magic
tech gf180mcuD
magscale 1 10
timestamp 1702237920
<< metal1 >>
rect 50082 329310 50094 329362
rect 50146 329359 50158 329362
rect 54786 329359 54798 329362
rect 50146 329313 54798 329359
rect 50146 329310 50158 329313
rect 54786 329310 54798 329313
rect 54850 329310 54862 329362
rect 109330 278910 109342 278962
rect 109394 278959 109406 278962
rect 113698 278959 113710 278962
rect 109394 278913 113710 278959
rect 109394 278910 109406 278913
rect 113698 278910 113710 278913
rect 113762 278910 113774 278962
rect 113586 270398 113598 270450
rect 113650 270447 113662 270450
rect 115826 270447 115838 270450
rect 113650 270401 115838 270447
rect 113650 270398 113662 270401
rect 115826 270398 115838 270401
rect 115890 270398 115902 270450
rect 43922 163102 43934 163154
rect 43986 163151 43998 163154
rect 45042 163151 45054 163154
rect 43986 163105 45054 163151
rect 43986 163102 43998 163105
rect 45042 163102 45054 163105
rect 45106 163102 45118 163154
rect 143714 161310 143726 161362
rect 143778 161359 143790 161362
rect 144386 161359 144398 161362
rect 143778 161313 144398 161359
rect 143778 161310 143790 161313
rect 144386 161310 144398 161313
rect 144450 161310 144462 161362
rect 373986 108334 373998 108386
rect 374050 108383 374062 108386
rect 374546 108383 374558 108386
rect 374050 108337 374558 108383
rect 374050 108334 374062 108337
rect 374546 108334 374558 108337
rect 374610 108334 374622 108386
rect 390450 45614 390462 45666
rect 390514 45663 390526 45666
rect 397842 45663 397854 45666
rect 390514 45617 397854 45663
rect 390514 45614 390526 45617
rect 397842 45614 397854 45617
rect 397906 45614 397918 45666
<< via1 >>
rect 50094 329310 50146 329362
rect 54798 329310 54850 329362
rect 109342 278910 109394 278962
rect 113710 278910 113762 278962
rect 113598 270398 113650 270450
rect 115838 270398 115890 270450
rect 43934 163102 43986 163154
rect 45054 163102 45106 163154
rect 143726 161310 143778 161362
rect 144398 161310 144450 161362
rect 373998 108334 374050 108386
rect 374558 108334 374610 108386
rect 390462 45614 390514 45666
rect 397854 45614 397906 45666
<< metal2 >>
rect 11032 595672 11256 597000
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 11032 595560 11284 595672
rect 11228 590772 11284 595560
rect 11228 590706 11284 590716
rect 33068 595560 33320 595672
rect 55132 595560 55384 595672
rect 77224 595672 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 143416 595672 143640 597000
rect 77224 595560 77476 595672
rect 99288 595560 99540 595672
rect 121352 595560 121604 595672
rect 33068 390628 33124 595560
rect 55132 511588 55188 595560
rect 77420 590884 77476 595560
rect 99484 590996 99540 595560
rect 99484 590930 99540 590940
rect 77420 590818 77476 590828
rect 118412 590884 118468 590894
rect 115052 588868 115108 588878
rect 55132 511522 55188 511532
rect 59612 548996 59668 549006
rect 33068 390562 33124 390572
rect 54572 509348 54628 509358
rect 1596 373716 1652 373726
rect 1484 308980 1540 308990
rect 28 304836 84 304846
rect 28 270340 84 304780
rect 28 270274 84 270284
rect 1484 164388 1540 308924
rect 1484 164322 1540 164332
rect 1596 148820 1652 373660
rect 25228 373268 25284 373278
rect 2492 368900 2548 368910
rect 2380 331044 2436 331054
rect 2268 317716 2324 317726
rect 2268 162148 2324 317660
rect 2380 162484 2436 330988
rect 2380 162418 2436 162428
rect 2268 162082 2324 162092
rect 1596 148754 1652 148764
rect 2492 148708 2548 368844
rect 23212 368116 23268 368126
rect 2940 364644 2996 364654
rect 2828 337204 2884 337214
rect 2716 337092 2772 337102
rect 2604 336980 2660 336990
rect 2604 313012 2660 336924
rect 2604 312946 2660 312956
rect 2716 310324 2772 337036
rect 2716 310258 2772 310268
rect 2716 305620 2772 305630
rect 2716 281428 2772 305564
rect 2828 304948 2884 337148
rect 2940 320404 2996 364588
rect 5628 363748 5684 363758
rect 4508 363636 4564 363646
rect 2940 320338 2996 320348
rect 3052 359604 3108 359614
rect 3052 315028 3108 359548
rect 3276 338548 3332 338558
rect 3052 314962 3108 314972
rect 3164 336868 3220 336878
rect 3164 312340 3220 336812
rect 3276 315700 3332 338492
rect 3276 315634 3332 315644
rect 4284 319060 4340 319070
rect 3164 312274 3220 312284
rect 3276 307636 3332 307646
rect 2828 304882 2884 304892
rect 2940 306292 2996 306302
rect 2716 281362 2772 281372
rect 2940 164276 2996 306236
rect 3276 194068 3332 307580
rect 3276 194002 3332 194012
rect 4172 273028 4228 273038
rect 2940 164210 2996 164220
rect 2492 148642 2548 148652
rect 4172 65268 4228 272972
rect 4284 268772 4340 319004
rect 4284 268706 4340 268716
rect 4508 162708 4564 363580
rect 4620 340228 4676 340238
rect 4620 313684 4676 340172
rect 4620 313618 4676 313628
rect 4732 338660 4788 338670
rect 4732 311668 4788 338604
rect 4732 311602 4788 311612
rect 4844 332724 4900 332734
rect 4732 309652 4788 309662
rect 4620 306964 4676 306974
rect 4620 280196 4676 306908
rect 4620 280130 4676 280140
rect 4732 279636 4788 309596
rect 4732 279570 4788 279580
rect 4844 164164 4900 332668
rect 5516 330372 5572 330382
rect 5516 320180 5572 330316
rect 5516 320114 5572 320124
rect 5628 304052 5684 363692
rect 18508 332724 18564 332734
rect 18508 329896 18564 332668
rect 19852 331044 19908 331054
rect 19852 329896 19908 330988
rect 23212 329896 23268 368060
rect 25228 329896 25284 373212
rect 27916 371364 27972 371374
rect 27916 329896 27972 371308
rect 37996 336084 38052 336094
rect 35980 335076 36036 335086
rect 28588 334852 28644 334862
rect 28588 329896 28644 334796
rect 35308 334516 35364 334526
rect 31948 333284 32004 333294
rect 31276 331604 31332 331614
rect 31052 330036 31108 330046
rect 31052 329924 31108 329980
rect 30632 329868 31108 329924
rect 31276 329896 31332 331548
rect 31948 329896 32004 333228
rect 35308 329896 35364 334460
rect 35980 329896 36036 335020
rect 36652 332948 36708 332958
rect 36652 329896 36708 332892
rect 37324 330708 37380 330718
rect 37324 329896 37380 330652
rect 37996 329896 38052 336028
rect 42700 333508 42756 333518
rect 38668 333396 38724 333406
rect 38668 329896 38724 333340
rect 41356 333060 41412 333070
rect 40012 332836 40068 332846
rect 40012 329896 40068 332780
rect 41356 329896 41412 333004
rect 42700 329896 42756 333452
rect 44716 333172 44772 333182
rect 43372 331716 43428 331726
rect 43372 329896 43428 331660
rect 44716 329896 44772 333116
rect 50092 329364 50148 329374
rect 49448 329362 50148 329364
rect 49448 329310 50094 329362
rect 50146 329310 50148 329362
rect 49448 329308 50148 329310
rect 50092 329298 50148 329308
rect 5628 303986 5684 303996
rect 54460 309204 54516 309214
rect 5516 283892 5572 283902
rect 5068 280532 5124 280542
rect 5068 280466 5124 280476
rect 5516 277844 5572 283836
rect 53452 281876 53508 281886
rect 13132 280644 13188 280654
rect 13132 280578 13188 280588
rect 23884 280644 23940 280654
rect 23884 280578 23940 280588
rect 40684 280644 40740 280654
rect 44716 280644 44772 280654
rect 40740 280588 41188 280644
rect 40684 280578 40740 280588
rect 25900 280532 25956 280542
rect 25900 280466 25956 280476
rect 26572 280532 26628 280542
rect 23212 280084 23268 280094
rect 5516 277778 5572 277788
rect 5740 276836 5796 280056
rect 6412 277060 6468 280056
rect 7084 277172 7140 280056
rect 7084 277106 7140 277116
rect 7756 277172 7812 280056
rect 7756 277106 7812 277116
rect 6412 276994 6468 277004
rect 5740 276770 5796 276780
rect 7980 276724 8036 276734
rect 7532 269668 7588 269678
rect 6748 264628 6804 264638
rect 6748 262836 6804 264572
rect 6748 262770 6804 262780
rect 4844 164098 4900 164108
rect 4508 162642 4564 162652
rect 4172 65202 4228 65212
rect 4284 158900 4340 158910
rect 4284 8820 4340 158844
rect 7532 121716 7588 269612
rect 7756 267988 7812 267998
rect 7644 266308 7700 266318
rect 7644 178052 7700 266252
rect 7756 220500 7812 267932
rect 7980 267092 8036 276668
rect 8428 274596 8484 280056
rect 9100 276388 9156 280056
rect 9100 276322 9156 276332
rect 9772 276276 9828 280056
rect 10444 276500 10500 280056
rect 11116 276948 11172 280056
rect 11116 276882 11172 276892
rect 10444 276434 10500 276444
rect 9772 276210 9828 276220
rect 11788 274708 11844 280056
rect 12460 278404 12516 280056
rect 12460 278338 12516 278348
rect 13804 276612 13860 280056
rect 13804 276546 13860 276556
rect 11788 274642 11844 274652
rect 8428 274530 8484 274540
rect 14476 270228 14532 280056
rect 15148 275492 15204 280056
rect 15148 275426 15204 275436
rect 14476 270162 14532 270172
rect 15820 269780 15876 280056
rect 16492 271908 16548 280056
rect 16828 278180 16884 278190
rect 16828 277060 16884 278124
rect 16828 276994 16884 277004
rect 16492 271842 16548 271852
rect 17164 271348 17220 280056
rect 17164 271282 17220 271292
rect 15820 269714 15876 269724
rect 7980 267026 8036 267036
rect 17836 266420 17892 280056
rect 18508 267876 18564 280056
rect 19180 273140 19236 280056
rect 19180 273074 19236 273084
rect 18508 267810 18564 267820
rect 17836 266354 17892 266364
rect 19852 264852 19908 280056
rect 20524 277956 20580 280056
rect 20524 277890 20580 277900
rect 21196 272804 21252 280056
rect 21868 274820 21924 280056
rect 21868 274754 21924 274764
rect 21196 272738 21252 272748
rect 22540 272692 22596 280056
rect 23212 280018 23268 280028
rect 24556 276724 24612 280056
rect 24556 276658 24612 276668
rect 22540 272626 22596 272636
rect 23436 276388 23492 276398
rect 23436 269892 23492 276332
rect 25228 273812 25284 280056
rect 26572 276612 26628 280476
rect 37996 280308 38052 280318
rect 37996 280242 38052 280252
rect 27244 279860 27300 280056
rect 27244 279794 27300 279804
rect 26908 278068 26964 278078
rect 26908 276836 26964 278012
rect 26908 276770 26964 276780
rect 26572 275604 26628 276556
rect 26572 275538 26628 275548
rect 25228 273746 25284 273756
rect 27916 272020 27972 280056
rect 28616 280028 29316 280084
rect 29260 276836 29316 280028
rect 29260 276770 29316 276780
rect 29932 276612 29988 280056
rect 31276 278628 31332 280056
rect 31276 278562 31332 278572
rect 29932 276546 29988 276556
rect 31948 273364 32004 280056
rect 34636 278852 34692 280056
rect 34636 278786 34692 278796
rect 35308 277172 35364 280056
rect 35308 277106 35364 277116
rect 31948 273298 32004 273308
rect 27916 271954 27972 271964
rect 35980 271796 36036 280056
rect 36680 280028 36932 280084
rect 36876 278516 36932 280028
rect 36876 275604 36932 278460
rect 38668 276164 38724 280056
rect 38668 276098 38724 276108
rect 36876 275538 36932 275548
rect 41132 275604 41188 280588
rect 44716 280578 44772 280588
rect 53452 280644 53508 281820
rect 53452 280578 53508 280588
rect 45388 280532 45444 280542
rect 45388 280466 45444 280476
rect 44044 280420 44100 280430
rect 44044 280354 44100 280364
rect 41132 275538 41188 275548
rect 35980 271730 36036 271740
rect 23436 269826 23492 269836
rect 42028 268436 42084 280056
rect 42700 278292 42756 280056
rect 42700 278226 42756 278236
rect 42028 268370 42084 268380
rect 43372 265188 43428 280056
rect 46060 266868 46116 280056
rect 46732 274932 46788 280056
rect 47404 276388 47460 280056
rect 48076 277060 48132 280056
rect 48748 277172 48804 280056
rect 48748 277106 48804 277116
rect 48076 276994 48132 277004
rect 47404 276322 47460 276332
rect 46732 274866 46788 274876
rect 49420 268324 49476 280056
rect 50092 277172 50148 280056
rect 54460 278740 54516 309148
rect 54572 280868 54628 509292
rect 54572 280802 54628 280812
rect 54684 416836 54740 416846
rect 54684 280420 54740 416780
rect 57036 361284 57092 361294
rect 55132 333396 55188 333406
rect 54796 329362 54852 329374
rect 54796 329310 54798 329362
rect 54850 329310 54852 329362
rect 54796 325948 54852 329310
rect 54796 325892 54964 325948
rect 54684 280354 54740 280364
rect 54908 280308 54964 325892
rect 55132 281540 55188 333340
rect 56700 333172 56756 333182
rect 56252 333060 56308 333070
rect 55132 281474 55188 281484
rect 56140 288148 56196 288158
rect 54908 280242 54964 280252
rect 54460 278674 54516 278684
rect 50092 277106 50148 277116
rect 56140 277172 56196 288092
rect 56140 277106 56196 277116
rect 56252 270116 56308 333004
rect 56476 332836 56532 332846
rect 56252 270050 56308 270060
rect 56364 319732 56420 319742
rect 56364 268548 56420 319676
rect 56476 273588 56532 332780
rect 56476 273522 56532 273532
rect 56588 312340 56644 312350
rect 56364 268482 56420 268492
rect 49420 268258 49476 268268
rect 56588 268212 56644 312284
rect 56700 275268 56756 333116
rect 56924 332836 56980 332846
rect 56812 302260 56868 302270
rect 56812 278908 56868 302204
rect 56924 280756 56980 332780
rect 57036 325108 57092 361228
rect 57932 339444 57988 339454
rect 57036 325042 57092 325052
rect 57148 327572 57204 327582
rect 57148 320964 57204 327516
rect 57932 326452 57988 339388
rect 57932 326386 57988 326396
rect 58716 331268 58772 331278
rect 57148 320898 57204 320908
rect 58156 324436 58212 324446
rect 58044 310324 58100 310334
rect 57932 307636 57988 307646
rect 57820 305620 57876 305630
rect 56924 280690 56980 280700
rect 57036 302932 57092 302942
rect 56812 278852 56980 278908
rect 56924 276388 56980 278852
rect 56924 276052 56980 276332
rect 57036 277060 57092 302876
rect 57820 280644 57876 305564
rect 57820 280578 57876 280588
rect 57036 276164 57092 277004
rect 57036 276098 57092 276108
rect 56924 275986 56980 275996
rect 56700 275202 56756 275212
rect 56588 268146 56644 268156
rect 46060 266802 46116 266812
rect 57932 265300 57988 307580
rect 58044 273476 58100 310268
rect 58156 281540 58212 324380
rect 58156 281474 58212 281484
rect 58268 322420 58324 322430
rect 58268 280532 58324 322364
rect 58716 314356 58772 331212
rect 58716 314290 58772 314300
rect 59500 319060 59556 319070
rect 58492 310996 58548 311006
rect 58268 280466 58324 280476
rect 58380 308308 58436 308318
rect 58380 275380 58436 308252
rect 58492 278628 58548 310940
rect 59388 302036 59444 302046
rect 58492 278562 58548 278572
rect 58604 289492 58660 289502
rect 58380 275314 58436 275324
rect 58044 273410 58100 273420
rect 58604 269556 58660 289436
rect 58716 284788 58772 284798
rect 58716 277732 58772 284732
rect 58716 277666 58772 277676
rect 58604 269490 58660 269500
rect 59388 266644 59444 301980
rect 59500 275156 59556 319004
rect 59612 281876 59668 548940
rect 60620 522564 60676 522574
rect 59836 378868 59892 378878
rect 59612 281810 59668 281820
rect 59724 333620 59780 333630
rect 59724 278516 59780 333564
rect 59836 288820 59892 378812
rect 59836 288754 59892 288764
rect 60060 332948 60116 332958
rect 60060 281764 60116 332892
rect 60620 327572 60676 522508
rect 113372 502516 113428 502526
rect 111692 460180 111748 460190
rect 88956 383908 89012 383918
rect 86492 364868 86548 364878
rect 78204 359268 78260 359278
rect 76188 349188 76244 349198
rect 70364 333844 70420 333854
rect 70364 333060 70420 333788
rect 73500 333732 73556 333742
rect 72828 333508 72884 333518
rect 70140 333004 70364 333060
rect 69468 332724 69524 332734
rect 69468 329896 69524 332668
rect 70140 329896 70196 333004
rect 70364 332994 70420 333004
rect 70476 333172 70532 333182
rect 70476 332724 70532 333116
rect 70476 332658 70532 332668
rect 72156 332948 72212 332958
rect 72156 329896 72212 332892
rect 72828 329896 72884 333452
rect 73500 330260 73556 333676
rect 75516 333620 75572 333630
rect 73500 329896 73556 330204
rect 74844 333396 74900 333406
rect 74844 332724 74900 333340
rect 74844 329896 74900 332668
rect 75516 329924 75572 333564
rect 76188 329896 76244 349132
rect 77532 332724 77588 332734
rect 76860 329924 76916 329934
rect 75516 329858 75572 329868
rect 77532 329896 77588 332668
rect 78204 329896 78260 359212
rect 86492 349468 86548 364812
rect 86492 349412 86996 349468
rect 84924 333844 84980 333854
rect 82908 333172 82964 333182
rect 78876 332948 78932 332958
rect 78876 329896 78932 332892
rect 79548 331268 79604 331278
rect 79548 329896 79604 331212
rect 82908 329896 82964 333116
rect 83580 331940 83636 331950
rect 83580 329896 83636 331884
rect 84252 331380 84308 331390
rect 84252 329896 84308 331324
rect 84924 329896 84980 333788
rect 86940 332836 86996 349412
rect 88284 333620 88340 333630
rect 86940 329896 86996 332780
rect 87612 333508 87668 333518
rect 87612 329896 87668 333452
rect 88284 329896 88340 333564
rect 88956 329896 89012 383852
rect 110012 375508 110068 375518
rect 93660 372148 93716 372158
rect 92988 331492 93044 331502
rect 92988 329896 93044 331436
rect 93660 329896 93716 372092
rect 110012 337708 110068 375452
rect 109788 337652 110068 337708
rect 110236 375508 110292 375518
rect 102396 334964 102452 334974
rect 101052 334404 101108 334414
rect 95004 332052 95060 332062
rect 95004 329896 95060 331996
rect 100380 331268 100436 331278
rect 100380 329896 100436 331212
rect 101052 329896 101108 334348
rect 101724 332836 101780 332846
rect 101724 329896 101780 332780
rect 102396 329896 102452 334908
rect 103740 331156 103796 331166
rect 103068 330260 103124 330270
rect 103068 329896 103124 330204
rect 103740 329896 103796 331100
rect 105084 331044 105140 331054
rect 104412 330484 104468 330494
rect 104412 329896 104468 330428
rect 105084 329896 105140 330988
rect 105756 330148 105812 330158
rect 105756 329896 105812 330092
rect 76860 329858 76916 329868
rect 60620 327506 60676 327516
rect 109788 320908 109844 337652
rect 109900 336084 109956 336094
rect 109900 332668 109956 336028
rect 109900 332612 110180 332668
rect 109788 320852 110068 320908
rect 60284 320180 60340 320190
rect 60060 281698 60116 281708
rect 60172 313012 60228 313022
rect 59724 278450 59780 278460
rect 60060 278180 60116 280056
rect 60060 276948 60116 278124
rect 60060 276882 60116 276892
rect 59500 275090 59556 275100
rect 59388 266578 59444 266588
rect 57932 265234 57988 265244
rect 43372 265122 43428 265132
rect 60172 265076 60228 312956
rect 60284 275044 60340 320124
rect 60396 315028 60452 315038
rect 60396 280420 60452 314972
rect 60396 280354 60452 280364
rect 60508 311668 60564 311678
rect 60284 274978 60340 274988
rect 60508 266756 60564 311612
rect 109340 303156 109396 303166
rect 70140 280756 70196 280766
rect 70140 280690 70196 280700
rect 74844 280756 74900 280766
rect 74844 280690 74900 280700
rect 87612 280756 87668 280766
rect 87612 280690 87668 280700
rect 89628 280756 89684 280766
rect 89628 280690 89684 280700
rect 74172 280084 74228 280094
rect 60732 276276 60788 280056
rect 60732 273252 60788 276220
rect 61404 277172 61460 280056
rect 61404 275604 61460 277116
rect 62076 278292 62132 280056
rect 62076 276724 62132 278236
rect 62076 276658 62132 276668
rect 62748 277956 62804 280056
rect 62748 276500 62804 277900
rect 63420 277060 63476 280056
rect 63420 276994 63476 277004
rect 62748 276434 62804 276444
rect 64092 276724 64148 280056
rect 61404 275538 61460 275548
rect 63868 276388 63924 276398
rect 63868 273812 63924 276332
rect 64092 275604 64148 276668
rect 64764 276388 64820 280056
rect 65436 277172 65492 280056
rect 65436 277106 65492 277116
rect 64764 276322 64820 276332
rect 64092 275538 64148 275548
rect 65548 275604 65604 275614
rect 65548 274708 65604 275548
rect 65548 274642 65604 274652
rect 63868 273746 63924 273756
rect 60732 273186 60788 273196
rect 66108 273140 66164 280056
rect 66780 275604 66836 280056
rect 67452 276948 67508 280056
rect 67452 276882 67508 276892
rect 68124 276500 68180 280056
rect 68796 278908 68852 280056
rect 68124 276434 68180 276444
rect 68684 278852 68852 278908
rect 66780 275538 66836 275548
rect 66108 273074 66164 273084
rect 68684 274708 68740 278852
rect 69468 276612 69524 280056
rect 70812 279860 70868 280056
rect 71512 280028 71988 280084
rect 70812 279794 70868 279804
rect 69468 276546 69524 276556
rect 71932 277172 71988 280028
rect 68684 269892 68740 274652
rect 68796 276500 68852 276510
rect 68796 274596 68852 276444
rect 68796 274530 68852 274540
rect 71932 271236 71988 277116
rect 72156 274596 72212 280056
rect 72828 278852 72884 280056
rect 73500 278908 73556 280056
rect 72828 278068 72884 278796
rect 72828 278002 72884 278012
rect 73052 278852 73556 278908
rect 72156 274530 72212 274540
rect 73052 276388 73108 278852
rect 74172 278516 74228 280028
rect 75516 280084 75572 280094
rect 77532 280084 77588 280094
rect 75516 280018 75572 280028
rect 74172 278450 74228 278460
rect 76188 279748 76244 280056
rect 71932 271170 71988 271180
rect 68684 269826 68740 269836
rect 60508 266690 60564 266700
rect 60172 265010 60228 265020
rect 19852 264786 19908 264796
rect 73052 264740 73108 276332
rect 75628 277172 75684 277182
rect 75628 271348 75684 277116
rect 76188 276836 76244 279692
rect 76860 277172 76916 280056
rect 77532 280018 77588 280028
rect 76860 277106 76916 277116
rect 78204 278404 78260 280056
rect 76188 276770 76244 276780
rect 78204 276388 78260 278348
rect 78204 276322 78260 276332
rect 75628 271282 75684 271292
rect 78876 271348 78932 280056
rect 79548 276724 79604 280056
rect 79548 276658 79604 276668
rect 80220 276052 80276 280056
rect 80892 276836 80948 280056
rect 80892 276500 80948 276780
rect 80892 276434 80948 276444
rect 81452 280028 81592 280084
rect 81676 280056 82264 280084
rect 81676 280028 82292 280056
rect 81452 277060 81508 280028
rect 81676 279972 81732 280028
rect 81676 279906 81732 279916
rect 82236 278404 82292 280028
rect 82236 278338 82292 278348
rect 80220 275986 80276 275996
rect 78876 271282 78932 271292
rect 81452 266420 81508 277004
rect 82236 276836 82292 276846
rect 82236 268100 82292 276780
rect 82908 276724 82964 280056
rect 83580 277172 83636 280056
rect 83580 277106 83636 277116
rect 84252 277060 84308 280056
rect 84252 276994 84308 277004
rect 84924 276948 84980 280056
rect 84924 276882 84980 276892
rect 82908 276658 82964 276668
rect 85596 273700 85652 280056
rect 85596 273634 85652 273644
rect 86268 273140 86324 280056
rect 86940 274820 86996 280056
rect 88284 276500 88340 280056
rect 88956 276612 89012 280056
rect 90300 277172 90356 280056
rect 90300 277106 90356 277116
rect 88956 276546 89012 276556
rect 88284 276434 88340 276444
rect 90972 276164 91028 280056
rect 90972 276098 91028 276108
rect 92988 276164 93044 280056
rect 93660 276948 93716 280056
rect 93660 276882 93716 276892
rect 94332 276948 94388 280056
rect 94332 276882 94388 276892
rect 92988 276098 93044 276108
rect 95676 276052 95732 280056
rect 97692 276836 97748 280056
rect 101052 277172 101108 280056
rect 101052 277106 101108 277116
rect 97692 276770 97748 276780
rect 95676 275986 95732 275996
rect 86940 274754 86996 274764
rect 100828 275604 100884 275614
rect 100828 273252 100884 275548
rect 101724 275604 101780 280056
rect 109340 278962 109396 303100
rect 109340 278910 109342 278962
rect 109394 278910 109396 278962
rect 109340 278908 109396 278910
rect 109228 278852 109396 278908
rect 109564 297332 109620 297342
rect 109564 282100 109620 297276
rect 109228 278786 109284 278796
rect 109564 278404 109620 282044
rect 109564 278338 109620 278348
rect 101724 275538 101780 275548
rect 106876 278068 106932 278078
rect 100828 273186 100884 273196
rect 86268 273074 86324 273084
rect 104972 273140 105028 273150
rect 82236 268034 82292 268044
rect 99932 269780 99988 269790
rect 81452 266354 81508 266364
rect 73052 264674 73108 264684
rect 7756 220434 7812 220444
rect 7644 177986 7700 177996
rect 10892 194068 10948 194078
rect 10892 162820 10948 194012
rect 20636 165732 20692 165742
rect 20440 165676 20636 165732
rect 20636 165666 20692 165676
rect 26684 165732 26740 165742
rect 26684 165666 26740 165676
rect 28028 165732 28084 165742
rect 39676 165732 39732 165742
rect 71708 165732 71764 165742
rect 38808 165676 39676 165732
rect 71512 165676 71708 165732
rect 28028 165666 28084 165676
rect 39676 165666 39732 165676
rect 71708 165666 71764 165676
rect 82236 165732 82292 165742
rect 82236 165666 82292 165676
rect 84028 165732 84084 165742
rect 84028 165666 84084 165676
rect 83804 165620 83860 165630
rect 83608 165564 83804 165620
rect 83804 165554 83860 165564
rect 45080 165116 45332 165172
rect 20860 162932 20916 165032
rect 20860 162866 20916 162876
rect 10892 162754 10948 162764
rect 21308 162596 21364 165032
rect 26236 162708 26292 165032
rect 27132 162932 27188 165032
rect 27608 165004 27860 165060
rect 27132 162866 27188 162876
rect 26236 162642 26292 162652
rect 21308 162530 21364 162540
rect 17948 159684 18004 159694
rect 17948 144900 18004 159628
rect 27804 159460 27860 165004
rect 28476 161140 28532 165032
rect 37884 164500 37940 165032
rect 37884 164434 37940 164444
rect 38332 164052 38388 165032
rect 43736 165004 43988 165060
rect 38332 163986 38388 163996
rect 43932 163154 43988 165004
rect 43932 163102 43934 163154
rect 43986 163102 43988 163154
rect 43932 163090 43988 163102
rect 44156 164164 44212 165032
rect 44156 163044 44212 164108
rect 44156 162978 44212 162988
rect 44380 165004 44632 165060
rect 44380 162484 44436 165004
rect 45052 163154 45108 163166
rect 45052 163102 45054 163154
rect 45106 163102 45108 163154
rect 44380 162418 44436 162428
rect 44940 163044 44996 163054
rect 28476 161074 28532 161084
rect 44828 162148 44884 162158
rect 27804 159394 27860 159404
rect 43484 159012 43540 159022
rect 38108 158788 38164 158798
rect 26460 158004 26516 158014
rect 18396 155428 18452 155438
rect 18396 144900 18452 155372
rect 17864 144844 18004 144900
rect 18312 144844 18452 144900
rect 18732 148932 18788 148942
rect 18732 144872 18788 148876
rect 25900 148820 25956 148830
rect 25900 144872 25956 148764
rect 26460 144900 26516 157948
rect 27356 157108 27412 157118
rect 26376 144844 26516 144900
rect 26796 150500 26852 150510
rect 26796 144872 26852 150444
rect 27356 144900 27412 157052
rect 27804 155540 27860 155550
rect 27804 144900 27860 155484
rect 37548 148932 37604 148942
rect 27272 144844 27412 144900
rect 27720 144844 27860 144900
rect 28140 148708 28196 148718
rect 28140 144872 28196 148652
rect 37548 144872 37604 148876
rect 38108 144900 38164 158732
rect 38024 144844 38164 144900
rect 38444 152852 38500 152862
rect 38444 144872 38500 152796
rect 43484 144900 43540 158956
rect 43932 157444 43988 157454
rect 43932 144900 43988 157388
rect 44380 155540 44436 155550
rect 44380 144900 44436 155484
rect 44828 144900 44884 162092
rect 44940 157332 44996 162988
rect 44940 157266 44996 157276
rect 45052 152068 45108 163102
rect 45276 162820 45332 165116
rect 45500 164276 45556 165032
rect 45976 165004 46228 165060
rect 53144 165004 53732 165060
rect 45500 163604 45556 164220
rect 45500 163538 45556 163548
rect 46172 164388 46228 165004
rect 45332 162764 45444 162820
rect 45276 162754 45332 162764
rect 45388 155652 45444 162764
rect 45388 155586 45444 155596
rect 45052 152002 45108 152012
rect 46172 148820 46228 164332
rect 46172 148754 46228 148764
rect 46396 163604 46452 163614
rect 46396 148708 46452 163548
rect 47852 162484 47908 162494
rect 46396 148642 46452 148652
rect 46620 157556 46676 157566
rect 43400 144844 43540 144900
rect 43848 144844 43988 144900
rect 44296 144844 44436 144900
rect 44744 144844 44884 144900
rect 45164 147924 45220 147934
rect 45164 144872 45220 147868
rect 46620 147924 46676 157500
rect 47852 152180 47908 162428
rect 53676 161028 53732 165004
rect 53676 160962 53732 160972
rect 63980 165004 64792 165060
rect 63980 163044 64036 165004
rect 63980 157556 64036 162988
rect 63980 157490 64036 157500
rect 64988 162260 65044 162270
rect 64988 157444 65044 162204
rect 65212 162148 65268 165032
rect 65212 162082 65268 162092
rect 65660 161476 65716 165032
rect 66108 162260 66164 165032
rect 66108 162194 66164 162204
rect 66332 165004 66584 165060
rect 65548 160468 65604 160478
rect 65548 159012 65604 160412
rect 65548 158946 65604 158956
rect 64988 157378 65044 157388
rect 47852 152114 47908 152124
rect 56924 157220 56980 157230
rect 46620 147858 46676 147868
rect 56924 144900 56980 157164
rect 64876 155652 64932 155662
rect 64876 149268 64932 155596
rect 65660 155540 65716 161420
rect 66332 160468 66388 165004
rect 71932 162484 71988 165032
rect 72380 163940 72436 165032
rect 72380 163874 72436 163884
rect 71932 162418 71988 162428
rect 81788 162372 81844 165032
rect 82684 162708 82740 165032
rect 82684 162642 82740 162652
rect 83132 162596 83188 165032
rect 91196 162932 91252 165032
rect 91196 162866 91252 162876
rect 91644 162820 91700 165032
rect 92092 164612 92148 165032
rect 92092 164546 92148 164556
rect 99932 162932 99988 269724
rect 99932 162866 99988 162876
rect 91644 162754 91700 162764
rect 83132 162530 83188 162540
rect 104972 162596 105028 273084
rect 105196 269892 105252 269902
rect 105196 162820 105252 269836
rect 105196 162754 105252 162764
rect 104972 162530 105028 162540
rect 106876 162484 106932 278012
rect 108332 276836 108388 276846
rect 108332 273364 108388 276780
rect 108332 273298 108388 273308
rect 110012 273364 110068 320852
rect 110124 305060 110180 332612
rect 110124 304994 110180 305004
rect 110236 277172 110292 375452
rect 110796 369908 110852 369918
rect 110684 362180 110740 362190
rect 110684 337092 110740 362124
rect 110684 336084 110740 337036
rect 110684 336018 110740 336028
rect 110796 335188 110852 369852
rect 110796 334628 110852 335132
rect 110796 334562 110852 334572
rect 110348 331268 110404 331278
rect 110348 301028 110404 331212
rect 110572 330148 110628 330158
rect 110348 300962 110404 300972
rect 110460 329588 110516 329598
rect 110236 277106 110292 277116
rect 110460 276948 110516 329532
rect 110572 309092 110628 330092
rect 110572 309026 110628 309036
rect 110908 304948 110964 304958
rect 110908 284564 110964 304892
rect 111132 284564 111188 284574
rect 110908 284508 111132 284564
rect 111132 284498 111188 284508
rect 110460 276882 110516 276892
rect 110012 273298 110068 273308
rect 111692 272132 111748 460124
rect 111804 389620 111860 389630
rect 111804 278404 111860 389564
rect 111916 341348 111972 341358
rect 111916 279860 111972 341292
rect 112252 336084 112308 336094
rect 112140 331044 112196 331054
rect 112028 330484 112084 330494
rect 112028 294308 112084 330428
rect 112140 302148 112196 330988
rect 112252 310772 112308 336028
rect 112252 310706 112308 310716
rect 112364 334628 112420 334638
rect 112364 308420 112420 334572
rect 112364 308354 112420 308364
rect 112588 317492 112644 317502
rect 112588 307412 112644 317436
rect 112588 307346 112644 307356
rect 112140 302082 112196 302092
rect 112028 294242 112084 294252
rect 112700 292180 112756 292190
rect 112700 290724 112756 292124
rect 111916 279794 111972 279804
rect 112588 288820 112644 288830
rect 112588 279076 112644 288764
rect 112700 279748 112756 290668
rect 112700 279682 112756 279692
rect 112588 279010 112644 279020
rect 111804 278338 111860 278348
rect 113372 273812 113428 502460
rect 113708 385588 113764 385598
rect 113484 374836 113540 374846
rect 113484 304948 113540 374780
rect 113484 304882 113540 304892
rect 113596 335748 113652 335758
rect 113372 273746 113428 273756
rect 113484 278964 113540 278974
rect 111692 272066 111748 272076
rect 113484 270452 113540 278908
rect 113596 277060 113652 335692
rect 113708 326452 113764 385532
rect 113708 326386 113764 326396
rect 113820 334404 113876 334414
rect 113820 287588 113876 334348
rect 114940 331492 114996 331502
rect 114268 331044 114324 331054
rect 114268 310996 114324 330988
rect 114940 317828 114996 331436
rect 115052 327124 115108 588812
rect 115836 372260 115892 372270
rect 115724 370020 115780 370030
rect 115612 368676 115668 368686
rect 115500 364756 115556 364766
rect 115052 327058 115108 327068
rect 115164 357028 115220 357038
rect 114940 317762 114996 317772
rect 115052 324212 115108 324222
rect 114268 310930 114324 310940
rect 113820 287522 113876 287532
rect 114044 279076 114100 279086
rect 113596 276994 113652 277004
rect 113708 278962 113764 278974
rect 113708 278910 113710 278962
rect 113762 278910 113764 278962
rect 113596 270452 113652 270462
rect 113484 270450 113652 270452
rect 113484 270398 113598 270450
rect 113650 270398 113652 270450
rect 113484 270396 113652 270398
rect 113596 270386 113652 270396
rect 113708 266196 113764 278910
rect 114044 276612 114100 279020
rect 115052 278180 115108 324156
rect 115052 278114 115108 278124
rect 114044 276546 114100 276556
rect 115164 274820 115220 356972
rect 115500 338660 115556 364700
rect 115612 340228 115668 368620
rect 115612 340162 115668 340172
rect 115500 338594 115556 338604
rect 115724 336980 115780 369964
rect 115724 336084 115780 336924
rect 115724 336018 115780 336028
rect 115164 274754 115220 274764
rect 115276 334628 115332 334638
rect 115276 273700 115332 334572
rect 115388 333284 115444 333294
rect 115388 279524 115444 333228
rect 115724 332836 115780 332846
rect 115612 331380 115668 331390
rect 115500 326788 115556 326798
rect 115500 312564 115556 326732
rect 115612 318948 115668 331324
rect 115724 324212 115780 332780
rect 115724 324146 115780 324156
rect 115612 318882 115668 318892
rect 115500 312498 115556 312508
rect 115500 307412 115556 307422
rect 115500 284228 115556 307356
rect 115836 300916 115892 372204
rect 117516 366996 117572 367006
rect 117516 339332 117572 366940
rect 117068 339108 117124 339118
rect 116732 336868 116788 336878
rect 116396 332052 116452 332062
rect 116396 308868 116452 331996
rect 116396 308802 116452 308812
rect 116620 331156 116676 331166
rect 116620 307748 116676 331100
rect 116620 307682 116676 307692
rect 115836 300850 115892 300860
rect 115500 284162 115556 284172
rect 115388 279458 115444 279468
rect 115276 273634 115332 273644
rect 116732 271348 116788 336812
rect 116956 333508 117012 333518
rect 116844 331940 116900 331950
rect 116844 280868 116900 331884
rect 116956 282884 117012 333452
rect 116956 282818 117012 282828
rect 117068 281652 117124 339052
rect 117516 338548 117572 339276
rect 117516 338482 117572 338492
rect 117292 337988 117348 337998
rect 117180 330260 117236 330270
rect 117180 285348 117236 330204
rect 117180 285282 117236 285292
rect 117292 281764 117348 337932
rect 117404 324212 117460 324222
rect 117404 286468 117460 324156
rect 117404 286402 117460 286412
rect 117516 309092 117572 309102
rect 117516 283108 117572 309036
rect 117516 283042 117572 283052
rect 117292 281698 117348 281708
rect 117068 281586 117124 281596
rect 116844 280802 116900 280812
rect 116732 271282 116788 271292
rect 118412 271236 118468 590828
rect 121548 590772 121604 595560
rect 121548 590706 121604 590716
rect 143388 595560 143640 595672
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 209608 595672 209832 597000
rect 231672 595672 231896 597000
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 319928 595672 320152 597000
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 386120 595672 386344 597000
rect 165480 595560 165732 595672
rect 118524 417844 118580 417854
rect 118524 273700 118580 417788
rect 143388 380548 143444 595560
rect 165676 590884 165732 595560
rect 165676 590818 165732 590828
rect 187516 595560 187768 595672
rect 209580 595560 209832 595672
rect 231644 595560 231896 595672
rect 253708 595560 253960 595672
rect 275772 595560 276024 595672
rect 297836 595560 298088 595672
rect 319900 595560 320152 595672
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386092 595560 386344 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 452312 595672 452536 597000
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 518504 595672 518728 597000
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 584696 595672 584920 597000
rect 430220 595560 430472 595672
rect 452284 595560 452536 595672
rect 474348 595560 474600 595672
rect 496412 595560 496664 595672
rect 518476 595560 518728 595672
rect 540540 595560 540792 595672
rect 562604 595560 562856 595672
rect 584668 595560 584920 595672
rect 143388 380482 143444 380492
rect 174188 376404 174244 376414
rect 167468 374948 167524 374958
rect 125132 374724 125188 374734
rect 119196 366436 119252 366446
rect 118636 361396 118692 361406
rect 118636 277956 118692 361340
rect 118860 347284 118916 347294
rect 118636 277890 118692 277900
rect 118748 336084 118804 336094
rect 118748 276276 118804 336028
rect 118860 278516 118916 347228
rect 118860 278450 118916 278460
rect 118972 331268 119028 331278
rect 118748 276210 118804 276220
rect 118972 276164 119028 331212
rect 119196 330372 119252 366380
rect 125132 364868 125188 374668
rect 149324 372036 149380 372046
rect 147980 371700 148036 371710
rect 133868 371588 133924 371598
rect 131180 368340 131236 368350
rect 125132 359912 125188 364812
rect 126476 367220 126532 367230
rect 125804 361284 125860 361294
rect 125804 359912 125860 361228
rect 126476 359912 126532 367164
rect 127820 363188 127876 363198
rect 127148 361396 127204 361406
rect 127148 359912 127204 361340
rect 127820 359912 127876 363132
rect 129164 363076 129220 363086
rect 128492 361508 128548 361518
rect 128492 359912 128548 361452
rect 129164 359912 129220 363020
rect 129836 360164 129892 360174
rect 129836 359912 129892 360108
rect 131180 359912 131236 368284
rect 132524 365092 132580 365102
rect 132300 360052 132356 360062
rect 132300 359940 132356 359996
rect 131880 359884 132356 359940
rect 132524 359912 132580 365036
rect 133196 359940 133252 359950
rect 133868 359912 133924 371532
rect 139244 371476 139300 371486
rect 137228 368452 137284 368462
rect 135884 368228 135940 368238
rect 134540 360276 134596 360286
rect 134540 359912 134596 360220
rect 135884 359912 135940 368172
rect 136556 361732 136612 361742
rect 136556 359912 136612 361676
rect 137228 359912 137284 368396
rect 138572 367108 138628 367118
rect 137900 364868 137956 364878
rect 137900 359912 137956 364812
rect 138572 359912 138628 367052
rect 139244 359912 139300 371420
rect 141932 370356 141988 370366
rect 139916 366548 139972 366558
rect 139916 359912 139972 366492
rect 140588 364980 140644 364990
rect 140588 359912 140644 364924
rect 141260 360500 141316 360510
rect 141260 359912 141316 360444
rect 141932 359912 141988 370300
rect 143948 369796 144004 369806
rect 143276 363972 143332 363982
rect 142604 361956 142660 361966
rect 142604 359912 142660 361900
rect 143276 359912 143332 363916
rect 143612 363188 143668 363198
rect 143612 362068 143668 363132
rect 143612 362002 143668 362012
rect 143948 359912 144004 369740
rect 144620 368564 144676 368574
rect 144620 359912 144676 368508
rect 146636 366772 146692 366782
rect 145964 363300 146020 363310
rect 145292 363188 145348 363198
rect 145292 359912 145348 363132
rect 145964 359912 146020 363244
rect 146636 359912 146692 366716
rect 147308 366660 147364 366670
rect 147308 359912 147364 366604
rect 147980 359912 148036 371644
rect 148652 361844 148708 361854
rect 148652 359912 148708 361788
rect 149324 359912 149380 371980
rect 162092 370020 162148 370030
rect 160076 369908 160132 369918
rect 149996 368788 150052 368798
rect 149996 359912 150052 368732
rect 159404 368676 159460 368686
rect 152684 366884 152740 366894
rect 151228 363076 151284 363086
rect 150668 361620 150724 361630
rect 150668 359912 150724 361564
rect 151228 360388 151284 363020
rect 151228 360322 151284 360332
rect 151340 362964 151396 362974
rect 151340 359912 151396 362908
rect 152012 362964 152068 362974
rect 152012 359912 152068 362908
rect 152684 359912 152740 366828
rect 154028 365428 154084 365438
rect 153356 362180 153412 362190
rect 153356 359912 153412 362124
rect 154028 359912 154084 365372
rect 156716 365316 156772 365326
rect 155372 365204 155428 365214
rect 154700 363524 154756 363534
rect 154700 359912 154756 363468
rect 155372 359912 155428 365148
rect 156156 362964 156212 362974
rect 155708 362180 155764 362190
rect 155708 361956 155764 362124
rect 155708 361890 155764 361900
rect 156156 359940 156212 362908
rect 156072 359884 156212 359940
rect 156716 359912 156772 365260
rect 158732 364756 158788 364766
rect 157836 362964 157892 362974
rect 157836 359940 157892 362908
rect 157416 359884 157892 359940
rect 158060 362180 158116 362190
rect 158060 359912 158116 362124
rect 158732 359912 158788 364700
rect 159404 359912 159460 368620
rect 160076 359912 160132 369852
rect 160748 363076 160804 363086
rect 160748 359912 160804 363020
rect 161420 361172 161476 361182
rect 133196 359874 133252 359884
rect 135212 359828 135268 359838
rect 135212 359762 135268 359772
rect 130508 359716 130564 359726
rect 130508 359650 130564 359660
rect 161420 359604 161476 361116
rect 162092 359912 162148 369964
rect 166796 368676 166852 368686
rect 165452 366996 165508 367006
rect 162764 366436 162820 366446
rect 162764 359912 162820 366380
rect 164108 363412 164164 363422
rect 163436 362180 163492 362190
rect 163436 359912 163492 362124
rect 164108 359912 164164 363356
rect 164668 363076 164724 363086
rect 164668 359940 164724 363020
rect 164668 359884 164808 359940
rect 165452 359912 165508 366940
rect 166124 364644 166180 364654
rect 161420 359538 161476 359548
rect 166124 359604 166180 364588
rect 166796 359912 166852 368620
rect 167468 359912 167524 374892
rect 168812 373268 168868 373278
rect 168140 370020 168196 370030
rect 168140 359912 168196 369964
rect 168812 362180 168868 373212
rect 169708 371924 169764 371934
rect 169708 371364 169764 371868
rect 168812 359912 168868 362124
rect 169484 369908 169540 369918
rect 169484 368116 169540 369852
rect 169484 359912 169540 368060
rect 169708 361228 169764 371308
rect 171500 371812 171556 371822
rect 170828 370132 170884 370142
rect 169708 361172 170212 361228
rect 170156 359912 170212 361172
rect 170828 359912 170884 370076
rect 171500 359912 171556 371756
rect 172172 366996 172228 367006
rect 172172 359912 172228 366940
rect 172844 363748 172900 363758
rect 172844 359912 172900 363692
rect 174188 359912 174244 376348
rect 174860 374836 174916 374846
rect 174860 359912 174916 374780
rect 187516 373828 187572 595560
rect 200732 590884 200788 590894
rect 200732 390740 200788 590828
rect 200732 390674 200788 390684
rect 187516 373762 187572 373772
rect 199948 374948 200004 374958
rect 176876 373604 176932 373614
rect 176204 372260 176260 372270
rect 175532 371364 175588 371374
rect 175532 359912 175588 371308
rect 176204 359912 176260 372204
rect 176876 359912 176932 373548
rect 180908 373492 180964 373502
rect 179564 373380 179620 373390
rect 177548 373268 177604 373278
rect 177548 359912 177604 373212
rect 178220 370244 178276 370254
rect 178220 359912 178276 370188
rect 178892 364644 178948 364654
rect 178892 359912 178948 364588
rect 179564 359912 179620 373324
rect 180236 366436 180292 366446
rect 180236 359912 180292 366380
rect 180908 359912 180964 373436
rect 181580 373044 181636 373054
rect 181580 359912 181636 372988
rect 199276 371364 199332 371374
rect 184268 369684 184324 369694
rect 183596 368116 183652 368126
rect 182924 363076 182980 363086
rect 182924 359912 182980 363020
rect 183596 359912 183652 368060
rect 184268 359912 184324 369628
rect 188972 368004 189028 368014
rect 186284 366324 186340 366334
rect 185612 364756 185668 364766
rect 184940 360612 184996 360622
rect 184940 359912 184996 360556
rect 185612 359912 185668 364700
rect 186284 359912 186340 366268
rect 187628 363412 187684 363422
rect 187628 359912 187684 363356
rect 188300 362964 188356 362974
rect 188300 359912 188356 362908
rect 188972 359912 189028 367948
rect 192556 360724 192612 360734
rect 192556 360164 192612 360668
rect 192556 360098 192612 360108
rect 192780 360164 192836 360174
rect 192780 359940 192836 360108
rect 192360 359884 192836 359940
rect 166124 359538 166180 359548
rect 173516 359604 173572 359614
rect 190764 359604 190820 359614
rect 190344 359548 190764 359604
rect 173516 359538 173572 359548
rect 190764 359538 190820 359548
rect 190988 359604 191044 359614
rect 192108 359604 192164 359614
rect 194012 359604 194068 359614
rect 195692 359604 195748 359614
rect 191688 359548 192108 359604
rect 193704 359548 194012 359604
rect 195048 359548 195692 359604
rect 190988 359538 191044 359548
rect 192108 359538 192164 359548
rect 194012 359538 194068 359548
rect 195692 359538 195748 359548
rect 182252 359492 182308 359502
rect 182252 359426 182308 359436
rect 186956 359492 187012 359502
rect 186956 359426 187012 359436
rect 189644 359492 189700 359502
rect 189644 359426 189700 359436
rect 193004 359492 193060 359502
rect 193004 359426 193060 359436
rect 194348 359492 194404 359502
rect 194348 359426 194404 359436
rect 120204 337540 120260 337550
rect 119196 329364 119252 330316
rect 119196 329298 119252 329308
rect 119980 334964 120036 334974
rect 119980 297108 120036 334908
rect 119980 297042 120036 297052
rect 120092 331716 120148 331726
rect 118972 276098 119028 276108
rect 119084 290724 119140 290734
rect 120092 290668 120148 331660
rect 118524 273634 118580 273644
rect 118412 271170 118468 271180
rect 113708 266130 113764 266140
rect 115836 270450 115892 270462
rect 115836 270398 115838 270450
rect 115890 270398 115892 270450
rect 115836 265412 115892 270398
rect 119084 268660 119140 290668
rect 119868 290612 120148 290668
rect 119868 281876 119924 290612
rect 119868 281810 119924 281820
rect 119980 282996 120036 283006
rect 119196 281540 119252 281550
rect 119196 279860 119252 281484
rect 119196 279794 119252 279804
rect 119980 279412 120036 282940
rect 119980 279346 120036 279356
rect 119084 268594 119140 268604
rect 119196 276724 119252 276734
rect 115836 265346 115892 265356
rect 119196 264964 119252 276668
rect 120204 274596 120260 337484
rect 120316 335076 120372 335086
rect 120316 276948 120372 335020
rect 120540 330708 120596 330718
rect 120540 277060 120596 330652
rect 121548 280756 121604 280766
rect 121548 280690 121604 280700
rect 141708 280644 141764 280654
rect 141708 280578 141764 280588
rect 127708 280532 127764 280542
rect 133644 280532 133700 280542
rect 127764 280476 128296 280532
rect 127708 280466 127764 280476
rect 133644 280466 133700 280476
rect 139692 280532 139748 280542
rect 139692 280466 139748 280476
rect 141036 280532 141092 280542
rect 141036 280466 141092 280476
rect 146412 280532 146468 280542
rect 163660 280532 163716 280542
rect 163240 280476 163660 280532
rect 146412 280466 146468 280476
rect 163660 280466 163716 280476
rect 198156 280532 198212 280542
rect 198156 280466 198212 280476
rect 151788 280420 151844 280430
rect 151788 280354 151844 280364
rect 153132 280308 153188 280318
rect 153132 280242 153188 280252
rect 166572 280196 166628 280206
rect 166572 280130 166628 280140
rect 121884 280084 121940 280094
rect 123004 280084 123060 280094
rect 137676 280084 137732 280094
rect 120540 276994 120596 277004
rect 120316 276882 120372 276892
rect 120876 276836 120932 280056
rect 121940 280028 122248 280084
rect 121884 280018 121940 280028
rect 120876 276770 120932 276780
rect 122892 276052 122948 280056
rect 123060 280028 123592 280084
rect 123676 280028 124264 280084
rect 124348 280028 124936 280084
rect 125020 280028 125608 280084
rect 123004 280018 123060 280028
rect 123676 279972 123732 280028
rect 123676 279906 123732 279916
rect 124348 277172 124404 280028
rect 125020 279748 125076 280028
rect 125020 279682 125076 279692
rect 125692 279972 125748 279982
rect 125692 279524 125748 279916
rect 125692 279458 125748 279468
rect 126252 277732 126308 280056
rect 126252 277666 126308 277676
rect 124348 277106 124404 277116
rect 122892 275986 122948 275996
rect 120204 274530 120260 274540
rect 126924 272692 126980 280056
rect 126924 272626 126980 272636
rect 127596 270228 127652 280056
rect 128940 272804 128996 280056
rect 128940 272738 128996 272748
rect 127596 270162 127652 270172
rect 129612 267876 129668 280056
rect 129612 267810 129668 267820
rect 119196 264898 119252 264908
rect 130284 264852 130340 280056
rect 130956 271908 131012 280056
rect 131628 277844 131684 280056
rect 132300 279860 132356 280056
rect 132300 279794 132356 279804
rect 131628 277778 131684 277788
rect 130956 271842 131012 271852
rect 132972 271124 133028 280056
rect 132972 271058 133028 271068
rect 134316 269556 134372 280056
rect 134988 279412 135044 280056
rect 134988 279346 135044 279356
rect 135660 274932 135716 280056
rect 135660 274866 135716 274876
rect 134316 269490 134372 269500
rect 136332 266868 136388 280056
rect 137004 278292 137060 280056
rect 159852 280084 159908 280094
rect 137676 280018 137732 280028
rect 137004 278226 137060 278236
rect 136332 266802 136388 266812
rect 138348 265188 138404 280056
rect 139020 268436 139076 280056
rect 139020 268370 139076 268380
rect 140364 266644 140420 280056
rect 142380 272020 142436 280056
rect 143052 275492 143108 280056
rect 143052 275426 143108 275436
rect 142380 271954 142436 271964
rect 143724 268324 143780 280056
rect 144396 271796 144452 280056
rect 145068 278628 145124 280056
rect 145068 278562 145124 278572
rect 145740 276948 145796 280056
rect 145740 276882 145796 276892
rect 144396 271730 144452 271740
rect 143724 268258 143780 268268
rect 147084 266756 147140 280056
rect 147756 268212 147812 280056
rect 147868 276836 147924 276846
rect 147868 273476 147924 276780
rect 147868 273410 147924 273420
rect 147756 268146 147812 268156
rect 147084 266690 147140 266700
rect 140364 266578 140420 266588
rect 138348 265122 138404 265132
rect 148428 265076 148484 280056
rect 149100 277060 149156 280056
rect 149100 276994 149156 277004
rect 149772 276276 149828 280056
rect 149772 276210 149828 276220
rect 150444 270004 150500 280056
rect 151116 277172 151172 280056
rect 151116 277106 151172 277116
rect 152460 275044 152516 280056
rect 152460 274978 152516 274988
rect 150444 269938 150500 269948
rect 153804 266980 153860 280056
rect 154476 270116 154532 280056
rect 155148 271572 155204 280056
rect 155820 271684 155876 280056
rect 156492 273588 156548 280056
rect 157164 275156 157220 280056
rect 157164 275090 157220 275100
rect 156492 273522 156548 273532
rect 155820 271618 155876 271628
rect 155148 271506 155204 271516
rect 154476 270050 154532 270060
rect 157052 270564 157108 270574
rect 153804 266914 153860 266924
rect 157052 265412 157108 270508
rect 157836 268548 157892 280056
rect 158508 275268 158564 280056
rect 159180 277172 159236 280056
rect 159852 280018 159908 280028
rect 159964 280028 160552 280084
rect 159180 277106 159236 277116
rect 159964 277172 160020 280028
rect 159964 277106 160020 277116
rect 161196 275380 161252 280056
rect 161196 275314 161252 275324
rect 158508 275202 158564 275212
rect 157836 268482 157892 268492
rect 157052 265346 157108 265356
rect 161868 265300 161924 280056
rect 162540 276836 162596 280056
rect 162540 276770 162596 276780
rect 163884 271460 163940 280056
rect 164556 278740 164612 280056
rect 164556 278674 164612 278684
rect 165228 277172 165284 280056
rect 165228 277106 165284 277116
rect 165900 277172 165956 280056
rect 167244 279636 167300 280056
rect 167244 279570 167300 279580
rect 165900 277106 165956 277116
rect 166236 277060 166292 277070
rect 166236 273028 166292 277004
rect 167916 276948 167972 280056
rect 167916 276882 167972 276892
rect 168140 280028 168616 280084
rect 168140 275604 168196 280028
rect 168140 275538 168196 275548
rect 169260 275604 169316 280056
rect 169260 275538 169316 275548
rect 169708 280028 169960 280084
rect 169708 275604 169764 280028
rect 169708 275538 169764 275548
rect 166236 272962 166292 272972
rect 163884 271394 163940 271404
rect 170604 266308 170660 280056
rect 171276 267988 171332 280056
rect 171276 267922 171332 267932
rect 170604 266242 170660 266252
rect 161868 265234 161924 265244
rect 148428 265010 148484 265020
rect 130284 264786 130340 264796
rect 171948 264628 172004 280056
rect 172620 270340 172676 280056
rect 173292 278516 173348 280056
rect 173292 278450 173348 278460
rect 173964 278404 174020 280056
rect 174636 278740 174692 280056
rect 174636 278674 174692 278684
rect 173964 278338 174020 278348
rect 175308 277172 175364 280056
rect 175308 277106 175364 277116
rect 175980 276276 176036 280056
rect 175980 276210 176036 276220
rect 176540 280028 176680 280084
rect 176540 275604 176596 280028
rect 176540 275538 176596 275548
rect 177324 275604 177380 280056
rect 177324 275538 177380 275548
rect 177996 271236 178052 280056
rect 178108 280028 178696 280084
rect 178108 275604 178164 280028
rect 179340 277060 179396 280056
rect 179340 276994 179396 277004
rect 179900 280028 180040 280084
rect 178108 275538 178164 275548
rect 179900 275604 179956 280028
rect 180684 275716 180740 280056
rect 181356 275828 181412 280056
rect 181356 275762 181412 275772
rect 181468 280028 182056 280084
rect 180684 275650 180740 275660
rect 179900 275538 179956 275548
rect 181468 275604 181524 280028
rect 181468 275538 181524 275548
rect 177996 271170 178052 271180
rect 172620 270274 172676 270284
rect 182700 267092 182756 280056
rect 183372 268772 183428 280056
rect 184044 277956 184100 280056
rect 184044 277890 184100 277900
rect 184716 275828 184772 280056
rect 184716 275762 184772 275772
rect 184828 280028 185416 280084
rect 184828 275604 184884 280028
rect 186060 275716 186116 280056
rect 186060 275650 186116 275660
rect 186396 276612 186452 276622
rect 184828 275538 184884 275548
rect 183372 268706 183428 268716
rect 182700 267026 182756 267036
rect 185612 268660 185668 268670
rect 181468 266196 181524 266206
rect 181468 265412 181524 266140
rect 185612 265524 185668 268604
rect 186396 268660 186452 276556
rect 186732 276276 186788 280056
rect 187404 278516 187460 280056
rect 187404 278450 187460 278460
rect 186732 276210 186788 276220
rect 188076 275940 188132 280056
rect 188076 275874 188132 275884
rect 188748 275604 188804 280056
rect 188748 275538 188804 275548
rect 189420 275604 189476 280056
rect 190092 276836 190148 280056
rect 190092 276770 190148 276780
rect 189420 275538 189476 275548
rect 186396 268594 186452 268604
rect 189084 275492 189140 275502
rect 185612 265458 185668 265468
rect 181468 265346 181524 265356
rect 171948 264562 172004 264572
rect 189084 264964 189140 275436
rect 190764 269668 190820 280056
rect 191436 275604 191492 280056
rect 191436 275538 191492 275548
rect 190764 269602 190820 269612
rect 192108 268100 192164 280056
rect 192780 276724 192836 280056
rect 192780 276658 192836 276668
rect 193452 270452 193508 280056
rect 194124 275716 194180 280056
rect 194124 275650 194180 275660
rect 194572 279972 194628 279982
rect 193452 270386 193508 270396
rect 192108 268034 192164 268044
rect 194572 270116 194628 279916
rect 194796 273364 194852 280056
rect 195468 273700 195524 280056
rect 195468 273634 195524 273644
rect 194796 273298 194852 273308
rect 196140 272132 196196 280056
rect 196812 273812 196868 280056
rect 197484 276164 197540 280056
rect 198828 278908 198884 280056
rect 198828 278852 199220 278908
rect 199164 278786 199220 278796
rect 197484 276098 197540 276108
rect 196812 273746 196868 273756
rect 196140 272066 196196 272076
rect 194572 267148 194628 270060
rect 194236 267092 194628 267148
rect 194236 266308 194292 267092
rect 194236 266242 194292 266252
rect 199276 265412 199332 371308
rect 199612 362964 199668 362974
rect 199388 301252 199444 301262
rect 199388 296436 199444 301196
rect 199388 296370 199444 296380
rect 199500 280756 199556 280766
rect 199500 280690 199556 280700
rect 199612 275492 199668 362908
rect 199612 275426 199668 275436
rect 199276 265346 199332 265356
rect 189084 264180 189140 264908
rect 189084 264114 189140 264124
rect 199388 168084 199444 168094
rect 199164 167524 199220 167534
rect 120092 165620 120148 165630
rect 122108 165620 122164 165630
rect 120148 165564 120456 165620
rect 121352 165564 122108 165620
rect 120092 165554 120148 165564
rect 122108 165554 122164 165564
rect 127596 165620 127652 165630
rect 154028 165620 154084 165630
rect 182476 165620 182532 165630
rect 183820 165620 183876 165630
rect 153160 165564 154028 165620
rect 182280 165564 182476 165620
rect 183624 165564 183820 165620
rect 127596 165554 127652 165564
rect 154028 165554 154084 165564
rect 182476 165554 182532 165564
rect 183820 165554 183876 165564
rect 184716 165620 184772 165630
rect 192332 165620 192388 165630
rect 192136 165564 192332 165620
rect 183708 165396 183764 165406
rect 120876 164164 120932 165032
rect 120876 164098 120932 164108
rect 126252 162932 126308 165032
rect 126728 165004 126980 165060
rect 126252 162866 126308 162876
rect 106876 162418 106932 162428
rect 81788 162306 81844 162316
rect 126924 160916 126980 165004
rect 127148 163828 127204 165032
rect 128072 165004 128324 165060
rect 127148 163762 127204 163772
rect 126924 160850 126980 160860
rect 128268 160804 128324 165004
rect 128492 164276 128548 165032
rect 128492 164210 128548 164220
rect 137900 162036 137956 165032
rect 138348 162820 138404 165032
rect 138796 164612 138852 165032
rect 138796 164546 138852 164556
rect 138348 162754 138404 162764
rect 137900 161970 137956 161980
rect 143724 161362 143780 165032
rect 144200 165004 144340 165060
rect 144648 165004 144900 165060
rect 144284 163044 144340 165004
rect 144172 162988 144340 163044
rect 143724 161310 143726 161362
rect 143778 161310 143780 161362
rect 143724 161298 143780 161310
rect 143836 162260 143892 162270
rect 143836 161588 143892 162204
rect 143836 161308 143892 161532
rect 144060 161476 144116 161486
rect 143836 161252 144004 161308
rect 128268 160738 128324 160748
rect 66332 160402 66388 160412
rect 143388 160468 143444 160478
rect 143388 159684 143444 160412
rect 127260 159012 127316 159022
rect 89852 157444 89908 157454
rect 65660 155474 65716 155484
rect 66108 157332 66164 157342
rect 56840 144844 56980 144900
rect 63980 148820 64036 148830
rect 63980 144872 64036 148764
rect 64428 148708 64484 148718
rect 64428 144872 64484 148652
rect 64876 144872 64932 149212
rect 65324 152180 65380 152190
rect 65324 149156 65380 152124
rect 65324 144872 65380 149100
rect 66108 149044 66164 157276
rect 82908 157332 82964 157342
rect 67116 152068 67172 152078
rect 67116 151172 67172 152012
rect 65436 148932 65492 148942
rect 65436 148708 65492 148876
rect 65436 148642 65492 148652
rect 66108 144900 66164 148988
rect 67004 151116 67116 151172
rect 67004 144900 67060 151116
rect 67116 151106 67172 151116
rect 71596 152068 71652 152078
rect 65800 144844 66164 144900
rect 66248 144844 67060 144900
rect 71148 150612 71204 150622
rect 71148 144872 71204 150556
rect 71596 144872 71652 152012
rect 81900 148708 81956 148718
rect 72044 147924 72100 147934
rect 72044 144872 72100 147868
rect 81452 147924 81508 147934
rect 81452 144872 81508 147868
rect 81900 144872 81956 148652
rect 82348 147924 82404 147934
rect 82348 144872 82404 147868
rect 82908 144900 82964 157276
rect 89180 155540 89236 155550
rect 83468 152180 83524 152190
rect 83468 149492 83524 152124
rect 83468 144900 83524 149436
rect 82824 144844 82964 144900
rect 83272 144844 83524 144900
rect 83692 152180 83748 152190
rect 83692 144872 83748 152124
rect 88620 148596 88676 148606
rect 88620 144872 88676 148540
rect 89180 144900 89236 155484
rect 89852 149380 89908 157388
rect 89852 144900 89908 149324
rect 126812 150724 126868 150734
rect 125916 148596 125972 148606
rect 118748 148148 118804 148158
rect 118300 148036 118356 148046
rect 89096 144844 89236 144900
rect 89544 144844 89908 144900
rect 117852 147924 117908 147934
rect 117852 144872 117908 147868
rect 118300 144872 118356 147980
rect 118748 144872 118804 148092
rect 125916 144872 125972 148540
rect 126364 147924 126420 147934
rect 126364 144872 126420 147868
rect 126812 144872 126868 150668
rect 127260 144872 127316 158956
rect 127708 155316 127764 155326
rect 127708 144872 127764 155260
rect 128156 152292 128212 152302
rect 128156 144872 128212 152236
rect 142828 151172 142884 151182
rect 138684 150388 138740 150398
rect 138012 149044 138068 149054
rect 137340 148484 137396 148494
rect 137340 144676 137396 148428
rect 138012 144872 138068 148988
rect 138684 144900 138740 150332
rect 142828 150388 142884 151116
rect 142828 150322 142884 150332
rect 142828 149044 142884 149054
rect 142828 148596 142884 148988
rect 142828 148530 142884 148540
rect 138488 144844 138740 144900
rect 143388 144872 143444 159628
rect 143948 156268 144004 161252
rect 143836 156212 144004 156268
rect 143836 144872 143892 156212
rect 144060 144900 144116 161420
rect 144172 149044 144228 162988
rect 144732 162148 144788 162158
rect 144284 161364 144340 161374
rect 144284 159684 144340 161308
rect 144284 159618 144340 159628
rect 144396 161362 144452 161374
rect 144396 161310 144398 161362
rect 144450 161310 144452 161362
rect 144396 150388 144452 161310
rect 144396 150322 144452 150332
rect 144172 148978 144228 148988
rect 144060 144844 144312 144900
rect 144732 144872 144788 162092
rect 144844 160692 144900 165004
rect 144844 160626 144900 160636
rect 145068 156324 145124 165032
rect 145404 165004 145544 165060
rect 145068 156258 145124 156268
rect 145180 162932 145236 162942
rect 145180 144872 145236 162876
rect 145404 160580 145460 165004
rect 145404 160524 145684 160580
rect 145628 148932 145684 160524
rect 145740 156324 145796 156334
rect 145740 149268 145796 156268
rect 145740 149202 145796 149212
rect 145628 148596 145684 148876
rect 145964 148820 146020 165032
rect 146076 162932 146132 162942
rect 146076 162148 146132 162876
rect 146076 162082 146132 162092
rect 164780 162148 164836 165032
rect 165228 162708 165284 165032
rect 165676 162932 165732 165032
rect 165676 162866 165732 162876
rect 166124 163044 166180 165032
rect 165228 162642 165284 162652
rect 164780 162082 164836 162092
rect 166124 161588 166180 162988
rect 166124 161522 166180 161532
rect 166236 162932 166292 162942
rect 166236 161476 166292 162876
rect 146076 160692 146132 160702
rect 146076 149156 146132 160636
rect 146076 148932 146132 149100
rect 146076 148866 146132 148876
rect 156828 160468 156884 160478
rect 145964 148754 146020 148764
rect 145628 148530 145684 148540
rect 156828 144872 156884 160412
rect 166236 152404 166292 161420
rect 166572 161364 166628 165032
rect 171500 164612 171556 165032
rect 171500 164546 171556 164556
rect 171948 162484 172004 165032
rect 172396 162596 172452 165032
rect 181804 163940 181860 165032
rect 181804 163874 181860 163884
rect 172396 162530 172452 162540
rect 171948 162418 172004 162428
rect 166572 161298 166628 161308
rect 167916 162372 167972 162382
rect 167916 161364 167972 162316
rect 182700 162260 182756 165032
rect 183148 162820 183204 165032
rect 183148 162754 183204 162764
rect 183260 164724 183316 164734
rect 182700 162194 182756 162204
rect 166236 152338 166292 152348
rect 166236 150388 166292 150398
rect 164892 149268 164948 149278
rect 164556 148820 164612 148830
rect 164556 148148 164612 148764
rect 164220 148092 164612 148148
rect 164220 144900 164276 148092
rect 164556 148036 164612 148092
rect 164556 147970 164612 147980
rect 164892 148260 164948 149212
rect 165788 149044 165844 149054
rect 164024 144844 164276 144900
rect 164444 147924 164500 147934
rect 164444 144872 164500 147868
rect 164892 144872 164948 148204
rect 165340 148932 165396 148942
rect 165340 148148 165396 148876
rect 165340 144872 165396 148092
rect 165788 147252 165844 148988
rect 165788 144872 165844 147196
rect 166236 144676 166292 150332
rect 167916 145572 167972 161308
rect 181916 160692 181972 160702
rect 181468 160580 181524 160590
rect 167916 145506 167972 145516
rect 171164 159236 171220 159246
rect 171164 144872 171220 159180
rect 172060 158900 172116 158910
rect 171612 150388 171668 150398
rect 171612 144872 171668 150332
rect 172060 144872 172116 158844
rect 181468 144872 181524 160524
rect 181916 144872 181972 160636
rect 182364 159124 182420 159134
rect 182364 144872 182420 159068
rect 182812 150836 182868 150846
rect 182812 144872 182868 150780
rect 183260 144872 183316 164668
rect 183708 144872 183764 165340
rect 184044 164612 184100 165032
rect 184716 164724 184772 165564
rect 192332 165554 192388 165564
rect 184716 164658 184772 164668
rect 184044 164546 184100 164556
rect 189420 164500 189476 164510
rect 189420 163380 189476 164444
rect 189420 161308 189476 163324
rect 191212 162932 191268 165032
rect 191660 164500 191716 165032
rect 191660 164434 191716 164444
rect 191212 162866 191268 162876
rect 199164 162484 199220 167468
rect 199276 164948 199332 164958
rect 199276 162820 199332 164892
rect 199276 162754 199332 162764
rect 199164 162418 199220 162428
rect 199164 162148 199220 162158
rect 189420 161252 189588 161308
rect 189084 148932 189140 148942
rect 188636 148596 188692 148606
rect 188636 144872 188692 148540
rect 189084 144872 189140 148876
rect 189532 144872 189588 161252
rect 137340 144620 137592 144676
rect 166236 144610 166292 144620
rect 166236 144564 166292 144574
rect 166236 144498 166292 144508
rect 199052 144564 199108 144574
rect 199052 129332 199108 144508
rect 199052 129266 199108 129276
rect 7532 121650 7588 121660
rect 199164 45332 199220 162092
rect 199276 161364 199332 161374
rect 199276 71988 199332 161308
rect 199388 148596 199444 168028
rect 199388 148530 199444 148540
rect 199948 148148 200004 374892
rect 202076 373716 202132 373726
rect 200620 373604 200676 373614
rect 199948 148082 200004 148092
rect 200060 366996 200116 367006
rect 200060 147924 200116 366940
rect 200172 347620 200228 347630
rect 200172 165508 200228 347564
rect 200172 165442 200228 165452
rect 200284 307300 200340 307310
rect 200284 150836 200340 307244
rect 200508 305060 200564 305070
rect 200508 297388 200564 305004
rect 200284 150770 200340 150780
rect 200396 297332 200564 297388
rect 200396 150388 200452 297332
rect 200508 290500 200564 290510
rect 200508 164164 200564 290444
rect 200620 278292 200676 373548
rect 201964 373156 202020 373166
rect 200844 371588 200900 371598
rect 200732 368340 200788 368350
rect 200732 303156 200788 368284
rect 200732 303090 200788 303100
rect 200620 278226 200676 278236
rect 200732 299124 200788 299134
rect 200508 164098 200564 164108
rect 200396 150322 200452 150332
rect 200732 148932 200788 299068
rect 200844 292404 200900 371532
rect 201628 368900 201684 368910
rect 200956 365092 201012 365102
rect 200956 297780 201012 365036
rect 201180 361508 201236 361518
rect 201068 360612 201124 360622
rect 201068 308532 201124 360556
rect 201180 313908 201236 361452
rect 201628 352100 201684 368844
rect 201628 352034 201684 352044
rect 201740 365540 201796 365550
rect 201740 340900 201796 365484
rect 201740 340834 201796 340844
rect 201852 363636 201908 363646
rect 201852 338660 201908 363580
rect 201964 353220 202020 373100
rect 201964 353154 202020 353164
rect 202076 350980 202132 373660
rect 208684 373492 208740 373502
rect 207452 373044 207508 373054
rect 203308 370020 203364 370030
rect 202076 350914 202132 350924
rect 202412 363300 202468 363310
rect 201852 338594 201908 338604
rect 202300 348740 202356 348750
rect 201180 313842 201236 313852
rect 201068 308466 201124 308476
rect 201740 308420 201796 308430
rect 201740 299124 201796 308364
rect 201740 299058 201796 299068
rect 200956 297714 201012 297724
rect 200844 292338 200900 292348
rect 201740 294980 201796 294990
rect 201628 287140 201684 287150
rect 200844 282660 200900 282670
rect 200844 164500 200900 282604
rect 201628 280644 201684 287084
rect 201628 280578 201684 280588
rect 201740 278068 201796 294924
rect 201740 278002 201796 278012
rect 201852 291620 201908 291630
rect 200844 164434 200900 164444
rect 201628 275604 201684 275614
rect 200732 148866 200788 148876
rect 201180 148148 201236 148158
rect 200060 147858 200116 147868
rect 200956 147924 201012 147934
rect 199276 71922 199332 71932
rect 199724 147476 199780 147486
rect 199724 66612 199780 147420
rect 200844 145572 200900 145582
rect 200732 129332 200788 129342
rect 200732 104132 200788 129276
rect 200732 104066 200788 104076
rect 200844 69300 200900 145516
rect 200844 69234 200900 69244
rect 199724 66546 199780 66556
rect 200956 61236 201012 147868
rect 201180 80052 201236 148092
rect 201628 147924 201684 275548
rect 201852 269892 201908 291564
rect 201852 269826 201908 269836
rect 201964 289380 202020 289390
rect 201964 163828 202020 289324
rect 202076 286020 202132 286030
rect 202076 167524 202132 285964
rect 202076 167458 202132 167468
rect 202188 283780 202244 283790
rect 202188 164948 202244 283724
rect 202300 168084 202356 348684
rect 202412 327572 202468 363244
rect 202636 363188 202692 363198
rect 202636 331828 202692 363132
rect 202636 331762 202692 331772
rect 202412 327506 202468 327516
rect 202524 329700 202580 329710
rect 202524 300804 202580 329644
rect 202524 300738 202580 300748
rect 202636 327460 202692 327470
rect 202636 297108 202692 327404
rect 202860 326340 202916 326350
rect 202860 310884 202916 326284
rect 202860 310818 202916 310828
rect 202636 297042 202692 297052
rect 202860 301700 202916 301710
rect 202524 292740 202580 292750
rect 202412 275828 202468 275838
rect 202412 206612 202468 275772
rect 202524 273140 202580 292684
rect 202524 273074 202580 273084
rect 202412 206546 202468 206556
rect 202524 266308 202580 266318
rect 202300 168018 202356 168028
rect 202188 164882 202244 164892
rect 201964 163762 202020 163772
rect 201628 147858 201684 147868
rect 201180 79986 201236 79996
rect 200956 61170 201012 61180
rect 202524 55860 202580 266252
rect 202748 152404 202804 152414
rect 202636 147924 202692 147934
rect 202636 63924 202692 147868
rect 202748 74676 202804 152348
rect 202860 150724 202916 301644
rect 203308 162708 203364 369964
rect 204988 369908 205044 369918
rect 204092 368116 204148 368126
rect 203308 155428 203364 162652
rect 203308 155362 203364 155372
rect 203420 343140 203476 343150
rect 203420 152292 203476 343084
rect 203532 320740 203588 320750
rect 203532 160468 203588 320684
rect 203644 284900 203700 284910
rect 203644 162260 203700 284844
rect 204092 187572 204148 368060
rect 204316 361732 204372 361742
rect 204092 187506 204148 187516
rect 204204 359604 204260 359614
rect 204204 182868 204260 359548
rect 204316 281652 204372 361676
rect 204316 281586 204372 281596
rect 204428 360500 204484 360510
rect 204428 262836 204484 360444
rect 204652 360276 204708 360286
rect 204652 289716 204708 360220
rect 204876 360052 204932 360062
rect 204876 300468 204932 359996
rect 204876 300402 204932 300412
rect 204652 289650 204708 289660
rect 204428 262770 204484 262780
rect 204204 182196 204260 182812
rect 204204 182130 204260 182140
rect 204988 163044 205044 369852
rect 205884 369684 205940 369694
rect 205772 364756 205828 364766
rect 204988 162978 205044 162988
rect 205100 346500 205156 346510
rect 203644 162194 203700 162204
rect 205100 160580 205156 346444
rect 205100 160514 205156 160524
rect 205212 306180 205268 306190
rect 203532 160402 203588 160412
rect 205212 159124 205268 306124
rect 205772 179508 205828 364700
rect 205884 184996 205940 369628
rect 205996 368788 206052 368798
rect 205996 227892 206052 368732
rect 206220 368452 206276 368462
rect 206108 366548 206164 366558
rect 206108 268212 206164 366492
rect 206220 278964 206276 368396
rect 207340 362068 207396 362078
rect 206332 359940 206388 359950
rect 206332 295092 206388 359884
rect 206556 359716 206612 359726
rect 206556 305844 206612 359660
rect 207340 316596 207396 362012
rect 207340 316530 207396 316540
rect 206556 305778 206612 305788
rect 206668 311780 206724 311790
rect 206332 295026 206388 295036
rect 206220 278898 206276 278908
rect 206108 268146 206164 268156
rect 205996 227826 206052 227836
rect 205884 184930 205940 184940
rect 205772 179442 205828 179452
rect 205212 159058 205268 159068
rect 204204 157556 204260 157566
rect 203420 152226 203476 152236
rect 204092 153860 204148 153870
rect 202860 150658 202916 150668
rect 203196 104132 203252 104142
rect 203196 99204 203252 104076
rect 204092 101556 204148 153804
rect 204204 109620 204260 157500
rect 204540 157444 204596 157454
rect 204428 153748 204484 153758
rect 204204 109554 204260 109564
rect 204316 147028 204372 147038
rect 204092 101490 204148 101500
rect 203196 99148 203364 99204
rect 203308 97524 203364 99148
rect 204316 98868 204372 146972
rect 204428 106932 204484 153692
rect 204540 112308 204596 157388
rect 206668 157108 206724 311724
rect 206780 310884 206836 310894
rect 206780 162596 206836 310828
rect 207452 195636 207508 372988
rect 208348 371924 208404 371934
rect 207900 369796 207956 369806
rect 207788 368564 207844 368574
rect 207676 366772 207732 366782
rect 207564 360388 207620 360398
rect 207564 311220 207620 360332
rect 207564 311154 207620 311164
rect 207452 195570 207508 195580
rect 207564 252084 207620 252094
rect 206780 162530 206836 162540
rect 206668 157042 206724 157052
rect 207452 155652 207508 155662
rect 204652 152180 204708 152190
rect 204652 117684 204708 152124
rect 206892 149380 206948 149390
rect 206780 148820 206836 148830
rect 206668 148708 206724 148718
rect 206668 147252 206724 148652
rect 206668 147186 206724 147196
rect 206780 144564 206836 148764
rect 206780 144498 206836 144508
rect 206892 141876 206948 149324
rect 206892 141810 206948 141820
rect 204652 117618 204708 117628
rect 207452 114996 207508 155596
rect 207452 114930 207508 114940
rect 204540 112242 204596 112252
rect 204428 106866 204484 106876
rect 204316 98802 204372 98812
rect 203420 97524 203476 97534
rect 203308 97468 203420 97524
rect 203420 97458 203476 97468
rect 202748 74610 202804 74620
rect 207452 97412 207508 97422
rect 202636 63858 202692 63868
rect 207452 57876 207508 97356
rect 207452 57810 207508 57820
rect 202524 55794 202580 55804
rect 207564 50484 207620 252028
rect 207676 241332 207732 366716
rect 207788 249396 207844 368508
rect 207900 252084 207956 369740
rect 208124 331828 208180 331838
rect 208012 325220 208068 325230
rect 208012 254772 208068 325164
rect 208012 254706 208068 254716
rect 207900 252018 207956 252028
rect 207788 249330 207844 249340
rect 208012 249508 208068 249518
rect 207676 241266 207732 241276
rect 207676 155428 207732 155438
rect 207676 77364 207732 155372
rect 207788 147364 207844 147374
rect 207788 88116 207844 147308
rect 207900 145460 207956 145470
rect 207900 93492 207956 145404
rect 208012 131124 208068 249452
rect 208124 246708 208180 331772
rect 208124 246642 208180 246652
rect 208236 327572 208292 327582
rect 208236 244020 208292 327516
rect 208236 243954 208292 243964
rect 208348 162372 208404 371868
rect 208460 366324 208516 366334
rect 208460 176820 208516 366268
rect 208460 176754 208516 176764
rect 208572 345380 208628 345390
rect 208348 162306 208404 162316
rect 208572 158900 208628 345324
rect 208684 199108 208740 373436
rect 209132 372036 209188 372046
rect 208684 199042 208740 199052
rect 208796 302820 208852 302830
rect 208796 159012 208852 302764
rect 209132 230580 209188 371980
rect 209244 367108 209300 367118
rect 209244 273588 209300 367052
rect 209580 360388 209636 595560
rect 210364 376404 210420 376414
rect 210028 368228 210084 368238
rect 209580 360322 209636 360332
rect 209916 364980 209972 364990
rect 209356 359828 209412 359838
rect 209356 287028 209412 359772
rect 209356 286962 209412 286972
rect 209244 273522 209300 273532
rect 209916 266084 209972 364924
rect 210028 285012 210084 368172
rect 210140 367220 210196 367230
rect 210140 322532 210196 367164
rect 210140 322466 210196 322476
rect 210252 361396 210308 361406
rect 210252 319956 210308 361340
rect 210252 319890 210308 319900
rect 210028 284946 210084 284956
rect 210140 297108 210196 297118
rect 209916 266018 209972 266028
rect 209132 230514 209188 230524
rect 210140 162036 210196 297052
rect 210364 277172 210420 376348
rect 211708 363972 211764 363982
rect 211708 325220 211764 363916
rect 211708 325154 211764 325164
rect 217196 343588 217252 343598
rect 217196 324968 217252 343532
rect 231644 336868 231700 595560
rect 231644 336802 231700 336812
rect 243628 589652 243684 589662
rect 230412 330148 230468 330158
rect 230412 324968 230468 330092
rect 243628 324968 243684 589596
rect 253708 589652 253764 595560
rect 253708 589586 253764 589596
rect 256844 373828 256900 373838
rect 256844 324968 256900 373772
rect 270060 341908 270116 341918
rect 270060 324968 270116 341852
rect 275772 330260 275828 595560
rect 296492 360388 296548 360398
rect 275772 330194 275828 330204
rect 283276 330260 283332 330270
rect 283276 324968 283332 330204
rect 296492 324968 296548 360332
rect 297836 357028 297892 595560
rect 297836 356962 297892 356972
rect 309708 380548 309764 380558
rect 309708 324968 309764 380492
rect 319900 330148 319956 595560
rect 319900 330082 319956 330092
rect 322924 590772 322980 590782
rect 322924 324968 322980 590716
rect 336140 357028 336196 357038
rect 336140 324968 336196 356972
rect 341964 341908 342020 595560
rect 364028 590772 364084 595560
rect 364028 590706 364084 590716
rect 341964 341842 342020 341852
rect 362572 390740 362628 390750
rect 349356 336868 349412 336878
rect 349356 324968 349412 336812
rect 362572 324968 362628 390684
rect 377132 361284 377188 361294
rect 375788 326340 375844 326350
rect 375564 326116 375620 326126
rect 373548 318724 373604 318734
rect 372764 317380 372820 317390
rect 371084 308644 371140 308654
rect 210364 277106 210420 277116
rect 370636 285796 370692 285806
rect 370076 265524 370132 265534
rect 370076 204036 370132 265468
rect 370412 262164 370468 262174
rect 370076 203970 370132 203980
rect 370300 206724 370356 206734
rect 210140 161970 210196 161980
rect 370076 171444 370132 171454
rect 208796 158946 208852 158956
rect 208572 158834 208628 158844
rect 208012 131058 208068 131068
rect 208124 147140 208180 147150
rect 207900 93426 207956 93436
rect 208124 90804 208180 147084
rect 208236 145348 208292 145358
rect 208236 96180 208292 145292
rect 208236 96114 208292 96124
rect 208124 90738 208180 90748
rect 207788 88050 207844 88060
rect 207676 77298 207732 77308
rect 207564 50418 207620 50428
rect 199164 45266 199220 45276
rect 370076 44436 370132 171388
rect 370188 161252 370244 161262
rect 370188 89460 370244 161196
rect 370300 147924 370356 206668
rect 370412 204708 370468 262108
rect 370412 204642 370468 204652
rect 370524 246036 370580 246046
rect 370300 147858 370356 147868
rect 370524 130788 370580 245980
rect 370636 234388 370692 285740
rect 370636 234322 370692 234332
rect 370748 273028 370804 273038
rect 370748 222628 370804 272972
rect 370972 269556 371028 269566
rect 370748 222562 370804 222572
rect 370860 239428 370916 239438
rect 370748 217812 370804 217822
rect 370748 209972 370804 217756
rect 370748 209906 370804 209916
rect 370748 202244 370804 202254
rect 370748 153860 370804 202188
rect 370860 165284 370916 239372
rect 370972 203140 371028 269500
rect 371084 240100 371140 308588
rect 372204 296884 372260 296894
rect 371980 285684 372036 285694
rect 371868 274708 371924 274718
rect 371196 263060 371252 263070
rect 371196 246036 371252 263004
rect 371196 245970 371252 245980
rect 371084 240034 371140 240044
rect 371196 234836 371252 234846
rect 371196 220108 371252 234780
rect 371868 233268 371924 274652
rect 371980 270340 372036 285628
rect 371980 270274 372036 270284
rect 372092 277844 372148 277854
rect 371868 233202 371924 233212
rect 371980 240660 372036 240670
rect 370972 203074 371028 203084
rect 371084 220052 371252 220108
rect 371868 231924 371924 231934
rect 370860 165218 370916 165228
rect 370972 173348 371028 173358
rect 370748 153794 370804 153804
rect 370524 130722 370580 130732
rect 370412 125524 370468 125534
rect 370188 89394 370244 89404
rect 370300 119924 370356 119934
rect 370300 78036 370356 119868
rect 370412 90132 370468 125468
rect 370972 90916 371028 173292
rect 371084 131012 371140 220052
rect 371756 218596 371812 218606
rect 371756 206724 371812 218540
rect 371756 206658 371812 206668
rect 371868 199556 371924 231868
rect 371868 199490 371924 199500
rect 371084 130946 371140 130956
rect 371980 130676 372036 240604
rect 372092 207172 372148 277788
rect 372204 273588 372260 296828
rect 372652 292516 372708 292526
rect 372204 273522 372260 273532
rect 372316 286804 372372 286814
rect 372316 270228 372372 286748
rect 372316 270162 372372 270172
rect 372428 271684 372484 271694
rect 372092 207106 372148 207116
rect 372204 264404 372260 264414
rect 372204 204820 372260 264348
rect 372428 239540 372484 271628
rect 372428 239474 372484 239484
rect 372540 257684 372596 257694
rect 372316 234164 372372 234174
rect 372316 205940 372372 234108
rect 372316 205874 372372 205884
rect 372428 225988 372484 225998
rect 372204 204754 372260 204764
rect 372204 202580 372260 202590
rect 371980 130610 372036 130620
rect 372092 163044 372148 163054
rect 372092 123508 372148 162988
rect 372204 157780 372260 202524
rect 372204 157714 372260 157724
rect 372316 174692 372372 174702
rect 372204 155540 372260 155550
rect 372204 137508 372260 155484
rect 372204 137442 372260 137452
rect 372092 123442 372148 123452
rect 372204 130676 372260 130686
rect 370972 90850 371028 90860
rect 372092 98868 372148 98878
rect 370412 90066 370468 90076
rect 370300 77970 370356 77980
rect 372092 68404 372148 98812
rect 372204 95060 372260 130620
rect 372316 125188 372372 174636
rect 372428 146804 372484 225932
rect 372540 204484 372596 257628
rect 372652 229348 372708 292460
rect 372652 229282 372708 229292
rect 372540 204418 372596 204428
rect 372652 222740 372708 222750
rect 372428 146738 372484 146748
rect 372540 180068 372596 180078
rect 372316 125122 372372 125132
rect 372204 94276 372260 95004
rect 372204 94210 372260 94220
rect 372428 109844 372484 109854
rect 372092 68338 372148 68348
rect 372428 67956 372484 109788
rect 372540 96628 372596 180012
rect 372652 132692 372708 222684
rect 372764 218708 372820 317324
rect 373324 271572 373380 271582
rect 373212 265412 373268 265422
rect 373100 265076 373156 265086
rect 372876 256116 372932 256126
rect 372876 240212 372932 256060
rect 372876 240146 372932 240156
rect 372988 240100 373044 240110
rect 372988 225092 373044 240044
rect 372988 225026 373044 225036
rect 372764 218642 372820 218652
rect 372988 224420 373044 224430
rect 372764 203028 372820 203038
rect 372764 153972 372820 202972
rect 372764 153906 372820 153916
rect 372988 150164 373044 224364
rect 373100 217924 373156 265020
rect 373212 248724 373268 265356
rect 373212 248658 373268 248668
rect 373100 217858 373156 217868
rect 373324 213220 373380 271516
rect 373436 246932 373492 246942
rect 373436 233492 373492 246876
rect 373436 233426 373492 233436
rect 373548 219156 373604 318668
rect 375452 317044 375508 317054
rect 374108 314020 374164 314030
rect 373996 271012 374052 271022
rect 373884 264740 373940 264750
rect 373884 243628 373940 264684
rect 373660 243572 373940 243628
rect 373660 240324 373716 243572
rect 373660 240258 373716 240268
rect 373884 242788 373940 242798
rect 373548 219090 373604 219100
rect 373772 240212 373828 240222
rect 373324 213154 373380 213164
rect 373436 211652 373492 211662
rect 373436 205604 373492 211596
rect 373436 205538 373492 205548
rect 373100 196756 373156 196766
rect 373100 194964 373156 196700
rect 373100 194898 373156 194908
rect 373212 196644 373268 196654
rect 373100 193284 373156 193294
rect 373100 189028 373156 193228
rect 373212 190484 373268 196588
rect 373212 190418 373268 190428
rect 373100 188962 373156 188972
rect 373324 175924 373380 175934
rect 373324 155428 373380 175868
rect 373324 155362 373380 155372
rect 372988 149156 373044 150108
rect 372988 149090 373044 149100
rect 372652 132626 372708 132636
rect 372764 147812 372820 147822
rect 372540 96562 372596 96572
rect 372652 122276 372708 122286
rect 372652 121044 372708 122220
rect 372540 95732 372596 95742
rect 372540 80052 372596 95676
rect 372652 80724 372708 120988
rect 372652 80658 372708 80668
rect 372540 79986 372596 79996
rect 372428 67890 372484 67900
rect 370076 44370 370132 44380
rect 372764 41860 372820 147756
rect 373100 132692 373156 132702
rect 372988 126644 373044 126654
rect 372988 124628 373044 126588
rect 372988 124562 373044 124572
rect 373100 108724 373156 132636
rect 373772 130900 373828 240156
rect 373884 238868 373940 242732
rect 373996 240436 374052 270956
rect 374108 263844 374164 313964
rect 374444 283108 374500 283118
rect 374332 271460 374388 271470
rect 374108 263778 374164 263788
rect 374220 270788 374276 270798
rect 373996 240370 374052 240380
rect 373884 238802 373940 238812
rect 373996 233492 374052 233502
rect 373884 233268 373940 233278
rect 373884 180068 373940 233212
rect 373996 231924 374052 233436
rect 373996 201460 374052 231868
rect 374108 217140 374164 217150
rect 374108 201572 374164 217084
rect 374220 215572 374276 270732
rect 374332 231868 374388 271404
rect 374444 263956 374500 283052
rect 375452 270116 375508 316988
rect 375564 304724 375620 326060
rect 375676 324436 375732 324446
rect 375676 310324 375732 324380
rect 375676 310258 375732 310268
rect 375788 305844 375844 326284
rect 377132 324324 377188 361228
rect 386092 343588 386148 595560
rect 408268 588868 408324 595560
rect 408268 588802 408324 588812
rect 430220 385588 430276 595560
rect 430220 385522 430276 385532
rect 452284 372148 452340 595560
rect 474348 375508 474404 595560
rect 494732 590212 494788 590222
rect 494732 383908 494788 590156
rect 496412 590212 496468 595560
rect 518476 590660 518532 595560
rect 518476 590594 518532 590604
rect 496412 590146 496468 590156
rect 494732 383842 494788 383852
rect 540540 378868 540596 595560
rect 562604 590548 562660 595560
rect 562604 590482 562660 590492
rect 584668 590212 584724 595560
rect 584668 590146 584724 590156
rect 590156 443268 590212 443278
rect 590156 437668 590212 443212
rect 590156 437602 590212 437612
rect 540540 378802 540596 378812
rect 474348 375442 474404 375452
rect 511532 377188 511588 377198
rect 452284 372082 452340 372092
rect 386092 343522 386148 343532
rect 408940 328132 408996 328142
rect 392812 327796 392868 327806
rect 389452 327684 389508 327694
rect 378588 326228 378644 326238
rect 377132 324258 377188 324268
rect 377916 324324 377972 324334
rect 375788 305778 375844 305788
rect 377692 314692 377748 314702
rect 375564 304658 375620 304668
rect 375564 303604 375620 303614
rect 375564 273364 375620 303548
rect 375788 298004 375844 298014
rect 375788 273476 375844 297948
rect 375788 273410 375844 273420
rect 376908 289828 376964 289838
rect 375564 273298 375620 273308
rect 375452 270050 375508 270060
rect 376236 271236 376292 271246
rect 374444 263890 374500 263900
rect 374556 268324 374612 268334
rect 374556 242228 374612 268268
rect 374668 267764 374724 267774
rect 374668 266868 374724 267708
rect 376012 267764 376068 267774
rect 374668 266802 374724 266812
rect 375228 267428 375284 267438
rect 375228 245476 375284 267372
rect 375676 266644 375732 266654
rect 375340 265636 375396 265646
rect 375340 255444 375396 265580
rect 375340 255378 375396 255388
rect 375452 265300 375508 265310
rect 375228 245410 375284 245420
rect 375340 250068 375396 250078
rect 374556 242162 374612 242172
rect 375228 235284 375284 235294
rect 374332 231812 374612 231868
rect 374220 215506 374276 215516
rect 374556 215460 374612 231812
rect 374668 221172 374724 221182
rect 374668 218596 374724 221116
rect 374668 218530 374724 218540
rect 374556 215394 374612 215404
rect 374556 215124 374612 215134
rect 374108 201506 374164 201516
rect 374332 202468 374388 202478
rect 373996 201394 374052 201404
rect 373884 180002 373940 180012
rect 373996 194852 374052 194862
rect 373996 178164 374052 194796
rect 374332 194516 374388 202412
rect 374556 201572 374612 215068
rect 374332 194450 374388 194460
rect 374444 195076 374500 195086
rect 374108 191716 374164 191726
rect 374108 181524 374164 191660
rect 374444 184884 374500 195020
rect 374444 184818 374500 184828
rect 374108 181458 374164 181468
rect 373996 178098 374052 178108
rect 374444 180740 374500 180750
rect 374332 176372 374388 176382
rect 374220 164612 374276 164622
rect 373772 130834 373828 130844
rect 373884 162596 373940 162606
rect 373772 124516 373828 124526
rect 373100 108658 373156 108668
rect 373212 124404 373268 124414
rect 373212 95732 373268 124348
rect 373772 116564 373828 124460
rect 373884 124404 373940 162540
rect 373996 156884 374052 156894
rect 373996 137284 374052 156828
rect 373996 137218 374052 137228
rect 374220 131124 374276 164556
rect 374332 136948 374388 176316
rect 374332 136882 374388 136892
rect 374220 131058 374276 131068
rect 374332 134596 374388 134606
rect 374108 130900 374164 130910
rect 374332 130900 374388 134540
rect 373884 124338 373940 124348
rect 373996 127204 374052 127214
rect 373772 116498 373828 116508
rect 373996 110964 374052 127148
rect 373996 110898 374052 110908
rect 373996 108388 374052 108398
rect 373212 95666 373268 95676
rect 373772 108386 374052 108388
rect 373772 108334 373998 108386
rect 374050 108334 374052 108386
rect 373772 108332 374052 108334
rect 372988 95508 373044 95518
rect 372876 94500 372932 94510
rect 372876 93828 372932 94444
rect 372876 93762 372932 93772
rect 372988 84084 373044 95452
rect 373772 94164 373828 108332
rect 373996 108322 374052 108332
rect 373772 94098 373828 94108
rect 373884 108164 373940 108174
rect 373212 90916 373268 90926
rect 372988 84018 373044 84028
rect 373100 85428 373156 85438
rect 373100 60564 373156 85372
rect 373212 70756 373268 90860
rect 373772 90692 373828 90702
rect 373212 70690 373268 70700
rect 373324 84084 373380 84094
rect 373100 60498 373156 60508
rect 373324 58324 373380 84028
rect 373772 69524 373828 90636
rect 373772 69458 373828 69468
rect 373884 67284 373940 108108
rect 374108 98644 374164 130844
rect 374220 130844 374388 130900
rect 374220 126028 374276 130844
rect 374332 130004 374388 130014
rect 374332 127988 374388 129948
rect 374332 127922 374388 127932
rect 374332 127764 374388 127774
rect 374332 127540 374388 127708
rect 374332 127474 374388 127484
rect 374220 125972 374388 126028
rect 374220 118804 374276 118814
rect 374220 116340 374276 118748
rect 374220 116274 374276 116284
rect 374332 109844 374388 125972
rect 374332 109778 374388 109788
rect 374108 98578 374164 98588
rect 374220 105364 374276 105374
rect 374108 95732 374164 95742
rect 374108 71316 374164 95676
rect 374108 71250 374164 71260
rect 373884 67218 373940 67228
rect 374220 62580 374276 105308
rect 374220 62514 374276 62524
rect 374332 104132 374388 104142
rect 374332 103124 374388 104076
rect 374332 61236 374388 103068
rect 374444 87332 374500 180684
rect 374556 152740 374612 201516
rect 375116 208516 375172 208526
rect 375116 197764 375172 208460
rect 375228 199444 375284 235228
rect 375340 235172 375396 250012
rect 375452 247604 375508 265244
rect 375452 247538 375508 247548
rect 375564 259924 375620 259934
rect 375340 235106 375396 235116
rect 375452 246932 375508 246942
rect 375452 213332 375508 246876
rect 375452 213266 375508 213276
rect 375228 199378 375284 199388
rect 375452 209524 375508 209534
rect 375116 197698 375172 197708
rect 375452 197652 375508 209468
rect 375564 204932 375620 259868
rect 375676 206052 375732 266588
rect 375900 261716 375956 261726
rect 375676 205986 375732 205996
rect 375788 256564 375844 256574
rect 375564 204866 375620 204876
rect 375788 204372 375844 256508
rect 375900 237748 375956 261660
rect 375900 237682 375956 237692
rect 375788 204306 375844 204316
rect 375900 237524 375956 237534
rect 375900 204148 375956 237468
rect 375788 204092 375956 204148
rect 375788 199332 375844 204092
rect 375900 203924 375956 203934
rect 375900 201012 375956 203868
rect 375900 200946 375956 200956
rect 375900 199332 375956 199342
rect 375788 199276 375900 199332
rect 375900 199266 375956 199276
rect 375452 197586 375508 197596
rect 375900 196084 375956 196094
rect 375788 195188 375844 195198
rect 375676 192500 375732 192510
rect 375452 190148 375508 190158
rect 375228 186564 375284 186574
rect 375228 160244 375284 186508
rect 375228 160178 375284 160188
rect 375340 164724 375396 164734
rect 374556 152674 374612 152684
rect 375228 155428 375284 155438
rect 374556 151172 374612 151182
rect 374556 115668 374612 151116
rect 375228 147140 375284 155372
rect 375228 145684 375284 147084
rect 375228 145618 375284 145628
rect 375228 131012 375284 131022
rect 375228 129332 375284 130956
rect 375228 129266 375284 129276
rect 375340 128884 375396 164668
rect 375452 151172 375508 190092
rect 375452 151106 375508 151116
rect 375564 170324 375620 170334
rect 375452 145684 375508 145694
rect 375452 137172 375508 145628
rect 375452 137106 375508 137116
rect 375340 128818 375396 128828
rect 374556 108386 374612 115612
rect 374556 108334 374558 108386
rect 374610 108334 374612 108386
rect 374556 108322 374612 108334
rect 374444 87266 374500 87276
rect 374556 107604 374612 107614
rect 374444 85652 374500 85662
rect 374444 84084 374500 85596
rect 374444 84018 374500 84028
rect 374332 61170 374388 61180
rect 374444 72212 374500 72222
rect 374444 59444 374500 72156
rect 374556 64596 374612 107548
rect 374556 64530 374612 64540
rect 375452 104244 375508 104254
rect 375452 61908 375508 104188
rect 375452 61842 375508 61852
rect 374444 59378 374500 59388
rect 373324 58258 373380 58268
rect 374556 52724 374612 52734
rect 374556 41972 374612 52668
rect 375564 44772 375620 170268
rect 375676 163940 375732 192444
rect 375676 163874 375732 163884
rect 375676 161924 375732 161934
rect 375676 137788 375732 161868
rect 375788 155428 375844 195132
rect 375788 155362 375844 155372
rect 375676 137732 375844 137788
rect 375788 123284 375844 137732
rect 375900 133924 375956 196028
rect 376012 173348 376068 267708
rect 376124 265524 376180 265534
rect 376124 253204 376180 265468
rect 376124 253138 376180 253148
rect 376012 173282 376068 173292
rect 376124 248948 376180 248958
rect 375900 133858 375956 133868
rect 376012 147924 376068 147934
rect 375676 110964 375732 110974
rect 375676 68628 375732 110908
rect 375788 82740 375844 123228
rect 375788 82674 375844 82684
rect 375900 106484 375956 106494
rect 375676 68562 375732 68572
rect 375900 63252 375956 106428
rect 376012 91476 376068 147868
rect 376124 132244 376180 248892
rect 376236 240324 376292 271180
rect 376236 240258 376292 240268
rect 376684 239540 376740 239550
rect 376684 239316 376740 239484
rect 376684 239250 376740 239260
rect 376236 225316 376292 225326
rect 376236 220500 376292 225260
rect 376236 220434 376292 220444
rect 376236 219156 376292 219166
rect 376236 213332 376292 219100
rect 376236 213266 376292 213276
rect 376236 205044 376292 205054
rect 376236 190148 376292 204988
rect 376908 202692 376964 289772
rect 377356 269780 377412 269790
rect 377356 243348 377412 269724
rect 377244 241332 377300 241342
rect 377132 239316 377188 239326
rect 376908 202626 376964 202636
rect 377020 236628 377076 236638
rect 376236 190082 376292 190092
rect 376124 97748 376180 132188
rect 376236 172004 376292 172014
rect 376236 98868 376292 171948
rect 377020 167300 377076 236572
rect 377020 167234 377076 167244
rect 377132 166628 377188 239260
rect 377132 166562 377188 166572
rect 377244 165956 377300 241276
rect 377244 164724 377300 165900
rect 377244 164658 377300 164668
rect 377356 164612 377412 243292
rect 377356 164546 377412 164556
rect 377468 246708 377524 246718
rect 377468 163268 377524 246652
rect 377468 163202 377524 163212
rect 377580 244020 377636 244030
rect 377580 160580 377636 243964
rect 377692 227892 377748 314636
rect 377916 303268 377972 324268
rect 377916 303202 377972 303212
rect 377692 227826 377748 227836
rect 377804 290500 377860 290510
rect 377804 202468 377860 290444
rect 377916 283780 377972 283790
rect 377916 276388 377972 283724
rect 377916 276322 377972 276332
rect 378028 235172 378084 235182
rect 376348 160244 376404 160254
rect 376348 156548 376404 160188
rect 377356 159908 377412 159918
rect 376348 156482 376404 156492
rect 377020 157892 377076 157902
rect 376796 153972 376852 153982
rect 376796 153188 376852 153916
rect 376796 153122 376852 153132
rect 377020 135604 377076 157836
rect 377132 155204 377188 155214
rect 377132 138964 377188 155148
rect 377244 153860 377300 153870
rect 377244 141092 377300 153804
rect 377244 140084 377300 141036
rect 377244 140018 377300 140028
rect 377132 138898 377188 138908
rect 377020 134708 377076 135548
rect 377020 134642 377076 134652
rect 377356 135940 377412 159852
rect 377468 159572 377524 159582
rect 377468 159124 377524 159516
rect 377468 154532 377524 159068
rect 377468 154466 377524 154476
rect 377468 153188 377524 153198
rect 377468 141204 377524 153132
rect 377468 141138 377524 141148
rect 377356 134484 377412 135884
rect 377356 134418 377412 134428
rect 377580 133476 377636 160524
rect 377580 133410 377636 133420
rect 377692 163268 377748 163278
rect 377468 132132 377524 132142
rect 376236 98802 376292 98812
rect 376348 130788 376404 130798
rect 376124 97682 376180 97692
rect 376348 95284 376404 130732
rect 377132 128884 377188 128894
rect 377020 98644 377076 98654
rect 376348 95218 376404 95228
rect 376460 96628 376516 96638
rect 376012 90692 376068 91420
rect 376012 90626 376068 90636
rect 376460 82964 376516 96572
rect 376460 82898 376516 82908
rect 375900 63186 375956 63196
rect 376236 70532 376292 70542
rect 376236 52724 376292 70476
rect 377020 65940 377076 98588
rect 377132 71988 377188 128828
rect 377244 128660 377300 128670
rect 377244 127204 377300 128604
rect 377244 127138 377300 127148
rect 377356 99764 377412 99774
rect 377356 99204 377412 99708
rect 377132 71922 377188 71932
rect 377244 84756 377300 84766
rect 377244 70532 377300 84700
rect 377244 70466 377300 70476
rect 377356 66612 377412 99148
rect 377468 96404 377524 132076
rect 377580 131684 377636 131694
rect 377580 130900 377636 131628
rect 377692 131572 377748 163212
rect 377804 157892 377860 202412
rect 377804 157220 377860 157836
rect 377804 157154 377860 157164
rect 377916 202692 377972 202702
rect 377916 202132 377972 202636
rect 377916 155876 377972 202076
rect 377916 136724 377972 155820
rect 377916 136658 377972 136668
rect 377916 135380 377972 135390
rect 377916 134372 377972 135324
rect 377916 134306 377972 134316
rect 378028 132132 378084 235116
rect 378588 222740 378644 326172
rect 389452 324968 389508 327628
rect 392140 326004 392196 326014
rect 392140 324968 392196 325948
rect 392812 324968 392868 327740
rect 408268 327796 408324 327806
rect 406252 326340 406308 326350
rect 397516 326228 397572 326238
rect 397516 324968 397572 326172
rect 398188 326004 398244 326014
rect 398188 324968 398244 325948
rect 406252 324968 406308 326284
rect 406924 326116 406980 326126
rect 406924 324968 406980 326060
rect 408268 324968 408324 327740
rect 408940 324968 408996 328076
rect 419692 328020 419748 328030
rect 409612 327908 409668 327918
rect 409612 324968 409668 327852
rect 417004 326228 417060 326238
rect 414306 324940 414316 324996
rect 414372 324940 414382 324996
rect 417004 324968 417060 326172
rect 417676 326116 417732 326126
rect 417676 324968 417732 326060
rect 419692 324968 419748 327964
rect 421036 327796 421092 327806
rect 421036 324968 421092 327740
rect 421708 327684 421764 327694
rect 421708 324968 421764 327628
rect 440300 326004 440356 326014
rect 423948 324996 424004 325006
rect 424004 324940 424424 324996
rect 423948 324930 424004 324940
rect 390124 324548 390180 324558
rect 390124 324482 390180 324492
rect 396844 324548 396900 324558
rect 396844 324482 396900 324492
rect 410956 324436 411012 324446
rect 410312 324380 410956 324436
rect 410956 324370 411012 324380
rect 418348 324436 418404 324446
rect 418348 324370 418404 324380
rect 418796 324436 418852 324446
rect 420812 324436 420868 324446
rect 418852 324380 419048 324436
rect 420392 324380 420812 324436
rect 418796 324370 418852 324380
rect 420812 324370 420868 324380
rect 422044 324436 422100 324446
rect 422604 324436 422660 324446
rect 424172 324436 424228 324446
rect 422100 324380 422408 324436
rect 422660 324380 423080 324436
rect 423752 324380 424172 324436
rect 422044 324370 422100 324380
rect 422604 324370 422660 324380
rect 424172 324370 424228 324380
rect 425068 324436 425124 324446
rect 426188 324436 426244 324446
rect 425768 324380 426188 324436
rect 425068 324370 425124 324380
rect 426188 324370 426244 324380
rect 426412 324436 426468 324446
rect 426412 324370 426468 324380
rect 440188 309988 440244 309998
rect 439292 305844 439348 305854
rect 379260 288484 379316 288494
rect 379148 287812 379204 287822
rect 378924 287140 378980 287150
rect 378812 261604 378868 261614
rect 378812 239428 378868 261548
rect 378812 239362 378868 239372
rect 378588 221844 378644 222684
rect 378812 227892 378868 227902
rect 378588 221778 378644 221788
rect 378700 222628 378756 222638
rect 378700 180740 378756 222572
rect 378700 180674 378756 180684
rect 378028 132066 378084 132076
rect 378140 163940 378196 163950
rect 377692 131506 377748 131516
rect 377804 132020 377860 132030
rect 377580 130834 377636 130844
rect 377804 130788 377860 131964
rect 377804 130722 377860 130732
rect 377916 131908 377972 131918
rect 377916 130676 377972 131852
rect 377916 130610 377972 130620
rect 377916 128772 377972 128782
rect 377916 127652 377972 128716
rect 377916 127586 377972 127596
rect 378028 127988 378084 127998
rect 377804 127540 377860 127550
rect 377692 124628 377748 124638
rect 377692 124404 377748 124572
rect 377468 96338 377524 96348
rect 377580 100884 377636 100894
rect 377356 66546 377412 66556
rect 377020 65874 377076 65884
rect 377580 65268 377636 100828
rect 377692 74004 377748 124348
rect 377692 73938 377748 73948
rect 377804 73332 377860 127484
rect 378028 127428 378084 127932
rect 377804 73266 377860 73276
rect 377916 127372 378084 127428
rect 377916 70644 377972 127372
rect 378140 122164 378196 163884
rect 378252 157780 378308 157790
rect 378252 157444 378308 157724
rect 378252 139412 378308 157388
rect 378252 139346 378308 139356
rect 378700 149380 378756 149390
rect 378700 149044 378756 149324
rect 378700 135492 378756 148988
rect 378812 145124 378868 227836
rect 378924 207396 378980 287084
rect 378924 207330 378980 207340
rect 379036 284452 379092 284462
rect 379036 204596 379092 284396
rect 379148 205380 379204 287756
rect 379148 205314 379204 205324
rect 379036 204530 379092 204540
rect 379260 204260 379316 288428
rect 379932 271796 379988 271806
rect 379484 264516 379540 264526
rect 379260 204194 379316 204204
rect 379372 263396 379428 263406
rect 379260 203924 379316 203934
rect 379036 197428 379092 197438
rect 378924 171444 378980 171454
rect 378924 147924 378980 171388
rect 379036 161252 379092 197372
rect 379036 161186 379092 161196
rect 379148 196308 379204 196318
rect 378924 147858 378980 147868
rect 378812 144564 378868 145068
rect 378812 144498 378868 144508
rect 378700 135426 378756 135436
rect 378812 141092 378868 141102
rect 378140 121044 378196 122108
rect 378140 120978 378196 120988
rect 378700 125300 378756 125310
rect 378700 107604 378756 125244
rect 378700 107538 378756 107548
rect 377916 70578 377972 70588
rect 377580 65202 377636 65212
rect 376236 52658 376292 52668
rect 375564 44706 375620 44716
rect 378812 43092 378868 141036
rect 378924 139412 378980 139422
rect 378924 137844 378980 139356
rect 378924 44884 378980 137788
rect 379148 134148 379204 196252
rect 379260 135268 379316 203868
rect 379372 172676 379428 263340
rect 379372 171444 379428 172620
rect 379484 172004 379540 264460
rect 379596 263620 379652 263630
rect 379596 246708 379652 263564
rect 379596 246642 379652 246652
rect 379820 263172 379876 263182
rect 379820 244020 379876 263116
rect 379820 243954 379876 243964
rect 379932 241220 379988 271740
rect 380044 271236 380100 275128
rect 380044 271170 380100 271180
rect 380716 271012 380772 275128
rect 381388 271460 381444 275128
rect 381388 271394 381444 271404
rect 380716 270946 380772 270956
rect 381388 271124 381444 271134
rect 381388 269892 381444 271068
rect 382060 270788 382116 275128
rect 382732 270900 382788 275128
rect 383404 271572 383460 275128
rect 383404 271506 383460 271516
rect 384076 271348 384132 275128
rect 384076 271282 384132 271292
rect 382732 270834 382788 270844
rect 382060 270722 382116 270732
rect 381388 269826 381444 269836
rect 384748 268436 384804 275128
rect 385420 272132 385476 275128
rect 385420 272066 385476 272076
rect 384748 268370 384804 268380
rect 386092 268212 386148 275128
rect 386764 268548 386820 275128
rect 387436 269556 387492 275128
rect 387436 269490 387492 269500
rect 386764 268482 386820 268492
rect 388108 268324 388164 275128
rect 388108 268258 388164 268268
rect 386092 268146 386148 268156
rect 379932 241154 379988 241164
rect 380044 267988 380100 267998
rect 379820 240324 379876 240334
rect 379708 234388 379764 234398
rect 379708 202244 379764 234332
rect 379820 205716 379876 240268
rect 380044 236852 380100 267932
rect 380268 266980 380324 266990
rect 380156 263508 380212 263518
rect 380156 243236 380212 263452
rect 380156 243170 380212 243180
rect 380268 237636 380324 266924
rect 388780 265076 388836 275128
rect 389452 271124 389508 275128
rect 390124 272132 390180 275128
rect 390124 271460 390180 272076
rect 394156 271572 394212 275128
rect 394156 271506 394212 271516
rect 390124 271394 390180 271404
rect 389452 271058 389508 271068
rect 401548 270116 401604 275128
rect 401548 270050 401604 270060
rect 404236 269892 404292 269902
rect 403564 267540 403620 267550
rect 403564 265748 403620 267484
rect 403564 265682 403620 265692
rect 388780 265010 388836 265020
rect 404236 264936 404292 269836
rect 405132 269892 405188 269902
rect 404908 264516 404964 264526
rect 405132 264516 405188 269836
rect 405580 267988 405636 275128
rect 406252 272020 406308 275128
rect 406252 271954 406308 271964
rect 406476 273252 406532 273262
rect 405580 267922 405636 267932
rect 405580 267428 405636 267438
rect 405580 264936 405636 267372
rect 406476 264516 406532 273196
rect 406924 268100 406980 275128
rect 407596 273364 407652 275128
rect 408268 273476 408324 275128
rect 408268 273410 408324 273420
rect 407596 273298 407652 273308
rect 408940 270228 408996 275128
rect 409612 271684 409668 275128
rect 409612 271618 409668 271628
rect 410060 275100 410312 275156
rect 410060 271124 410116 275100
rect 410060 271058 410116 271068
rect 410284 273364 410340 273374
rect 408940 270162 408996 270172
rect 409836 271012 409892 271022
rect 406924 268034 406980 268044
rect 409612 267988 409668 267998
rect 408716 267764 408772 267774
rect 407596 265412 407652 265422
rect 407596 264936 407652 265356
rect 408716 264964 408772 267708
rect 408296 264908 408772 264964
rect 408940 267316 408996 267326
rect 408940 264936 408996 267260
rect 409612 264936 409668 267932
rect 409836 267764 409892 270956
rect 409836 267698 409892 267708
rect 410284 265412 410340 273308
rect 410956 271236 411012 275128
rect 410956 271170 411012 271180
rect 410956 270340 411012 270350
rect 410956 265748 411012 270284
rect 411628 269780 411684 275128
rect 412300 271124 412356 275128
rect 412972 271908 413028 275128
rect 413644 273588 413700 275128
rect 413644 273522 413700 273532
rect 412972 271842 413028 271852
rect 412300 271058 412356 271068
rect 414316 271124 414372 275128
rect 414316 271058 414372 271068
rect 414988 270228 415044 275128
rect 415660 271124 415716 275128
rect 416332 271684 416388 275128
rect 417004 271796 417060 275128
rect 417004 271730 417060 271740
rect 417452 271796 417508 271806
rect 416332 271618 416388 271628
rect 415660 271058 415716 271068
rect 414988 270162 415044 270172
rect 411628 269714 411684 269724
rect 415660 270004 415716 270014
rect 414988 267764 415044 267774
rect 410956 265682 411012 265692
rect 412972 266868 413028 266878
rect 410284 264936 410340 265356
rect 412300 265636 412356 265646
rect 411628 265300 411684 265310
rect 411628 264936 411684 265244
rect 412300 264936 412356 265580
rect 412972 264936 413028 266812
rect 414316 265524 414372 265534
rect 414316 264936 414372 265468
rect 414988 264936 415044 267708
rect 415660 264936 415716 269948
rect 417452 267652 417508 271740
rect 416332 267204 416388 267214
rect 416332 264936 416388 267148
rect 417452 264964 417508 267596
rect 417676 266980 417732 275128
rect 419692 271124 419748 275128
rect 419692 271058 419748 271068
rect 419916 271684 419972 271694
rect 417676 266914 417732 266924
rect 418348 268100 418404 268110
rect 417452 264908 417704 264964
rect 418348 264936 418404 268044
rect 419916 267988 419972 271628
rect 420364 270340 420420 270350
rect 419916 267922 419972 267932
rect 420028 268772 420084 268782
rect 420028 266644 420084 268716
rect 420028 266578 420084 266588
rect 420364 267204 420420 270284
rect 423052 267540 423108 275128
rect 430444 268772 430500 268782
rect 423052 267474 423108 267484
rect 429772 267876 429828 267886
rect 420364 264936 420420 267148
rect 423388 267428 423444 267438
rect 404964 264460 405188 264516
rect 406280 264488 406532 264516
rect 406252 264460 406532 264488
rect 417004 264516 417060 264526
rect 404908 264450 404964 264460
rect 406252 264404 406308 264460
rect 417004 264450 417060 264460
rect 423388 264516 423444 267372
rect 429772 264936 429828 267820
rect 430444 264936 430500 268716
rect 439292 264740 439348 305788
rect 440188 273028 440244 309932
rect 440188 272962 440244 272972
rect 439292 264674 439348 264684
rect 440188 268100 440244 268110
rect 423388 264450 423444 264460
rect 406252 264338 406308 264348
rect 403564 264292 403620 264302
rect 403564 264226 403620 264236
rect 406252 264292 406308 264302
rect 406252 264226 406308 264236
rect 406924 264292 406980 264302
rect 406924 264226 406980 264236
rect 410956 264292 411012 264302
rect 410956 264226 411012 264236
rect 413644 264292 413700 264302
rect 413644 264226 413700 264236
rect 380268 237570 380324 237580
rect 380492 242228 380548 242238
rect 380044 236786 380100 236796
rect 379932 221732 379988 221742
rect 379932 218372 379988 221676
rect 379932 218306 379988 218316
rect 380380 215348 380436 215358
rect 379820 205688 380072 205716
rect 379820 205660 380100 205688
rect 379708 202178 379764 202188
rect 379484 171938 379540 171948
rect 379596 198548 379652 198558
rect 379372 171378 379428 171388
rect 379260 135202 379316 135212
rect 379484 159236 379540 159246
rect 379148 134082 379204 134092
rect 378924 44818 378980 44828
rect 379036 132356 379092 132366
rect 379036 93044 379092 132300
rect 379372 131796 379428 131806
rect 379148 123956 379204 123966
rect 379148 99204 379204 123900
rect 379260 122052 379316 122062
rect 379260 104132 379316 121996
rect 379260 104066 379316 104076
rect 379148 99138 379204 99148
rect 379260 96404 379316 96414
rect 378812 43026 378868 43036
rect 379036 42756 379092 92988
rect 379148 95060 379204 95070
rect 379148 44324 379204 95004
rect 379260 46340 379316 96348
rect 379260 46274 379316 46284
rect 379372 91924 379428 131740
rect 379484 125524 379540 159180
rect 379596 134260 379652 198492
rect 379932 196196 379988 196206
rect 379932 176372 379988 196140
rect 379932 176306 379988 176316
rect 379596 134194 379652 134204
rect 379708 167300 379764 167310
rect 379708 127540 379764 167244
rect 379708 127474 379764 127484
rect 379820 165284 379876 165294
rect 379484 125458 379540 125468
rect 379820 124404 379876 165228
rect 380044 161308 380100 205660
rect 379932 161252 380100 161308
rect 380268 198436 380324 198446
rect 379932 155540 379988 161252
rect 379932 155474 379988 155484
rect 380156 146244 380212 146254
rect 380156 138964 380212 146188
rect 380268 144508 380324 198380
rect 380380 197540 380436 215292
rect 380492 201460 380548 242172
rect 380604 240436 380660 240446
rect 380604 215068 380660 240380
rect 380604 215012 380884 215068
rect 380828 211708 380884 215012
rect 380828 211652 380996 211708
rect 380940 205380 380996 211652
rect 381836 205716 381892 205726
rect 381836 205380 381892 205660
rect 382060 205716 382116 205726
rect 382060 205650 382116 205660
rect 383404 205716 383460 205726
rect 384748 205716 384804 205726
rect 383460 205660 383684 205716
rect 383404 205650 383460 205660
rect 380744 205352 380996 205380
rect 381416 205352 381892 205380
rect 380492 201394 380548 201404
rect 380716 205324 380996 205352
rect 381388 205324 381892 205352
rect 380380 197474 380436 197484
rect 380716 196588 380772 205324
rect 381388 203028 381444 205324
rect 382620 203252 382676 203262
rect 382732 203252 382788 205128
rect 382676 203196 382788 203252
rect 383628 203252 383684 205660
rect 384748 205650 384804 205660
rect 384076 205492 384132 205502
rect 384076 205426 384132 205436
rect 417004 205492 417060 205502
rect 417004 205426 417060 205436
rect 419244 205380 419300 205390
rect 419300 205352 419720 205380
rect 419300 205324 419748 205352
rect 419244 205314 419300 205324
rect 385420 205268 385476 205278
rect 382620 203186 382676 203196
rect 383628 203186 383684 203196
rect 384972 205212 385420 205268
rect 381388 202962 381444 202972
rect 384188 202804 384244 202814
rect 384636 202804 384692 202814
rect 384244 202748 384636 202804
rect 384188 202738 384244 202748
rect 384636 202738 384692 202748
rect 384636 202468 384692 202478
rect 384636 202132 384692 202412
rect 384636 202066 384692 202076
rect 384972 198436 385028 205212
rect 385420 205202 385476 205212
rect 386092 205268 386148 205278
rect 386092 198548 386148 205212
rect 386764 205268 386820 205278
rect 386092 198482 386148 198492
rect 386428 203140 386484 203150
rect 384972 198370 385028 198380
rect 380604 196532 380772 196588
rect 380604 144508 380660 196532
rect 386428 196084 386484 203084
rect 386764 198324 386820 205212
rect 389452 205268 389508 205278
rect 387436 203140 387492 205128
rect 387436 203074 387492 203084
rect 388108 201460 388164 205128
rect 388108 201394 388164 201404
rect 388220 203252 388276 203262
rect 386764 198258 386820 198268
rect 388220 196308 388276 203196
rect 388444 201348 388500 201358
rect 388444 196420 388500 201292
rect 388780 201348 388836 205128
rect 389452 203252 389508 205212
rect 399532 205156 399588 205166
rect 389452 203186 389508 203196
rect 389788 205100 390152 205156
rect 403340 205156 403396 205166
rect 388780 201282 388836 201292
rect 388444 196354 388500 196364
rect 389788 198100 389844 205100
rect 399532 205090 399588 205100
rect 391468 205044 391524 205054
rect 390460 202804 390516 202814
rect 390908 202804 390964 202814
rect 390516 202748 390908 202804
rect 390460 202738 390516 202748
rect 390908 202738 390964 202748
rect 391468 201236 391524 204988
rect 402220 203924 402276 205128
rect 400204 202804 400260 202814
rect 391468 201170 391524 201180
rect 398188 201684 398244 201694
rect 388220 196242 388276 196252
rect 389788 196196 389844 198044
rect 389788 196130 389844 196140
rect 386428 196018 386484 196028
rect 398188 194628 398244 201628
rect 400204 194936 400260 202748
rect 402220 201908 402276 203868
rect 402220 201842 402276 201852
rect 410956 205156 411012 205166
rect 403340 197092 403396 205100
rect 404908 201684 404964 205128
rect 406924 204484 406980 205128
rect 406924 204418 406980 204428
rect 407596 205044 407652 205054
rect 404908 201460 404964 201628
rect 404908 201394 404964 201404
rect 403340 197026 403396 197036
rect 403564 197876 403620 197886
rect 403564 194936 403620 197820
rect 405580 197764 405636 197774
rect 405580 194936 405636 197708
rect 407596 194936 407652 204988
rect 408268 204932 408324 205128
rect 408268 204866 408324 204876
rect 408940 204372 408996 205128
rect 410284 204708 410340 205128
rect 410284 204642 410340 204652
rect 413644 205156 413700 205166
rect 408940 204306 408996 204316
rect 408940 199556 408996 199566
rect 408940 194936 408996 199500
rect 410284 199444 410340 199454
rect 409612 197652 409668 197662
rect 409612 194936 409668 197596
rect 410284 194936 410340 199388
rect 410956 199444 411012 205100
rect 411628 202692 411684 205128
rect 412300 204820 412356 205128
rect 412300 204754 412356 204764
rect 412972 202916 413028 205128
rect 413644 205090 413700 205100
rect 412972 202850 413028 202860
rect 414316 204596 414372 205128
rect 411628 202626 411684 202636
rect 414316 202468 414372 204540
rect 414316 202402 414372 202412
rect 414764 205044 414820 205054
rect 410956 199378 411012 199388
rect 411628 201236 411684 201246
rect 410956 197092 411012 197102
rect 410956 194936 411012 197036
rect 411628 194936 411684 201180
rect 413420 201012 413476 201022
rect 412300 197988 412356 197998
rect 412300 194936 412356 197932
rect 413420 194852 413476 200956
rect 414764 199556 414820 204988
rect 414988 202916 415044 205128
rect 415660 204036 415716 205128
rect 415660 203970 415716 203980
rect 416332 203028 416388 205128
rect 416332 202962 416388 202972
rect 416668 204260 416724 204270
rect 416668 203028 416724 204204
rect 416668 202962 416724 202972
rect 414988 202850 415044 202860
rect 416556 202916 416612 202926
rect 416556 199668 416612 202860
rect 417676 202580 417732 205128
rect 418348 204372 418404 205128
rect 418572 205044 418628 205054
rect 418348 204316 418516 204372
rect 418348 204148 418404 204158
rect 418348 203252 418404 204092
rect 418348 203186 418404 203196
rect 417676 202514 417732 202524
rect 418460 202356 418516 204316
rect 418572 203140 418628 204988
rect 418572 203074 418628 203084
rect 418460 202290 418516 202300
rect 419020 202244 419076 205128
rect 419692 204260 419748 205324
rect 419692 204194 419748 204204
rect 423052 203028 423108 205128
rect 423052 202692 423108 202972
rect 423052 202626 423108 202636
rect 427084 203252 427140 205128
rect 427084 202580 427140 203196
rect 427084 202514 427140 202524
rect 429772 203140 429828 205128
rect 419020 202178 419076 202188
rect 429772 201684 429828 203084
rect 429772 201618 429828 201628
rect 416556 199602 416612 199612
rect 417676 201124 417732 201134
rect 414764 199490 414820 199500
rect 417004 199332 417060 199342
rect 416332 197540 416388 197550
rect 416332 194936 416388 197484
rect 417004 194936 417060 199276
rect 417676 194936 417732 201068
rect 439404 199444 439460 199454
rect 418348 198212 418404 198222
rect 418348 194936 418404 198156
rect 423500 194852 423556 194862
rect 413420 194796 413672 194852
rect 398188 194562 398244 194572
rect 423500 194628 423556 194796
rect 423500 194562 423556 194572
rect 380268 144452 380436 144508
rect 380604 144452 380884 144508
rect 380156 138908 380324 138964
rect 380044 137508 380100 137518
rect 380044 132468 380100 137452
rect 380044 132402 380100 132412
rect 380268 126028 380324 138908
rect 380380 136724 380436 144452
rect 380828 141148 380884 144452
rect 380828 141092 380996 141148
rect 380380 136658 380436 136668
rect 380492 138964 380548 138974
rect 379820 124338 379876 124348
rect 380156 125972 380324 126028
rect 380380 127204 380436 127214
rect 379484 123844 379540 123854
rect 379484 105364 379540 123788
rect 379484 105298 379540 105308
rect 379596 121044 379652 121054
rect 379148 44258 379204 44268
rect 379372 43204 379428 91868
rect 379484 95284 379540 95294
rect 379484 46228 379540 95228
rect 379596 82068 379652 120988
rect 379596 82002 379652 82012
rect 380156 67228 380212 125972
rect 380268 123732 380324 123742
rect 380268 106484 380324 123676
rect 380268 106418 380324 106428
rect 380380 100884 380436 127148
rect 380380 100818 380436 100828
rect 380380 97748 380436 97758
rect 380156 67172 380324 67228
rect 379484 46162 379540 46172
rect 379820 65604 379876 65614
rect 379820 45780 379876 65548
rect 379820 45724 380072 45780
rect 380268 44660 380324 67172
rect 380268 44594 380324 44604
rect 379372 43138 379428 43148
rect 380380 42980 380436 97692
rect 380492 46004 380548 138908
rect 380716 135716 380772 135726
rect 380716 135650 380772 135660
rect 380940 135716 380996 141092
rect 380940 129388 380996 135660
rect 381388 136052 381444 136062
rect 381388 132692 381444 135996
rect 382060 135716 382116 135726
rect 381388 132626 381444 132636
rect 381836 135660 382060 135716
rect 381836 132692 381892 135660
rect 382060 135650 382116 135660
rect 383628 135716 383684 135726
rect 385420 135716 385476 135726
rect 383628 135268 383684 135660
rect 384972 135660 385420 135716
rect 383432 135240 383684 135268
rect 383404 135212 383684 135240
rect 384748 135268 384804 135278
rect 382732 134820 382788 135128
rect 382732 134754 382788 134764
rect 381836 132626 381892 132636
rect 383404 132692 383460 135212
rect 384748 135202 384804 135212
rect 383404 132626 383460 132636
rect 384076 132580 384132 135128
rect 384076 132514 384132 132524
rect 384972 132580 385028 135660
rect 385420 135650 385476 135660
rect 388780 135716 388836 135726
rect 388780 135650 388836 135660
rect 396844 135716 396900 135726
rect 396844 135650 396900 135660
rect 397516 135716 397572 135726
rect 397516 135650 397572 135660
rect 398188 135156 398244 135166
rect 384972 132514 385028 132524
rect 385644 134260 385700 134270
rect 385644 132580 385700 134204
rect 386092 134260 386148 135128
rect 386092 134194 386148 134204
rect 385644 132514 385700 132524
rect 386428 134148 386484 134158
rect 381724 132468 381780 132478
rect 381724 132132 381780 132412
rect 381724 132066 381780 132076
rect 384524 132244 384580 132254
rect 384524 131684 384580 132188
rect 384524 131618 384580 131628
rect 386428 131684 386484 134092
rect 386764 134148 386820 135128
rect 386764 134082 386820 134092
rect 386540 133924 386596 133934
rect 386540 132580 386596 133868
rect 387436 133924 387492 135128
rect 387436 133858 387492 133868
rect 388108 134372 388164 135128
rect 386540 132514 386596 132524
rect 386428 131618 386484 131628
rect 380716 129332 380996 129388
rect 380716 126028 380772 129332
rect 388108 129220 388164 134316
rect 389452 134036 389508 135128
rect 389452 131460 389508 133980
rect 389452 131394 389508 131404
rect 398188 134932 398244 135100
rect 398188 131124 398244 134876
rect 398188 131058 398244 131068
rect 404236 131796 404292 135128
rect 388108 129154 388164 129164
rect 380604 125972 380772 126028
rect 382172 129108 382228 129118
rect 380604 67508 380660 125972
rect 382172 122276 382228 129052
rect 404236 129108 404292 131740
rect 409612 129332 409668 135128
rect 410284 132132 410340 135128
rect 410956 132244 411012 135128
rect 410956 132178 411012 132188
rect 410284 132066 410340 132076
rect 411628 132020 411684 135128
rect 412300 132468 412356 135128
rect 412300 132402 412356 132412
rect 412972 132356 413028 135128
rect 412972 132290 413028 132300
rect 411628 131954 411684 131964
rect 413644 131908 413700 135128
rect 414316 132580 414372 135128
rect 414316 132514 414372 132524
rect 414876 132692 414932 132702
rect 413644 131842 413700 131852
rect 409612 129266 409668 129276
rect 411516 131684 411572 131694
rect 404236 129042 404292 129052
rect 411516 127204 411572 131628
rect 411516 127138 411572 127148
rect 414092 131236 414148 131246
rect 414092 123956 414148 131180
rect 414876 128996 414932 132636
rect 414988 132468 415044 135128
rect 414988 131236 415044 132412
rect 415660 132580 415716 135128
rect 415660 131684 415716 132524
rect 415660 131618 415716 131628
rect 416332 132244 416388 135128
rect 414988 131170 415044 131180
rect 414876 128930 414932 128940
rect 414092 123890 414148 123900
rect 382172 122210 382228 122220
rect 416332 122052 416388 132188
rect 417004 132132 417060 135128
rect 417004 132066 417060 132076
rect 417452 135100 417704 135156
rect 417452 132356 417508 135100
rect 418348 132692 418404 135128
rect 418348 132626 418404 132636
rect 419020 134260 419076 135128
rect 417452 123844 417508 132300
rect 417900 132132 417956 132142
rect 417900 125412 417956 132076
rect 419020 126028 419076 134204
rect 419244 135100 419720 135156
rect 419244 132020 419300 135100
rect 439404 132580 439460 199388
rect 439404 132514 439460 132524
rect 419020 125972 419188 126028
rect 417900 125346 417956 125356
rect 417452 123778 417508 123788
rect 419132 123732 419188 125972
rect 419244 125300 419300 131964
rect 440188 131796 440244 268044
rect 440300 201460 440356 325948
rect 441980 310660 442036 310670
rect 441868 307300 441924 307310
rect 440524 276388 440580 276398
rect 440300 201394 440356 201404
rect 440412 267988 440468 267998
rect 440188 131730 440244 131740
rect 440300 196756 440356 196766
rect 419244 125234 419300 125244
rect 419132 123666 419188 123676
rect 416332 121986 416388 121996
rect 440300 83412 440356 196700
rect 440412 161924 440468 267932
rect 440524 202916 440580 276332
rect 441868 270452 441924 307244
rect 441980 274708 442036 310604
rect 442092 309316 442148 309326
rect 442092 275604 442148 309260
rect 442092 275538 442148 275548
rect 441980 274642 442036 274652
rect 441868 270386 441924 270396
rect 445228 267764 445284 267774
rect 442316 267316 442372 267326
rect 441980 265412 442036 265422
rect 440524 202850 440580 202860
rect 440636 205604 440692 205614
rect 440412 161858 440468 161868
rect 440524 202580 440580 202590
rect 440300 83346 440356 83356
rect 440412 136948 440468 136958
rect 440412 81396 440468 136892
rect 440524 134260 440580 202524
rect 440636 172004 440692 205548
rect 441868 194516 441924 194526
rect 441868 177380 441924 194460
rect 441868 177314 441924 177324
rect 440636 171938 440692 171948
rect 441980 163268 442036 265356
rect 442204 228564 442260 228574
rect 442092 226548 442148 226558
rect 442092 201572 442148 226492
rect 442204 206612 442260 228508
rect 442316 208348 442372 267260
rect 443660 266868 443716 266878
rect 443548 263396 443604 263406
rect 442316 208292 442596 208348
rect 442204 206546 442260 206556
rect 442092 201506 442148 201516
rect 442316 193396 442372 193406
rect 442204 191828 442260 191838
rect 442092 191772 442204 191828
rect 442092 170660 442148 191772
rect 442204 191762 442260 191772
rect 442316 191604 442372 193340
rect 442204 191548 442372 191604
rect 442204 172676 442260 191548
rect 442540 190596 442596 208292
rect 442204 172610 442260 172620
rect 442316 190540 442596 190596
rect 442092 170594 442148 170604
rect 441980 163202 442036 163212
rect 442316 162932 442372 190540
rect 442652 164612 442708 164622
rect 442316 162866 442372 162876
rect 442540 163940 442596 163950
rect 442204 161252 442260 161262
rect 442092 159908 442148 159918
rect 441868 157892 441924 157902
rect 441868 135044 441924 157836
rect 442092 137396 442148 159852
rect 442092 137330 442148 137340
rect 442092 137060 442148 137070
rect 441868 134978 441924 134988
rect 441980 135492 442036 135502
rect 441980 134820 442036 135436
rect 440524 134194 440580 134204
rect 441868 134764 442036 134820
rect 440412 81330 440468 81340
rect 380604 67228 380660 67452
rect 380604 67172 380772 67228
rect 380492 45938 380548 45948
rect 380716 45752 380772 67172
rect 441868 66612 441924 134764
rect 442092 126028 442148 137004
rect 442204 134372 442260 161196
rect 442428 160580 442484 160590
rect 442204 134306 442260 134316
rect 442316 159236 442372 159246
rect 442316 130228 442372 159180
rect 442428 135380 442484 160524
rect 442428 135314 442484 135324
rect 442316 130162 442372 130172
rect 441980 125972 442148 126028
rect 442540 125972 442596 163884
rect 442652 137788 442708 164556
rect 442652 137732 443044 137788
rect 442652 137396 442708 137406
rect 442652 128660 442708 137340
rect 442876 135604 442932 135614
rect 442652 128594 442708 128604
rect 442764 133700 442820 133710
rect 441980 69300 442036 125972
rect 442540 125906 442596 125916
rect 442316 125188 442372 125198
rect 442316 87444 442372 125132
rect 442428 123508 442484 123518
rect 442428 89460 442484 123452
rect 442428 89394 442484 89404
rect 442316 87378 442372 87388
rect 441980 69234 442036 69244
rect 442764 68628 442820 133644
rect 442876 69972 442932 135548
rect 442988 128772 443044 137732
rect 442988 128706 443044 128716
rect 443548 124292 443604 263340
rect 443660 137284 443716 266812
rect 443660 137218 443716 137228
rect 443772 191716 443828 191726
rect 443548 124226 443604 124236
rect 443660 128548 443716 128558
rect 443660 75348 443716 128492
rect 443772 76020 443828 191660
rect 445228 135156 445284 267708
rect 445340 263060 445396 263070
rect 445340 137172 445396 263004
rect 448588 196644 448644 196654
rect 446908 195076 446964 195086
rect 445340 137106 445396 137116
rect 445452 194628 445508 194638
rect 445228 135090 445284 135100
rect 445452 77364 445508 194572
rect 445564 193284 445620 193294
rect 445564 78036 445620 193228
rect 446908 78708 446964 195020
rect 448588 84756 448644 196588
rect 448588 84690 448644 84700
rect 446908 78642 446964 78652
rect 445564 77970 445620 77980
rect 445452 77298 445508 77308
rect 443772 75954 443828 75964
rect 443660 75282 443716 75292
rect 442876 69906 442932 69916
rect 457772 69972 457828 69982
rect 442764 68562 442820 68572
rect 441868 66546 441924 66556
rect 457772 47012 457828 69916
rect 457772 46946 457828 46956
rect 381388 45780 381444 45790
rect 381388 45714 381444 45724
rect 382060 45780 382116 45790
rect 382060 45714 382116 45724
rect 384076 45780 384132 45790
rect 384076 45714 384132 45724
rect 384748 45780 384804 45790
rect 384748 45714 384804 45724
rect 388108 45780 388164 45790
rect 388108 45714 388164 45724
rect 396844 45780 396900 45790
rect 396844 45714 396900 45724
rect 398188 45780 398244 45790
rect 398188 45714 398244 45724
rect 403564 45780 403620 45790
rect 403564 45714 403620 45724
rect 417676 45780 417732 45790
rect 417676 45714 417732 45724
rect 390460 45668 390516 45678
rect 390460 45574 390516 45612
rect 397852 45668 397908 45678
rect 397852 45574 397908 45612
rect 418348 45668 418404 45678
rect 418348 45602 418404 45612
rect 382732 45556 382788 45566
rect 383852 45556 383908 45566
rect 383432 45500 383852 45556
rect 382732 45490 382788 45500
rect 383852 45490 383908 45500
rect 384972 45556 385028 45566
rect 386428 45556 386484 45566
rect 386988 45556 387044 45566
rect 389004 45556 389060 45566
rect 391916 45556 391972 45566
rect 412972 45556 413028 45566
rect 385028 45500 385448 45556
rect 386484 45500 386792 45556
rect 387044 45500 387464 45556
rect 389060 45500 389480 45556
rect 391972 45500 392840 45556
rect 384972 45490 385028 45500
rect 386428 45490 386484 45500
rect 386988 45490 387044 45500
rect 389004 45490 389060 45500
rect 391916 45490 391972 45500
rect 412972 45490 413028 45500
rect 388332 45444 388388 45454
rect 407596 45444 407652 45454
rect 388388 45388 388808 45444
rect 388332 45378 388388 45388
rect 407596 45378 407652 45388
rect 386092 45220 386148 45230
rect 386092 45154 386148 45164
rect 405580 45220 405636 45230
rect 405580 45154 405636 45164
rect 402892 45108 402948 45118
rect 380380 42914 380436 42924
rect 396172 42980 396228 45080
rect 398860 44324 398916 45080
rect 398860 44258 398916 44268
rect 396172 42914 396228 42924
rect 379036 42690 379092 42700
rect 399532 42756 399588 45080
rect 400204 43204 400260 45080
rect 400876 43652 400932 45080
rect 416332 45108 416388 45118
rect 402892 45042 402948 45052
rect 400876 43586 400932 43596
rect 404236 43540 404292 45080
rect 406252 44772 406308 45080
rect 406252 44706 406308 44716
rect 406924 44436 406980 45080
rect 406924 44370 406980 44380
rect 404236 43474 404292 43484
rect 400204 43138 400260 43148
rect 399532 42690 399588 42700
rect 374556 41906 374612 41916
rect 372764 41794 372820 41804
rect 408940 40292 408996 45080
rect 409612 41748 409668 45080
rect 410284 42868 410340 45080
rect 410956 44884 411012 45080
rect 410956 44818 411012 44828
rect 413644 42980 413700 45080
rect 414316 43092 414372 45080
rect 415660 43540 415716 45080
rect 485548 45108 485604 45118
rect 416332 45042 416388 45052
rect 415660 43474 415716 43484
rect 417004 43204 417060 45080
rect 419692 43652 419748 45080
rect 419692 43586 419748 43596
rect 420364 43652 420420 45080
rect 420364 43586 420420 43596
rect 421036 43428 421092 45080
rect 421036 43362 421092 43372
rect 422380 43316 422436 45080
rect 423052 44660 423108 45080
rect 423052 44594 423108 44604
rect 422380 43250 422436 43260
rect 417004 43138 417060 43148
rect 414316 43026 414372 43036
rect 413644 42914 413700 42924
rect 410284 42802 410340 42812
rect 423724 41860 423780 45080
rect 484204 43540 484260 45080
rect 484876 43652 484932 45080
rect 485548 45042 485604 45052
rect 484876 43586 484932 43596
rect 484204 43474 484260 43484
rect 511532 43540 511588 377132
rect 540092 350756 540148 350766
rect 511532 43474 511588 43484
rect 512428 69972 512484 69982
rect 512428 41972 512484 69916
rect 512540 69300 512596 69310
rect 512540 45332 512596 69244
rect 512540 45266 512596 45276
rect 540092 43652 540148 350700
rect 573692 337540 573748 337550
rect 573692 45108 573748 337484
rect 573692 45042 573748 45052
rect 540092 43586 540148 43596
rect 512428 41906 512484 41916
rect 423724 41794 423780 41804
rect 409612 41682 409668 41692
rect 408940 40226 408996 40236
rect 4284 8754 4340 8764
rect 396396 5572 396452 5582
rect 395976 5516 396396 5572
rect 396396 5506 396452 5516
rect 437612 5572 437668 5582
rect 483084 5572 483140 5582
rect 437668 5516 437892 5572
rect 437612 5506 437668 5516
rect 401324 5460 401380 5470
rect 400680 5404 401324 5460
rect 401324 5394 401380 5404
rect 382508 5348 382564 5358
rect 420140 5348 420196 5358
rect 381864 5292 382508 5348
rect 419496 5292 420140 5348
rect 382508 5282 382564 5292
rect 420140 5282 420196 5292
rect 353612 5236 353668 5246
rect 353612 5170 353668 5180
rect 386652 5236 386708 5246
rect 429548 5236 429604 5246
rect 428904 5180 429548 5236
rect 15372 5124 15428 5134
rect 47852 5124 47908 5134
rect 91756 5124 91812 5134
rect 333228 5124 333284 5134
rect 361676 5124 361732 5134
rect 367724 5124 367780 5134
rect 11564 480 11732 532
rect 13468 480 13636 532
rect 15372 480 15428 5068
rect 28700 5012 28756 5022
rect 21084 3444 21140 3454
rect 19180 2660 19236 2670
rect 17276 2548 17332 2558
rect 17276 480 17332 2492
rect 19180 480 19236 2604
rect 21084 480 21140 3388
rect 26796 2884 26852 2894
rect 24892 2772 24948 2782
rect 22988 480 23156 532
rect 24892 480 24948 2716
rect 26796 480 26852 2828
rect 28700 480 28756 4956
rect 30604 4900 30660 4910
rect 30604 480 30660 4844
rect 40124 4788 40180 4798
rect 36316 3220 36372 3230
rect 34412 3108 34468 3118
rect 32508 2996 32564 3006
rect 32508 480 32564 2940
rect 34412 480 34468 3052
rect 36316 480 36372 3164
rect 38220 2212 38276 2222
rect 38220 480 38276 2156
rect 40124 480 40180 4732
rect 43932 4676 43988 4686
rect 41916 2436 41972 2446
rect 41916 480 41972 2380
rect 43932 480 43988 4620
rect 11368 476 11732 480
rect 11368 392 11620 476
rect 11368 -960 11592 392
rect 11676 84 11732 476
rect 11676 18 11732 28
rect 13272 476 13636 480
rect 13272 392 13524 476
rect 13272 -960 13496 392
rect 13580 196 13636 476
rect 13580 130 13636 140
rect 15176 392 15428 480
rect 17080 392 17332 480
rect 18984 392 19236 480
rect 20888 392 21140 480
rect 22792 476 23156 480
rect 22792 392 23044 476
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 18984 -960 19208 392
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 23100 308 23156 476
rect 23100 242 23156 252
rect 24696 392 24948 480
rect 26600 392 26852 480
rect 28504 392 28756 480
rect 30408 392 30660 480
rect 32312 392 32564 480
rect 34216 392 34468 480
rect 36120 392 36372 480
rect 38024 392 38276 480
rect 39928 392 40180 480
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 392
rect 30408 -960 30632 392
rect 32312 -960 32536 392
rect 34216 -960 34440 392
rect 36120 -960 36344 392
rect 38024 -960 38248 392
rect 39928 -960 40152 392
rect 41832 -960 42056 480
rect 43736 392 43988 480
rect 43736 -960 43960 392
rect 44716 84 44772 5096
rect 45836 4564 45892 4574
rect 45836 480 45892 4508
rect 44716 18 44772 28
rect 45640 392 45892 480
rect 45640 -960 45864 392
rect 46284 196 46340 5096
rect 47852 5058 47908 5068
rect 47740 4452 47796 4462
rect 47740 480 47796 4396
rect 49420 2548 49476 5096
rect 50988 2660 51044 5096
rect 51996 5068 52584 5124
rect 50988 2594 51044 2604
rect 51548 4340 51604 4350
rect 49420 2482 49476 2492
rect 49644 2324 49700 2334
rect 49644 480 49700 2268
rect 51548 480 51604 4284
rect 51996 3444 52052 5068
rect 51996 3378 52052 3388
rect 53452 4228 53508 4238
rect 53452 480 53508 4172
rect 46284 130 46340 140
rect 47544 392 47796 480
rect 49448 392 49700 480
rect 51352 392 51604 480
rect 53256 392 53508 480
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51352 -960 51576 392
rect 53256 -960 53480 392
rect 54124 308 54180 5096
rect 55692 2772 55748 5096
rect 57260 2884 57316 5096
rect 58856 5068 58996 5124
rect 58940 5012 58996 5068
rect 58940 4946 58996 4956
rect 60396 4900 60452 5096
rect 60396 4834 60452 4844
rect 57260 2818 57316 2828
rect 57372 4116 57428 4126
rect 55692 2706 55748 2716
rect 55356 2548 55412 2558
rect 55356 480 55412 2492
rect 57372 2100 57428 4060
rect 61068 4004 61124 4014
rect 57260 2044 57428 2100
rect 59164 2660 59220 2670
rect 57260 480 57316 2044
rect 59164 480 59220 2604
rect 61068 480 61124 3948
rect 61964 2996 62020 5096
rect 63532 3108 63588 5096
rect 63532 3042 63588 3052
rect 64876 4900 64932 4910
rect 61964 2930 62020 2940
rect 62972 2772 63028 2782
rect 62972 480 63028 2716
rect 64876 480 64932 4844
rect 65100 3220 65156 5096
rect 65100 3154 65156 3164
rect 66668 2212 66724 5096
rect 68236 4788 68292 5096
rect 68236 4722 68292 4732
rect 68684 5012 68740 5022
rect 66668 2146 66724 2156
rect 66780 2884 66836 2894
rect 66780 480 66836 2828
rect 68684 480 68740 4956
rect 69804 2436 69860 5096
rect 69804 2370 69860 2380
rect 70476 4788 70532 4798
rect 70476 480 70532 4732
rect 71372 4676 71428 5096
rect 71372 4610 71428 4620
rect 72492 4676 72548 4686
rect 72492 480 72548 4620
rect 72940 4564 72996 5096
rect 72940 4498 72996 4508
rect 73052 5012 73108 5022
rect 73052 4004 73108 4956
rect 73052 3938 73108 3948
rect 74396 4564 74452 4574
rect 74396 480 74452 4508
rect 74508 4452 74564 5096
rect 74508 4386 74564 4396
rect 76076 2324 76132 5096
rect 76076 2258 76132 2268
rect 76300 4452 76356 4462
rect 76300 480 76356 4396
rect 77644 4340 77700 5096
rect 77644 4274 77700 4284
rect 78204 4340 78260 4350
rect 78204 480 78260 4284
rect 79212 4228 79268 5096
rect 79212 4162 79268 4172
rect 80108 2996 80164 3006
rect 80108 480 80164 2940
rect 80780 2548 80836 5096
rect 80780 2482 80836 2492
rect 82012 4228 82068 4238
rect 82012 480 82068 4172
rect 82348 4116 82404 5096
rect 82348 4050 82404 4060
rect 83244 5068 83944 5124
rect 84812 5068 85512 5124
rect 83244 2660 83300 5068
rect 84812 5012 84868 5068
rect 84812 4946 84868 4956
rect 85820 5012 85876 5022
rect 83244 2594 83300 2604
rect 83916 4116 83972 4126
rect 83916 480 83972 4060
rect 85820 480 85876 4956
rect 87052 2772 87108 5096
rect 88620 4900 88676 5096
rect 88620 4834 88676 4844
rect 89628 4900 89684 4910
rect 87052 2706 87108 2716
rect 87724 2548 87780 2558
rect 87724 480 87780 2492
rect 89628 480 89684 4844
rect 90188 2884 90244 5096
rect 91756 5058 91812 5068
rect 93324 4788 93380 5096
rect 93324 4722 93380 4732
rect 94892 4676 94948 5096
rect 94892 4610 94948 4620
rect 95340 4788 95396 4798
rect 90188 2818 90244 2828
rect 93436 2772 93492 2782
rect 91532 2660 91588 2670
rect 91532 480 91588 2604
rect 93436 480 93492 2716
rect 95340 480 95396 4732
rect 96460 4564 96516 5096
rect 96460 4498 96516 4508
rect 98028 4452 98084 5096
rect 98028 4386 98084 4396
rect 99036 4676 99092 4686
rect 97244 2884 97300 2894
rect 97244 480 97300 2828
rect 99036 480 99092 4620
rect 99596 4340 99652 5096
rect 99596 4274 99652 4284
rect 101052 4564 101108 4574
rect 101052 480 101108 4508
rect 101164 2996 101220 5096
rect 102732 4228 102788 5096
rect 102732 4162 102788 4172
rect 102956 4452 103012 4462
rect 101164 2930 101220 2940
rect 102956 480 103012 4396
rect 104300 4116 104356 5096
rect 105896 5068 106036 5124
rect 105980 5012 106036 5068
rect 105980 4946 106036 4956
rect 106764 5012 106820 5022
rect 104300 4050 104356 4060
rect 104860 4340 104916 4350
rect 104860 480 104916 4284
rect 106764 480 106820 4956
rect 107436 2548 107492 5096
rect 109004 4900 109060 5096
rect 109004 4834 109060 4844
rect 109900 5068 110600 5124
rect 107436 2482 107492 2492
rect 108668 4228 108724 4238
rect 108668 480 108724 4172
rect 109900 2660 109956 5068
rect 109900 2594 109956 2604
rect 110572 4900 110628 4910
rect 110572 480 110628 4844
rect 112140 2772 112196 5096
rect 113708 4788 113764 5096
rect 113708 4722 113764 4732
rect 112140 2706 112196 2716
rect 112476 4116 112532 4126
rect 112476 480 112532 4060
rect 115276 2884 115332 5096
rect 116844 4676 116900 5096
rect 116844 4610 116900 4620
rect 118412 4564 118468 5096
rect 118412 4498 118468 4508
rect 119980 4452 120036 5096
rect 119980 4386 120036 4396
rect 120092 4788 120148 4798
rect 115276 2818 115332 2828
rect 118188 2772 118244 2782
rect 116284 2660 116340 2670
rect 114380 2548 114436 2558
rect 114380 480 114436 2492
rect 116284 480 116340 2604
rect 118188 480 118244 2716
rect 120092 480 120148 4732
rect 121548 4340 121604 5096
rect 122668 5068 123144 5124
rect 122668 5012 122724 5068
rect 122668 4946 122724 4956
rect 123900 5012 123956 5022
rect 121548 4274 121604 4284
rect 121996 2884 122052 2894
rect 121996 480 122052 2828
rect 123900 480 123956 4956
rect 124684 4228 124740 5096
rect 126252 4900 126308 5096
rect 126252 4834 126308 4844
rect 127596 4900 127652 4910
rect 124684 4162 124740 4172
rect 125804 4676 125860 4686
rect 125804 480 125860 4620
rect 127596 480 127652 4844
rect 127820 4116 127876 5096
rect 127820 4050 127876 4060
rect 129388 2548 129444 5096
rect 129388 2482 129444 2492
rect 129612 4564 129668 4574
rect 129612 480 129668 4508
rect 130956 2660 131012 5096
rect 130956 2594 131012 2604
rect 131516 4452 131572 4462
rect 131516 480 131572 4396
rect 132524 2772 132580 5096
rect 134092 4788 134148 5096
rect 134092 4722 134148 4732
rect 135660 2884 135716 5096
rect 136556 5068 137256 5124
rect 136556 5012 136612 5068
rect 136556 4946 136612 4956
rect 138796 4676 138852 5096
rect 138796 4610 138852 4620
rect 139132 5012 139188 5022
rect 135660 2818 135716 2828
rect 132524 2706 132580 2716
rect 137228 2772 137284 2782
rect 135324 2660 135380 2670
rect 133420 2548 133476 2558
rect 133420 480 133476 2492
rect 135324 480 135380 2604
rect 137228 480 137284 2716
rect 139132 480 139188 4956
rect 140364 4900 140420 5096
rect 140364 4834 140420 4844
rect 141036 4900 141092 4910
rect 141036 480 141092 4844
rect 141932 4564 141988 5096
rect 141932 4498 141988 4508
rect 142940 4788 142996 4798
rect 142940 480 142996 4732
rect 143500 4452 143556 5096
rect 143500 4386 143556 4396
rect 144844 4676 144900 4686
rect 144844 480 144900 4620
rect 145068 2548 145124 5096
rect 146636 2660 146692 5096
rect 146636 2594 146692 2604
rect 146748 4564 146804 4574
rect 145068 2482 145124 2492
rect 146748 480 146804 4508
rect 148204 2772 148260 5096
rect 149548 5068 149800 5124
rect 149548 5012 149604 5068
rect 149548 4946 149604 4956
rect 151340 4900 151396 5096
rect 151340 4834 151396 4844
rect 152908 4788 152964 5096
rect 152908 4722 152964 4732
rect 154476 4676 154532 5096
rect 154476 4610 154532 4620
rect 156044 4564 156100 5096
rect 156044 4498 156100 4508
rect 148204 2706 148260 2716
rect 148652 4452 148708 4462
rect 148652 480 148708 4396
rect 157612 4452 157668 5096
rect 157612 4386 157668 4396
rect 158172 4676 158228 4686
rect 150556 3780 150612 3790
rect 150556 480 150612 3724
rect 152460 3668 152516 3678
rect 152460 480 152516 3612
rect 154364 3556 154420 3566
rect 154364 480 154420 3500
rect 156156 3444 156212 3454
rect 156156 480 156212 3388
rect 158172 480 158228 4620
rect 159180 3780 159236 5096
rect 159180 3714 159236 3724
rect 160076 5012 160132 5022
rect 160076 480 160132 4956
rect 160748 3668 160804 5096
rect 160748 3602 160804 3612
rect 161980 3892 162036 3902
rect 161980 480 162036 3836
rect 162316 3556 162372 5096
rect 162316 3490 162372 3500
rect 163884 3444 163940 5096
rect 165452 4676 165508 5096
rect 166348 5068 167048 5124
rect 166348 5012 166404 5068
rect 166348 4946 166404 4956
rect 165452 4610 165508 4620
rect 168588 3892 168644 5096
rect 168588 3826 168644 3836
rect 163884 3378 163940 3388
rect 164108 3780 164164 3790
rect 164108 532 164164 3724
rect 170156 3780 170212 5096
rect 170156 3714 170212 3724
rect 163884 480 164164 532
rect 165788 3668 165844 3678
rect 165788 480 165844 3612
rect 171724 3668 171780 5096
rect 171724 3602 171780 3612
rect 167692 3556 167748 3566
rect 167692 480 167748 3500
rect 173292 3556 173348 5096
rect 173292 3490 173348 3500
rect 169596 3444 169652 3454
rect 169596 480 169652 3388
rect 174860 3444 174916 5096
rect 174860 3378 174916 3388
rect 175308 2772 175364 2782
rect 173404 2660 173460 2670
rect 171500 2548 171556 2558
rect 171500 480 171556 2492
rect 173404 480 173460 2604
rect 175308 480 175364 2716
rect 176428 2548 176484 5096
rect 177996 2660 178052 5096
rect 179564 2772 179620 5096
rect 179564 2706 179620 2716
rect 177996 2594 178052 2604
rect 179116 2660 179172 2670
rect 176428 2482 176484 2492
rect 177212 2436 177268 2446
rect 177212 480 177268 2380
rect 179116 480 179172 2604
rect 181020 2548 181076 2558
rect 181020 480 181076 2492
rect 181132 2436 181188 5096
rect 182700 2660 182756 5096
rect 182700 2594 182756 2604
rect 182924 2660 182980 2670
rect 181132 2370 181188 2380
rect 182924 480 182980 2604
rect 184268 2548 184324 5096
rect 185836 2660 185892 5096
rect 185836 2594 185892 2604
rect 186732 3556 186788 3566
rect 184268 2482 184324 2492
rect 184716 2548 184772 2558
rect 184716 480 184772 2492
rect 186732 480 186788 3500
rect 187404 2548 187460 5096
rect 188972 3556 189028 5096
rect 188972 3490 189028 3500
rect 187404 2482 187460 2492
rect 188636 3444 188692 3454
rect 188636 480 188692 3388
rect 190540 3444 190596 5096
rect 190540 3378 190596 3388
rect 191436 5068 192136 5124
rect 193116 5068 193704 5124
rect 194796 5068 195272 5124
rect 196476 5068 196840 5124
rect 198156 5068 198408 5124
rect 190540 480 190708 532
rect 54124 242 54180 252
rect 55160 392 55412 480
rect 57064 392 57316 480
rect 58968 392 59220 480
rect 60872 392 61124 480
rect 62776 392 63028 480
rect 64680 392 64932 480
rect 66584 392 66836 480
rect 68488 392 68740 480
rect 55160 -960 55384 392
rect 57064 -960 57288 392
rect 58968 -960 59192 392
rect 60872 -960 61096 392
rect 62776 -960 63000 392
rect 64680 -960 64904 392
rect 66584 -960 66808 392
rect 68488 -960 68712 392
rect 70392 -960 70616 480
rect 72296 392 72548 480
rect 74200 392 74452 480
rect 76104 392 76356 480
rect 78008 392 78260 480
rect 79912 392 80164 480
rect 81816 392 82068 480
rect 83720 392 83972 480
rect 85624 392 85876 480
rect 87528 392 87780 480
rect 89432 392 89684 480
rect 91336 392 91588 480
rect 93240 392 93492 480
rect 95144 392 95396 480
rect 97048 392 97300 480
rect 72296 -960 72520 392
rect 74200 -960 74424 392
rect 76104 -960 76328 392
rect 78008 -960 78232 392
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 83720 -960 83944 392
rect 85624 -960 85848 392
rect 87528 -960 87752 392
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 -960 97272 392
rect 98952 -960 99176 480
rect 100856 392 101108 480
rect 102760 392 103012 480
rect 104664 392 104916 480
rect 106568 392 106820 480
rect 108472 392 108724 480
rect 110376 392 110628 480
rect 112280 392 112532 480
rect 114184 392 114436 480
rect 116088 392 116340 480
rect 117992 392 118244 480
rect 119896 392 120148 480
rect 121800 392 122052 480
rect 123704 392 123956 480
rect 125608 392 125860 480
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104664 -960 104888 392
rect 106568 -960 106792 392
rect 108472 -960 108696 392
rect 110376 -960 110600 392
rect 112280 -960 112504 392
rect 114184 -960 114408 392
rect 116088 -960 116312 392
rect 117992 -960 118216 392
rect 119896 -960 120120 392
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 -960 125832 392
rect 127512 -960 127736 480
rect 129416 392 129668 480
rect 131320 392 131572 480
rect 133224 392 133476 480
rect 135128 392 135380 480
rect 137032 392 137284 480
rect 138936 392 139188 480
rect 140840 392 141092 480
rect 142744 392 142996 480
rect 144648 392 144900 480
rect 146552 392 146804 480
rect 148456 392 148708 480
rect 150360 392 150612 480
rect 152264 392 152516 480
rect 154168 392 154420 480
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 -960 135352 392
rect 137032 -960 137256 392
rect 138936 -960 139160 392
rect 140840 -960 141064 392
rect 142744 -960 142968 392
rect 144648 -960 144872 392
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 -960 150584 392
rect 152264 -960 152488 392
rect 154168 -960 154392 392
rect 156072 -960 156296 480
rect 157976 392 158228 480
rect 159880 392 160132 480
rect 161784 392 162036 480
rect 163688 476 164164 480
rect 163688 392 163940 476
rect 165592 392 165844 480
rect 167496 392 167748 480
rect 169400 392 169652 480
rect 171304 392 171556 480
rect 173208 392 173460 480
rect 175112 392 175364 480
rect 177016 392 177268 480
rect 178920 392 179172 480
rect 180824 392 181076 480
rect 182728 392 182980 480
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 -960 162008 392
rect 163688 -960 163912 392
rect 165592 -960 165816 392
rect 167496 -960 167720 392
rect 169400 -960 169624 392
rect 171304 -960 171528 392
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 -960 177240 392
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 480
rect 186536 392 186788 480
rect 188440 392 188692 480
rect 190344 476 190708 480
rect 190344 392 190596 476
rect 190652 420 190708 476
rect 191436 420 191492 5068
rect 192444 480 192612 532
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 -960 190568 392
rect 190652 364 191492 420
rect 192248 476 192612 480
rect 192248 392 192500 476
rect 192556 420 192612 476
rect 193116 420 193172 5068
rect 194348 480 194516 532
rect 192248 -960 192472 392
rect 192556 364 193172 420
rect 194152 476 194516 480
rect 194152 392 194404 476
rect 194460 420 194516 476
rect 194796 420 194852 5068
rect 196476 2548 196532 5068
rect 196252 2492 196532 2548
rect 196252 480 196308 2492
rect 198156 480 198212 5068
rect 199948 480 200004 5096
rect 201544 5068 201796 5124
rect 203112 5068 203700 5124
rect 204680 5068 205044 5124
rect 206248 5068 206836 5124
rect 207816 5068 208404 5124
rect 201740 480 201796 5068
rect 203644 480 203700 5068
rect 194152 -960 194376 392
rect 194460 364 194852 420
rect 196056 392 196308 480
rect 197960 392 198212 480
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199864 -960 200088 480
rect 201740 392 201992 480
rect 203644 392 203896 480
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 204988 420 205044 5068
rect 205436 480 205604 532
rect 205436 476 205800 480
rect 205436 420 205492 476
rect 204988 364 205492 420
rect 205548 392 205800 476
rect 205576 -960 205800 392
rect 206780 420 206836 5068
rect 207340 480 207508 532
rect 207340 476 207704 480
rect 207340 420 207396 476
rect 206780 364 207396 420
rect 207452 392 207704 476
rect 207480 -960 207704 392
rect 208348 420 208404 5068
rect 209356 3444 209412 5096
rect 210924 3556 210980 5096
rect 210924 3490 210980 3500
rect 209356 3378 209412 3388
rect 211260 3444 211316 3454
rect 209244 480 209412 532
rect 211260 480 211316 3388
rect 212492 3444 212548 5096
rect 212492 3378 212548 3388
rect 213164 3556 213220 3566
rect 213164 480 213220 3500
rect 214060 3556 214116 5096
rect 214060 3490 214116 3500
rect 215068 3444 215124 3454
rect 215068 480 215124 3388
rect 215628 3444 215684 5096
rect 215628 3378 215684 3388
rect 216972 3556 217028 3566
rect 216972 480 217028 3500
rect 217196 3556 217252 5096
rect 218764 3668 218820 5096
rect 218764 3602 218820 3612
rect 217196 3490 217252 3500
rect 218876 3444 218932 3454
rect 218876 480 218932 3388
rect 220332 3444 220388 5096
rect 220332 3378 220388 3388
rect 220780 3556 220836 3566
rect 220780 480 220836 3500
rect 221900 3556 221956 5096
rect 221900 3490 221956 3500
rect 222684 3668 222740 3678
rect 222684 480 222740 3612
rect 223468 3668 223524 5096
rect 223468 3602 223524 3612
rect 224588 3444 224644 3454
rect 224588 480 224644 3388
rect 225036 2548 225092 5096
rect 225036 2482 225092 2492
rect 226492 3556 226548 3566
rect 226492 480 226548 3500
rect 226604 2660 226660 5096
rect 226604 2594 226660 2604
rect 228172 2436 228228 5096
rect 228172 2370 228228 2380
rect 228508 3668 228564 3678
rect 228508 480 228564 3612
rect 229740 2884 229796 5096
rect 229740 2818 229796 2828
rect 231308 2772 231364 5096
rect 231308 2706 231364 2716
rect 232204 2660 232260 2670
rect 230300 2548 230356 2558
rect 230300 480 230356 2492
rect 232204 480 232260 2604
rect 232876 2548 232932 5096
rect 234444 2660 234500 5096
rect 236012 3444 236068 5096
rect 237580 3556 237636 5096
rect 239148 4452 239204 5096
rect 240716 4564 240772 5096
rect 242284 4676 242340 5096
rect 242284 4610 242340 4620
rect 240716 4498 240772 4508
rect 239148 4386 239204 4396
rect 243852 3668 243908 5096
rect 245420 3780 245476 5096
rect 245420 3714 245476 3724
rect 243852 3602 243908 3612
rect 237580 3490 237636 3500
rect 245532 3556 245588 3566
rect 236012 3378 236068 3388
rect 243628 3444 243684 3454
rect 234444 2594 234500 2604
rect 236012 2884 236068 2894
rect 232876 2482 232932 2492
rect 234108 2436 234164 2446
rect 234108 480 234164 2380
rect 236012 480 236068 2828
rect 237916 2772 237972 2782
rect 237916 480 237972 2716
rect 241724 2660 241780 2670
rect 239820 2548 239876 2558
rect 239820 480 239876 2492
rect 241724 480 241780 2604
rect 243628 480 243684 3388
rect 245532 480 245588 3500
rect 246988 3444 247044 5096
rect 246988 3378 247044 3388
rect 247436 4452 247492 4462
rect 247436 480 247492 4396
rect 248556 2772 248612 5096
rect 248556 2706 248612 2716
rect 249340 4564 249396 4574
rect 249340 480 249396 4508
rect 250124 2548 250180 5096
rect 250124 2482 250180 2492
rect 251244 4676 251300 4686
rect 251244 480 251300 4620
rect 251692 2436 251748 5096
rect 251692 2370 251748 2380
rect 253148 3668 253204 3678
rect 253148 480 253204 3612
rect 253260 3332 253316 5096
rect 253260 3266 253316 3276
rect 254828 3220 254884 5096
rect 254828 3154 254884 3164
rect 255052 3780 255108 3790
rect 255052 480 255108 3724
rect 256396 3108 256452 5096
rect 256396 3042 256452 3052
rect 257068 3444 257124 3454
rect 257068 480 257124 3388
rect 257964 2660 258020 5096
rect 259532 2996 259588 5096
rect 259532 2930 259588 2940
rect 257964 2594 258020 2604
rect 258860 2772 258916 2782
rect 258860 480 258916 2716
rect 260764 2548 260820 2558
rect 260764 480 260820 2492
rect 261100 2548 261156 5096
rect 262668 2884 262724 5096
rect 262668 2818 262724 2828
rect 264236 2772 264292 5096
rect 264236 2706 264292 2716
rect 264572 3332 264628 3342
rect 261100 2482 261156 2492
rect 262668 2436 262724 2446
rect 262668 480 262724 2380
rect 264572 480 264628 3276
rect 265804 2324 265860 5096
rect 265804 2258 265860 2268
rect 266476 3220 266532 3230
rect 266476 480 266532 3164
rect 267372 2436 267428 5096
rect 268940 3332 268996 5096
rect 268940 3266 268996 3276
rect 267372 2370 267428 2380
rect 268380 3108 268436 3118
rect 268380 480 268436 3052
rect 270284 2660 270340 2670
rect 270284 480 270340 2604
rect 270508 2660 270564 5096
rect 272076 3220 272132 5096
rect 272076 3154 272132 3164
rect 273644 3108 273700 5096
rect 273644 3042 273700 3052
rect 270508 2594 270564 2604
rect 272188 2996 272244 3006
rect 272188 480 272244 2940
rect 274092 2548 274148 2558
rect 274092 480 274148 2492
rect 275212 2548 275268 5096
rect 276780 2996 276836 5096
rect 276780 2930 276836 2940
rect 275212 2482 275268 2492
rect 275996 2884 276052 2894
rect 275996 480 276052 2828
rect 278348 2884 278404 5096
rect 278348 2818 278404 2828
rect 277900 2772 277956 2782
rect 277900 480 277956 2716
rect 279916 2772 279972 5096
rect 281484 4004 281540 5096
rect 283052 4788 283108 5096
rect 284620 4900 284676 5096
rect 284620 4834 284676 4844
rect 283052 4722 283108 4732
rect 281484 3938 281540 3948
rect 279916 2706 279972 2716
rect 283612 3332 283668 3342
rect 281708 2436 281764 2446
rect 279804 2324 279860 2334
rect 279804 480 279860 2268
rect 281708 480 281764 2380
rect 283612 480 283668 3276
rect 285628 2660 285684 2670
rect 285628 480 285684 2604
rect 286188 2660 286244 5096
rect 287756 4116 287812 5096
rect 289324 4228 289380 5096
rect 290892 4340 290948 5096
rect 290892 4274 290948 4284
rect 289324 4162 289380 4172
rect 287756 4050 287812 4060
rect 286188 2594 286244 2604
rect 287420 3220 287476 3230
rect 287420 480 287476 3164
rect 289324 3108 289380 3118
rect 289324 480 289380 3052
rect 291228 2548 291284 2558
rect 291228 480 291284 2492
rect 292460 2548 292516 5096
rect 294056 5068 294756 5124
rect 294700 5012 294756 5068
rect 294700 4946 294756 4956
rect 295596 4452 295652 5096
rect 297164 4564 297220 5096
rect 298732 4676 298788 5096
rect 298732 4610 298788 4620
rect 297164 4498 297220 4508
rect 295596 4386 295652 4396
rect 298844 4004 298900 4014
rect 292460 2482 292516 2492
rect 293132 2996 293188 3006
rect 293132 480 293188 2940
rect 295036 2884 295092 2894
rect 295036 480 295092 2828
rect 296940 2772 296996 2782
rect 296940 480 296996 2716
rect 298844 480 298900 3948
rect 300300 3220 300356 5096
rect 300300 3154 300356 3164
rect 300748 4788 300804 4798
rect 300748 480 300804 4732
rect 301868 4788 301924 5096
rect 301868 4722 301924 4732
rect 302652 4900 302708 4910
rect 302652 480 302708 4844
rect 303436 3108 303492 5096
rect 305004 4900 305060 5096
rect 305004 4834 305060 4844
rect 303436 3042 303492 3052
rect 306460 4116 306516 4126
rect 304556 2660 304612 2670
rect 304556 480 304612 2604
rect 306460 480 306516 4060
rect 306572 2996 306628 5096
rect 306572 2930 306628 2940
rect 308140 2660 308196 5096
rect 308140 2594 308196 2604
rect 308364 4228 308420 4238
rect 308364 480 308420 4172
rect 309708 2884 309764 5096
rect 309708 2818 309764 2828
rect 310268 4340 310324 4350
rect 310268 480 310324 4284
rect 311276 2772 311332 5096
rect 311276 2706 311332 2716
rect 312172 2548 312228 2558
rect 312172 480 312228 2492
rect 312844 2548 312900 5096
rect 312844 2482 312900 2492
rect 314188 5012 314244 5022
rect 314188 480 314244 4956
rect 314412 4004 314468 5096
rect 316008 5068 316708 5124
rect 316652 5012 316708 5068
rect 316652 4946 316708 4956
rect 314412 3938 314468 3948
rect 315980 4452 316036 4462
rect 315980 480 316036 4396
rect 317548 4116 317604 5096
rect 317548 4050 317604 4060
rect 317884 4564 317940 4574
rect 317884 480 317940 4508
rect 319116 4228 319172 5096
rect 319116 4162 319172 4172
rect 319788 4676 319844 4686
rect 319788 480 319844 4620
rect 320684 4340 320740 5096
rect 322252 4452 322308 5096
rect 322252 4386 322308 4396
rect 323596 4788 323652 4798
rect 320684 4274 320740 4284
rect 321692 3220 321748 3230
rect 321692 480 321748 3164
rect 323596 480 323652 4732
rect 323820 3332 323876 5096
rect 323820 3266 323876 3276
rect 325388 3220 325444 5096
rect 326956 4564 327012 5096
rect 326956 4498 327012 4508
rect 327404 4900 327460 4910
rect 325388 3154 325444 3164
rect 325500 3108 325556 3118
rect 325500 480 325556 3052
rect 327404 480 327460 4844
rect 328524 4676 328580 5096
rect 328524 4610 328580 4620
rect 330092 3108 330148 5096
rect 330092 3042 330148 3052
rect 329308 2996 329364 3006
rect 329308 480 329364 2940
rect 331212 2660 331268 2670
rect 331212 480 331268 2604
rect 331660 2660 331716 5096
rect 333228 5058 333284 5068
rect 334796 2996 334852 5096
rect 336364 4788 336420 5096
rect 337932 4900 337988 5096
rect 337932 4834 337988 4844
rect 336364 4722 336420 4732
rect 334796 2930 334852 2940
rect 338828 4004 338884 4014
rect 331660 2594 331716 2604
rect 333116 2884 333172 2894
rect 333116 480 333172 2828
rect 335020 2772 335076 2782
rect 335020 480 335076 2716
rect 336924 2548 336980 2558
rect 336924 480 336980 2492
rect 338828 480 338884 3948
rect 339500 2884 339556 5096
rect 341096 5068 341796 5124
rect 339500 2818 339556 2828
rect 340732 5012 340788 5022
rect 340732 480 340788 4956
rect 341740 5012 341796 5068
rect 341740 4946 341796 4956
rect 342524 5068 342664 5124
rect 342524 532 342580 5068
rect 209244 476 209608 480
rect 209244 420 209300 476
rect 208348 364 209300 420
rect 209356 392 209608 476
rect 211260 392 211512 480
rect 213164 392 213416 480
rect 215068 392 215320 480
rect 216972 392 217224 480
rect 218876 392 219128 480
rect 220780 392 221032 480
rect 222684 392 222936 480
rect 224588 392 224840 480
rect 226492 392 226744 480
rect 209384 -960 209608 392
rect 211288 -960 211512 392
rect 213192 -960 213416 392
rect 215096 -960 215320 392
rect 217000 -960 217224 392
rect 218904 -960 219128 392
rect 220808 -960 221032 392
rect 222712 -960 222936 392
rect 224616 -960 224840 392
rect 226520 -960 226744 392
rect 228424 -960 228648 480
rect 230300 392 230552 480
rect 232204 392 232456 480
rect 234108 392 234360 480
rect 236012 392 236264 480
rect 237916 392 238168 480
rect 239820 392 240072 480
rect 241724 392 241976 480
rect 243628 392 243880 480
rect 245532 392 245784 480
rect 247436 392 247688 480
rect 249340 392 249592 480
rect 251244 392 251496 480
rect 253148 392 253400 480
rect 255052 392 255304 480
rect 230328 -960 230552 392
rect 232232 -960 232456 392
rect 234136 -960 234360 392
rect 236040 -960 236264 392
rect 237944 -960 238168 392
rect 239848 -960 240072 392
rect 241752 -960 241976 392
rect 243656 -960 243880 392
rect 245560 -960 245784 392
rect 247464 -960 247688 392
rect 249368 -960 249592 392
rect 251272 -960 251496 392
rect 253176 -960 253400 392
rect 255080 -960 255304 392
rect 256984 -960 257208 480
rect 258860 392 259112 480
rect 260764 392 261016 480
rect 262668 392 262920 480
rect 264572 392 264824 480
rect 266476 392 266728 480
rect 268380 392 268632 480
rect 270284 392 270536 480
rect 272188 392 272440 480
rect 274092 392 274344 480
rect 275996 392 276248 480
rect 277900 392 278152 480
rect 279804 392 280056 480
rect 281708 392 281960 480
rect 283612 392 283864 480
rect 258888 -960 259112 392
rect 260792 -960 261016 392
rect 262696 -960 262920 392
rect 264600 -960 264824 392
rect 266504 -960 266728 392
rect 268408 -960 268632 392
rect 270312 -960 270536 392
rect 272216 -960 272440 392
rect 274120 -960 274344 392
rect 276024 -960 276248 392
rect 277928 -960 278152 392
rect 279832 -960 280056 392
rect 281736 -960 281960 392
rect 283640 -960 283864 392
rect 285544 -960 285768 480
rect 287420 392 287672 480
rect 289324 392 289576 480
rect 291228 392 291480 480
rect 293132 392 293384 480
rect 295036 392 295288 480
rect 296940 392 297192 480
rect 298844 392 299096 480
rect 300748 392 301000 480
rect 302652 392 302904 480
rect 304556 392 304808 480
rect 306460 392 306712 480
rect 308364 392 308616 480
rect 310268 392 310520 480
rect 312172 392 312424 480
rect 287448 -960 287672 392
rect 289352 -960 289576 392
rect 291256 -960 291480 392
rect 293160 -960 293384 392
rect 295064 -960 295288 392
rect 296968 -960 297192 392
rect 298872 -960 299096 392
rect 300776 -960 301000 392
rect 302680 -960 302904 392
rect 304584 -960 304808 392
rect 306488 -960 306712 392
rect 308392 -960 308616 392
rect 310296 -960 310520 392
rect 312200 -960 312424 392
rect 314104 -960 314328 480
rect 315980 392 316232 480
rect 317884 392 318136 480
rect 319788 392 320040 480
rect 321692 392 321944 480
rect 323596 392 323848 480
rect 325500 392 325752 480
rect 327404 392 327656 480
rect 329308 392 329560 480
rect 331212 392 331464 480
rect 333116 392 333368 480
rect 335020 392 335272 480
rect 336924 392 337176 480
rect 338828 392 339080 480
rect 340732 392 340984 480
rect 342748 4116 342804 4126
rect 342748 480 342804 4060
rect 344204 2548 344260 5096
rect 344204 2482 344260 2492
rect 344540 4228 344596 4238
rect 344540 480 344596 4172
rect 345772 2324 345828 5096
rect 347368 5068 347732 5124
rect 345772 2258 345828 2268
rect 346444 4340 346500 4350
rect 346444 480 346500 4284
rect 347676 1764 347732 5068
rect 348348 4452 348404 4462
rect 347676 1708 347844 1764
rect 347788 756 347844 1708
rect 347788 690 347844 700
rect 348348 480 348404 4396
rect 348908 2772 348964 5096
rect 350504 5068 351092 5124
rect 351036 3892 351092 5068
rect 351036 3826 351092 3836
rect 348908 2706 348964 2716
rect 350252 3332 350308 3342
rect 350252 480 350308 3276
rect 352044 868 352100 5096
rect 354060 4564 354116 4574
rect 352044 802 352100 812
rect 352156 3220 352212 3230
rect 352156 480 352212 3164
rect 354060 480 354116 4508
rect 355180 3220 355236 5096
rect 355180 3154 355236 3164
rect 355964 4676 356020 4686
rect 355964 480 356020 4620
rect 356748 532 356804 5096
rect 342524 466 342580 476
rect 316008 -960 316232 392
rect 317912 -960 318136 392
rect 319816 -960 320040 392
rect 321720 -960 321944 392
rect 323624 -960 323848 392
rect 325528 -960 325752 392
rect 327432 -960 327656 392
rect 329336 -960 329560 392
rect 331240 -960 331464 392
rect 333144 -960 333368 392
rect 335048 -960 335272 392
rect 336952 -960 337176 392
rect 338856 -960 339080 392
rect 340760 -960 340984 392
rect 342664 -960 342888 480
rect 344540 392 344792 480
rect 346444 392 346696 480
rect 348348 392 348600 480
rect 350252 392 350504 480
rect 352156 392 352408 480
rect 354060 392 354312 480
rect 355964 392 356216 480
rect 356748 466 356804 476
rect 357868 3108 357924 3118
rect 357868 480 357924 3052
rect 358316 2436 358372 5096
rect 358316 2370 358372 2380
rect 359548 3556 359604 3566
rect 359548 2324 359604 3500
rect 359884 3332 359940 5096
rect 359884 3266 359940 3276
rect 359548 2258 359604 2268
rect 359772 2660 359828 2670
rect 359772 480 359828 2604
rect 361452 1876 361508 5096
rect 361452 1810 361508 1820
rect 361676 480 361732 5068
rect 363020 2660 363076 5096
rect 363020 2594 363076 2604
rect 363580 2996 363636 3006
rect 363580 480 363636 2940
rect 364588 2212 364644 5096
rect 366044 5068 366184 5124
rect 369320 5068 369572 5124
rect 364588 2146 364644 2156
rect 365484 4788 365540 4798
rect 364476 1876 364532 1886
rect 364476 644 364532 1820
rect 364476 578 364532 588
rect 365484 480 365540 4732
rect 366044 1764 366100 5068
rect 367724 5058 367780 5068
rect 367388 4900 367444 4910
rect 366156 3668 366212 3678
rect 366156 3332 366212 3612
rect 366156 3266 366212 3276
rect 366044 1708 366324 1764
rect 357868 392 358120 480
rect 359772 392 360024 480
rect 361676 392 361928 480
rect 363580 392 363832 480
rect 365484 392 365736 480
rect 344568 -960 344792 392
rect 346472 -960 346696 392
rect 348376 -960 348600 392
rect 350280 -960 350504 392
rect 352184 -960 352408 392
rect 354088 -960 354312 392
rect 355992 -960 356216 392
rect 357896 -960 358120 392
rect 359800 -960 360024 392
rect 361704 -960 361928 392
rect 363608 -960 363832 392
rect 365512 -960 365736 392
rect 366268 420 366324 1708
rect 367388 480 367444 4844
rect 369292 2884 369348 2894
rect 369292 480 369348 2828
rect 369516 2324 369572 5068
rect 369516 2258 369572 2268
rect 366380 420 366436 430
rect 366268 364 366380 420
rect 367388 392 367640 480
rect 369292 392 369544 480
rect 366380 354 366436 364
rect 367416 -960 367640 392
rect 369320 -960 369544 392
rect 370860 308 370916 5096
rect 371308 5012 371364 5022
rect 371308 480 371364 4956
rect 372428 3220 372484 5096
rect 373996 3332 374052 5096
rect 375592 5068 376292 5124
rect 373996 3266 374052 3276
rect 372428 3154 372484 3164
rect 375004 2548 375060 2558
rect 372988 480 373156 532
rect 375004 480 375060 2492
rect 370860 242 370916 252
rect 371224 -960 371448 480
rect 372988 476 373352 480
rect 372988 196 373044 476
rect 373100 392 373352 476
rect 375004 392 375256 480
rect 372988 130 373044 140
rect 373128 -960 373352 392
rect 375032 -960 375256 392
rect 376236 196 376292 5068
rect 376908 3556 376964 3566
rect 376908 480 376964 3500
rect 377132 2548 377188 5096
rect 377916 3556 377972 3566
rect 377916 3332 377972 3500
rect 377916 3266 377972 3276
rect 378700 2996 378756 5096
rect 378700 2930 378756 2940
rect 380044 5068 380296 5124
rect 377132 2482 377188 2492
rect 378812 756 378868 766
rect 378812 480 378868 700
rect 376908 392 377160 480
rect 378812 392 379064 480
rect 376236 130 376292 140
rect 376936 -960 377160 392
rect 378840 -960 379064 392
rect 380044 84 380100 5068
rect 382620 3892 382676 3902
rect 381388 3780 381444 3790
rect 381388 3220 381444 3724
rect 381388 3154 381444 3164
rect 380716 2772 380772 2782
rect 380716 480 380772 2716
rect 382620 480 382676 3836
rect 383404 3332 383460 5096
rect 383404 3266 383460 3276
rect 384972 1540 385028 5096
rect 386540 3108 386596 5096
rect 386540 3042 386596 3052
rect 384972 1474 385028 1484
rect 384524 868 384580 878
rect 384524 480 384580 812
rect 386652 480 386708 5180
rect 429548 5170 429604 5180
rect 403116 5124 403172 5134
rect 420364 5124 420420 5134
rect 434252 5124 434308 5134
rect 387996 3892 388052 3902
rect 387996 3332 388052 3836
rect 387996 3266 388052 3276
rect 388108 1988 388164 5096
rect 389564 4004 389620 4014
rect 388108 1922 388164 1932
rect 388332 3444 388388 3454
rect 380716 392 380968 480
rect 382620 392 382872 480
rect 384524 392 384776 480
rect 380044 18 380100 28
rect 380744 -960 380968 392
rect 382648 -960 382872 392
rect 384552 -960 384776 392
rect 386456 392 386708 480
rect 388332 480 388388 3388
rect 389564 2212 389620 3948
rect 389676 2772 389732 5096
rect 389676 2706 389732 2716
rect 389564 2146 389620 2156
rect 391244 2212 391300 5096
rect 392840 5068 393092 5124
rect 393036 5012 393092 5068
rect 393036 4946 393092 4956
rect 394044 3668 394100 3678
rect 391244 2146 391300 2156
rect 392140 2436 392196 2446
rect 390124 532 390180 542
rect 388332 392 388584 480
rect 390180 480 390292 532
rect 392140 480 392196 2380
rect 394044 480 394100 3612
rect 394380 1652 394436 5096
rect 397516 2100 397572 5096
rect 397516 2034 397572 2044
rect 397852 2660 397908 2670
rect 394380 1586 394436 1596
rect 395948 644 396004 654
rect 395948 480 396004 588
rect 397852 480 397908 2604
rect 399084 756 399140 5096
rect 401436 4116 401492 4126
rect 399084 690 399140 700
rect 399868 4004 399924 4014
rect 399868 480 399924 3948
rect 401436 2996 401492 4060
rect 401436 2930 401492 2940
rect 402220 2884 402276 5096
rect 403172 5068 403284 5124
rect 403116 5058 403172 5068
rect 402220 2818 402276 2828
rect 401660 644 401716 654
rect 401660 480 401716 588
rect 390180 476 390488 480
rect 390124 466 390180 476
rect 390236 392 390488 476
rect 392140 392 392392 480
rect 394044 392 394296 480
rect 395948 392 396200 480
rect 397852 392 398104 480
rect 386456 -960 386680 392
rect 388360 -960 388584 392
rect 390264 -960 390488 392
rect 392168 -960 392392 392
rect 394072 -960 394296 392
rect 395976 -960 396200 392
rect 397880 -960 398104 392
rect 399784 -960 400008 480
rect 401660 392 401912 480
rect 401688 -960 401912 392
rect 403228 420 403284 5068
rect 403788 868 403844 5096
rect 405356 2996 405412 5096
rect 406952 5068 407652 5124
rect 407596 3668 407652 5068
rect 407596 3602 407652 3612
rect 405356 2930 405412 2940
rect 403788 802 403844 812
rect 405468 2324 405524 2334
rect 403452 480 403620 532
rect 405468 480 405524 2268
rect 408492 644 408548 5096
rect 408492 578 408548 588
rect 409276 3780 409332 3790
rect 407260 480 407428 532
rect 409276 480 409332 3724
rect 410060 3220 410116 5096
rect 411656 5068 412356 5124
rect 411516 4228 411572 4238
rect 410060 3154 410116 3164
rect 411180 3556 411236 3566
rect 411180 480 411236 3500
rect 411516 2772 411572 4172
rect 412300 4004 412356 5068
rect 412300 3938 412356 3948
rect 411516 2706 411572 2716
rect 413196 1204 413252 5096
rect 414764 2772 414820 5096
rect 414764 2706 414820 2716
rect 413196 1138 413252 1148
rect 414988 2548 415044 2558
rect 412972 480 413140 532
rect 414988 480 415044 2492
rect 416332 2212 416388 5096
rect 416892 4116 416948 4126
rect 416332 2146 416388 2156
rect 416668 3780 416724 3790
rect 416668 1988 416724 3724
rect 416668 1922 416724 1932
rect 416892 480 416948 4060
rect 417900 532 417956 5096
rect 403452 476 403816 480
rect 403452 420 403508 476
rect 403228 364 403508 420
rect 403564 392 403816 476
rect 405468 392 405720 480
rect 403592 -960 403816 392
rect 405496 -960 405720 392
rect 407260 476 407624 480
rect 407260 308 407316 476
rect 407372 392 407624 476
rect 409276 392 409528 480
rect 411180 392 411432 480
rect 407260 242 407316 252
rect 407400 -960 407624 392
rect 409304 -960 409528 392
rect 411208 -960 411432 392
rect 412972 476 413336 480
rect 412972 196 413028 476
rect 413084 392 413336 476
rect 414988 392 415240 480
rect 416892 392 417144 480
rect 417900 466 417956 476
rect 418684 480 418852 532
rect 418684 476 419048 480
rect 412972 130 413028 140
rect 413112 -960 413336 392
rect 415016 -960 415240 392
rect 416920 -960 417144 392
rect 418684 84 418740 476
rect 418796 392 419048 476
rect 418684 18 418740 28
rect 418824 -960 419048 392
rect 420364 420 420420 5068
rect 421036 2324 421092 5096
rect 422632 5068 423332 5124
rect 421036 2258 421092 2268
rect 422604 3892 422660 3902
rect 420588 480 420756 532
rect 422604 480 422660 3836
rect 423276 1428 423332 5068
rect 424172 2660 424228 5096
rect 425740 4900 425796 5096
rect 425740 4834 425796 4844
rect 424172 2594 424228 2604
rect 426412 3108 426468 3118
rect 423276 1362 423332 1372
rect 424508 1540 424564 1550
rect 424508 480 424564 1484
rect 426412 480 426468 3052
rect 420588 476 420952 480
rect 420588 420 420644 476
rect 420364 364 420644 420
rect 420700 392 420952 476
rect 422604 392 422856 480
rect 424508 392 424760 480
rect 426412 392 426664 480
rect 420728 -960 420952 392
rect 422632 -960 422856 392
rect 424536 -960 424760 392
rect 426440 -960 426664 392
rect 427308 420 427364 5096
rect 430220 4228 430276 4238
rect 428428 3892 428484 3902
rect 428428 2100 428484 3836
rect 428428 2034 428484 2044
rect 428540 3780 428596 3790
rect 428540 480 428596 3724
rect 427308 354 427364 364
rect 428344 392 428596 480
rect 430220 480 430276 4172
rect 430444 1988 430500 5096
rect 432040 5068 433076 5124
rect 433608 5068 434252 5124
rect 435176 5068 435876 5124
rect 430444 1922 430500 1932
rect 432124 2436 432180 2446
rect 432124 480 432180 2380
rect 430220 392 430472 480
rect 432124 392 432376 480
rect 428344 -960 428568 392
rect 430248 -960 430472 392
rect 432152 -960 432376 392
rect 433020 308 433076 5068
rect 434252 5058 434308 5068
rect 434364 5012 434420 5022
rect 434364 4900 434420 4956
rect 434252 4844 434420 4900
rect 434252 480 434308 4844
rect 435820 3780 435876 5068
rect 435820 3714 435876 3724
rect 435036 3444 435092 3454
rect 435036 2884 435092 3388
rect 435036 2818 435092 2828
rect 436716 1876 436772 5096
rect 436716 1810 436772 1820
rect 433020 242 433076 252
rect 434056 392 434308 480
rect 435932 1652 435988 1662
rect 435932 480 435988 1596
rect 437836 480 437892 5516
rect 443548 5460 443604 5470
rect 442988 5124 443044 5134
rect 438284 2548 438340 5096
rect 438284 2482 438340 2492
rect 439740 3892 439796 3902
rect 439740 480 439796 3836
rect 439852 2884 439908 5096
rect 440188 3556 440244 3566
rect 440188 2996 440244 3500
rect 441420 3108 441476 5096
rect 442988 5058 443044 5068
rect 441420 3042 441476 3052
rect 440188 2930 440244 2940
rect 439852 2818 439908 2828
rect 441644 756 441700 766
rect 441644 480 441700 700
rect 443548 480 443604 5404
rect 462476 5460 462532 5470
rect 444556 4340 444612 5096
rect 444556 4274 444612 4284
rect 445452 3444 445508 3454
rect 445452 480 445508 3388
rect 446124 756 446180 5096
rect 447692 3332 447748 5096
rect 447692 3266 447748 3276
rect 449260 1876 449316 5096
rect 450268 3668 450324 3678
rect 449260 1810 449316 1820
rect 449372 3556 449428 3566
rect 446124 690 446180 700
rect 447356 868 447412 878
rect 447356 480 447412 812
rect 449372 480 449428 3500
rect 450268 2212 450324 3612
rect 450268 2146 450324 2156
rect 450828 868 450884 5096
rect 450828 802 450884 812
rect 451164 3556 451220 3566
rect 451164 480 451220 3500
rect 452396 3220 452452 5096
rect 453992 5068 454692 5124
rect 454636 5012 454692 5068
rect 454636 4946 454692 4956
rect 452396 3154 452452 3164
rect 454972 3444 455028 3454
rect 453068 644 453124 654
rect 453068 480 453124 588
rect 454972 480 455028 3388
rect 455532 1316 455588 5096
rect 456988 4004 457044 4014
rect 456876 3556 456932 3566
rect 456876 2324 456932 3500
rect 456876 2258 456932 2268
rect 455532 1250 455588 1260
rect 456988 480 457044 3948
rect 457100 2996 457156 5096
rect 457100 2930 457156 2940
rect 458668 2212 458724 5096
rect 458668 2146 458724 2156
rect 460236 1540 460292 5096
rect 460236 1474 460292 1484
rect 460684 2772 460740 2782
rect 458780 980 458836 990
rect 458780 480 458836 924
rect 460684 480 460740 2716
rect 461804 2100 461860 5096
rect 462476 3220 462532 5404
rect 465724 5348 465780 5358
rect 463372 4452 463428 5096
rect 463372 4386 463428 4396
rect 462476 3154 462532 3164
rect 462588 3668 462644 3678
rect 461804 2034 461860 2044
rect 462588 480 462644 3612
rect 464940 644 464996 5096
rect 464940 578 464996 588
rect 464380 532 464436 542
rect 435932 392 436184 480
rect 437836 392 438088 480
rect 439740 392 439992 480
rect 441644 392 441896 480
rect 443548 392 443800 480
rect 445452 392 445704 480
rect 447356 392 447608 480
rect 434056 -960 434280 392
rect 435960 -960 436184 392
rect 437864 -960 438088 392
rect 439768 -960 439992 392
rect 441672 -960 441896 392
rect 443576 -960 443800 392
rect 445480 -960 445704 392
rect 447384 -960 447608 392
rect 449288 -960 449512 480
rect 451164 392 451416 480
rect 453068 392 453320 480
rect 454972 392 455224 480
rect 451192 -960 451416 392
rect 453096 -960 453320 392
rect 455000 -960 455224 392
rect 456904 -960 457128 480
rect 458780 392 459032 480
rect 460684 392 460936 480
rect 462588 392 462840 480
rect 464436 480 464548 532
rect 464436 476 464744 480
rect 464380 466 464436 476
rect 464492 392 464744 476
rect 458808 -960 459032 392
rect 460712 -960 460936 392
rect 462616 -960 462840 392
rect 464520 -960 464744 392
rect 465724 420 465780 5292
rect 474348 5348 474404 5358
rect 474348 5282 474404 5292
rect 478156 5236 478212 5246
rect 478044 5180 478156 5236
rect 466508 3220 466564 5096
rect 468076 4564 468132 5096
rect 468076 4498 468132 4508
rect 466508 3154 466564 3164
rect 468300 3556 468356 3566
rect 466284 480 466452 532
rect 468300 480 468356 3500
rect 469644 532 469700 5096
rect 471212 3332 471268 5096
rect 471212 3266 471268 3276
rect 471996 3444 472052 3454
rect 471996 1988 472052 3388
rect 471996 1922 472052 1932
rect 472108 2660 472164 2670
rect 466284 476 466648 480
rect 466284 420 466340 476
rect 465724 364 466340 420
rect 466396 392 466648 476
rect 468300 392 468552 480
rect 469644 466 469700 476
rect 470204 1428 470260 1438
rect 470204 480 470260 1372
rect 472108 480 472164 2604
rect 472780 2436 472836 5096
rect 472780 2370 472836 2380
rect 474012 4900 474068 4910
rect 474012 480 474068 4844
rect 475916 2660 475972 5096
rect 477484 4676 477540 5096
rect 477484 4610 477540 4620
rect 475916 2594 475972 2604
rect 475804 480 475972 532
rect 478044 480 478100 5180
rect 478156 5170 478212 5180
rect 482860 5124 482916 5134
rect 470204 392 470456 480
rect 472108 392 472360 480
rect 474012 392 474264 480
rect 466424 -960 466648 392
rect 468328 -960 468552 392
rect 470232 -960 470456 392
rect 472136 -960 472360 392
rect 474040 -960 474264 392
rect 475804 476 476168 480
rect 475804 420 475860 476
rect 475916 392 476168 476
rect 475804 354 475860 364
rect 475944 -960 476168 392
rect 477848 392 478100 480
rect 477848 -960 478072 392
rect 479052 84 479108 5096
rect 480396 3668 480452 3678
rect 479724 3444 479780 3454
rect 479724 480 479780 3388
rect 480396 2884 480452 3612
rect 480396 2818 480452 2828
rect 480620 2324 480676 5096
rect 480620 2258 480676 2268
rect 482188 1988 482244 5096
rect 482188 1922 482244 1932
rect 481516 480 481684 532
rect 479724 392 479976 480
rect 479052 18 479108 28
rect 479752 -960 479976 392
rect 481516 476 481880 480
rect 481516 308 481572 476
rect 481628 392 481880 476
rect 481516 242 481572 252
rect 481656 -960 481880 392
rect 482860 420 482916 5068
rect 483084 3220 483140 5516
rect 523516 5572 523572 5582
rect 506380 5460 506436 5470
rect 493164 5236 493220 5246
rect 493164 5170 493220 5180
rect 495404 5124 495460 5134
rect 483084 3154 483140 3164
rect 483756 1204 483812 5096
rect 485324 3108 485380 5096
rect 486892 4788 486948 5096
rect 486892 4722 486948 4732
rect 485324 3042 485380 3052
rect 485548 3780 485604 3790
rect 483756 1138 483812 1148
rect 483420 480 483588 532
rect 485548 480 485604 3724
rect 487228 480 487396 532
rect 483420 476 483784 480
rect 483420 420 483476 476
rect 482860 364 483476 420
rect 483532 392 483784 476
rect 483560 -960 483784 392
rect 485464 -960 485688 480
rect 487228 476 487592 480
rect 487228 196 487284 476
rect 487340 392 487592 476
rect 487228 130 487284 140
rect 487368 -960 487592 392
rect 488460 196 488516 5096
rect 490028 2996 490084 5096
rect 490028 2930 490084 2940
rect 491148 3668 491204 3678
rect 489244 2548 489300 2558
rect 489244 480 489300 2492
rect 491148 480 491204 3612
rect 491596 2884 491652 5096
rect 494760 5068 495404 5124
rect 495404 5058 495460 5068
rect 496300 4900 496356 5096
rect 496300 4834 496356 4844
rect 496860 4340 496916 4350
rect 491596 2818 491652 2828
rect 492156 3556 492212 3566
rect 492156 1876 492212 3500
rect 492156 1810 492212 1820
rect 493052 3444 493108 3454
rect 493052 480 493108 3388
rect 494956 3444 495012 3454
rect 494956 480 495012 3388
rect 496860 480 496916 4284
rect 497868 1652 497924 5096
rect 499436 3332 499492 5096
rect 499436 3266 499492 3276
rect 500668 3444 500724 3454
rect 497868 1586 497924 1596
rect 498764 756 498820 766
rect 498764 480 498820 700
rect 500668 480 500724 3388
rect 501004 3332 501060 5096
rect 502600 5068 503412 5124
rect 501004 3266 501060 3276
rect 502572 3556 502628 3566
rect 502572 480 502628 3500
rect 489244 392 489496 480
rect 491148 392 491400 480
rect 493052 392 493304 480
rect 494956 392 495208 480
rect 496860 392 497112 480
rect 498764 392 499016 480
rect 500668 392 500920 480
rect 502572 392 502824 480
rect 488460 130 488516 140
rect 489272 -960 489496 392
rect 491176 -960 491400 392
rect 493080 -960 493304 392
rect 494984 -960 495208 392
rect 496888 -960 497112 392
rect 498792 -960 499016 392
rect 500696 -960 500920 392
rect 502600 -960 502824 392
rect 503356 84 503412 5068
rect 503804 3780 503860 3790
rect 503804 2212 503860 3724
rect 503804 2146 503860 2156
rect 503916 3444 503972 3454
rect 503916 1316 503972 3388
rect 504140 2548 504196 5096
rect 504140 2482 504196 2492
rect 505708 2548 505764 5096
rect 505708 2482 505764 2492
rect 503916 1250 503972 1260
rect 504476 868 504532 878
rect 504476 480 504532 812
rect 506380 480 506436 5404
rect 507276 5124 507332 5134
rect 507276 5058 507332 5068
rect 508284 5012 508340 5022
rect 507276 2660 507332 2670
rect 507276 980 507332 2604
rect 507276 914 507332 924
rect 508284 480 508340 4956
rect 508844 2772 508900 5096
rect 508844 2706 508900 2716
rect 510188 3444 510244 3454
rect 509068 2324 509124 2334
rect 509068 868 509124 2268
rect 509068 802 509124 812
rect 510188 480 510244 3388
rect 510412 2660 510468 5096
rect 512008 5068 512484 5124
rect 512428 3668 512484 5068
rect 512428 3602 512484 3612
rect 510412 2594 510468 2604
rect 510524 3444 510580 3454
rect 510524 1540 510580 3388
rect 513548 2548 513604 5096
rect 515144 5068 515732 5124
rect 515676 5012 515732 5068
rect 515676 4946 515732 4956
rect 519708 4452 519764 4462
rect 513548 2482 513604 2492
rect 514108 3780 514164 3790
rect 510524 1474 510580 1484
rect 512092 756 512148 766
rect 512092 480 512148 700
rect 514108 480 514164 3724
rect 515900 3444 515956 3454
rect 515900 480 515956 3388
rect 517804 2100 517860 2110
rect 517804 480 517860 2044
rect 519708 480 519764 4396
rect 521612 644 521668 654
rect 521612 480 521668 588
rect 523516 480 523572 5516
rect 533036 5348 533092 5358
rect 525420 4564 525476 4574
rect 524188 3556 524244 3566
rect 524188 2436 524244 3500
rect 524188 2370 524244 2380
rect 525420 480 525476 4508
rect 531132 3556 531188 3566
rect 529228 3444 529284 3454
rect 527212 532 527268 542
rect 504476 392 504728 480
rect 506380 392 506632 480
rect 508284 392 508536 480
rect 510188 392 510440 480
rect 512092 392 512344 480
rect 503468 84 503524 94
rect 503356 28 503468 84
rect 503468 18 503524 28
rect 504504 -960 504728 392
rect 506408 -960 506632 392
rect 508312 -960 508536 392
rect 510216 -960 510440 392
rect 512120 -960 512344 392
rect 514024 -960 514248 480
rect 515900 392 516152 480
rect 517804 392 518056 480
rect 519708 392 519960 480
rect 521612 392 521864 480
rect 523516 392 523768 480
rect 525420 392 525672 480
rect 527268 480 527380 532
rect 529228 480 529284 3388
rect 531132 480 531188 3500
rect 533036 480 533092 5292
rect 555884 5236 555940 5246
rect 548268 4788 548324 4798
rect 536844 4676 536900 4686
rect 534940 868 534996 878
rect 534940 480 534996 812
rect 536844 480 536900 4620
rect 546364 3108 546420 3118
rect 542556 1764 542612 1774
rect 542612 1708 542724 1764
rect 542556 1698 542612 1708
rect 540652 756 540708 766
rect 538748 644 538804 654
rect 538748 480 538804 588
rect 540652 480 540708 700
rect 542668 480 542724 1708
rect 544348 480 544516 532
rect 546364 480 546420 3052
rect 548268 480 548324 4732
rect 552076 2996 552132 3006
rect 550060 480 550228 532
rect 552076 480 552132 2940
rect 553980 2884 554036 2894
rect 553980 480 554036 2828
rect 555884 480 555940 5180
rect 573020 5124 573076 5134
rect 559692 4900 559748 4910
rect 557788 3444 557844 3454
rect 557788 480 557844 3388
rect 559692 480 559748 4844
rect 565404 3444 565460 3454
rect 563500 1764 563556 1774
rect 561596 1652 561652 1662
rect 561596 480 561652 1596
rect 563500 480 563556 1708
rect 565404 480 565460 3388
rect 569212 644 569268 654
rect 567196 480 567364 532
rect 569212 480 569268 588
rect 571228 644 571284 654
rect 571228 480 571284 588
rect 573020 480 573076 5068
rect 584444 5012 584500 5022
rect 580636 3668 580692 3678
rect 574924 2772 574980 2782
rect 574924 480 574980 2716
rect 576828 2660 576884 2670
rect 576828 480 576884 2604
rect 580636 480 580692 3612
rect 582540 2548 582596 2558
rect 582540 480 582596 2492
rect 584444 480 584500 4956
rect 527268 476 527576 480
rect 527212 466 527268 476
rect 527324 392 527576 476
rect 529228 392 529480 480
rect 531132 392 531384 480
rect 533036 392 533288 480
rect 534940 392 535192 480
rect 536844 392 537096 480
rect 538748 392 539000 480
rect 540652 392 540904 480
rect 515928 -960 516152 392
rect 517832 -960 518056 392
rect 519736 -960 519960 392
rect 521640 -960 521864 392
rect 523544 -960 523768 392
rect 525448 -960 525672 392
rect 527352 -960 527576 392
rect 529256 -960 529480 392
rect 531160 -960 531384 392
rect 533064 -960 533288 392
rect 534968 -960 535192 392
rect 536872 -960 537096 392
rect 538776 -960 539000 392
rect 540680 -960 540904 392
rect 542584 -960 542808 480
rect 544348 476 544712 480
rect 544348 308 544404 476
rect 544460 392 544712 476
rect 546364 392 546616 480
rect 548268 392 548520 480
rect 544348 242 544404 252
rect 544488 -960 544712 392
rect 546392 -960 546616 392
rect 548296 -960 548520 392
rect 550060 476 550424 480
rect 550060 196 550116 476
rect 550172 392 550424 476
rect 552076 392 552328 480
rect 553980 392 554232 480
rect 555884 392 556136 480
rect 557788 392 558040 480
rect 559692 392 559944 480
rect 561596 392 561848 480
rect 563500 392 563752 480
rect 565404 392 565656 480
rect 550060 130 550116 140
rect 550200 -960 550424 392
rect 552104 -960 552328 392
rect 554008 -960 554232 392
rect 555912 -960 556136 392
rect 557816 -960 558040 392
rect 559720 -960 559944 392
rect 561624 -960 561848 392
rect 563528 -960 563752 392
rect 565432 -960 565656 392
rect 567196 476 567560 480
rect 567196 84 567252 476
rect 567308 392 567560 476
rect 569212 392 569464 480
rect 567196 18 567252 28
rect 567336 -960 567560 392
rect 569240 -960 569464 392
rect 571144 -960 571368 480
rect 573020 392 573272 480
rect 574924 392 575176 480
rect 576828 392 577080 480
rect 573048 -960 573272 392
rect 574952 -960 575176 392
rect 576856 -960 577080 392
rect 578760 -960 578984 480
rect 580636 392 580888 480
rect 582540 392 582792 480
rect 584444 392 584696 480
rect 580664 -960 580888 392
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 11228 590716 11284 590772
rect 99484 590940 99540 590996
rect 77420 590828 77476 590884
rect 118412 590828 118468 590884
rect 115052 588812 115108 588868
rect 55132 511532 55188 511588
rect 59612 548940 59668 548996
rect 33068 390572 33124 390628
rect 54572 509292 54628 509348
rect 1596 373660 1652 373716
rect 1484 308924 1540 308980
rect 28 304780 84 304836
rect 28 270284 84 270340
rect 1484 164332 1540 164388
rect 25228 373212 25284 373268
rect 2492 368844 2548 368900
rect 2380 330988 2436 331044
rect 2268 317660 2324 317716
rect 2380 162428 2436 162484
rect 2268 162092 2324 162148
rect 1596 148764 1652 148820
rect 23212 368060 23268 368116
rect 2940 364588 2996 364644
rect 2828 337148 2884 337204
rect 2716 337036 2772 337092
rect 2604 336924 2660 336980
rect 2604 312956 2660 313012
rect 2716 310268 2772 310324
rect 2716 305564 2772 305620
rect 5628 363692 5684 363748
rect 4508 363580 4564 363636
rect 2940 320348 2996 320404
rect 3052 359548 3108 359604
rect 3276 338492 3332 338548
rect 3052 314972 3108 315028
rect 3164 336812 3220 336868
rect 3276 315644 3332 315700
rect 4284 319004 4340 319060
rect 3164 312284 3220 312340
rect 3276 307580 3332 307636
rect 2828 304892 2884 304948
rect 2940 306236 2996 306292
rect 2716 281372 2772 281428
rect 3276 194012 3332 194068
rect 4172 272972 4228 273028
rect 2940 164220 2996 164276
rect 2492 148652 2548 148708
rect 4284 268716 4340 268772
rect 4620 340172 4676 340228
rect 4620 313628 4676 313684
rect 4732 338604 4788 338660
rect 4732 311612 4788 311668
rect 4844 332668 4900 332724
rect 4732 309596 4788 309652
rect 4620 306908 4676 306964
rect 4620 280140 4676 280196
rect 4732 279580 4788 279636
rect 5516 330316 5572 330372
rect 5516 320124 5572 320180
rect 18508 332668 18564 332724
rect 19852 330988 19908 331044
rect 27916 371308 27972 371364
rect 37996 336028 38052 336084
rect 35980 335020 36036 335076
rect 28588 334796 28644 334852
rect 35308 334460 35364 334516
rect 31948 333228 32004 333284
rect 31276 331548 31332 331604
rect 31052 329980 31108 330036
rect 36652 332892 36708 332948
rect 37324 330652 37380 330708
rect 42700 333452 42756 333508
rect 38668 333340 38724 333396
rect 41356 333004 41412 333060
rect 40012 332780 40068 332836
rect 44716 333116 44772 333172
rect 43372 331660 43428 331716
rect 5628 303996 5684 304052
rect 54460 309148 54516 309204
rect 5516 283836 5572 283892
rect 5068 280476 5124 280532
rect 53452 281820 53508 281876
rect 13132 280588 13188 280644
rect 23884 280588 23940 280644
rect 40684 280588 40740 280644
rect 25900 280476 25956 280532
rect 26572 280476 26628 280532
rect 5516 277788 5572 277844
rect 7084 277116 7140 277172
rect 7756 277116 7812 277172
rect 6412 277004 6468 277060
rect 5740 276780 5796 276836
rect 7980 276668 8036 276724
rect 7532 269612 7588 269668
rect 6748 264572 6804 264628
rect 6748 262780 6804 262836
rect 4844 164108 4900 164164
rect 4508 162652 4564 162708
rect 4172 65212 4228 65268
rect 4284 158844 4340 158900
rect 7756 267932 7812 267988
rect 7644 266252 7700 266308
rect 9100 276332 9156 276388
rect 11116 276892 11172 276948
rect 10444 276444 10500 276500
rect 9772 276220 9828 276276
rect 12460 278348 12516 278404
rect 13804 276556 13860 276612
rect 11788 274652 11844 274708
rect 8428 274540 8484 274596
rect 15148 275436 15204 275492
rect 14476 270172 14532 270228
rect 16828 278124 16884 278180
rect 16828 277004 16884 277060
rect 16492 271852 16548 271908
rect 17164 271292 17220 271348
rect 15820 269724 15876 269780
rect 7980 267036 8036 267092
rect 19180 273084 19236 273140
rect 18508 267820 18564 267876
rect 17836 266364 17892 266420
rect 20524 277900 20580 277956
rect 21868 274764 21924 274820
rect 21196 272748 21252 272804
rect 23212 280028 23268 280084
rect 24556 276668 24612 276724
rect 22540 272636 22596 272692
rect 23436 276332 23492 276388
rect 37996 280252 38052 280308
rect 27244 279804 27300 279860
rect 26908 278012 26964 278068
rect 26908 276780 26964 276836
rect 26572 276556 26628 276612
rect 26572 275548 26628 275604
rect 25228 273756 25284 273812
rect 29260 276780 29316 276836
rect 31276 278572 31332 278628
rect 29932 276556 29988 276612
rect 34636 278796 34692 278852
rect 35308 277116 35364 277172
rect 31948 273308 32004 273364
rect 27916 271964 27972 272020
rect 36876 278460 36932 278516
rect 38668 276108 38724 276164
rect 36876 275548 36932 275604
rect 44716 280588 44772 280644
rect 53452 280588 53508 280644
rect 45388 280476 45444 280532
rect 44044 280364 44100 280420
rect 41132 275548 41188 275604
rect 35980 271740 36036 271796
rect 23436 269836 23492 269892
rect 42700 278236 42756 278292
rect 42028 268380 42084 268436
rect 48748 277116 48804 277172
rect 48076 277004 48132 277060
rect 47404 276332 47460 276388
rect 46732 274876 46788 274932
rect 54572 280812 54628 280868
rect 54684 416780 54740 416836
rect 57036 361228 57092 361284
rect 55132 333340 55188 333396
rect 54684 280364 54740 280420
rect 56700 333116 56756 333172
rect 56252 333004 56308 333060
rect 55132 281484 55188 281540
rect 56140 288092 56196 288148
rect 54908 280252 54964 280308
rect 54460 278684 54516 278740
rect 50092 277116 50148 277172
rect 56140 277116 56196 277172
rect 56476 332780 56532 332836
rect 56252 270060 56308 270116
rect 56364 319676 56420 319732
rect 56476 273532 56532 273588
rect 56588 312284 56644 312340
rect 56364 268492 56420 268548
rect 49420 268268 49476 268324
rect 56924 332780 56980 332836
rect 56812 302204 56868 302260
rect 57932 339388 57988 339444
rect 57036 325052 57092 325108
rect 57148 327516 57204 327572
rect 57932 326396 57988 326452
rect 58716 331212 58772 331268
rect 57148 320908 57204 320964
rect 58156 324380 58212 324436
rect 58044 310268 58100 310324
rect 57932 307580 57988 307636
rect 57820 305564 57876 305620
rect 56924 280700 56980 280756
rect 57036 302876 57092 302932
rect 56924 276332 56980 276388
rect 57820 280588 57876 280644
rect 57036 277004 57092 277060
rect 57036 276108 57092 276164
rect 56924 275996 56980 276052
rect 56700 275212 56756 275268
rect 56588 268156 56644 268212
rect 46060 266812 46116 266868
rect 58156 281484 58212 281540
rect 58268 322364 58324 322420
rect 58716 314300 58772 314356
rect 59500 319004 59556 319060
rect 58492 310940 58548 310996
rect 58268 280476 58324 280532
rect 58380 308252 58436 308308
rect 59388 301980 59444 302036
rect 58492 278572 58548 278628
rect 58604 289436 58660 289492
rect 58380 275324 58436 275380
rect 58044 273420 58100 273476
rect 58716 284732 58772 284788
rect 58716 277676 58772 277732
rect 58604 269500 58660 269556
rect 60620 522508 60676 522564
rect 59836 378812 59892 378868
rect 59612 281820 59668 281876
rect 59724 333564 59780 333620
rect 59836 288764 59892 288820
rect 60060 332892 60116 332948
rect 113372 502460 113428 502516
rect 111692 460124 111748 460180
rect 88956 383852 89012 383908
rect 86492 364812 86548 364868
rect 78204 359212 78260 359268
rect 76188 349132 76244 349188
rect 70364 333788 70420 333844
rect 73500 333676 73556 333732
rect 72828 333452 72884 333508
rect 70364 333004 70420 333060
rect 69468 332668 69524 332724
rect 70476 333116 70532 333172
rect 70476 332668 70532 332724
rect 72156 332892 72212 332948
rect 75516 333564 75572 333620
rect 73500 330204 73556 330260
rect 74844 333340 74900 333396
rect 74844 332668 74900 332724
rect 75516 329868 75572 329924
rect 77532 332668 77588 332724
rect 76860 329868 76916 329924
rect 84924 333788 84980 333844
rect 82908 333116 82964 333172
rect 78876 332892 78932 332948
rect 79548 331212 79604 331268
rect 83580 331884 83636 331940
rect 84252 331324 84308 331380
rect 88284 333564 88340 333620
rect 86940 332780 86996 332836
rect 87612 333452 87668 333508
rect 110012 375452 110068 375508
rect 93660 372092 93716 372148
rect 92988 331436 93044 331492
rect 110236 375452 110292 375508
rect 102396 334908 102452 334964
rect 101052 334348 101108 334404
rect 95004 331996 95060 332052
rect 100380 331212 100436 331268
rect 101724 332780 101780 332836
rect 103740 331100 103796 331156
rect 103068 330204 103124 330260
rect 105084 330988 105140 331044
rect 104412 330428 104468 330484
rect 105756 330092 105812 330148
rect 60620 327516 60676 327572
rect 109900 336028 109956 336084
rect 60284 320124 60340 320180
rect 60060 281708 60116 281764
rect 60172 312956 60228 313012
rect 59724 278460 59780 278516
rect 60060 278124 60116 278180
rect 60060 276892 60116 276948
rect 59500 275100 59556 275156
rect 59388 266588 59444 266644
rect 57932 265244 57988 265300
rect 43372 265132 43428 265188
rect 60396 314972 60452 315028
rect 60396 280364 60452 280420
rect 60508 311612 60564 311668
rect 60284 274988 60340 275044
rect 109340 303100 109396 303156
rect 70140 280700 70196 280756
rect 74844 280700 74900 280756
rect 87612 280700 87668 280756
rect 89628 280700 89684 280756
rect 60732 276220 60788 276276
rect 61404 277116 61460 277172
rect 62076 278236 62132 278292
rect 62076 276668 62132 276724
rect 62748 277900 62804 277956
rect 63420 277004 63476 277060
rect 62748 276444 62804 276500
rect 64092 276668 64148 276724
rect 61404 275548 61460 275604
rect 63868 276332 63924 276388
rect 65436 277116 65492 277172
rect 64764 276332 64820 276388
rect 64092 275548 64148 275604
rect 65548 275548 65604 275604
rect 65548 274652 65604 274708
rect 63868 273756 63924 273812
rect 60732 273196 60788 273252
rect 67452 276892 67508 276948
rect 68124 276444 68180 276500
rect 66780 275548 66836 275604
rect 66108 273084 66164 273140
rect 70812 279804 70868 279860
rect 69468 276556 69524 276612
rect 71932 277116 71988 277172
rect 68684 274652 68740 274708
rect 68796 276444 68852 276500
rect 68796 274540 68852 274596
rect 72828 278796 72884 278852
rect 72828 278012 72884 278068
rect 74172 280028 74228 280084
rect 72156 274540 72212 274596
rect 75516 280028 75572 280084
rect 74172 278460 74228 278516
rect 76188 279692 76244 279748
rect 73052 276332 73108 276388
rect 71932 271180 71988 271236
rect 68684 269836 68740 269892
rect 60508 266700 60564 266756
rect 60172 265020 60228 265076
rect 19852 264796 19908 264852
rect 75628 277116 75684 277172
rect 77532 280028 77588 280084
rect 76860 277116 76916 277172
rect 78204 278348 78260 278404
rect 76188 276780 76244 276836
rect 78204 276332 78260 276388
rect 75628 271292 75684 271348
rect 79548 276668 79604 276724
rect 80892 276780 80948 276836
rect 80892 276444 80948 276500
rect 81676 279916 81732 279972
rect 82236 278348 82292 278404
rect 81452 277004 81508 277060
rect 80220 275996 80276 276052
rect 78876 271292 78932 271348
rect 82236 276780 82292 276836
rect 83580 277116 83636 277172
rect 84252 277004 84308 277060
rect 84924 276892 84980 276948
rect 82908 276668 82964 276724
rect 85596 273644 85652 273700
rect 90300 277116 90356 277172
rect 88956 276556 89012 276612
rect 88284 276444 88340 276500
rect 90972 276108 91028 276164
rect 93660 276892 93716 276948
rect 94332 276892 94388 276948
rect 92988 276108 93044 276164
rect 101052 277116 101108 277172
rect 97692 276780 97748 276836
rect 95676 275996 95732 276052
rect 86940 274764 86996 274820
rect 100828 275548 100884 275604
rect 109564 297276 109620 297332
rect 109564 282044 109620 282100
rect 109228 278796 109284 278852
rect 109564 278348 109620 278404
rect 101724 275548 101780 275604
rect 106876 278012 106932 278068
rect 100828 273196 100884 273252
rect 86268 273084 86324 273140
rect 104972 273084 105028 273140
rect 82236 268044 82292 268100
rect 99932 269724 99988 269780
rect 81452 266364 81508 266420
rect 73052 264684 73108 264740
rect 7756 220444 7812 220500
rect 7644 177996 7700 178052
rect 10892 194012 10948 194068
rect 20636 165676 20692 165732
rect 26684 165676 26740 165732
rect 28028 165676 28084 165732
rect 39676 165676 39732 165732
rect 71708 165676 71764 165732
rect 82236 165676 82292 165732
rect 84028 165676 84084 165732
rect 83804 165564 83860 165620
rect 20860 162876 20916 162932
rect 10892 162764 10948 162820
rect 27132 162876 27188 162932
rect 26236 162652 26292 162708
rect 21308 162540 21364 162596
rect 17948 159628 18004 159684
rect 37884 164444 37940 164500
rect 38332 163996 38388 164052
rect 44156 164108 44212 164164
rect 44156 162988 44212 163044
rect 44380 162428 44436 162484
rect 44940 162988 44996 163044
rect 28476 161084 28532 161140
rect 44828 162092 44884 162148
rect 27804 159404 27860 159460
rect 43484 158956 43540 159012
rect 38108 158732 38164 158788
rect 26460 157948 26516 158004
rect 18396 155372 18452 155428
rect 18732 148876 18788 148932
rect 25900 148764 25956 148820
rect 27356 157052 27412 157108
rect 26796 150444 26852 150500
rect 27804 155484 27860 155540
rect 37548 148876 37604 148932
rect 28140 148652 28196 148708
rect 38444 152796 38500 152852
rect 43932 157388 43988 157444
rect 44380 155484 44436 155540
rect 44940 157276 44996 157332
rect 45500 164220 45556 164276
rect 45500 163548 45556 163604
rect 46172 164332 46228 164388
rect 45276 162764 45332 162820
rect 45388 155596 45444 155652
rect 45052 152012 45108 152068
rect 46172 148764 46228 148820
rect 46396 163548 46452 163604
rect 47852 162428 47908 162484
rect 46396 148652 46452 148708
rect 46620 157500 46676 157556
rect 45164 147868 45220 147924
rect 53676 160972 53732 161028
rect 63980 162988 64036 163044
rect 63980 157500 64036 157556
rect 64988 162204 65044 162260
rect 65212 162092 65268 162148
rect 66108 162204 66164 162260
rect 65660 161420 65716 161476
rect 65548 160412 65604 160468
rect 65548 158956 65604 159012
rect 64988 157388 65044 157444
rect 47852 152124 47908 152180
rect 56924 157164 56980 157220
rect 46620 147868 46676 147924
rect 64876 155596 64932 155652
rect 72380 163884 72436 163940
rect 71932 162428 71988 162484
rect 82684 162652 82740 162708
rect 91196 162876 91252 162932
rect 92092 164556 92148 164612
rect 99932 162876 99988 162932
rect 91644 162764 91700 162820
rect 83132 162540 83188 162596
rect 105196 269836 105252 269892
rect 105196 162764 105252 162820
rect 104972 162540 105028 162596
rect 108332 276780 108388 276836
rect 108332 273308 108388 273364
rect 110124 305004 110180 305060
rect 110796 369852 110852 369908
rect 110684 362124 110740 362180
rect 110684 337036 110740 337092
rect 110684 336028 110740 336084
rect 110796 335132 110852 335188
rect 110796 334572 110852 334628
rect 110348 331212 110404 331268
rect 110572 330092 110628 330148
rect 110348 300972 110404 301028
rect 110460 329532 110516 329588
rect 110236 277116 110292 277172
rect 110572 309036 110628 309092
rect 110908 304892 110964 304948
rect 111132 284508 111188 284564
rect 110460 276892 110516 276948
rect 110012 273308 110068 273364
rect 111804 389564 111860 389620
rect 111916 341292 111972 341348
rect 112252 336028 112308 336084
rect 112140 330988 112196 331044
rect 112028 330428 112084 330484
rect 112252 310716 112308 310772
rect 112364 334572 112420 334628
rect 112364 308364 112420 308420
rect 112588 317436 112644 317492
rect 112588 307356 112644 307412
rect 112140 302092 112196 302148
rect 112028 294252 112084 294308
rect 112700 292124 112756 292180
rect 112700 290668 112756 290724
rect 111916 279804 111972 279860
rect 112588 288764 112644 288820
rect 112700 279692 112756 279748
rect 112588 279020 112644 279076
rect 111804 278348 111860 278404
rect 113708 385532 113764 385588
rect 113484 374780 113540 374836
rect 113484 304892 113540 304948
rect 113596 335692 113652 335748
rect 113372 273756 113428 273812
rect 113484 278908 113540 278964
rect 111692 272076 111748 272132
rect 113708 326396 113764 326452
rect 113820 334348 113876 334404
rect 114940 331436 114996 331492
rect 114268 330988 114324 331044
rect 115836 372204 115892 372260
rect 115724 369964 115780 370020
rect 115612 368620 115668 368676
rect 115500 364700 115556 364756
rect 115052 327068 115108 327124
rect 115164 356972 115220 357028
rect 114940 317772 114996 317828
rect 115052 324156 115108 324212
rect 114268 310940 114324 310996
rect 113820 287532 113876 287588
rect 114044 279020 114100 279076
rect 113596 277004 113652 277060
rect 115052 278124 115108 278180
rect 114044 276556 114100 276612
rect 115612 340172 115668 340228
rect 115500 338604 115556 338660
rect 115724 336924 115780 336980
rect 115724 336028 115780 336084
rect 115164 274764 115220 274820
rect 115276 334572 115332 334628
rect 115388 333228 115444 333284
rect 115724 332780 115780 332836
rect 115612 331324 115668 331380
rect 115500 326732 115556 326788
rect 115724 324156 115780 324212
rect 115612 318892 115668 318948
rect 115500 312508 115556 312564
rect 115500 307356 115556 307412
rect 117516 366940 117572 366996
rect 117516 339276 117572 339332
rect 117068 339052 117124 339108
rect 116732 336812 116788 336868
rect 116396 331996 116452 332052
rect 116396 308812 116452 308868
rect 116620 331100 116676 331156
rect 116620 307692 116676 307748
rect 115836 300860 115892 300916
rect 115500 284172 115556 284228
rect 115388 279468 115444 279524
rect 115276 273644 115332 273700
rect 116956 333452 117012 333508
rect 116844 331884 116900 331940
rect 116956 282828 117012 282884
rect 117516 338492 117572 338548
rect 117292 337932 117348 337988
rect 117180 330204 117236 330260
rect 117180 285292 117236 285348
rect 117404 324156 117460 324212
rect 117404 286412 117460 286468
rect 117516 309036 117572 309092
rect 117516 283052 117572 283108
rect 117292 281708 117348 281764
rect 117068 281596 117124 281652
rect 116844 280812 116900 280868
rect 116732 271292 116788 271348
rect 121548 590716 121604 590772
rect 118524 417788 118580 417844
rect 165676 590828 165732 590884
rect 143388 380492 143444 380548
rect 174188 376348 174244 376404
rect 167468 374892 167524 374948
rect 125132 374668 125188 374724
rect 119196 366380 119252 366436
rect 118636 361340 118692 361396
rect 118860 347228 118916 347284
rect 118636 277900 118692 277956
rect 118748 336028 118804 336084
rect 118860 278460 118916 278516
rect 118972 331212 119028 331268
rect 118748 276220 118804 276276
rect 149324 371980 149380 372036
rect 147980 371644 148036 371700
rect 133868 371532 133924 371588
rect 131180 368284 131236 368340
rect 125132 364812 125188 364868
rect 126476 367164 126532 367220
rect 125804 361228 125860 361284
rect 127820 363132 127876 363188
rect 127148 361340 127204 361396
rect 129164 363020 129220 363076
rect 128492 361452 128548 361508
rect 129836 360108 129892 360164
rect 132524 365036 132580 365092
rect 132300 359996 132356 360052
rect 133196 359884 133252 359940
rect 139244 371420 139300 371476
rect 137228 368396 137284 368452
rect 135884 368172 135940 368228
rect 134540 360220 134596 360276
rect 136556 361676 136612 361732
rect 138572 367052 138628 367108
rect 137900 364812 137956 364868
rect 141932 370300 141988 370356
rect 139916 366492 139972 366548
rect 140588 364924 140644 364980
rect 141260 360444 141316 360500
rect 143948 369740 144004 369796
rect 143276 363916 143332 363972
rect 142604 361900 142660 361956
rect 143612 363132 143668 363188
rect 143612 362012 143668 362068
rect 144620 368508 144676 368564
rect 146636 366716 146692 366772
rect 145964 363244 146020 363300
rect 145292 363132 145348 363188
rect 147308 366604 147364 366660
rect 148652 361788 148708 361844
rect 162092 369964 162148 370020
rect 160076 369852 160132 369908
rect 149996 368732 150052 368788
rect 159404 368620 159460 368676
rect 152684 366828 152740 366884
rect 151228 363020 151284 363076
rect 150668 361564 150724 361620
rect 151228 360332 151284 360388
rect 151340 362908 151396 362964
rect 152012 362908 152068 362964
rect 154028 365372 154084 365428
rect 153356 362124 153412 362180
rect 156716 365260 156772 365316
rect 155372 365148 155428 365204
rect 154700 363468 154756 363524
rect 156156 362908 156212 362964
rect 155708 362124 155764 362180
rect 155708 361900 155764 361956
rect 158732 364700 158788 364756
rect 157836 362908 157892 362964
rect 158060 362124 158116 362180
rect 160748 363020 160804 363076
rect 161420 361116 161476 361172
rect 135212 359772 135268 359828
rect 130508 359660 130564 359716
rect 166796 368620 166852 368676
rect 165452 366940 165508 366996
rect 162764 366380 162820 366436
rect 164108 363356 164164 363412
rect 163436 362124 163492 362180
rect 164668 363020 164724 363076
rect 166124 364588 166180 364644
rect 161420 359548 161476 359604
rect 168812 373212 168868 373268
rect 168140 369964 168196 370020
rect 169708 371868 169764 371924
rect 169708 371308 169764 371364
rect 168812 362124 168868 362180
rect 169484 369852 169540 369908
rect 169484 368060 169540 368116
rect 171500 371756 171556 371812
rect 170828 370076 170884 370132
rect 172172 366940 172228 366996
rect 172844 363692 172900 363748
rect 174860 374780 174916 374836
rect 200732 590828 200788 590884
rect 200732 390684 200788 390740
rect 187516 373772 187572 373828
rect 199948 374892 200004 374948
rect 176876 373548 176932 373604
rect 176204 372204 176260 372260
rect 175532 371308 175588 371364
rect 180908 373436 180964 373492
rect 179564 373324 179620 373380
rect 177548 373212 177604 373268
rect 178220 370188 178276 370244
rect 178892 364588 178948 364644
rect 180236 366380 180292 366436
rect 181580 372988 181636 373044
rect 199276 371308 199332 371364
rect 184268 369628 184324 369684
rect 183596 368060 183652 368116
rect 182924 363020 182980 363076
rect 188972 367948 189028 368004
rect 186284 366268 186340 366324
rect 185612 364700 185668 364756
rect 184940 360556 184996 360612
rect 187628 363356 187684 363412
rect 188300 362908 188356 362964
rect 192556 360668 192612 360724
rect 192556 360108 192612 360164
rect 192780 360108 192836 360164
rect 166124 359548 166180 359604
rect 173516 359548 173572 359604
rect 190764 359548 190820 359604
rect 190988 359548 191044 359604
rect 192108 359548 192164 359604
rect 194012 359548 194068 359604
rect 195692 359548 195748 359604
rect 182252 359436 182308 359492
rect 186956 359436 187012 359492
rect 189644 359436 189700 359492
rect 193004 359436 193060 359492
rect 194348 359436 194404 359492
rect 120204 337484 120260 337540
rect 119196 330316 119252 330372
rect 119196 329308 119252 329364
rect 119980 334908 120036 334964
rect 119980 297052 120036 297108
rect 120092 331660 120148 331716
rect 118972 276108 119028 276164
rect 119084 290668 119140 290724
rect 118524 273644 118580 273700
rect 118412 271180 118468 271236
rect 113708 266140 113764 266196
rect 119868 281820 119924 281876
rect 119980 282940 120036 282996
rect 119196 281484 119252 281540
rect 119196 279804 119252 279860
rect 119980 279356 120036 279412
rect 119084 268604 119140 268660
rect 119196 276668 119252 276724
rect 115836 265356 115892 265412
rect 120316 335020 120372 335076
rect 120540 330652 120596 330708
rect 121548 280700 121604 280756
rect 141708 280588 141764 280644
rect 127708 280476 127764 280532
rect 133644 280476 133700 280532
rect 139692 280476 139748 280532
rect 141036 280476 141092 280532
rect 146412 280476 146468 280532
rect 163660 280476 163716 280532
rect 198156 280476 198212 280532
rect 151788 280364 151844 280420
rect 153132 280252 153188 280308
rect 166572 280140 166628 280196
rect 120540 277004 120596 277060
rect 120316 276892 120372 276948
rect 121884 280028 121940 280084
rect 120876 276780 120932 276836
rect 123004 280028 123060 280084
rect 123676 279916 123732 279972
rect 125020 279692 125076 279748
rect 125692 279916 125748 279972
rect 125692 279468 125748 279524
rect 126252 277676 126308 277732
rect 124348 277116 124404 277172
rect 122892 275996 122948 276052
rect 120204 274540 120260 274596
rect 126924 272636 126980 272692
rect 128940 272748 128996 272804
rect 127596 270172 127652 270228
rect 129612 267820 129668 267876
rect 119196 264908 119252 264964
rect 132300 279804 132356 279860
rect 131628 277788 131684 277844
rect 130956 271852 131012 271908
rect 132972 271068 133028 271124
rect 134988 279356 135044 279412
rect 135660 274876 135716 274932
rect 134316 269500 134372 269556
rect 137676 280028 137732 280084
rect 137004 278236 137060 278292
rect 136332 266812 136388 266868
rect 139020 268380 139076 268436
rect 143052 275436 143108 275492
rect 142380 271964 142436 272020
rect 145068 278572 145124 278628
rect 145740 276892 145796 276948
rect 144396 271740 144452 271796
rect 143724 268268 143780 268324
rect 147868 276780 147924 276836
rect 147868 273420 147924 273476
rect 147756 268156 147812 268212
rect 147084 266700 147140 266756
rect 140364 266588 140420 266644
rect 138348 265132 138404 265188
rect 149100 277004 149156 277060
rect 149772 276220 149828 276276
rect 151116 277116 151172 277172
rect 152460 274988 152516 275044
rect 150444 269948 150500 270004
rect 157164 275100 157220 275156
rect 156492 273532 156548 273588
rect 155820 271628 155876 271684
rect 155148 271516 155204 271572
rect 154476 270060 154532 270116
rect 157052 270508 157108 270564
rect 153804 266924 153860 266980
rect 159852 280028 159908 280084
rect 159180 277116 159236 277172
rect 159964 277116 160020 277172
rect 161196 275324 161252 275380
rect 158508 275212 158564 275268
rect 157836 268492 157892 268548
rect 157052 265356 157108 265412
rect 162540 276780 162596 276836
rect 164556 278684 164612 278740
rect 165228 277116 165284 277172
rect 167244 279580 167300 279636
rect 165900 277116 165956 277172
rect 166236 277004 166292 277060
rect 167916 276892 167972 276948
rect 168140 275548 168196 275604
rect 169260 275548 169316 275604
rect 169708 275548 169764 275604
rect 166236 272972 166292 273028
rect 163884 271404 163940 271460
rect 171276 267932 171332 267988
rect 170604 266252 170660 266308
rect 161868 265244 161924 265300
rect 148428 265020 148484 265076
rect 130284 264796 130340 264852
rect 173292 278460 173348 278516
rect 174636 278684 174692 278740
rect 173964 278348 174020 278404
rect 175308 277116 175364 277172
rect 175980 276220 176036 276276
rect 176540 275548 176596 275604
rect 177324 275548 177380 275604
rect 179340 277004 179396 277060
rect 178108 275548 178164 275604
rect 181356 275772 181412 275828
rect 180684 275660 180740 275716
rect 179900 275548 179956 275604
rect 181468 275548 181524 275604
rect 177996 271180 178052 271236
rect 172620 270284 172676 270340
rect 184044 277900 184100 277956
rect 184716 275772 184772 275828
rect 186060 275660 186116 275716
rect 186396 276556 186452 276612
rect 184828 275548 184884 275604
rect 183372 268716 183428 268772
rect 182700 267036 182756 267092
rect 185612 268604 185668 268660
rect 181468 266140 181524 266196
rect 187404 278460 187460 278516
rect 186732 276220 186788 276276
rect 188076 275884 188132 275940
rect 188748 275548 188804 275604
rect 190092 276780 190148 276836
rect 189420 275548 189476 275604
rect 186396 268604 186452 268660
rect 189084 275436 189140 275492
rect 185612 265468 185668 265524
rect 181468 265356 181524 265412
rect 171948 264572 172004 264628
rect 191436 275548 191492 275604
rect 190764 269612 190820 269668
rect 192780 276668 192836 276724
rect 194124 275660 194180 275716
rect 194572 279916 194628 279972
rect 193452 270396 193508 270452
rect 192108 268044 192164 268100
rect 195468 273644 195524 273700
rect 194796 273308 194852 273364
rect 199164 278796 199220 278852
rect 197484 276108 197540 276164
rect 196812 273756 196868 273812
rect 196140 272076 196196 272132
rect 194572 270060 194628 270116
rect 194236 266252 194292 266308
rect 199612 362908 199668 362964
rect 199388 301196 199444 301252
rect 199388 296380 199444 296436
rect 199500 280700 199556 280756
rect 199612 275436 199668 275492
rect 199276 265356 199332 265412
rect 189084 264908 189140 264964
rect 189084 264124 189140 264180
rect 199388 168028 199444 168084
rect 199164 167468 199220 167524
rect 120092 165564 120148 165620
rect 122108 165564 122164 165620
rect 127596 165564 127652 165620
rect 154028 165564 154084 165620
rect 182476 165564 182532 165620
rect 183820 165564 183876 165620
rect 184716 165564 184772 165620
rect 192332 165564 192388 165620
rect 183708 165340 183764 165396
rect 120876 164108 120932 164164
rect 126252 162876 126308 162932
rect 106876 162428 106932 162484
rect 81788 162316 81844 162372
rect 127148 163772 127204 163828
rect 126924 160860 126980 160916
rect 128492 164220 128548 164276
rect 138796 164556 138852 164612
rect 138348 162764 138404 162820
rect 137900 161980 137956 162036
rect 143836 162204 143892 162260
rect 143836 161532 143892 161588
rect 144060 161420 144116 161476
rect 128268 160748 128324 160804
rect 66332 160412 66388 160468
rect 143388 160412 143444 160468
rect 143388 159628 143444 159684
rect 127260 158956 127316 159012
rect 89852 157388 89908 157444
rect 65660 155484 65716 155540
rect 66108 157276 66164 157332
rect 64876 149212 64932 149268
rect 63980 148764 64036 148820
rect 64428 148652 64484 148708
rect 65324 152124 65380 152180
rect 65324 149100 65380 149156
rect 82908 157276 82964 157332
rect 67116 152012 67172 152068
rect 66108 148988 66164 149044
rect 65436 148876 65492 148932
rect 65436 148652 65492 148708
rect 67116 151116 67172 151172
rect 71596 152012 71652 152068
rect 71148 150556 71204 150612
rect 81900 148652 81956 148708
rect 72044 147868 72100 147924
rect 81452 147868 81508 147924
rect 82348 147868 82404 147924
rect 89180 155484 89236 155540
rect 83468 152124 83524 152180
rect 83468 149436 83524 149492
rect 83692 152124 83748 152180
rect 88620 148540 88676 148596
rect 89852 149324 89908 149380
rect 126812 150668 126868 150724
rect 125916 148540 125972 148596
rect 118748 148092 118804 148148
rect 118300 147980 118356 148036
rect 117852 147868 117908 147924
rect 126364 147868 126420 147924
rect 127708 155260 127764 155316
rect 128156 152236 128212 152292
rect 142828 151116 142884 151172
rect 138684 150332 138740 150388
rect 138012 148988 138068 149044
rect 137340 148428 137396 148484
rect 142828 150332 142884 150388
rect 142828 148988 142884 149044
rect 142828 148540 142884 148596
rect 144732 162092 144788 162148
rect 144284 161308 144340 161364
rect 144284 159628 144340 159684
rect 144396 150332 144452 150388
rect 144172 148988 144228 149044
rect 144844 160636 144900 160692
rect 145068 156268 145124 156324
rect 145180 162876 145236 162932
rect 145740 156268 145796 156324
rect 145740 149212 145796 149268
rect 145628 148876 145684 148932
rect 146076 162876 146132 162932
rect 146076 162092 146132 162148
rect 165676 162876 165732 162932
rect 166124 162988 166180 163044
rect 165228 162652 165284 162708
rect 164780 162092 164836 162148
rect 166124 161532 166180 161588
rect 166236 162876 166292 162932
rect 166236 161420 166292 161476
rect 146076 160636 146132 160692
rect 146076 149100 146132 149156
rect 146076 148876 146132 148932
rect 156828 160412 156884 160468
rect 145964 148764 146020 148820
rect 145628 148540 145684 148596
rect 171500 164556 171556 164612
rect 181804 163884 181860 163940
rect 172396 162540 172452 162596
rect 171948 162428 172004 162484
rect 166572 161308 166628 161364
rect 167916 162316 167972 162372
rect 183148 162764 183204 162820
rect 183260 164668 183316 164724
rect 182700 162204 182756 162260
rect 167916 161308 167972 161364
rect 166236 152348 166292 152404
rect 166236 150332 166292 150388
rect 164892 149212 164948 149268
rect 164556 148764 164612 148820
rect 164556 147980 164612 148036
rect 165788 148988 165844 149044
rect 164892 148204 164948 148260
rect 164444 147868 164500 147924
rect 165340 148876 165396 148932
rect 165340 148092 165396 148148
rect 165788 147196 165844 147252
rect 181916 160636 181972 160692
rect 181468 160524 181524 160580
rect 167916 145516 167972 145572
rect 171164 159180 171220 159236
rect 172060 158844 172116 158900
rect 171612 150332 171668 150388
rect 182364 159068 182420 159124
rect 182812 150780 182868 150836
rect 184716 164668 184772 164724
rect 184044 164556 184100 164612
rect 189420 164444 189476 164500
rect 189420 163324 189476 163380
rect 191660 164444 191716 164500
rect 191212 162876 191268 162932
rect 199276 164892 199332 164948
rect 199276 162764 199332 162820
rect 199164 162428 199220 162484
rect 199164 162092 199220 162148
rect 189084 148876 189140 148932
rect 188636 148540 188692 148596
rect 166236 144620 166292 144676
rect 166236 144508 166292 144564
rect 199052 144508 199108 144564
rect 199052 129276 199108 129332
rect 7532 121660 7588 121716
rect 199276 161308 199332 161364
rect 199388 148540 199444 148596
rect 202076 373660 202132 373716
rect 200620 373548 200676 373604
rect 199948 148092 200004 148148
rect 200060 366940 200116 366996
rect 200172 347564 200228 347620
rect 200172 165452 200228 165508
rect 200284 307244 200340 307300
rect 200508 305004 200564 305060
rect 200284 150780 200340 150836
rect 200508 290444 200564 290500
rect 201964 373100 202020 373156
rect 200844 371532 200900 371588
rect 200732 368284 200788 368340
rect 200732 303100 200788 303156
rect 200620 278236 200676 278292
rect 200732 299068 200788 299124
rect 200508 164108 200564 164164
rect 200396 150332 200452 150388
rect 201628 368844 201684 368900
rect 200956 365036 201012 365092
rect 201180 361452 201236 361508
rect 201068 360556 201124 360612
rect 201628 352044 201684 352100
rect 201740 365484 201796 365540
rect 201740 340844 201796 340900
rect 201852 363580 201908 363636
rect 201964 353164 202020 353220
rect 208684 373436 208740 373492
rect 207452 372988 207508 373044
rect 203308 369964 203364 370020
rect 202076 350924 202132 350980
rect 202412 363244 202468 363300
rect 201852 338604 201908 338660
rect 202300 348684 202356 348740
rect 201180 313852 201236 313908
rect 201068 308476 201124 308532
rect 201740 308364 201796 308420
rect 201740 299068 201796 299124
rect 200956 297724 201012 297780
rect 200844 292348 200900 292404
rect 201740 294924 201796 294980
rect 201628 287084 201684 287140
rect 200844 282604 200900 282660
rect 201628 280588 201684 280644
rect 201740 278012 201796 278068
rect 201852 291564 201908 291620
rect 200844 164444 200900 164500
rect 201628 275548 201684 275604
rect 200732 148876 200788 148932
rect 201180 148092 201236 148148
rect 200060 147868 200116 147924
rect 200956 147868 201012 147924
rect 199276 71932 199332 71988
rect 199724 147420 199780 147476
rect 200844 145516 200900 145572
rect 200732 129276 200788 129332
rect 200732 104076 200788 104132
rect 200844 69244 200900 69300
rect 199724 66556 199780 66612
rect 201852 269836 201908 269892
rect 201964 289324 202020 289380
rect 202076 285964 202132 286020
rect 202076 167468 202132 167524
rect 202188 283724 202244 283780
rect 202636 363132 202692 363188
rect 202636 331772 202692 331828
rect 202412 327516 202468 327572
rect 202524 329644 202580 329700
rect 202524 300748 202580 300804
rect 202636 327404 202692 327460
rect 202860 326284 202916 326340
rect 202860 310828 202916 310884
rect 202636 297052 202692 297108
rect 202860 301644 202916 301700
rect 202524 292684 202580 292740
rect 202412 275772 202468 275828
rect 202524 273084 202580 273140
rect 202412 206556 202468 206612
rect 202524 266252 202580 266308
rect 202300 168028 202356 168084
rect 202188 164892 202244 164948
rect 201964 163772 202020 163828
rect 201628 147868 201684 147924
rect 201180 79996 201236 80052
rect 200956 61180 201012 61236
rect 202748 152348 202804 152404
rect 202636 147868 202692 147924
rect 204988 369852 205044 369908
rect 204092 368060 204148 368116
rect 203308 162652 203364 162708
rect 203308 155372 203364 155428
rect 203420 343084 203476 343140
rect 203532 320684 203588 320740
rect 203644 284844 203700 284900
rect 204316 361676 204372 361732
rect 204092 187516 204148 187572
rect 204204 359548 204260 359604
rect 204316 281596 204372 281652
rect 204428 360444 204484 360500
rect 204652 360220 204708 360276
rect 204876 359996 204932 360052
rect 204876 300412 204932 300468
rect 204652 289660 204708 289716
rect 204428 262780 204484 262836
rect 204204 182812 204260 182868
rect 204204 182140 204260 182196
rect 205884 369628 205940 369684
rect 205772 364700 205828 364756
rect 204988 162988 205044 163044
rect 205100 346444 205156 346500
rect 203644 162204 203700 162260
rect 205100 160524 205156 160580
rect 205212 306124 205268 306180
rect 203532 160412 203588 160468
rect 205996 368732 206052 368788
rect 206220 368396 206276 368452
rect 206108 366492 206164 366548
rect 207340 362012 207396 362068
rect 206332 359884 206388 359940
rect 206556 359660 206612 359716
rect 207340 316540 207396 316596
rect 206556 305788 206612 305844
rect 206668 311724 206724 311780
rect 206332 295036 206388 295092
rect 206220 278908 206276 278964
rect 206108 268156 206164 268212
rect 205996 227836 206052 227892
rect 205884 184940 205940 184996
rect 205772 179452 205828 179508
rect 205212 159068 205268 159124
rect 204204 157500 204260 157556
rect 203420 152236 203476 152292
rect 204092 153804 204148 153860
rect 202860 150668 202916 150724
rect 203196 104076 203252 104132
rect 204540 157388 204596 157444
rect 204428 153692 204484 153748
rect 204204 109564 204260 109620
rect 204316 146972 204372 147028
rect 204092 101500 204148 101556
rect 206780 310828 206836 310884
rect 208348 371868 208404 371924
rect 207900 369740 207956 369796
rect 207788 368508 207844 368564
rect 207676 366716 207732 366772
rect 207564 360332 207620 360388
rect 207564 311164 207620 311220
rect 207452 195580 207508 195636
rect 207564 252028 207620 252084
rect 206780 162540 206836 162596
rect 206668 157052 206724 157108
rect 207452 155596 207508 155652
rect 204652 152124 204708 152180
rect 206892 149324 206948 149380
rect 206780 148764 206836 148820
rect 206668 148652 206724 148708
rect 206668 147196 206724 147252
rect 206780 144508 206836 144564
rect 206892 141820 206948 141876
rect 204652 117628 204708 117684
rect 207452 114940 207508 114996
rect 204540 112252 204596 112308
rect 204428 106876 204484 106932
rect 204316 98812 204372 98868
rect 203420 97468 203476 97524
rect 202748 74620 202804 74676
rect 207452 97356 207508 97412
rect 202636 63868 202692 63924
rect 207452 57820 207508 57876
rect 202524 55804 202580 55860
rect 208124 331772 208180 331828
rect 208012 325164 208068 325220
rect 208012 254716 208068 254772
rect 207900 252028 207956 252084
rect 207788 249340 207844 249396
rect 208012 249452 208068 249508
rect 207676 241276 207732 241332
rect 207676 155372 207732 155428
rect 207788 147308 207844 147364
rect 207900 145404 207956 145460
rect 208124 246652 208180 246708
rect 208236 327516 208292 327572
rect 208236 243964 208292 244020
rect 208460 366268 208516 366324
rect 208460 176764 208516 176820
rect 208572 345324 208628 345380
rect 208348 162316 208404 162372
rect 209132 371980 209188 372036
rect 208684 199052 208740 199108
rect 208796 302764 208852 302820
rect 209244 367052 209300 367108
rect 210364 376348 210420 376404
rect 210028 368172 210084 368228
rect 209580 360332 209636 360388
rect 209916 364924 209972 364980
rect 209356 359772 209412 359828
rect 209356 286972 209412 287028
rect 209244 273532 209300 273588
rect 210140 367164 210196 367220
rect 210140 322476 210196 322532
rect 210252 361340 210308 361396
rect 210252 319900 210308 319956
rect 210028 284956 210084 285012
rect 210140 297052 210196 297108
rect 209916 266028 209972 266084
rect 209132 230524 209188 230580
rect 211708 363916 211764 363972
rect 211708 325164 211764 325220
rect 217196 343532 217252 343588
rect 231644 336812 231700 336868
rect 243628 589596 243684 589652
rect 230412 330092 230468 330148
rect 253708 589596 253764 589652
rect 256844 373772 256900 373828
rect 270060 341852 270116 341908
rect 296492 360332 296548 360388
rect 275772 330204 275828 330260
rect 283276 330204 283332 330260
rect 297836 356972 297892 357028
rect 309708 380492 309764 380548
rect 319900 330092 319956 330148
rect 322924 590716 322980 590772
rect 336140 356972 336196 357028
rect 364028 590716 364084 590772
rect 341964 341852 342020 341908
rect 362572 390684 362628 390740
rect 349356 336812 349412 336868
rect 377132 361228 377188 361284
rect 375788 326284 375844 326340
rect 375564 326060 375620 326116
rect 373548 318668 373604 318724
rect 372764 317324 372820 317380
rect 371084 308588 371140 308644
rect 210364 277116 210420 277172
rect 370636 285740 370692 285796
rect 370076 265468 370132 265524
rect 370412 262108 370468 262164
rect 370076 203980 370132 204036
rect 370300 206668 370356 206724
rect 210140 161980 210196 162036
rect 370076 171388 370132 171444
rect 208796 158956 208852 159012
rect 208572 158844 208628 158900
rect 208012 131068 208068 131124
rect 208124 147084 208180 147140
rect 207900 93436 207956 93492
rect 208236 145292 208292 145348
rect 208236 96124 208292 96180
rect 208124 90748 208180 90804
rect 207788 88060 207844 88116
rect 207676 77308 207732 77364
rect 207564 50428 207620 50484
rect 199164 45276 199220 45332
rect 370188 161196 370244 161252
rect 370412 204652 370468 204708
rect 370524 245980 370580 246036
rect 370300 147868 370356 147924
rect 370636 234332 370692 234388
rect 370748 272972 370804 273028
rect 370972 269500 371028 269556
rect 370748 222572 370804 222628
rect 370860 239372 370916 239428
rect 370748 217756 370804 217812
rect 370748 209916 370804 209972
rect 370748 202188 370804 202244
rect 372204 296828 372260 296884
rect 371980 285628 372036 285684
rect 371868 274652 371924 274708
rect 371196 263004 371252 263060
rect 371196 245980 371252 246036
rect 371084 240044 371140 240100
rect 371196 234780 371252 234836
rect 371980 270284 372036 270340
rect 372092 277788 372148 277844
rect 371868 233212 371924 233268
rect 371980 240604 372036 240660
rect 370972 203084 371028 203140
rect 371868 231868 371924 231924
rect 370860 165228 370916 165284
rect 370972 173292 371028 173348
rect 370748 153804 370804 153860
rect 370524 130732 370580 130788
rect 370412 125468 370468 125524
rect 370188 89404 370244 89460
rect 370300 119868 370356 119924
rect 371756 218540 371812 218596
rect 371756 206668 371812 206724
rect 371868 199500 371924 199556
rect 371084 130956 371140 131012
rect 372652 292460 372708 292516
rect 372204 273532 372260 273588
rect 372316 286748 372372 286804
rect 372316 270172 372372 270228
rect 372428 271628 372484 271684
rect 372092 207116 372148 207172
rect 372204 264348 372260 264404
rect 372428 239484 372484 239540
rect 372540 257628 372596 257684
rect 372316 234108 372372 234164
rect 372316 205884 372372 205940
rect 372428 225932 372484 225988
rect 372204 204764 372260 204820
rect 372204 202524 372260 202580
rect 371980 130620 372036 130676
rect 372092 162988 372148 163044
rect 372204 157724 372260 157780
rect 372316 174636 372372 174692
rect 372204 155484 372260 155540
rect 372204 137452 372260 137508
rect 372092 123452 372148 123508
rect 372204 130620 372260 130676
rect 370972 90860 371028 90916
rect 372092 98812 372148 98868
rect 370412 90076 370468 90132
rect 370300 77980 370356 78036
rect 372652 229292 372708 229348
rect 372540 204428 372596 204484
rect 372652 222684 372708 222740
rect 372428 146748 372484 146804
rect 372540 180012 372596 180068
rect 372316 125132 372372 125188
rect 372204 95004 372260 95060
rect 372204 94220 372260 94276
rect 372428 109788 372484 109844
rect 372092 68348 372148 68404
rect 373324 271516 373380 271572
rect 373212 265356 373268 265412
rect 373100 265020 373156 265076
rect 372876 256060 372932 256116
rect 372876 240156 372932 240212
rect 372988 240044 373044 240100
rect 372988 225036 373044 225092
rect 372764 218652 372820 218708
rect 372988 224364 373044 224420
rect 372764 202972 372820 203028
rect 372764 153916 372820 153972
rect 373212 248668 373268 248724
rect 373100 217868 373156 217924
rect 373436 246876 373492 246932
rect 373436 233436 373492 233492
rect 375452 316988 375508 317044
rect 374108 313964 374164 314020
rect 373996 270956 374052 271012
rect 373884 264684 373940 264740
rect 373660 240268 373716 240324
rect 373884 242732 373940 242788
rect 373548 219100 373604 219156
rect 373772 240156 373828 240212
rect 373324 213164 373380 213220
rect 373436 211596 373492 211652
rect 373436 205548 373492 205604
rect 373100 196700 373156 196756
rect 373100 194908 373156 194964
rect 373212 196588 373268 196644
rect 373100 193228 373156 193284
rect 373212 190428 373268 190484
rect 373100 188972 373156 189028
rect 373324 175868 373380 175924
rect 373324 155372 373380 155428
rect 372988 150108 373044 150164
rect 372988 149100 373044 149156
rect 372652 132636 372708 132692
rect 372764 147756 372820 147812
rect 372540 96572 372596 96628
rect 372652 122220 372708 122276
rect 372652 120988 372708 121044
rect 372540 95676 372596 95732
rect 372652 80668 372708 80724
rect 372540 79996 372596 80052
rect 372428 67900 372484 67956
rect 370076 44380 370132 44436
rect 373100 132636 373156 132692
rect 372988 126588 373044 126644
rect 372988 124572 373044 124628
rect 374444 283052 374500 283108
rect 374332 271404 374388 271460
rect 374108 263788 374164 263844
rect 374220 270732 374276 270788
rect 373996 240380 374052 240436
rect 373884 238812 373940 238868
rect 373996 233436 374052 233492
rect 373884 233212 373940 233268
rect 373996 231868 374052 231924
rect 374108 217084 374164 217140
rect 375676 324380 375732 324436
rect 375676 310268 375732 310324
rect 408268 588812 408324 588868
rect 430220 385532 430276 385588
rect 494732 590156 494788 590212
rect 518476 590604 518532 590660
rect 496412 590156 496468 590212
rect 494732 383852 494788 383908
rect 562604 590492 562660 590548
rect 584668 590156 584724 590212
rect 590156 443212 590212 443268
rect 590156 437612 590212 437668
rect 540540 378812 540596 378868
rect 474348 375452 474404 375508
rect 511532 377132 511588 377188
rect 452284 372092 452340 372148
rect 386092 343532 386148 343588
rect 408940 328076 408996 328132
rect 392812 327740 392868 327796
rect 389452 327628 389508 327684
rect 378588 326172 378644 326228
rect 377132 324268 377188 324324
rect 377916 324268 377972 324324
rect 375788 305788 375844 305844
rect 377692 314636 377748 314692
rect 375564 304668 375620 304724
rect 375564 303548 375620 303604
rect 375788 297948 375844 298004
rect 375788 273420 375844 273476
rect 376908 289772 376964 289828
rect 375564 273308 375620 273364
rect 375452 270060 375508 270116
rect 376236 271180 376292 271236
rect 374444 263900 374500 263956
rect 374556 268268 374612 268324
rect 374668 267708 374724 267764
rect 376012 267708 376068 267764
rect 374668 266812 374724 266868
rect 375228 267372 375284 267428
rect 375676 266588 375732 266644
rect 375340 265580 375396 265636
rect 375340 255388 375396 255444
rect 375452 265244 375508 265300
rect 375228 245420 375284 245476
rect 375340 250012 375396 250068
rect 374556 242172 374612 242228
rect 375228 235228 375284 235284
rect 374220 215516 374276 215572
rect 374668 221116 374724 221172
rect 374668 218540 374724 218596
rect 374556 215404 374612 215460
rect 374556 215068 374612 215124
rect 374108 201516 374164 201572
rect 374332 202412 374388 202468
rect 373996 201404 374052 201460
rect 373884 180012 373940 180068
rect 373996 194796 374052 194852
rect 374556 201516 374612 201572
rect 374332 194460 374388 194516
rect 374444 195020 374500 195076
rect 374108 191660 374164 191716
rect 374444 184828 374500 184884
rect 374108 181468 374164 181524
rect 373996 178108 374052 178164
rect 374444 180684 374500 180740
rect 374332 176316 374388 176372
rect 374220 164556 374276 164612
rect 373772 130844 373828 130900
rect 373884 162540 373940 162596
rect 373772 124460 373828 124516
rect 373100 108668 373156 108724
rect 373212 124348 373268 124404
rect 373996 156828 374052 156884
rect 373996 137228 374052 137284
rect 374332 136892 374388 136948
rect 374220 131068 374276 131124
rect 374332 134540 374388 134596
rect 374108 130844 374164 130900
rect 373884 124348 373940 124404
rect 373996 127148 374052 127204
rect 373772 116508 373828 116564
rect 373996 110908 374052 110964
rect 373212 95676 373268 95732
rect 372988 95452 373044 95508
rect 372876 94444 372932 94500
rect 372876 93772 372932 93828
rect 373772 94108 373828 94164
rect 373884 108108 373940 108164
rect 373212 90860 373268 90916
rect 372988 84028 373044 84084
rect 373100 85372 373156 85428
rect 373772 90636 373828 90692
rect 373212 70700 373268 70756
rect 373324 84028 373380 84084
rect 373100 60508 373156 60564
rect 373772 69468 373828 69524
rect 374332 129948 374388 130004
rect 374332 127932 374388 127988
rect 374332 127708 374388 127764
rect 374332 127484 374388 127540
rect 374220 118748 374276 118804
rect 374220 116284 374276 116340
rect 374332 109788 374388 109844
rect 374108 98588 374164 98644
rect 374220 105308 374276 105364
rect 374108 95676 374164 95732
rect 374108 71260 374164 71316
rect 373884 67228 373940 67284
rect 374220 62524 374276 62580
rect 374332 104076 374388 104132
rect 374332 103068 374388 103124
rect 375116 208460 375172 208516
rect 375452 247548 375508 247604
rect 375564 259868 375620 259924
rect 375340 235116 375396 235172
rect 375452 246876 375508 246932
rect 375452 213276 375508 213332
rect 375228 199388 375284 199444
rect 375452 209468 375508 209524
rect 375116 197708 375172 197764
rect 375900 261660 375956 261716
rect 375676 205996 375732 206052
rect 375788 256508 375844 256564
rect 375564 204876 375620 204932
rect 375900 237692 375956 237748
rect 375788 204316 375844 204372
rect 375900 237468 375956 237524
rect 375900 203868 375956 203924
rect 375900 200956 375956 201012
rect 375900 199276 375956 199332
rect 375452 197596 375508 197652
rect 375900 196028 375956 196084
rect 375788 195132 375844 195188
rect 375676 192444 375732 192500
rect 375452 190092 375508 190148
rect 375228 186508 375284 186564
rect 375228 160188 375284 160244
rect 375340 164668 375396 164724
rect 374556 152684 374612 152740
rect 375228 155372 375284 155428
rect 374556 151116 374612 151172
rect 375228 147084 375284 147140
rect 375228 145628 375284 145684
rect 375228 130956 375284 131012
rect 375228 129276 375284 129332
rect 375452 151116 375508 151172
rect 375564 170268 375620 170324
rect 375452 145628 375508 145684
rect 375452 137116 375508 137172
rect 375340 128828 375396 128884
rect 374556 115612 374612 115668
rect 374444 87276 374500 87332
rect 374556 107548 374612 107604
rect 374444 85596 374500 85652
rect 374444 84028 374500 84084
rect 374332 61180 374388 61236
rect 374444 72156 374500 72212
rect 374556 64540 374612 64596
rect 375452 104188 375508 104244
rect 375452 61852 375508 61908
rect 374444 59388 374500 59444
rect 373324 58268 373380 58324
rect 374556 52668 374612 52724
rect 375676 163884 375732 163940
rect 375676 161868 375732 161924
rect 375788 155372 375844 155428
rect 376124 265468 376180 265524
rect 376124 253148 376180 253204
rect 376012 173292 376068 173348
rect 376124 248892 376180 248948
rect 375900 133868 375956 133924
rect 376012 147868 376068 147924
rect 375788 123228 375844 123284
rect 375676 110908 375732 110964
rect 375788 82684 375844 82740
rect 375900 106428 375956 106484
rect 375676 68572 375732 68628
rect 376236 240268 376292 240324
rect 376684 239484 376740 239540
rect 376684 239260 376740 239316
rect 376236 225260 376292 225316
rect 376236 220444 376292 220500
rect 376236 219100 376292 219156
rect 376236 213276 376292 213332
rect 376236 204988 376292 205044
rect 377356 269724 377412 269780
rect 377356 243292 377412 243348
rect 377244 241276 377300 241332
rect 377132 239260 377188 239316
rect 376908 202636 376964 202692
rect 377020 236572 377076 236628
rect 376236 190092 376292 190148
rect 376124 132188 376180 132244
rect 376236 171948 376292 172004
rect 377020 167244 377076 167300
rect 377132 166572 377188 166628
rect 377244 165900 377300 165956
rect 377244 164668 377300 164724
rect 377356 164556 377412 164612
rect 377468 246652 377524 246708
rect 377468 163212 377524 163268
rect 377580 243964 377636 244020
rect 377916 303212 377972 303268
rect 377692 227836 377748 227892
rect 377804 290444 377860 290500
rect 377916 283724 377972 283780
rect 377916 276332 377972 276388
rect 378028 235116 378084 235172
rect 377804 202412 377860 202468
rect 377580 160524 377636 160580
rect 376348 160188 376404 160244
rect 377356 159852 377412 159908
rect 376348 156492 376404 156548
rect 377020 157836 377076 157892
rect 376796 153916 376852 153972
rect 376796 153132 376852 153188
rect 377132 155148 377188 155204
rect 377244 153804 377300 153860
rect 377244 141036 377300 141092
rect 377244 140028 377300 140084
rect 377132 138908 377188 138964
rect 377020 135548 377076 135604
rect 377020 134652 377076 134708
rect 377468 159516 377524 159572
rect 377468 159068 377524 159124
rect 377468 154476 377524 154532
rect 377468 153132 377524 153188
rect 377468 141148 377524 141204
rect 377356 135884 377412 135940
rect 377356 134428 377412 134484
rect 377580 133420 377636 133476
rect 377692 163212 377748 163268
rect 377468 132076 377524 132132
rect 376236 98812 376292 98868
rect 376348 130732 376404 130788
rect 376124 97692 376180 97748
rect 377132 128828 377188 128884
rect 377020 98588 377076 98644
rect 376348 95228 376404 95284
rect 376460 96572 376516 96628
rect 376012 91420 376068 91476
rect 376012 90636 376068 90692
rect 376460 82908 376516 82964
rect 375900 63196 375956 63252
rect 376236 70476 376292 70532
rect 377244 128604 377300 128660
rect 377244 127148 377300 127204
rect 377356 99708 377412 99764
rect 377356 99148 377412 99204
rect 377132 71932 377188 71988
rect 377244 84700 377300 84756
rect 377244 70476 377300 70532
rect 377580 131628 377636 131684
rect 377804 157836 377860 157892
rect 377804 157164 377860 157220
rect 377916 202636 377972 202692
rect 377916 202076 377972 202132
rect 377916 155820 377972 155876
rect 377916 136668 377972 136724
rect 377916 135324 377972 135380
rect 377916 134316 377972 134372
rect 392140 325948 392196 326004
rect 408268 327740 408324 327796
rect 406252 326284 406308 326340
rect 397516 326172 397572 326228
rect 398188 325948 398244 326004
rect 406924 326060 406980 326116
rect 419692 327964 419748 328020
rect 409612 327852 409668 327908
rect 417004 326172 417060 326228
rect 414316 324940 414372 324996
rect 417676 326060 417732 326116
rect 421036 327740 421092 327796
rect 421708 327628 421764 327684
rect 440300 325948 440356 326004
rect 423948 324940 424004 324996
rect 390124 324492 390180 324548
rect 396844 324492 396900 324548
rect 410956 324380 411012 324436
rect 418348 324380 418404 324436
rect 418796 324380 418852 324436
rect 420812 324380 420868 324436
rect 422044 324380 422100 324436
rect 422604 324380 422660 324436
rect 424172 324380 424228 324436
rect 425068 324380 425124 324436
rect 426188 324380 426244 324436
rect 426412 324380 426468 324436
rect 440188 309932 440244 309988
rect 439292 305788 439348 305844
rect 379260 288428 379316 288484
rect 379148 287756 379204 287812
rect 378924 287084 378980 287140
rect 378812 261548 378868 261604
rect 378812 239372 378868 239428
rect 378588 222684 378644 222740
rect 378812 227836 378868 227892
rect 378588 221788 378644 221844
rect 378700 222572 378756 222628
rect 378700 180684 378756 180740
rect 378028 132076 378084 132132
rect 378140 163884 378196 163940
rect 377692 131516 377748 131572
rect 377804 131964 377860 132020
rect 377580 130844 377636 130900
rect 377804 130732 377860 130788
rect 377916 131852 377972 131908
rect 377916 130620 377972 130676
rect 377916 128716 377972 128772
rect 377916 127596 377972 127652
rect 378028 127932 378084 127988
rect 377804 127484 377860 127540
rect 377692 124572 377748 124628
rect 377692 124348 377748 124404
rect 377468 96348 377524 96404
rect 377580 100828 377636 100884
rect 377356 66556 377412 66612
rect 377020 65884 377076 65940
rect 377692 73948 377748 74004
rect 377804 73276 377860 73332
rect 378252 157724 378308 157780
rect 378252 157388 378308 157444
rect 378252 139356 378308 139412
rect 378700 149324 378756 149380
rect 378700 148988 378756 149044
rect 378924 207340 378980 207396
rect 379036 284396 379092 284452
rect 379148 205324 379204 205380
rect 379036 204540 379092 204596
rect 379932 271740 379988 271796
rect 379484 264460 379540 264516
rect 379260 204204 379316 204260
rect 379372 263340 379428 263396
rect 379260 203868 379316 203924
rect 379036 197372 379092 197428
rect 378924 171388 378980 171444
rect 379036 161196 379092 161252
rect 379148 196252 379204 196308
rect 378924 147868 378980 147924
rect 378812 145068 378868 145124
rect 378812 144508 378868 144564
rect 378700 135436 378756 135492
rect 378812 141036 378868 141092
rect 378140 122108 378196 122164
rect 378140 120988 378196 121044
rect 378700 125244 378756 125300
rect 378700 107548 378756 107604
rect 377916 70588 377972 70644
rect 377580 65212 377636 65268
rect 376236 52668 376292 52724
rect 375564 44716 375620 44772
rect 378924 139356 378980 139412
rect 378924 137788 378980 137844
rect 379372 172620 379428 172676
rect 379596 263564 379652 263620
rect 379596 246652 379652 246708
rect 379820 263116 379876 263172
rect 379820 243964 379876 244020
rect 380044 271180 380100 271236
rect 381388 271404 381444 271460
rect 380716 270956 380772 271012
rect 381388 271068 381444 271124
rect 383404 271516 383460 271572
rect 384076 271292 384132 271348
rect 382732 270844 382788 270900
rect 382060 270732 382116 270788
rect 381388 269836 381444 269892
rect 385420 272076 385476 272132
rect 384748 268380 384804 268436
rect 387436 269500 387492 269556
rect 386764 268492 386820 268548
rect 388108 268268 388164 268324
rect 386092 268156 386148 268212
rect 379932 241164 379988 241220
rect 380044 267932 380100 267988
rect 379820 240268 379876 240324
rect 379708 234332 379764 234388
rect 380268 266924 380324 266980
rect 380156 263452 380212 263508
rect 380156 243180 380212 243236
rect 390124 272076 390180 272132
rect 394156 271516 394212 271572
rect 390124 271404 390180 271460
rect 389452 271068 389508 271124
rect 401548 270060 401604 270116
rect 404236 269836 404292 269892
rect 403564 267484 403620 267540
rect 403564 265692 403620 265748
rect 388780 265020 388836 265076
rect 405132 269836 405188 269892
rect 406252 271964 406308 272020
rect 406476 273196 406532 273252
rect 405580 267932 405636 267988
rect 405580 267372 405636 267428
rect 408268 273420 408324 273476
rect 407596 273308 407652 273364
rect 409612 271628 409668 271684
rect 410060 271068 410116 271124
rect 410284 273308 410340 273364
rect 408940 270172 408996 270228
rect 409836 270956 409892 271012
rect 406924 268044 406980 268100
rect 409612 267932 409668 267988
rect 408716 267708 408772 267764
rect 407596 265356 407652 265412
rect 408940 267260 408996 267316
rect 409836 267708 409892 267764
rect 410956 271180 411012 271236
rect 410956 270284 411012 270340
rect 413644 273532 413700 273588
rect 412972 271852 413028 271908
rect 412300 271068 412356 271124
rect 414316 271068 414372 271124
rect 417004 271740 417060 271796
rect 417452 271740 417508 271796
rect 416332 271628 416388 271684
rect 415660 271068 415716 271124
rect 414988 270172 415044 270228
rect 411628 269724 411684 269780
rect 415660 269948 415716 270004
rect 414988 267708 415044 267764
rect 410956 265692 411012 265748
rect 412972 266812 413028 266868
rect 410284 265356 410340 265412
rect 412300 265580 412356 265636
rect 411628 265244 411684 265300
rect 414316 265468 414372 265524
rect 417452 267596 417508 267652
rect 416332 267148 416388 267204
rect 419692 271068 419748 271124
rect 419916 271628 419972 271684
rect 417676 266924 417732 266980
rect 418348 268044 418404 268100
rect 420364 270284 420420 270340
rect 419916 267932 419972 267988
rect 420028 268716 420084 268772
rect 420028 266588 420084 266644
rect 430444 268716 430500 268772
rect 423052 267484 423108 267540
rect 429772 267820 429828 267876
rect 420364 267148 420420 267204
rect 423388 267372 423444 267428
rect 404908 264460 404964 264516
rect 417004 264460 417060 264516
rect 440188 272972 440244 273028
rect 439292 264684 439348 264740
rect 440188 268044 440244 268100
rect 423388 264460 423444 264516
rect 406252 264348 406308 264404
rect 403564 264236 403620 264292
rect 406252 264236 406308 264292
rect 406924 264236 406980 264292
rect 410956 264236 411012 264292
rect 413644 264236 413700 264292
rect 380268 237580 380324 237636
rect 380492 242172 380548 242228
rect 380044 236796 380100 236852
rect 379932 221676 379988 221732
rect 379932 218316 379988 218372
rect 380380 215292 380436 215348
rect 379708 202188 379764 202244
rect 379484 171948 379540 172004
rect 379596 198492 379652 198548
rect 379372 171388 379428 171444
rect 379260 135212 379316 135268
rect 379484 159180 379540 159236
rect 379148 134092 379204 134148
rect 378924 44828 378980 44884
rect 379036 132300 379092 132356
rect 379372 131740 379428 131796
rect 379148 123900 379204 123956
rect 379260 121996 379316 122052
rect 379260 104076 379316 104132
rect 379148 99148 379204 99204
rect 379260 96348 379316 96404
rect 379036 92988 379092 93044
rect 378812 43036 378868 43092
rect 379148 95004 379204 95060
rect 379260 46284 379316 46340
rect 379932 196140 379988 196196
rect 379932 176316 379988 176372
rect 379596 134204 379652 134260
rect 379708 167244 379764 167300
rect 379708 127484 379764 127540
rect 379820 165228 379876 165284
rect 379484 125468 379540 125524
rect 380268 198380 380324 198436
rect 379932 155484 379988 155540
rect 380156 146188 380212 146244
rect 380604 240380 380660 240436
rect 381836 205660 381892 205716
rect 382060 205660 382116 205716
rect 383404 205660 383460 205716
rect 380492 201404 380548 201460
rect 380380 197484 380436 197540
rect 382620 203196 382676 203252
rect 384748 205660 384804 205716
rect 384076 205436 384132 205492
rect 417004 205436 417060 205492
rect 419244 205324 419300 205380
rect 383628 203196 383684 203252
rect 385420 205212 385476 205268
rect 381388 202972 381444 203028
rect 384188 202748 384244 202804
rect 384636 202748 384692 202804
rect 384636 202412 384692 202468
rect 384636 202076 384692 202132
rect 386092 205212 386148 205268
rect 386764 205212 386820 205268
rect 386092 198492 386148 198548
rect 386428 203084 386484 203140
rect 384972 198380 385028 198436
rect 389452 205212 389508 205268
rect 387436 203084 387492 203140
rect 388108 201404 388164 201460
rect 388220 203196 388276 203252
rect 386764 198268 386820 198324
rect 388444 201292 388500 201348
rect 389452 203196 389508 203252
rect 399532 205100 399588 205156
rect 388780 201292 388836 201348
rect 388444 196364 388500 196420
rect 391468 204988 391524 205044
rect 390460 202748 390516 202804
rect 390908 202748 390964 202804
rect 402220 203868 402276 203924
rect 400204 202748 400260 202804
rect 391468 201180 391524 201236
rect 398188 201628 398244 201684
rect 389788 198044 389844 198100
rect 388220 196252 388276 196308
rect 389788 196140 389844 196196
rect 386428 196028 386484 196084
rect 402220 201852 402276 201908
rect 403340 205100 403396 205156
rect 406924 204428 406980 204484
rect 407596 204988 407652 205044
rect 404908 201628 404964 201684
rect 404908 201404 404964 201460
rect 403340 197036 403396 197092
rect 403564 197820 403620 197876
rect 405580 197708 405636 197764
rect 408268 204876 408324 204932
rect 410284 204652 410340 204708
rect 410956 205100 411012 205156
rect 408940 204316 408996 204372
rect 408940 199500 408996 199556
rect 410284 199388 410340 199444
rect 409612 197596 409668 197652
rect 412300 204764 412356 204820
rect 413644 205100 413700 205156
rect 412972 202860 413028 202916
rect 414316 204540 414372 204596
rect 411628 202636 411684 202692
rect 414316 202412 414372 202468
rect 414764 204988 414820 205044
rect 410956 199388 411012 199444
rect 411628 201180 411684 201236
rect 410956 197036 411012 197092
rect 413420 200956 413476 201012
rect 412300 197932 412356 197988
rect 415660 203980 415716 204036
rect 416332 202972 416388 203028
rect 416668 204204 416724 204260
rect 416668 202972 416724 203028
rect 414988 202860 415044 202916
rect 416556 202860 416612 202916
rect 418572 204988 418628 205044
rect 418348 204092 418404 204148
rect 418348 203196 418404 203252
rect 417676 202524 417732 202580
rect 418572 203084 418628 203140
rect 418460 202300 418516 202356
rect 419692 204204 419748 204260
rect 423052 202972 423108 203028
rect 423052 202636 423108 202692
rect 427084 203196 427140 203252
rect 427084 202524 427140 202580
rect 429772 203084 429828 203140
rect 419020 202188 419076 202244
rect 429772 201628 429828 201684
rect 416556 199612 416612 199668
rect 417676 201068 417732 201124
rect 414764 199500 414820 199556
rect 417004 199276 417060 199332
rect 416332 197484 416388 197540
rect 439404 199388 439460 199444
rect 418348 198156 418404 198212
rect 423500 194796 423556 194852
rect 398188 194572 398244 194628
rect 423500 194572 423556 194628
rect 380044 137452 380100 137508
rect 380044 132412 380100 132468
rect 380380 136668 380436 136724
rect 380492 138908 380548 138964
rect 379820 124348 379876 124404
rect 380380 127148 380436 127204
rect 379484 123788 379540 123844
rect 379484 105308 379540 105364
rect 379596 120988 379652 121044
rect 379372 91868 379428 91924
rect 379148 44268 379204 44324
rect 379484 95228 379540 95284
rect 379596 82012 379652 82068
rect 380268 123676 380324 123732
rect 380268 106428 380324 106484
rect 380380 100828 380436 100884
rect 380380 97692 380436 97748
rect 379484 46172 379540 46228
rect 379820 65548 379876 65604
rect 380268 44604 380324 44660
rect 379372 43148 379428 43204
rect 380716 135660 380772 135716
rect 380940 135660 380996 135716
rect 381388 135996 381444 136052
rect 381388 132636 381444 132692
rect 382060 135660 382116 135716
rect 383628 135660 383684 135716
rect 385420 135660 385476 135716
rect 384748 135212 384804 135268
rect 382732 134764 382788 134820
rect 381836 132636 381892 132692
rect 383404 132636 383460 132692
rect 384076 132524 384132 132580
rect 388780 135660 388836 135716
rect 396844 135660 396900 135716
rect 397516 135660 397572 135716
rect 384972 132524 385028 132580
rect 385644 134204 385700 134260
rect 386092 134204 386148 134260
rect 385644 132524 385700 132580
rect 386428 134092 386484 134148
rect 381724 132412 381780 132468
rect 381724 132076 381780 132132
rect 384524 132188 384580 132244
rect 384524 131628 384580 131684
rect 386764 134092 386820 134148
rect 386540 133868 386596 133924
rect 387436 133868 387492 133924
rect 388108 134316 388164 134372
rect 386540 132524 386596 132580
rect 386428 131628 386484 131684
rect 389452 133980 389508 134036
rect 389452 131404 389508 131460
rect 398188 135100 398244 135156
rect 398188 134876 398244 134932
rect 398188 131068 398244 131124
rect 404236 131740 404292 131796
rect 388108 129164 388164 129220
rect 382172 129052 382228 129108
rect 410956 132188 411012 132244
rect 410284 132076 410340 132132
rect 412300 132412 412356 132468
rect 412972 132300 413028 132356
rect 411628 131964 411684 132020
rect 414316 132524 414372 132580
rect 414876 132636 414932 132692
rect 413644 131852 413700 131908
rect 409612 129276 409668 129332
rect 411516 131628 411572 131684
rect 404236 129052 404292 129108
rect 411516 127148 411572 127204
rect 414092 131180 414148 131236
rect 414988 132412 415044 132468
rect 415660 132524 415716 132580
rect 415660 131628 415716 131684
rect 416332 132188 416388 132244
rect 414988 131180 415044 131236
rect 414876 128940 414932 128996
rect 414092 123900 414148 123956
rect 382172 122220 382228 122276
rect 417004 132076 417060 132132
rect 418348 132636 418404 132692
rect 419020 134204 419076 134260
rect 417452 132300 417508 132356
rect 417900 132076 417956 132132
rect 439404 132524 439460 132580
rect 419244 131964 419300 132020
rect 417900 125356 417956 125412
rect 417452 123788 417508 123844
rect 441980 310604 442036 310660
rect 441868 307244 441924 307300
rect 440524 276332 440580 276388
rect 440300 201404 440356 201460
rect 440412 267932 440468 267988
rect 440188 131740 440244 131796
rect 440300 196700 440356 196756
rect 419244 125244 419300 125300
rect 419132 123676 419188 123732
rect 416332 121996 416388 122052
rect 442092 309260 442148 309316
rect 442092 275548 442148 275604
rect 441980 274652 442036 274708
rect 441868 270396 441924 270452
rect 445228 267708 445284 267764
rect 442316 267260 442372 267316
rect 441980 265356 442036 265412
rect 440524 202860 440580 202916
rect 440636 205548 440692 205604
rect 440412 161868 440468 161924
rect 440524 202524 440580 202580
rect 440300 83356 440356 83412
rect 440412 136892 440468 136948
rect 441868 194460 441924 194516
rect 441868 177324 441924 177380
rect 440636 171948 440692 172004
rect 442204 228508 442260 228564
rect 442092 226492 442148 226548
rect 443660 266812 443716 266868
rect 443548 263340 443604 263396
rect 442204 206556 442260 206612
rect 442092 201516 442148 201572
rect 442316 193340 442372 193396
rect 442204 191772 442260 191828
rect 442204 172620 442260 172676
rect 442092 170604 442148 170660
rect 441980 163212 442036 163268
rect 442652 164556 442708 164612
rect 442316 162876 442372 162932
rect 442540 163884 442596 163940
rect 442204 161196 442260 161252
rect 442092 159852 442148 159908
rect 441868 157836 441924 157892
rect 442092 137340 442148 137396
rect 442092 137004 442148 137060
rect 441868 134988 441924 135044
rect 441980 135436 442036 135492
rect 440524 134204 440580 134260
rect 440412 81340 440468 81396
rect 380604 67452 380660 67508
rect 380492 45948 380548 46004
rect 442428 160524 442484 160580
rect 442204 134316 442260 134372
rect 442316 159180 442372 159236
rect 442428 135324 442484 135380
rect 442316 130172 442372 130228
rect 442652 137340 442708 137396
rect 442876 135548 442932 135604
rect 442652 128604 442708 128660
rect 442764 133644 442820 133700
rect 442540 125916 442596 125972
rect 442316 125132 442372 125188
rect 442428 123452 442484 123508
rect 442428 89404 442484 89460
rect 442316 87388 442372 87444
rect 441980 69244 442036 69300
rect 442988 128716 443044 128772
rect 443660 137228 443716 137284
rect 443772 191660 443828 191716
rect 443548 124236 443604 124292
rect 443660 128492 443716 128548
rect 445340 263004 445396 263060
rect 448588 196588 448644 196644
rect 446908 195020 446964 195076
rect 445340 137116 445396 137172
rect 445452 194572 445508 194628
rect 445228 135100 445284 135156
rect 445564 193228 445620 193284
rect 448588 84700 448644 84756
rect 446908 78652 446964 78708
rect 445564 77980 445620 78036
rect 445452 77308 445508 77364
rect 443772 75964 443828 76020
rect 443660 75292 443716 75348
rect 442876 69916 442932 69972
rect 457772 69916 457828 69972
rect 442764 68572 442820 68628
rect 441868 66556 441924 66612
rect 457772 46956 457828 47012
rect 381388 45724 381444 45780
rect 382060 45724 382116 45780
rect 384076 45724 384132 45780
rect 384748 45724 384804 45780
rect 388108 45724 388164 45780
rect 396844 45724 396900 45780
rect 398188 45724 398244 45780
rect 403564 45724 403620 45780
rect 417676 45724 417732 45780
rect 390460 45666 390516 45668
rect 390460 45614 390462 45666
rect 390462 45614 390514 45666
rect 390514 45614 390516 45666
rect 390460 45612 390516 45614
rect 397852 45666 397908 45668
rect 397852 45614 397854 45666
rect 397854 45614 397906 45666
rect 397906 45614 397908 45666
rect 397852 45612 397908 45614
rect 418348 45612 418404 45668
rect 382732 45500 382788 45556
rect 383852 45500 383908 45556
rect 384972 45500 385028 45556
rect 386428 45500 386484 45556
rect 386988 45500 387044 45556
rect 389004 45500 389060 45556
rect 391916 45500 391972 45556
rect 412972 45500 413028 45556
rect 388332 45388 388388 45444
rect 407596 45388 407652 45444
rect 386092 45164 386148 45220
rect 405580 45164 405636 45220
rect 380380 42924 380436 42980
rect 398860 44268 398916 44324
rect 396172 42924 396228 42980
rect 379036 42700 379092 42756
rect 402892 45052 402948 45108
rect 400876 43596 400932 43652
rect 406252 44716 406308 44772
rect 406924 44380 406980 44436
rect 404236 43484 404292 43540
rect 400204 43148 400260 43204
rect 399532 42700 399588 42756
rect 374556 41916 374612 41972
rect 372764 41804 372820 41860
rect 410956 44828 411012 44884
rect 416332 45052 416388 45108
rect 415660 43484 415716 43540
rect 419692 43596 419748 43652
rect 420364 43596 420420 43652
rect 421036 43372 421092 43428
rect 423052 44604 423108 44660
rect 422380 43260 422436 43316
rect 417004 43148 417060 43204
rect 414316 43036 414372 43092
rect 413644 42924 413700 42980
rect 410284 42812 410340 42868
rect 485548 45052 485604 45108
rect 484876 43596 484932 43652
rect 484204 43484 484260 43540
rect 540092 350700 540148 350756
rect 511532 43484 511588 43540
rect 512428 69916 512484 69972
rect 512540 69244 512596 69300
rect 512540 45276 512596 45332
rect 573692 337484 573748 337540
rect 573692 45052 573748 45108
rect 540092 43596 540148 43652
rect 512428 41916 512484 41972
rect 423724 41804 423780 41860
rect 409612 41692 409668 41748
rect 408940 40236 408996 40292
rect 4284 8764 4340 8820
rect 396396 5516 396452 5572
rect 437612 5516 437668 5572
rect 401324 5404 401380 5460
rect 382508 5292 382564 5348
rect 420140 5292 420196 5348
rect 353612 5180 353668 5236
rect 386652 5180 386708 5236
rect 429548 5180 429604 5236
rect 15372 5068 15428 5124
rect 28700 4956 28756 5012
rect 21084 3388 21140 3444
rect 19180 2604 19236 2660
rect 17276 2492 17332 2548
rect 26796 2828 26852 2884
rect 24892 2716 24948 2772
rect 30604 4844 30660 4900
rect 40124 4732 40180 4788
rect 36316 3164 36372 3220
rect 34412 3052 34468 3108
rect 32508 2940 32564 2996
rect 38220 2156 38276 2212
rect 43932 4620 43988 4676
rect 41916 2380 41972 2436
rect 11676 28 11732 84
rect 13580 140 13636 196
rect 23100 252 23156 308
rect 45836 4508 45892 4564
rect 44716 28 44772 84
rect 47852 5068 47908 5124
rect 47740 4396 47796 4452
rect 50988 2604 51044 2660
rect 51548 4284 51604 4340
rect 49420 2492 49476 2548
rect 49644 2268 49700 2324
rect 51996 3388 52052 3444
rect 53452 4172 53508 4228
rect 46284 140 46340 196
rect 58940 4956 58996 5012
rect 60396 4844 60452 4900
rect 57260 2828 57316 2884
rect 57372 4060 57428 4116
rect 55692 2716 55748 2772
rect 55356 2492 55412 2548
rect 61068 3948 61124 4004
rect 59164 2604 59220 2660
rect 63532 3052 63588 3108
rect 64876 4844 64932 4900
rect 61964 2940 62020 2996
rect 62972 2716 63028 2772
rect 65100 3164 65156 3220
rect 68236 4732 68292 4788
rect 68684 4956 68740 5012
rect 66668 2156 66724 2212
rect 66780 2828 66836 2884
rect 69804 2380 69860 2436
rect 70476 4732 70532 4788
rect 71372 4620 71428 4676
rect 72492 4620 72548 4676
rect 72940 4508 72996 4564
rect 73052 4956 73108 5012
rect 73052 3948 73108 4004
rect 74396 4508 74452 4564
rect 74508 4396 74564 4452
rect 76076 2268 76132 2324
rect 76300 4396 76356 4452
rect 77644 4284 77700 4340
rect 78204 4284 78260 4340
rect 79212 4172 79268 4228
rect 80108 2940 80164 2996
rect 80780 2492 80836 2548
rect 82012 4172 82068 4228
rect 82348 4060 82404 4116
rect 84812 4956 84868 5012
rect 85820 4956 85876 5012
rect 83244 2604 83300 2660
rect 83916 4060 83972 4116
rect 88620 4844 88676 4900
rect 89628 4844 89684 4900
rect 87052 2716 87108 2772
rect 87724 2492 87780 2548
rect 91756 5068 91812 5124
rect 93324 4732 93380 4788
rect 94892 4620 94948 4676
rect 95340 4732 95396 4788
rect 90188 2828 90244 2884
rect 93436 2716 93492 2772
rect 91532 2604 91588 2660
rect 96460 4508 96516 4564
rect 98028 4396 98084 4452
rect 99036 4620 99092 4676
rect 97244 2828 97300 2884
rect 99596 4284 99652 4340
rect 101052 4508 101108 4564
rect 102732 4172 102788 4228
rect 102956 4396 103012 4452
rect 101164 2940 101220 2996
rect 105980 4956 106036 5012
rect 106764 4956 106820 5012
rect 104300 4060 104356 4116
rect 104860 4284 104916 4340
rect 109004 4844 109060 4900
rect 107436 2492 107492 2548
rect 108668 4172 108724 4228
rect 109900 2604 109956 2660
rect 110572 4844 110628 4900
rect 113708 4732 113764 4788
rect 112140 2716 112196 2772
rect 112476 4060 112532 4116
rect 116844 4620 116900 4676
rect 118412 4508 118468 4564
rect 119980 4396 120036 4452
rect 120092 4732 120148 4788
rect 115276 2828 115332 2884
rect 118188 2716 118244 2772
rect 116284 2604 116340 2660
rect 114380 2492 114436 2548
rect 122668 4956 122724 5012
rect 123900 4956 123956 5012
rect 121548 4284 121604 4340
rect 121996 2828 122052 2884
rect 126252 4844 126308 4900
rect 127596 4844 127652 4900
rect 124684 4172 124740 4228
rect 125804 4620 125860 4676
rect 127820 4060 127876 4116
rect 129388 2492 129444 2548
rect 129612 4508 129668 4564
rect 130956 2604 131012 2660
rect 131516 4396 131572 4452
rect 134092 4732 134148 4788
rect 136556 4956 136612 5012
rect 138796 4620 138852 4676
rect 139132 4956 139188 5012
rect 135660 2828 135716 2884
rect 132524 2716 132580 2772
rect 137228 2716 137284 2772
rect 135324 2604 135380 2660
rect 133420 2492 133476 2548
rect 140364 4844 140420 4900
rect 141036 4844 141092 4900
rect 141932 4508 141988 4564
rect 142940 4732 142996 4788
rect 143500 4396 143556 4452
rect 144844 4620 144900 4676
rect 146636 2604 146692 2660
rect 146748 4508 146804 4564
rect 145068 2492 145124 2548
rect 149548 4956 149604 5012
rect 151340 4844 151396 4900
rect 152908 4732 152964 4788
rect 154476 4620 154532 4676
rect 156044 4508 156100 4564
rect 148204 2716 148260 2772
rect 148652 4396 148708 4452
rect 157612 4396 157668 4452
rect 158172 4620 158228 4676
rect 150556 3724 150612 3780
rect 152460 3612 152516 3668
rect 154364 3500 154420 3556
rect 156156 3388 156212 3444
rect 159180 3724 159236 3780
rect 160076 4956 160132 5012
rect 160748 3612 160804 3668
rect 161980 3836 162036 3892
rect 162316 3500 162372 3556
rect 166348 4956 166404 5012
rect 165452 4620 165508 4676
rect 168588 3836 168644 3892
rect 163884 3388 163940 3444
rect 164108 3724 164164 3780
rect 170156 3724 170212 3780
rect 165788 3612 165844 3668
rect 171724 3612 171780 3668
rect 167692 3500 167748 3556
rect 173292 3500 173348 3556
rect 169596 3388 169652 3444
rect 174860 3388 174916 3444
rect 175308 2716 175364 2772
rect 173404 2604 173460 2660
rect 171500 2492 171556 2548
rect 179564 2716 179620 2772
rect 177996 2604 178052 2660
rect 179116 2604 179172 2660
rect 176428 2492 176484 2548
rect 177212 2380 177268 2436
rect 181020 2492 181076 2548
rect 182700 2604 182756 2660
rect 182924 2604 182980 2660
rect 181132 2380 181188 2436
rect 185836 2604 185892 2660
rect 186732 3500 186788 3556
rect 184268 2492 184324 2548
rect 184716 2492 184772 2548
rect 188972 3500 189028 3556
rect 187404 2492 187460 2548
rect 188636 3388 188692 3444
rect 190540 3388 190596 3444
rect 54124 252 54180 308
rect 210924 3500 210980 3556
rect 209356 3388 209412 3444
rect 211260 3388 211316 3444
rect 212492 3388 212548 3444
rect 213164 3500 213220 3556
rect 214060 3500 214116 3556
rect 215068 3388 215124 3444
rect 215628 3388 215684 3444
rect 216972 3500 217028 3556
rect 218764 3612 218820 3668
rect 217196 3500 217252 3556
rect 218876 3388 218932 3444
rect 220332 3388 220388 3444
rect 220780 3500 220836 3556
rect 221900 3500 221956 3556
rect 222684 3612 222740 3668
rect 223468 3612 223524 3668
rect 224588 3388 224644 3444
rect 225036 2492 225092 2548
rect 226492 3500 226548 3556
rect 226604 2604 226660 2660
rect 228172 2380 228228 2436
rect 228508 3612 228564 3668
rect 229740 2828 229796 2884
rect 231308 2716 231364 2772
rect 232204 2604 232260 2660
rect 230300 2492 230356 2548
rect 242284 4620 242340 4676
rect 240716 4508 240772 4564
rect 239148 4396 239204 4452
rect 245420 3724 245476 3780
rect 243852 3612 243908 3668
rect 237580 3500 237636 3556
rect 245532 3500 245588 3556
rect 236012 3388 236068 3444
rect 243628 3388 243684 3444
rect 234444 2604 234500 2660
rect 236012 2828 236068 2884
rect 232876 2492 232932 2548
rect 234108 2380 234164 2436
rect 237916 2716 237972 2772
rect 241724 2604 241780 2660
rect 239820 2492 239876 2548
rect 246988 3388 247044 3444
rect 247436 4396 247492 4452
rect 248556 2716 248612 2772
rect 249340 4508 249396 4564
rect 250124 2492 250180 2548
rect 251244 4620 251300 4676
rect 251692 2380 251748 2436
rect 253148 3612 253204 3668
rect 253260 3276 253316 3332
rect 254828 3164 254884 3220
rect 255052 3724 255108 3780
rect 256396 3052 256452 3108
rect 257068 3388 257124 3444
rect 259532 2940 259588 2996
rect 257964 2604 258020 2660
rect 258860 2716 258916 2772
rect 260764 2492 260820 2548
rect 262668 2828 262724 2884
rect 264236 2716 264292 2772
rect 264572 3276 264628 3332
rect 261100 2492 261156 2548
rect 262668 2380 262724 2436
rect 265804 2268 265860 2324
rect 266476 3164 266532 3220
rect 268940 3276 268996 3332
rect 267372 2380 267428 2436
rect 268380 3052 268436 3108
rect 270284 2604 270340 2660
rect 272076 3164 272132 3220
rect 273644 3052 273700 3108
rect 270508 2604 270564 2660
rect 272188 2940 272244 2996
rect 274092 2492 274148 2548
rect 276780 2940 276836 2996
rect 275212 2492 275268 2548
rect 275996 2828 276052 2884
rect 278348 2828 278404 2884
rect 277900 2716 277956 2772
rect 284620 4844 284676 4900
rect 283052 4732 283108 4788
rect 281484 3948 281540 4004
rect 279916 2716 279972 2772
rect 283612 3276 283668 3332
rect 281708 2380 281764 2436
rect 279804 2268 279860 2324
rect 285628 2604 285684 2660
rect 290892 4284 290948 4340
rect 289324 4172 289380 4228
rect 287756 4060 287812 4116
rect 286188 2604 286244 2660
rect 287420 3164 287476 3220
rect 289324 3052 289380 3108
rect 291228 2492 291284 2548
rect 294700 4956 294756 5012
rect 298732 4620 298788 4676
rect 297164 4508 297220 4564
rect 295596 4396 295652 4452
rect 298844 3948 298900 4004
rect 292460 2492 292516 2548
rect 293132 2940 293188 2996
rect 295036 2828 295092 2884
rect 296940 2716 296996 2772
rect 300300 3164 300356 3220
rect 300748 4732 300804 4788
rect 301868 4732 301924 4788
rect 302652 4844 302708 4900
rect 305004 4844 305060 4900
rect 303436 3052 303492 3108
rect 306460 4060 306516 4116
rect 304556 2604 304612 2660
rect 306572 2940 306628 2996
rect 308140 2604 308196 2660
rect 308364 4172 308420 4228
rect 309708 2828 309764 2884
rect 310268 4284 310324 4340
rect 311276 2716 311332 2772
rect 312172 2492 312228 2548
rect 312844 2492 312900 2548
rect 314188 4956 314244 5012
rect 316652 4956 316708 5012
rect 314412 3948 314468 4004
rect 315980 4396 316036 4452
rect 317548 4060 317604 4116
rect 317884 4508 317940 4564
rect 319116 4172 319172 4228
rect 319788 4620 319844 4676
rect 322252 4396 322308 4452
rect 323596 4732 323652 4788
rect 320684 4284 320740 4340
rect 321692 3164 321748 3220
rect 323820 3276 323876 3332
rect 326956 4508 327012 4564
rect 327404 4844 327460 4900
rect 325388 3164 325444 3220
rect 325500 3052 325556 3108
rect 328524 4620 328580 4676
rect 330092 3052 330148 3108
rect 329308 2940 329364 2996
rect 331212 2604 331268 2660
rect 333228 5068 333284 5124
rect 337932 4844 337988 4900
rect 336364 4732 336420 4788
rect 334796 2940 334852 2996
rect 338828 3948 338884 4004
rect 331660 2604 331716 2660
rect 333116 2828 333172 2884
rect 335020 2716 335076 2772
rect 336924 2492 336980 2548
rect 339500 2828 339556 2884
rect 340732 4956 340788 5012
rect 341740 4956 341796 5012
rect 342524 476 342580 532
rect 342748 4060 342804 4116
rect 344204 2492 344260 2548
rect 344540 4172 344596 4228
rect 345772 2268 345828 2324
rect 346444 4284 346500 4340
rect 348348 4396 348404 4452
rect 347788 700 347844 756
rect 351036 3836 351092 3892
rect 348908 2716 348964 2772
rect 350252 3276 350308 3332
rect 354060 4508 354116 4564
rect 352044 812 352100 868
rect 352156 3164 352212 3220
rect 355180 3164 355236 3220
rect 355964 4620 356020 4676
rect 356748 476 356804 532
rect 357868 3052 357924 3108
rect 358316 2380 358372 2436
rect 359548 3500 359604 3556
rect 359884 3276 359940 3332
rect 359548 2268 359604 2324
rect 359772 2604 359828 2660
rect 361452 1820 361508 1876
rect 361676 5068 361732 5124
rect 363020 2604 363076 2660
rect 363580 2940 363636 2996
rect 367724 5068 367780 5124
rect 364588 2156 364644 2212
rect 365484 4732 365540 4788
rect 364476 1820 364532 1876
rect 364476 588 364532 644
rect 367388 4844 367444 4900
rect 366156 3612 366212 3668
rect 366156 3276 366212 3332
rect 369292 2828 369348 2884
rect 369516 2268 369572 2324
rect 366380 364 366436 420
rect 371308 4956 371364 5012
rect 373996 3276 374052 3332
rect 372428 3164 372484 3220
rect 375004 2492 375060 2548
rect 370860 252 370916 308
rect 372988 140 373044 196
rect 376908 3500 376964 3556
rect 377916 3500 377972 3556
rect 377916 3276 377972 3332
rect 378700 2940 378756 2996
rect 377132 2492 377188 2548
rect 378812 700 378868 756
rect 376236 140 376292 196
rect 382620 3836 382676 3892
rect 381388 3724 381444 3780
rect 381388 3164 381444 3220
rect 380716 2716 380772 2772
rect 383404 3276 383460 3332
rect 386540 3052 386596 3108
rect 384972 1484 385028 1540
rect 384524 812 384580 868
rect 387996 3836 388052 3892
rect 387996 3276 388052 3332
rect 389564 3948 389620 4004
rect 388108 1932 388164 1988
rect 388332 3388 388388 3444
rect 380044 28 380100 84
rect 389676 2716 389732 2772
rect 389564 2156 389620 2212
rect 393036 4956 393092 5012
rect 394044 3612 394100 3668
rect 391244 2156 391300 2212
rect 392140 2380 392196 2436
rect 390124 476 390180 532
rect 397516 2044 397572 2100
rect 397852 2604 397908 2660
rect 394380 1596 394436 1652
rect 395948 588 396004 644
rect 401436 4060 401492 4116
rect 399084 700 399140 756
rect 399868 3948 399924 4004
rect 401436 2940 401492 2996
rect 403116 5068 403172 5124
rect 402220 2828 402276 2884
rect 401660 588 401716 644
rect 407596 3612 407652 3668
rect 405356 2940 405412 2996
rect 403788 812 403844 868
rect 405468 2268 405524 2324
rect 408492 588 408548 644
rect 409276 3724 409332 3780
rect 411516 4172 411572 4228
rect 410060 3164 410116 3220
rect 411180 3500 411236 3556
rect 412300 3948 412356 4004
rect 411516 2716 411572 2772
rect 414764 2716 414820 2772
rect 413196 1148 413252 1204
rect 414988 2492 415044 2548
rect 416892 4060 416948 4116
rect 416332 2156 416388 2212
rect 416668 3724 416724 3780
rect 416668 1932 416724 1988
rect 420364 5068 420420 5124
rect 407260 252 407316 308
rect 417900 476 417956 532
rect 412972 140 413028 196
rect 418684 28 418740 84
rect 421036 2268 421092 2324
rect 422604 3836 422660 3892
rect 425740 4844 425796 4900
rect 424172 2604 424228 2660
rect 426412 3052 426468 3108
rect 423276 1372 423332 1428
rect 424508 1484 424564 1540
rect 430220 4172 430276 4228
rect 428428 3836 428484 3892
rect 428428 2044 428484 2100
rect 428540 3724 428596 3780
rect 427308 364 427364 420
rect 434252 5068 434308 5124
rect 430444 1932 430500 1988
rect 432124 2380 432180 2436
rect 434364 4956 434420 5012
rect 435820 3724 435876 3780
rect 435036 3388 435092 3444
rect 435036 2828 435092 2884
rect 436716 1820 436772 1876
rect 433020 252 433076 308
rect 435932 1596 435988 1652
rect 483084 5516 483140 5572
rect 443548 5404 443604 5460
rect 438284 2492 438340 2548
rect 439740 3836 439796 3892
rect 440188 3500 440244 3556
rect 442988 5068 443044 5124
rect 441420 3052 441476 3108
rect 440188 2940 440244 2996
rect 439852 2828 439908 2884
rect 441644 700 441700 756
rect 462476 5404 462532 5460
rect 444556 4284 444612 4340
rect 445452 3388 445508 3444
rect 447692 3276 447748 3332
rect 450268 3612 450324 3668
rect 449260 1820 449316 1876
rect 449372 3500 449428 3556
rect 446124 700 446180 756
rect 447356 812 447412 868
rect 450268 2156 450324 2212
rect 450828 812 450884 868
rect 451164 3500 451220 3556
rect 454636 4956 454692 5012
rect 452396 3164 452452 3220
rect 454972 3388 455028 3444
rect 453068 588 453124 644
rect 456988 3948 457044 4004
rect 456876 3500 456932 3556
rect 456876 2268 456932 2324
rect 455532 1260 455588 1316
rect 457100 2940 457156 2996
rect 458668 2156 458724 2212
rect 460236 1484 460292 1540
rect 460684 2716 460740 2772
rect 458780 924 458836 980
rect 465724 5292 465780 5348
rect 463372 4396 463428 4452
rect 462476 3164 462532 3220
rect 462588 3612 462644 3668
rect 461804 2044 461860 2100
rect 464940 588 464996 644
rect 464380 476 464436 532
rect 474348 5292 474404 5348
rect 478156 5180 478212 5236
rect 468076 4508 468132 4564
rect 466508 3164 466564 3220
rect 468300 3500 468356 3556
rect 471212 3276 471268 3332
rect 471996 3388 472052 3444
rect 471996 1932 472052 1988
rect 472108 2604 472164 2660
rect 469644 476 469700 532
rect 470204 1372 470260 1428
rect 472780 2380 472836 2436
rect 474012 4844 474068 4900
rect 477484 4620 477540 4676
rect 475916 2604 475972 2660
rect 475804 364 475860 420
rect 480396 3612 480452 3668
rect 479724 3388 479780 3444
rect 480396 2828 480452 2884
rect 480620 2268 480676 2324
rect 482188 1932 482244 1988
rect 482860 5068 482916 5124
rect 479052 28 479108 84
rect 481516 252 481572 308
rect 523516 5516 523572 5572
rect 506380 5404 506436 5460
rect 493164 5180 493220 5236
rect 483084 3164 483140 3220
rect 486892 4732 486948 4788
rect 485324 3052 485380 3108
rect 485548 3724 485604 3780
rect 483756 1148 483812 1204
rect 487228 140 487284 196
rect 490028 2940 490084 2996
rect 491148 3612 491204 3668
rect 489244 2492 489300 2548
rect 495404 5068 495460 5124
rect 496300 4844 496356 4900
rect 496860 4284 496916 4340
rect 491596 2828 491652 2884
rect 492156 3500 492212 3556
rect 492156 1820 492212 1876
rect 493052 3388 493108 3444
rect 494956 3388 495012 3444
rect 499436 3276 499492 3332
rect 500668 3388 500724 3444
rect 497868 1596 497924 1652
rect 498764 700 498820 756
rect 501004 3276 501060 3332
rect 502572 3500 502628 3556
rect 488460 140 488516 196
rect 503804 3724 503860 3780
rect 503804 2156 503860 2212
rect 503916 3388 503972 3444
rect 504140 2492 504196 2548
rect 505708 2492 505764 2548
rect 503916 1260 503972 1316
rect 504476 812 504532 868
rect 507276 5068 507332 5124
rect 508284 4956 508340 5012
rect 507276 2604 507332 2660
rect 507276 924 507332 980
rect 508844 2716 508900 2772
rect 510188 3388 510244 3444
rect 509068 2268 509124 2324
rect 509068 812 509124 868
rect 512428 3612 512484 3668
rect 510412 2604 510468 2660
rect 510524 3388 510580 3444
rect 515676 4956 515732 5012
rect 519708 4396 519764 4452
rect 513548 2492 513604 2548
rect 514108 3724 514164 3780
rect 510524 1484 510580 1540
rect 512092 700 512148 756
rect 515900 3388 515956 3444
rect 517804 2044 517860 2100
rect 521612 588 521668 644
rect 533036 5292 533092 5348
rect 525420 4508 525476 4564
rect 524188 3500 524244 3556
rect 524188 2380 524244 2436
rect 531132 3500 531188 3556
rect 529228 3388 529284 3444
rect 503468 28 503524 84
rect 527212 476 527268 532
rect 555884 5180 555940 5236
rect 548268 4732 548324 4788
rect 536844 4620 536900 4676
rect 534940 812 534996 868
rect 546364 3052 546420 3108
rect 542556 1708 542612 1764
rect 540652 700 540708 756
rect 538748 588 538804 644
rect 552076 2940 552132 2996
rect 553980 2828 554036 2884
rect 573020 5068 573076 5124
rect 559692 4844 559748 4900
rect 557788 3388 557844 3444
rect 565404 3388 565460 3444
rect 563500 1708 563556 1764
rect 561596 1596 561652 1652
rect 569212 588 569268 644
rect 571228 588 571284 644
rect 584444 4956 584500 5012
rect 580636 3612 580692 3668
rect 574924 2716 574980 2772
rect 576828 2604 576884 2660
rect 582540 2492 582596 2548
rect 544348 252 544404 308
rect 550060 140 550116 196
rect 567196 28 567252 84
<< metal3 >>
rect 99474 590940 99484 590996
rect 99540 590940 111692 590996
rect 111748 590940 111758 590996
rect 77410 590828 77420 590884
rect 77476 590828 118412 590884
rect 118468 590828 118478 590884
rect 165666 590828 165676 590884
rect 165732 590828 200732 590884
rect 200788 590828 200798 590884
rect 11218 590716 11228 590772
rect 11284 590716 120092 590772
rect 120148 590716 120158 590772
rect 121538 590716 121548 590772
rect 121604 590716 199948 590772
rect 200004 590716 200014 590772
rect 322914 590716 322924 590772
rect 322980 590716 364028 590772
rect 364084 590716 364094 590772
rect 106642 590604 106652 590660
rect 106708 590604 518476 590660
rect 518532 590604 518542 590660
rect 52882 590492 52892 590548
rect 52948 590492 562604 590548
rect 562660 590492 562670 590548
rect 494722 590156 494732 590212
rect 494788 590156 496412 590212
rect 496468 590156 496478 590212
rect 584658 590156 584668 590212
rect 584724 590156 584762 590212
rect 243618 589596 243628 589652
rect 243684 589596 253708 589652
rect 253764 589596 253774 589652
rect 115042 588812 115052 588868
rect 115108 588812 408268 588868
rect 408324 588812 408334 588868
rect 595560 588644 597000 588840
rect 590482 588588 590492 588644
rect 590548 588616 597000 588644
rect 590548 588588 595672 588616
rect -960 587188 480 587384
rect -960 587160 199836 587188
rect 392 587132 199836 587160
rect 199892 587132 199902 587188
rect 595560 575428 597000 575624
rect 54562 575372 54572 575428
rect 54628 575400 597000 575428
rect 54628 575372 595672 575400
rect -960 573076 480 573272
rect -960 573048 120204 573076
rect 392 573020 120204 573048
rect 120260 573020 120270 573076
rect 595560 562212 597000 562408
rect 590594 562156 590604 562212
rect 590660 562184 597000 562212
rect 590660 562156 595672 562184
rect -960 558964 480 559160
rect -960 558936 111804 558964
rect 392 558908 111804 558936
rect 111860 558908 111870 558964
rect 595560 548996 597000 549192
rect 59602 548940 59612 548996
rect 59668 548968 597000 548996
rect 59668 548940 595672 548968
rect -960 544852 480 545048
rect -960 544824 108332 544852
rect 392 544796 108332 544824
rect 108388 544796 108398 544852
rect 595560 535780 597000 535976
rect 59826 535724 59836 535780
rect 59892 535752 597000 535780
rect 59892 535724 595672 535752
rect -960 530740 480 530936
rect -960 530712 2492 530740
rect 392 530684 2492 530712
rect 2548 530684 2558 530740
rect 54450 523292 54460 523348
rect 54516 523292 590604 523348
rect 590660 523292 590670 523348
rect 595560 522564 597000 522760
rect 60610 522508 60620 522564
rect 60676 522536 597000 522564
rect 60676 522508 595672 522536
rect -960 516628 480 516824
rect -960 516600 532 516628
rect 392 516572 532 516600
rect 476 516516 532 516572
rect 18 516460 28 516516
rect 84 516460 532 516516
rect 55122 511532 55132 511588
rect 55188 511532 200060 511588
rect 200116 511532 200126 511588
rect 595560 509348 597000 509544
rect 54562 509292 54572 509348
rect 54628 509320 597000 509348
rect 54628 509292 595672 509320
rect -960 502516 480 502712
rect -960 502488 113372 502516
rect 392 502460 113372 502488
rect 113428 502460 113438 502516
rect 595560 496132 597000 496328
rect 49522 496076 49532 496132
rect 49588 496104 597000 496132
rect 49588 496076 595672 496104
rect -960 488404 480 488600
rect -960 488376 4172 488404
rect 392 488348 4172 488376
rect 4228 488348 4238 488404
rect 59602 482972 59612 483028
rect 59668 482972 590492 483028
rect 590548 482972 590558 483028
rect 595560 482916 597000 483112
rect 62962 482860 62972 482916
rect 63028 482888 597000 482916
rect 63028 482860 595672 482888
rect -960 474292 480 474488
rect -960 474264 114268 474292
rect 392 474236 114268 474264
rect 114324 474236 114334 474292
rect 595560 469700 597000 469896
rect 1474 469644 1484 469700
rect 1540 469672 597000 469700
rect 1540 469644 595672 469672
rect -960 460180 480 460376
rect -960 460152 111692 460180
rect 392 460124 111692 460152
rect 111748 460124 111758 460180
rect 595560 456484 597000 456680
rect 60610 456428 60620 456484
rect 60676 456456 597000 456484
rect 60676 456428 595672 456456
rect -960 446068 480 446264
rect -960 446040 4396 446068
rect 392 446012 4396 446040
rect 4452 446012 4462 446068
rect 595560 443268 597000 443464
rect 590146 443212 590156 443268
rect 590212 443240 597000 443268
rect 590212 443212 595672 443240
rect 60498 437612 60508 437668
rect 60564 437612 590156 437668
rect 590212 437612 590222 437668
rect -960 431956 480 432152
rect -960 431928 110012 431956
rect 392 431900 110012 431928
rect 110068 431900 110078 431956
rect 595560 430164 597000 430248
rect 57922 430108 57932 430164
rect 57988 430108 597000 430164
rect 595560 430024 597000 430108
rect -960 417844 480 418040
rect -960 417816 118524 417844
rect 392 417788 118524 417816
rect 118580 417788 118590 417844
rect 595560 416836 597000 417032
rect 54674 416780 54684 416836
rect 54740 416808 597000 416836
rect 54740 416780 595672 416808
rect -960 403732 480 403928
rect -960 403704 532 403732
rect 392 403676 532 403704
rect 476 403620 532 403676
rect 595560 403620 597000 403816
rect 130 403564 140 403620
rect 196 403564 532 403620
rect 3154 403564 3164 403620
rect 3220 403592 597000 403620
rect 3220 403564 595672 403592
rect 200722 390684 200732 390740
rect 200788 390684 362572 390740
rect 362628 390684 362638 390740
rect 33058 390572 33068 390628
rect 33124 390572 203420 390628
rect 203476 390572 203486 390628
rect 595560 390404 597000 390600
rect 513202 390348 513212 390404
rect 513268 390376 597000 390404
rect 513268 390348 595672 390376
rect -960 389620 480 389816
rect -960 389592 111804 389620
rect 392 389564 111804 389592
rect 111860 389564 111870 389620
rect 113698 385532 113708 385588
rect 113764 385532 430220 385588
rect 430276 385532 430286 385588
rect 88946 383852 88956 383908
rect 89012 383852 494732 383908
rect 494788 383852 494798 383908
rect 143378 380492 143388 380548
rect 143444 380492 309708 380548
rect 309764 380492 309774 380548
rect 59826 378812 59836 378868
rect 59892 378812 540540 378868
rect 540596 378812 540606 378868
rect 595560 377188 597000 377384
rect 511522 377132 511532 377188
rect 511588 377160 597000 377188
rect 511588 377132 595672 377160
rect 174178 376348 174188 376404
rect 174244 376348 210364 376404
rect 210420 376348 210430 376404
rect -960 375508 480 375704
rect -960 375480 110012 375508
rect 392 375452 110012 375480
rect 110068 375452 110078 375508
rect 110226 375452 110236 375508
rect 110292 375452 474348 375508
rect 474404 375452 474414 375508
rect 167458 374892 167468 374948
rect 167524 374892 199948 374948
rect 200004 374892 200014 374948
rect 113474 374780 113484 374836
rect 113540 374780 174860 374836
rect 174916 374780 174926 374836
rect 125122 374668 125132 374724
rect 125188 374668 387212 374724
rect 387268 374668 387278 374724
rect 187506 373772 187516 373828
rect 187572 373772 256844 373828
rect 256900 373772 256910 373828
rect 1586 373660 1596 373716
rect 1652 373660 202076 373716
rect 202132 373660 202142 373716
rect 176866 373548 176876 373604
rect 176932 373548 200620 373604
rect 200676 373548 200686 373604
rect 180898 373436 180908 373492
rect 180964 373436 208684 373492
rect 208740 373436 208750 373492
rect 179554 373324 179564 373380
rect 179620 373324 212156 373380
rect 212212 373324 212222 373380
rect 25218 373212 25228 373268
rect 25284 373212 168812 373268
rect 168868 373212 168878 373268
rect 177538 373212 177548 373268
rect 177604 373212 211932 373268
rect 211988 373212 211998 373268
rect 54674 373100 54684 373156
rect 54740 373100 201964 373156
rect 202020 373100 202030 373156
rect 181570 372988 181580 373044
rect 181636 372988 207452 373044
rect 207508 372988 207518 373044
rect 115826 372204 115836 372260
rect 115892 372204 176204 372260
rect 176260 372204 176270 372260
rect 93650 372092 93660 372148
rect 93716 372092 452284 372148
rect 452340 372092 452350 372148
rect 149314 371980 149324 372036
rect 149380 371980 209132 372036
rect 209188 371980 209198 372036
rect 169698 371868 169708 371924
rect 169764 371868 208348 371924
rect 208404 371868 208414 371924
rect 171490 371756 171500 371812
rect 171556 371756 197708 371812
rect 197764 371756 197774 371812
rect 147970 371644 147980 371700
rect 148036 371644 211708 371700
rect 211764 371644 211774 371700
rect 133858 371532 133868 371588
rect 133924 371532 200844 371588
rect 200900 371532 200910 371588
rect 139234 371420 139244 371476
rect 139300 371420 210252 371476
rect 210308 371420 210318 371476
rect 27906 371308 27916 371364
rect 27972 371308 169708 371364
rect 169764 371308 169774 371364
rect 175522 371308 175532 371364
rect 175588 371308 199276 371364
rect 199332 371308 199342 371364
rect 141922 370300 141932 370356
rect 141988 370300 210140 370356
rect 210196 370300 210206 370356
rect 178210 370188 178220 370244
rect 178276 370188 196588 370244
rect 196644 370188 196654 370244
rect 170818 370076 170828 370132
rect 170884 370076 194908 370132
rect 194964 370076 194974 370132
rect 115714 369964 115724 370020
rect 115780 369964 162092 370020
rect 162148 369964 162158 370020
rect 168130 369964 168140 370020
rect 168196 369964 203308 370020
rect 203364 369964 203374 370020
rect 110786 369852 110796 369908
rect 110852 369852 160076 369908
rect 160132 369852 160142 369908
rect 169474 369852 169484 369908
rect 169540 369852 204988 369908
rect 205044 369852 205054 369908
rect 143938 369740 143948 369796
rect 144004 369740 207900 369796
rect 207956 369740 207966 369796
rect 184258 369628 184268 369684
rect 184324 369628 205884 369684
rect 205940 369628 205950 369684
rect 2482 368844 2492 368900
rect 2548 368844 201628 368900
rect 201684 368844 201694 368900
rect 149986 368732 149996 368788
rect 150052 368732 205996 368788
rect 206052 368732 206062 368788
rect 115602 368620 115612 368676
rect 115668 368620 159404 368676
rect 159460 368620 159470 368676
rect 166786 368620 166796 368676
rect 166852 368620 199500 368676
rect 199556 368620 199566 368676
rect 144610 368508 144620 368564
rect 144676 368508 207788 368564
rect 207844 368508 207854 368564
rect 137218 368396 137228 368452
rect 137284 368396 206220 368452
rect 206276 368396 206286 368452
rect 131170 368284 131180 368340
rect 131236 368284 200732 368340
rect 200788 368284 200798 368340
rect 135874 368172 135884 368228
rect 135940 368172 210028 368228
rect 210084 368172 210094 368228
rect 23202 368060 23212 368116
rect 23268 368060 169484 368116
rect 169540 368060 169550 368116
rect 183586 368060 183596 368116
rect 183652 368060 204092 368116
rect 204148 368060 204158 368116
rect 188962 367948 188972 368004
rect 189028 367948 213388 368004
rect 213444 367948 213454 368004
rect 126466 367164 126476 367220
rect 126532 367164 210140 367220
rect 210196 367164 210206 367220
rect 138562 367052 138572 367108
rect 138628 367052 209244 367108
rect 209300 367052 209310 367108
rect 117506 366940 117516 366996
rect 117572 366940 165452 366996
rect 165508 366940 165518 366996
rect 172162 366940 172172 366996
rect 172228 366940 200060 366996
rect 200116 366940 200126 366996
rect 152674 366828 152684 366884
rect 152740 366828 204204 366884
rect 204260 366828 204270 366884
rect 146626 366716 146636 366772
rect 146692 366716 207676 366772
rect 207732 366716 207742 366772
rect 147298 366604 147308 366660
rect 147364 366604 210028 366660
rect 210084 366604 210094 366660
rect 139906 366492 139916 366548
rect 139972 366492 206108 366548
rect 206164 366492 206174 366548
rect 119186 366380 119196 366436
rect 119252 366380 162764 366436
rect 162820 366380 162830 366436
rect 180226 366380 180236 366436
rect 180292 366380 195020 366436
rect 195076 366380 195086 366436
rect 186274 366268 186284 366324
rect 186340 366268 208460 366324
rect 208516 366268 208526 366324
rect 112466 365484 112476 365540
rect 112532 365484 201740 365540
rect 201796 365484 201806 365540
rect 154018 365372 154028 365428
rect 154084 365372 209692 365428
rect 209748 365372 209758 365428
rect 156706 365260 156716 365316
rect 156772 365260 209244 365316
rect 209300 365260 209310 365316
rect 155362 365148 155372 365204
rect 155428 365148 209468 365204
rect 209524 365148 209534 365204
rect 132514 365036 132524 365092
rect 132580 365036 200956 365092
rect 201012 365036 201022 365092
rect 140578 364924 140588 364980
rect 140644 364924 209916 364980
rect 209972 364924 209982 364980
rect 86482 364812 86492 364868
rect 86548 364812 125132 364868
rect 125188 364812 125198 364868
rect 137890 364812 137900 364868
rect 137956 364812 213500 364868
rect 213556 364812 213566 364868
rect 115490 364700 115500 364756
rect 115556 364700 158732 364756
rect 158788 364700 158798 364756
rect 185602 364700 185612 364756
rect 185668 364700 205772 364756
rect 205828 364700 205838 364756
rect 2930 364588 2940 364644
rect 2996 364588 166124 364644
rect 166180 364588 166190 364644
rect 178882 364588 178892 364644
rect 178948 364588 199724 364644
rect 199780 364588 199790 364644
rect 595560 363972 597000 364168
rect 143266 363916 143276 363972
rect 143332 363916 211708 363972
rect 211764 363916 211774 363972
rect 590482 363916 590492 363972
rect 590548 363944 597000 363972
rect 590548 363916 595672 363944
rect 5618 363692 5628 363748
rect 5684 363692 171276 363748
rect 171332 363692 172844 363748
rect 172900 363692 172910 363748
rect 4498 363580 4508 363636
rect 4564 363580 201852 363636
rect 201908 363580 201918 363636
rect 154690 363468 154700 363524
rect 154756 363468 204316 363524
rect 204372 363468 204382 363524
rect 114146 363356 114156 363412
rect 114212 363356 164108 363412
rect 164164 363356 164174 363412
rect 187618 363356 187628 363412
rect 187684 363356 196700 363412
rect 196756 363356 196766 363412
rect 145954 363244 145964 363300
rect 146020 363244 202412 363300
rect 202468 363244 202478 363300
rect 127810 363132 127820 363188
rect 127876 363132 143612 363188
rect 143668 363132 143678 363188
rect 145282 363132 145292 363188
rect 145348 363132 202636 363188
rect 202692 363132 202702 363188
rect 129154 363020 129164 363076
rect 129220 363020 151228 363076
rect 151284 363020 151294 363076
rect 160710 363020 160748 363076
rect 160804 363020 160814 363076
rect 164630 363020 164668 363076
rect 164724 363020 164734 363076
rect 182914 363020 182924 363076
rect 182980 363020 194572 363076
rect 194628 363020 194638 363076
rect 151302 362908 151340 362964
rect 151396 362908 151406 362964
rect 151974 362908 152012 362964
rect 152068 362908 152078 362964
rect 156118 362908 156156 362964
rect 156212 362908 156222 362964
rect 157798 362908 157836 362964
rect 157892 362908 157902 362964
rect 188290 362908 188300 362964
rect 188356 362908 199612 362964
rect 199668 362908 199678 362964
rect 149492 362236 158116 362292
rect 149492 362180 149548 362236
rect 158060 362180 158116 362236
rect 110674 362124 110684 362180
rect 110740 362124 149548 362180
rect 153346 362124 153356 362180
rect 153412 362124 155708 362180
rect 155764 362124 155774 362180
rect 158050 362124 158060 362180
rect 158116 362124 158126 362180
rect 163398 362124 163436 362180
rect 163492 362124 163502 362180
rect 168802 362124 168812 362180
rect 168868 362124 193340 362180
rect 193396 362124 193406 362180
rect 199938 362124 199948 362180
rect 200004 362124 200284 362180
rect 200340 362124 200350 362180
rect 143602 362012 143612 362068
rect 143668 362012 207340 362068
rect 207396 362012 207406 362068
rect 142594 361900 142604 361956
rect 142660 361900 155372 361956
rect 155428 361900 155438 361956
rect 155698 361900 155708 361956
rect 155764 361900 205996 361956
rect 206052 361900 206062 361956
rect 148642 361788 148652 361844
rect 148708 361788 207564 361844
rect 207620 361788 207630 361844
rect 136546 361676 136556 361732
rect 136612 361676 204316 361732
rect 204372 361676 204382 361732
rect -960 361396 480 361592
rect 150630 361564 150668 361620
rect 150724 361564 150734 361620
rect 155362 361564 155372 361620
rect 155428 361564 211820 361620
rect 211876 361564 211886 361620
rect 128482 361452 128492 361508
rect 128548 361452 201180 361508
rect 201236 361452 201246 361508
rect -960 361368 118636 361396
rect 392 361340 118636 361368
rect 118692 361340 118702 361396
rect 127138 361340 127148 361396
rect 127204 361340 210252 361396
rect 210308 361340 210318 361396
rect 57026 361228 57036 361284
rect 57092 361228 125804 361284
rect 125860 361228 377132 361284
rect 377188 361228 377198 361284
rect 161382 361116 161420 361172
rect 161476 361116 161486 361172
rect 184940 360668 191548 360724
rect 192546 360668 192556 360724
rect 192612 360668 201124 360724
rect 184940 360612 184996 360668
rect 191492 360612 191548 360668
rect 201068 360612 201124 360668
rect 184930 360556 184940 360612
rect 184996 360556 185006 360612
rect 191492 360556 197372 360612
rect 197428 360556 197438 360612
rect 201058 360556 201068 360612
rect 201124 360556 201134 360612
rect 141250 360444 141260 360500
rect 141316 360444 204428 360500
rect 204484 360444 204494 360500
rect 151218 360332 151228 360388
rect 151284 360332 207564 360388
rect 207620 360332 207630 360388
rect 209570 360332 209580 360388
rect 209636 360332 296492 360388
rect 296548 360332 296558 360388
rect 134530 360220 134540 360276
rect 134596 360220 204652 360276
rect 204708 360220 204718 360276
rect 129826 360108 129836 360164
rect 129892 360108 192556 360164
rect 192612 360108 192622 360164
rect 192770 360108 192780 360164
rect 192836 360108 194684 360164
rect 194740 360108 194750 360164
rect 132290 359996 132300 360052
rect 132356 359996 204876 360052
rect 204932 359996 204942 360052
rect 133186 359884 133196 359940
rect 133252 359884 206332 359940
rect 206388 359884 206398 359940
rect 135202 359772 135212 359828
rect 135268 359772 209356 359828
rect 209412 359772 209422 359828
rect 130498 359660 130508 359716
rect 130564 359660 206556 359716
rect 206612 359660 206622 359716
rect 3042 359548 3052 359604
rect 3108 359548 161420 359604
rect 161476 359548 161486 359604
rect 166086 359548 166124 359604
rect 166180 359548 166190 359604
rect 173478 359548 173516 359604
rect 173572 359548 173582 359604
rect 190726 359548 190764 359604
rect 190820 359548 190830 359604
rect 190978 359548 190988 359604
rect 191044 359548 191082 359604
rect 192098 359548 192108 359604
rect 192164 359548 192556 359604
rect 192612 359548 192622 359604
rect 194002 359548 194012 359604
rect 194068 359548 194236 359604
rect 194292 359548 194302 359604
rect 195654 359548 195692 359604
rect 195748 359548 195758 359604
rect 197362 359548 197372 359604
rect 197428 359548 204204 359604
rect 204260 359548 204270 359604
rect 182214 359436 182252 359492
rect 182308 359436 182318 359492
rect 186918 359436 186956 359492
rect 187012 359436 187022 359492
rect 189522 359436 189532 359492
rect 189588 359436 189644 359492
rect 189700 359436 189710 359492
rect 192966 359436 193004 359492
rect 193060 359436 193070 359492
rect 194310 359436 194348 359492
rect 194404 359436 194414 359492
rect 78194 359212 78204 359268
rect 78260 359212 120120 359268
rect 200050 358652 200060 358708
rect 200116 358652 200396 358708
rect 200452 358652 200462 358708
rect 63746 358092 63756 358148
rect 63812 358092 120120 358148
rect 199266 357644 199276 357700
rect 199332 357644 199342 357700
rect 199266 357084 199276 357140
rect 199332 357084 199342 357140
rect 115154 356972 115164 357028
rect 115220 356972 120120 357028
rect 199276 356552 199332 357084
rect 297826 356972 297836 357028
rect 297892 356972 336140 357028
rect 336196 356972 336206 357028
rect 199378 355964 199388 356020
rect 199444 355964 199454 356020
rect 117394 355852 117404 355908
rect 117460 355852 120120 355908
rect 199388 355432 199444 355964
rect 58258 354732 58268 354788
rect 58324 354732 120120 354788
rect 199864 354284 202076 354340
rect 202132 354284 202142 354340
rect 58594 353612 58604 353668
rect 58660 353612 120120 353668
rect 199864 353164 201964 353220
rect 202020 353164 202030 353220
rect 117170 352492 117180 352548
rect 117236 352492 120120 352548
rect 199864 352044 201628 352100
rect 201684 352044 201694 352100
rect 91522 351372 91532 351428
rect 91588 351372 120120 351428
rect 199864 350924 202076 350980
rect 202132 350924 202142 350980
rect 595560 350756 597000 350952
rect 540082 350700 540092 350756
rect 540148 350728 597000 350756
rect 540148 350700 595672 350728
rect 116610 350252 116620 350308
rect 116676 350252 120120 350308
rect 199864 349804 201852 349860
rect 201908 349804 201918 349860
rect 76178 349132 76188 349188
rect 76244 349132 120120 349188
rect 199864 348684 202300 348740
rect 202356 348684 202366 348740
rect 61282 348012 61292 348068
rect 61348 348012 120120 348068
rect 199864 347564 200172 347620
rect 200228 347564 200238 347620
rect -960 347284 480 347480
rect -960 347256 118860 347284
rect 392 347228 118860 347256
rect 118916 347228 118926 347284
rect 112578 346892 112588 346948
rect 112644 346892 120120 346948
rect 199864 346444 205100 346500
rect 205156 346444 205166 346500
rect 107426 345772 107436 345828
rect 107492 345772 120120 345828
rect 199864 345324 208572 345380
rect 208628 345324 208638 345380
rect 64642 344652 64652 344708
rect 64708 344652 120120 344708
rect 199864 344204 200620 344260
rect 200676 344204 200686 344260
rect 58482 343532 58492 343588
rect 58548 343532 120120 343588
rect 217186 343532 217196 343588
rect 217252 343532 386092 343588
rect 386148 343532 386158 343588
rect 199864 343084 203420 343140
rect 203476 343084 203486 343140
rect 57810 342412 57820 342468
rect 57876 342412 120120 342468
rect 199864 341964 202188 342020
rect 202244 341964 202254 342020
rect 270050 341852 270060 341908
rect 270116 341852 341964 341908
rect 342020 341852 342030 341908
rect 111906 341292 111916 341348
rect 111972 341292 120120 341348
rect 199864 340844 201740 340900
rect 201796 340844 201806 340900
rect 56578 340284 56588 340340
rect 56644 340284 107436 340340
rect 107492 340284 107502 340340
rect 4610 340172 4620 340228
rect 4676 340172 115612 340228
rect 115668 340172 116732 340228
rect 116788 340172 116798 340228
rect 117058 340172 117068 340228
rect 117124 340172 120120 340228
rect 199864 339724 201964 339780
rect 202020 339724 202030 339780
rect 57922 339388 57932 339444
rect 57988 339388 108668 339444
rect 108724 339388 108734 339444
rect 117506 339276 117516 339332
rect 117572 339276 118636 339332
rect 118692 339276 118702 339332
rect 117058 339052 117068 339108
rect 117124 339052 120120 339108
rect 60050 338828 60060 338884
rect 60116 338828 116620 338884
rect 116676 338828 116686 338884
rect 56802 338716 56812 338772
rect 56868 338716 112588 338772
rect 112644 338716 112654 338772
rect 4722 338604 4732 338660
rect 4788 338604 115500 338660
rect 115556 338604 116844 338660
rect 116900 338604 116910 338660
rect 199864 338604 201852 338660
rect 201908 338604 201918 338660
rect 3266 338492 3276 338548
rect 3332 338492 117516 338548
rect 117572 338492 117582 338548
rect 117282 337932 117292 337988
rect 117348 337932 120120 337988
rect 595560 337540 597000 337736
rect 119186 337484 119196 337540
rect 119252 337484 120204 337540
rect 120260 337484 120270 337540
rect 199864 337484 210364 337540
rect 210420 337484 210430 337540
rect 573682 337484 573692 337540
rect 573748 337512 597000 337540
rect 573748 337484 595672 337512
rect 58706 337260 58716 337316
rect 58772 337260 117180 337316
rect 117236 337260 117246 337316
rect 2818 337148 2828 337204
rect 2884 337148 109116 337204
rect 109172 337148 109182 337204
rect 2706 337036 2716 337092
rect 2772 337036 110684 337092
rect 110740 337036 110750 337092
rect 2594 336924 2604 336980
rect 2660 336924 115724 336980
rect 115780 336924 115790 336980
rect 116508 336924 119196 336980
rect 119252 336924 119262 336980
rect 116508 336868 116564 336924
rect 3154 336812 3164 336868
rect 3220 336812 116564 336868
rect 116722 336812 116732 336868
rect 116788 336812 120120 336868
rect 231634 336812 231644 336868
rect 231700 336812 349356 336868
rect 349412 336812 349422 336868
rect 199266 336364 199276 336420
rect 199332 336364 199342 336420
rect 102452 336140 118804 336196
rect 102452 336084 102508 336140
rect 118748 336084 118804 336140
rect 37986 336028 37996 336084
rect 38052 336028 102508 336084
rect 109106 336028 109116 336084
rect 109172 336028 109900 336084
rect 109956 336028 109966 336084
rect 110674 336028 110684 336084
rect 110740 336028 112252 336084
rect 112308 336028 112318 336084
rect 115714 336028 115724 336084
rect 115780 336028 116956 336084
rect 117012 336028 117022 336084
rect 118738 336028 118748 336084
rect 118804 336028 118814 336084
rect 113586 335692 113596 335748
rect 113652 335692 120120 335748
rect 199864 335244 206892 335300
rect 206948 335244 206958 335300
rect 7522 335132 7532 335188
rect 7588 335132 110796 335188
rect 110852 335132 110862 335188
rect 35970 335020 35980 335076
rect 36036 335020 120316 335076
rect 120372 335020 120382 335076
rect 102386 334908 102396 334964
rect 102452 334908 119980 334964
rect 120036 334908 120046 334964
rect 28578 334796 28588 334852
rect 28644 334796 118748 334852
rect 118804 334796 118814 334852
rect 110786 334572 110796 334628
rect 110852 334572 112364 334628
rect 112420 334572 112430 334628
rect 115266 334572 115276 334628
rect 115332 334572 120120 334628
rect 35298 334460 35308 334516
rect 35364 334460 120540 334516
rect 120596 334460 120606 334516
rect 56914 334348 56924 334404
rect 56980 334348 64652 334404
rect 64708 334348 64718 334404
rect 101042 334348 101052 334404
rect 101108 334348 113820 334404
rect 113876 334348 113886 334404
rect 199864 334124 202076 334180
rect 202132 334124 202142 334180
rect 70354 333788 70364 333844
rect 70420 333788 84924 333844
rect 84980 333788 84990 333844
rect 73490 333676 73500 333732
rect 73556 333676 75796 333732
rect 75740 333620 75796 333676
rect 59714 333564 59724 333620
rect 59780 333564 75516 333620
rect 75572 333564 75582 333620
rect 75740 333564 88284 333620
rect 88340 333564 88350 333620
rect 42690 333452 42700 333508
rect 42756 333452 51212 333508
rect 51268 333452 51278 333508
rect 63522 333452 63532 333508
rect 63588 333452 72828 333508
rect 72884 333452 87612 333508
rect 87668 333452 87678 333508
rect 116946 333452 116956 333508
rect 117012 333452 120120 333508
rect -960 333172 480 333368
rect 38658 333340 38668 333396
rect 38724 333340 51436 333396
rect 51492 333340 51502 333396
rect 55122 333340 55132 333396
rect 55188 333340 74844 333396
rect 74900 333340 74910 333396
rect 31938 333228 31948 333284
rect 32004 333228 115388 333284
rect 115444 333228 115454 333284
rect -960 333144 4284 333172
rect 392 333116 4284 333144
rect 4340 333116 4350 333172
rect 44706 333116 44716 333172
rect 44772 333116 56700 333172
rect 56756 333116 56766 333172
rect 70466 333116 70476 333172
rect 70532 333116 82908 333172
rect 82964 333116 82974 333172
rect 41346 333004 41356 333060
rect 41412 333004 56252 333060
rect 56308 333004 56318 333060
rect 60386 333004 60396 333060
rect 60452 333004 70364 333060
rect 70420 333004 70430 333060
rect 199864 333004 203308 333060
rect 203364 333004 203374 333060
rect 36642 332892 36652 332948
rect 36708 332892 53004 332948
rect 53060 332892 53070 332948
rect 60050 332892 60060 332948
rect 60116 332892 72156 332948
rect 72212 332892 78876 332948
rect 78932 332892 78942 332948
rect 40002 332780 40012 332836
rect 40068 332780 56476 332836
rect 56532 332780 56542 332836
rect 56914 332780 56924 332836
rect 56980 332780 86940 332836
rect 86996 332780 87006 332836
rect 101714 332780 101724 332836
rect 101780 332780 115724 332836
rect 115780 332780 115790 332836
rect 4834 332668 4844 332724
rect 4900 332668 18508 332724
rect 18564 332668 18574 332724
rect 63634 332668 63644 332724
rect 63700 332668 69468 332724
rect 69524 332668 70476 332724
rect 70532 332668 70542 332724
rect 74834 332668 74844 332724
rect 74900 332668 77532 332724
rect 77588 332668 77598 332724
rect 94994 331996 95004 332052
rect 95060 331996 116396 332052
rect 116452 331996 116462 332052
rect 83570 331884 83580 331940
rect 83636 331884 116844 331940
rect 116900 331884 116910 331940
rect 56690 331772 56700 331828
rect 56756 331772 91532 331828
rect 91588 331772 91598 331828
rect 120092 331716 120148 332360
rect 199864 331884 201964 331940
rect 202020 331884 202030 331940
rect 202626 331772 202636 331828
rect 202692 331772 208124 331828
rect 208180 331772 208190 331828
rect 43362 331660 43372 331716
rect 43428 331660 119196 331716
rect 119252 331660 119262 331716
rect 120082 331660 120092 331716
rect 120148 331660 120158 331716
rect 31266 331548 31276 331604
rect 31332 331548 119868 331604
rect 119924 331548 119934 331604
rect 92978 331436 92988 331492
rect 93044 331436 114940 331492
rect 114996 331436 115006 331492
rect 84242 331324 84252 331380
rect 84308 331324 115612 331380
rect 115668 331324 115678 331380
rect 58706 331212 58716 331268
rect 58772 331212 79548 331268
rect 79604 331212 79614 331268
rect 100370 331212 100380 331268
rect 100436 331212 110348 331268
rect 110404 331212 110414 331268
rect 118962 331212 118972 331268
rect 119028 331212 120120 331268
rect 103730 331100 103740 331156
rect 103796 331100 116620 331156
rect 116676 331100 116686 331156
rect 2370 330988 2380 331044
rect 2436 330988 19852 331044
rect 19908 330988 19918 331044
rect 105074 330988 105084 331044
rect 105140 330988 112140 331044
rect 112196 330988 112206 331044
rect 114146 330988 114156 331044
rect 114212 330988 114268 331044
rect 114324 330988 114334 331044
rect 57698 330876 57708 330932
rect 57764 330876 62972 330932
rect 63028 330876 63038 330932
rect 56466 330764 56476 330820
rect 56532 330764 61292 330820
rect 61348 330764 61358 330820
rect 37314 330652 37324 330708
rect 37380 330652 120540 330708
rect 120596 330652 120606 330708
rect 104402 330428 104412 330484
rect 104468 330428 112028 330484
rect 112084 330428 112094 330484
rect 5506 330316 5516 330372
rect 5572 330316 119196 330372
rect 119252 330316 119262 330372
rect 199276 330260 199332 330792
rect 58034 330204 58044 330260
rect 58100 330204 73500 330260
rect 73556 330204 73566 330260
rect 103058 330204 103068 330260
rect 103124 330204 117180 330260
rect 117236 330204 117246 330260
rect 199266 330204 199276 330260
rect 199332 330204 199342 330260
rect 275762 330204 275772 330260
rect 275828 330204 283276 330260
rect 283332 330204 283342 330260
rect 105746 330092 105756 330148
rect 105812 330092 110572 330148
rect 110628 330092 110638 330148
rect 31042 329980 31052 330036
rect 31108 329980 119644 330036
rect 119700 329980 119710 330036
rect 75506 329868 75516 329924
rect 75572 329868 76860 329924
rect 76916 329868 76926 329924
rect 109928 329756 115052 329812
rect 115108 329756 115118 329812
rect 120092 329588 120148 330120
rect 230402 330092 230412 330148
rect 230468 330092 319900 330148
rect 319956 330092 319966 330148
rect 199864 329644 202524 329700
rect 202580 329644 202590 329700
rect 110450 329532 110460 329588
rect 110516 329532 120148 329588
rect 119186 329308 119196 329364
rect 119252 329308 120316 329364
rect 120372 329308 120382 329364
rect 200050 329252 200060 329308
rect 200116 329252 200126 329308
rect 200060 329196 200284 329252
rect 200340 329196 200350 329252
rect 109928 329084 118860 329140
rect 118916 329084 118926 329140
rect 115938 328972 115948 329028
rect 116004 328972 120120 329028
rect 199864 328524 210476 328580
rect 210532 328524 210542 328580
rect 109928 328412 111916 328468
rect 111972 328412 111982 328468
rect 408930 328076 408940 328132
rect 408996 328076 423948 328132
rect 424004 328076 424014 328132
rect 419682 327964 419692 328020
rect 419748 327964 431788 328020
rect 431844 327964 431854 328020
rect 112242 327852 112252 327908
rect 112308 327852 120120 327908
rect 409602 327852 409612 327908
rect 409668 327852 420140 327908
rect 420196 327852 420206 327908
rect 109928 327740 112588 327796
rect 112644 327740 112654 327796
rect 380258 327740 380268 327796
rect 380324 327740 392812 327796
rect 392868 327740 392878 327796
rect 408258 327740 408268 327796
rect 408324 327740 420028 327796
rect 420084 327740 420094 327796
rect 421026 327740 421036 327796
rect 421092 327740 426860 327796
rect 426916 327740 426926 327796
rect 370626 327628 370636 327684
rect 370692 327628 389452 327684
rect 389508 327628 389518 327684
rect 421698 327628 421708 327684
rect 421764 327628 426748 327684
rect 426804 327628 426814 327684
rect 57138 327516 57148 327572
rect 57204 327516 60620 327572
rect 60676 327516 60686 327572
rect 202402 327516 202412 327572
rect 202468 327516 208236 327572
rect 208292 327516 208302 327572
rect 199864 327404 202636 327460
rect 202692 327404 202702 327460
rect 109928 327068 115052 327124
rect 115108 327068 115118 327124
rect 115490 326732 115500 326788
rect 115556 326732 120120 326788
rect 54936 326396 57932 326452
rect 57988 326396 57998 326452
rect 109928 326396 113708 326452
rect 113764 326396 113774 326452
rect 199864 326284 202860 326340
rect 202916 326284 202926 326340
rect 375778 326284 375788 326340
rect 375844 326284 406252 326340
rect 406308 326284 406318 326340
rect 378578 326172 378588 326228
rect 378644 326172 397516 326228
rect 397572 326172 397582 326228
rect 416994 326172 417004 326228
rect 417060 326172 428428 326228
rect 428484 326172 428494 326228
rect 375554 326060 375564 326116
rect 375620 326060 406924 326116
rect 406980 326060 406990 326116
rect 417666 326060 417676 326116
rect 417732 326060 433468 326116
rect 433524 326060 433534 326116
rect 379698 325948 379708 326004
rect 379764 325948 392140 326004
rect 392196 325948 392206 326004
rect 398178 325948 398188 326004
rect 398244 325948 440300 326004
rect 440356 325948 440366 326004
rect 54936 325724 57932 325780
rect 57988 325724 57998 325780
rect 109928 325724 113484 325780
rect 113540 325724 113550 325780
rect 115266 325612 115276 325668
rect 115332 325612 120120 325668
rect 199266 325164 199276 325220
rect 199332 325164 199342 325220
rect 208002 325164 208012 325220
rect 208068 325164 211708 325220
rect 211764 325164 211774 325220
rect 5068 324660 5124 325080
rect 5282 324828 5292 324884
rect 5348 324828 5358 324884
rect 4946 324604 4956 324660
rect 5012 324604 5124 324660
rect 5292 324408 5348 324828
rect 54908 324660 54964 325080
rect 56998 325052 57036 325108
rect 57092 325052 60088 325108
rect 109928 325052 113820 325108
rect 113876 325052 113886 325108
rect 208114 325052 208124 325108
rect 208180 325052 212268 325108
rect 212324 325052 212334 325108
rect 410722 324940 410732 324996
rect 410788 324940 414316 324996
rect 414372 324940 414382 324996
rect 423378 324940 423388 324996
rect 423444 324940 423948 324996
rect 424004 324940 424014 324996
rect 377570 324828 377580 324884
rect 377636 324828 442092 324884
rect 442148 324828 442158 324884
rect 376114 324716 376124 324772
rect 376180 324716 441868 324772
rect 441924 324716 441934 324772
rect 54908 324604 58380 324660
rect 58436 324604 58446 324660
rect 373874 324604 373884 324660
rect 373940 324604 440300 324660
rect 440356 324604 440366 324660
rect 115490 324492 115500 324548
rect 115556 324492 120120 324548
rect 380370 324492 380380 324548
rect 380436 324492 390124 324548
rect 390180 324492 390190 324548
rect 396834 324492 396844 324548
rect 396900 324492 432124 324548
rect 432180 324492 432190 324548
rect 54936 324380 58156 324436
rect 58212 324380 58222 324436
rect 109928 324380 112028 324436
rect 112084 324380 112094 324436
rect 375666 324380 375676 324436
rect 375732 324380 410732 324436
rect 410788 324380 410798 324436
rect 410946 324380 410956 324436
rect 411012 324380 411404 324436
rect 411460 324380 411470 324436
rect 418310 324380 418348 324436
rect 418404 324380 418414 324436
rect 418758 324380 418796 324436
rect 418852 324380 418862 324436
rect 420802 324380 420812 324436
rect 420868 324380 421260 324436
rect 421316 324380 421326 324436
rect 422006 324380 422044 324436
rect 422100 324380 422110 324436
rect 422566 324380 422604 324436
rect 422660 324380 422670 324436
rect 424134 324380 424172 324436
rect 424228 324380 424238 324436
rect 425030 324380 425068 324436
rect 425124 324380 425134 324436
rect 426150 324380 426188 324436
rect 426244 324380 426254 324436
rect 426402 324380 426412 324436
rect 426468 324380 426506 324436
rect 595560 324324 597000 324520
rect 377122 324268 377132 324324
rect 377188 324268 377916 324324
rect 377972 324296 597000 324324
rect 377972 324268 595672 324296
rect 114258 324156 114268 324212
rect 114324 324156 115052 324212
rect 115108 324156 115118 324212
rect 115714 324156 115724 324212
rect 115780 324156 117404 324212
rect 117460 324156 117470 324212
rect 199378 324044 199388 324100
rect 199444 324044 199454 324100
rect 54936 323708 57932 323764
rect 57988 323708 57998 323764
rect 109928 323708 113708 323764
rect 113764 323708 113774 323764
rect 113250 323372 113260 323428
rect 113316 323372 120120 323428
rect 426402 323372 426412 323428
rect 426468 323372 436828 323428
rect 436884 323372 436894 323428
rect 54936 323036 58156 323092
rect 58212 323036 58222 323092
rect 109928 323036 113036 323092
rect 113092 323036 113102 323092
rect 379026 323036 379036 323092
rect 379092 323036 442316 323092
rect 442372 323036 442382 323092
rect 199864 322924 201852 322980
rect 201908 322924 201918 322980
rect 378802 322924 378812 322980
rect 378868 322924 442204 322980
rect 442260 322924 442270 322980
rect 375442 322812 375452 322868
rect 375508 322812 441980 322868
rect 442036 322812 442046 322868
rect 373650 322700 373660 322756
rect 373716 322700 440412 322756
rect 440468 322700 440478 322756
rect 373762 322588 373772 322644
rect 373828 322588 440188 322644
rect 440244 322588 440254 322644
rect 210130 322476 210140 322532
rect 210196 322476 210206 322532
rect 54936 322364 58268 322420
rect 58324 322364 58334 322420
rect 58594 322364 58604 322420
rect 58660 322364 60088 322420
rect 109928 322364 113596 322420
rect 113652 322364 113662 322420
rect 115602 322252 115612 322308
rect 115668 322252 120120 322308
rect 210140 321944 210196 322476
rect 199864 321804 206668 321860
rect 206724 321804 206734 321860
rect 54908 321076 54964 321720
rect 58706 321692 58716 321748
rect 58772 321692 60088 321748
rect 109928 321692 113372 321748
rect 113428 321692 113438 321748
rect 55412 321132 60228 321188
rect 114818 321132 114828 321188
rect 114884 321132 120120 321188
rect 55412 321076 55468 321132
rect 60172 321076 60228 321132
rect 54908 321020 55468 321076
rect 56130 321020 56140 321076
rect 56196 321020 57820 321076
rect 57876 321020 57886 321076
rect 60162 321020 60172 321076
rect 60228 321020 60238 321076
rect 109928 321020 117404 321076
rect 117460 321020 117470 321076
rect 57110 320908 57148 320964
rect 57204 320908 57214 320964
rect 199864 320684 203532 320740
rect 203588 320684 203598 320740
rect 2930 320348 2940 320404
rect 2996 320348 5096 320404
rect 54908 320180 54964 320376
rect 56690 320348 56700 320404
rect 56756 320348 60088 320404
rect 109928 320348 117292 320404
rect 117348 320348 117358 320404
rect 5506 320124 5516 320180
rect 5572 320124 5582 320180
rect 54908 320124 60284 320180
rect 60340 320124 60350 320180
rect 5516 319704 5572 320124
rect 115378 320012 115388 320068
rect 115444 320012 120120 320068
rect 199836 320012 210588 320068
rect 210644 320012 210654 320068
rect 54936 319676 56364 319732
rect 56420 319676 56430 319732
rect 60050 319676 60060 319732
rect 60116 319676 60126 319732
rect 109928 319676 113148 319732
rect 113204 319676 113214 319732
rect 199836 319592 199892 320012
rect 210242 319900 210252 319956
rect 210308 319900 210318 319956
rect 210252 319256 210308 319900
rect -960 319060 480 319256
rect -960 319032 4284 319060
rect 392 319004 4284 319032
rect 4340 319004 4350 319060
rect 54936 319004 59500 319060
rect 59556 319004 59566 319060
rect 109928 319004 116620 319060
rect 116676 319004 116686 319060
rect 115602 318892 115612 318948
rect 115668 318892 120120 318948
rect 373538 318668 373548 318724
rect 373604 318668 380072 318724
rect 5058 318332 5068 318388
rect 5124 318332 5134 318388
rect 109928 318332 117180 318388
rect 117236 318332 117246 318388
rect 199276 317828 199332 318472
rect 369880 318108 373884 318164
rect 373940 318108 373950 318164
rect 114930 317772 114940 317828
rect 114996 317772 120120 317828
rect 199266 317772 199276 317828
rect 199332 317772 199342 317828
rect 2258 317660 2268 317716
rect 2324 317660 5096 317716
rect 109928 317660 115164 317716
rect 115220 317660 115230 317716
rect 58258 317436 58268 317492
rect 58324 317436 60116 317492
rect 112550 317436 112588 317492
rect 112644 317436 112654 317492
rect 60060 317016 60116 317436
rect 199864 317324 202300 317380
rect 202356 317324 202366 317380
rect 372754 317324 372764 317380
rect 372820 317324 380072 317380
rect 109928 316988 115948 317044
rect 116004 316988 116014 317044
rect 369880 316988 375452 317044
rect 375508 316988 375518 317044
rect 115826 316652 115836 316708
rect 115892 316652 120120 316708
rect 376002 316652 376012 316708
rect 376068 316652 380072 316708
rect 207330 316540 207340 316596
rect 207396 316540 210056 316596
rect 56466 316316 56476 316372
rect 56532 316316 60088 316372
rect 109928 316316 113932 316372
rect 113988 316316 113998 316372
rect 199864 316204 200172 316260
rect 200228 316204 200238 316260
rect 377458 315980 377468 316036
rect 377524 315980 380072 316036
rect 369880 315868 377580 315924
rect 377636 315868 377646 315924
rect 3266 315644 3276 315700
rect 3332 315644 5096 315700
rect 109928 315644 115724 315700
rect 115780 315644 115790 315700
rect 117170 315532 117180 315588
rect 117236 315532 120120 315588
rect 376786 315308 376796 315364
rect 376852 315308 380072 315364
rect 199602 315084 199612 315140
rect 199668 315084 199678 315140
rect 3042 314972 3052 315028
rect 3108 314972 5096 315028
rect 54936 314972 60396 315028
rect 60452 314972 60462 315028
rect 109928 314972 117180 315028
rect 117236 314972 117246 315028
rect 369880 314748 373772 314804
rect 373828 314748 373838 314804
rect 377682 314636 377692 314692
rect 377748 314636 380072 314692
rect 117282 314412 117292 314468
rect 117348 314412 120120 314468
rect 54936 314300 58268 314356
rect 58324 314300 58334 314356
rect 58706 314300 58716 314356
rect 58772 314300 60088 314356
rect 109928 314300 115836 314356
rect 115892 314300 115902 314356
rect 58716 314244 58772 314300
rect 56242 314188 56252 314244
rect 56308 314188 58772 314244
rect 116946 313964 116956 314020
rect 117012 313964 120428 314020
rect 120484 313964 120494 314020
rect 199864 313964 202524 314020
rect 202580 313964 202590 314020
rect 374098 313964 374108 314020
rect 374164 313964 380072 314020
rect 201170 313852 201180 313908
rect 201236 313852 210056 313908
rect 4610 313628 4620 313684
rect 4676 313628 5096 313684
rect 54908 313460 54964 313656
rect 56802 313628 56812 313684
rect 56868 313628 60088 313684
rect 369880 313628 379036 313684
rect 379092 313628 379102 313684
rect 54908 313404 55468 313460
rect 55412 313012 55468 313404
rect 116610 313292 116620 313348
rect 116676 313292 120120 313348
rect 2594 312956 2604 313012
rect 2660 312956 5096 313012
rect 55412 312956 60172 313012
rect 60228 312956 60238 313012
rect 199864 312844 200508 312900
rect 200564 312844 200574 312900
rect 439880 312620 443548 312676
rect 443604 312620 443614 312676
rect 114034 312508 114044 312564
rect 114100 312508 115500 312564
rect 115556 312508 115566 312564
rect 369880 312508 373772 312564
rect 373828 312508 373838 312564
rect 3154 312284 3164 312340
rect 3220 312284 5096 312340
rect 54936 312284 56588 312340
rect 56644 312284 56654 312340
rect 113138 312172 113148 312228
rect 113204 312172 120120 312228
rect 439880 311948 441868 312004
rect 441924 311948 441934 312004
rect 199864 311724 206668 311780
rect 206724 311724 206734 311780
rect 4722 311612 4732 311668
rect 4788 311612 5096 311668
rect 54936 311612 60508 311668
rect 60564 311612 60574 311668
rect 369880 311388 378812 311444
rect 378868 311388 378878 311444
rect 439880 311276 445228 311332
rect 445284 311276 445294 311332
rect 207554 311164 207564 311220
rect 207620 311164 210056 311220
rect 595560 311108 597000 311304
rect 113362 311052 113372 311108
rect 113428 311052 120120 311108
rect 543442 311052 543452 311108
rect 543508 311080 597000 311108
rect 543508 311052 595672 311080
rect 3042 310940 3052 310996
rect 3108 310940 5096 310996
rect 54936 310940 58492 310996
rect 58548 310940 58558 310996
rect 114258 310940 114268 310996
rect 114324 310940 114362 310996
rect 202850 310828 202860 310884
rect 202916 310828 206780 310884
rect 206836 310828 206846 310884
rect 112242 310716 112252 310772
rect 112308 310716 116956 310772
rect 117012 310716 117022 310772
rect 199864 310604 200284 310660
rect 200340 310604 200350 310660
rect 377346 310604 377356 310660
rect 377412 310604 380072 310660
rect 439880 310604 441980 310660
rect 442036 310604 442046 310660
rect 2706 310268 2716 310324
rect 2772 310268 5096 310324
rect 54936 310268 58044 310324
rect 58100 310268 58110 310324
rect 369880 310268 375676 310324
rect 375732 310268 375742 310324
rect 115938 309932 115948 309988
rect 116004 309932 120120 309988
rect 439880 309932 440188 309988
rect 440244 309932 440254 309988
rect 4722 309596 4732 309652
rect 4788 309596 5096 309652
rect 54460 309204 54516 309624
rect 199864 309484 200396 309540
rect 200452 309484 200462 309540
rect 439880 309260 442092 309316
rect 442148 309260 442158 309316
rect 54450 309148 54460 309204
rect 54516 309148 54526 309204
rect 57026 309148 57036 309204
rect 57092 309148 58492 309204
rect 58548 309148 58558 309204
rect 369880 309148 375452 309204
rect 375508 309148 375518 309204
rect 110562 309036 110572 309092
rect 110628 309036 117516 309092
rect 117572 309036 117582 309092
rect 1474 308924 1484 308980
rect 1540 308924 5096 308980
rect 54936 308924 58716 308980
rect 58772 308924 58782 308980
rect 116386 308812 116396 308868
rect 116452 308812 120120 308868
rect 5282 308700 5292 308756
rect 5348 308700 5358 308756
rect 5292 308280 5348 308700
rect 371074 308588 371084 308644
rect 371140 308588 380072 308644
rect 439880 308588 445340 308644
rect 445396 308588 445406 308644
rect 201058 308476 201068 308532
rect 201124 308476 210056 308532
rect 112354 308364 112364 308420
rect 112420 308364 118524 308420
rect 118580 308364 118590 308420
rect 199864 308364 201740 308420
rect 201796 308364 201806 308420
rect 54936 308252 58380 308308
rect 58436 308252 58446 308308
rect 369880 308028 373884 308084
rect 373940 308028 373950 308084
rect 439880 307916 442540 307972
rect 442596 307916 442606 307972
rect 116610 307692 116620 307748
rect 116676 307692 120120 307748
rect 3266 307580 3276 307636
rect 3332 307580 5096 307636
rect 54936 307580 57932 307636
rect 57988 307580 57998 307636
rect 112578 307356 112588 307412
rect 112644 307356 115500 307412
rect 115556 307356 115566 307412
rect 199864 307244 200284 307300
rect 200340 307244 200350 307300
rect 439880 307244 441868 307300
rect 441924 307244 441934 307300
rect 4610 306908 4620 306964
rect 4676 306908 5096 306964
rect 369880 306908 373660 306964
rect 373716 306908 373726 306964
rect 117282 306572 117292 306628
rect 117348 306572 120120 306628
rect 439880 306572 443660 306628
rect 443716 306572 443726 306628
rect 2930 306236 2940 306292
rect 2996 306236 5096 306292
rect 109928 306236 114828 306292
rect 114884 306236 114894 306292
rect 199864 306124 205212 306180
rect 205268 306124 205278 306180
rect 439292 305844 439348 305928
rect 206546 305788 206556 305844
rect 206612 305788 210056 305844
rect 369880 305788 375788 305844
rect 375844 305788 375854 305844
rect 439282 305788 439292 305844
rect 439348 305788 439358 305844
rect 2706 305564 2716 305620
rect 2772 305564 5096 305620
rect 54936 305564 57820 305620
rect 57876 305564 57886 305620
rect 115042 305452 115052 305508
rect 115108 305452 120120 305508
rect 439880 305228 440860 305284
rect 440916 305228 440926 305284
rect -960 304948 480 305144
rect 110114 305004 110124 305060
rect 110180 305004 118412 305060
rect 118468 305004 118478 305060
rect 199864 305004 200508 305060
rect 200564 305004 200574 305060
rect -960 304920 532 304948
rect 392 304892 532 304920
rect 2818 304892 2828 304948
rect 2884 304892 5096 304948
rect 54936 304892 57708 304948
rect 57764 304892 57774 304948
rect 109928 304892 110908 304948
rect 110964 304892 113484 304948
rect 113540 304892 113550 304948
rect 476 304836 532 304892
rect 18 304780 28 304836
rect 84 304780 532 304836
rect 54908 304668 57148 304724
rect 57204 304668 57214 304724
rect 369880 304668 375564 304724
rect 375620 304668 375630 304724
rect 54908 304248 54964 304668
rect 439880 304556 442652 304612
rect 442708 304556 442718 304612
rect 115714 304332 115724 304388
rect 115780 304332 120120 304388
rect 56578 304220 56588 304276
rect 56644 304220 60088 304276
rect 5618 303996 5628 304052
rect 5684 303996 5694 304052
rect 5628 303576 5684 303996
rect 199826 303884 199836 303940
rect 199892 303884 199902 303940
rect 439880 303884 442204 303940
rect 442260 303884 442270 303940
rect 54936 303548 58492 303604
rect 58548 303548 58558 303604
rect 109340 303156 109396 303576
rect 369880 303548 375564 303604
rect 375620 303548 375630 303604
rect 118850 303212 118860 303268
rect 118916 303212 120120 303268
rect 376226 303212 376236 303268
rect 376292 303212 377916 303268
rect 377972 303212 380072 303268
rect 439880 303212 441980 303268
rect 442036 303212 442046 303268
rect 109330 303100 109340 303156
rect 109396 303100 109406 303156
rect 200722 303100 200732 303156
rect 200788 303100 210056 303156
rect 54936 302876 56364 302932
rect 56420 302876 56430 302932
rect 57026 302876 57036 302932
rect 57092 302876 60088 302932
rect 109928 302876 115612 302932
rect 115668 302876 115678 302932
rect 199864 302764 208796 302820
rect 208852 302764 208862 302820
rect 439880 302540 441084 302596
rect 441140 302540 441150 302596
rect 369880 302428 377244 302484
rect 377300 302428 377310 302484
rect 54796 302036 54852 302232
rect 56802 302204 56812 302260
rect 56868 302204 60088 302260
rect 112130 302092 112140 302148
rect 112196 302092 120120 302148
rect 54796 301980 59388 302036
rect 59444 301980 59454 302036
rect 376450 301868 376460 301924
rect 376516 301868 380072 301924
rect 439880 301868 440972 301924
rect 441028 301868 441038 301924
rect 199864 301644 202860 301700
rect 202916 301644 202926 301700
rect 54450 301532 54460 301588
rect 54516 301532 54526 301588
rect 56914 301532 56924 301588
rect 56980 301532 60088 301588
rect 369880 301308 380100 301364
rect 199266 301196 199276 301252
rect 199332 301196 199388 301252
rect 199444 301196 199454 301252
rect 380044 301224 380100 301308
rect 439880 301196 440300 301252
rect 440356 301196 440366 301252
rect 110338 300972 110348 301028
rect 110404 300972 120120 301028
rect 54936 300860 59724 300916
rect 59780 300860 59790 300916
rect 109928 300860 110908 300916
rect 110964 300860 115836 300916
rect 115892 300860 115902 300916
rect 202514 300748 202524 300804
rect 202580 300748 206780 300804
rect 206836 300748 206846 300804
rect 113810 300524 113820 300580
rect 113876 300524 115836 300580
rect 115892 300524 115902 300580
rect 199266 300524 199276 300580
rect 199332 300524 199342 300580
rect 204866 300412 204876 300468
rect 204932 300412 210056 300468
rect 54936 300188 56476 300244
rect 56532 300188 56542 300244
rect 109928 300188 113260 300244
rect 113316 300188 113326 300244
rect 369880 300188 376460 300244
rect 376516 300188 376526 300244
rect 380044 300132 380100 300552
rect 439880 300524 442204 300580
rect 442260 300524 442270 300580
rect 372932 300076 380100 300132
rect 111906 299964 111916 300020
rect 111972 299964 120148 300020
rect 120092 299880 120148 299964
rect 199864 299404 202188 299460
rect 202244 299404 202254 299460
rect 372932 299124 372988 300076
rect 377234 299852 377244 299908
rect 377300 299852 380072 299908
rect 439880 299852 440412 299908
rect 440468 299852 440478 299908
rect 373650 299180 373660 299236
rect 373716 299180 380072 299236
rect 439880 299180 442316 299236
rect 442372 299180 442382 299236
rect 112242 299068 112252 299124
rect 112308 299068 112700 299124
rect 112756 299068 112766 299124
rect 200722 299068 200732 299124
rect 200788 299068 201740 299124
rect 201796 299068 201806 299124
rect 369880 299068 372988 299124
rect 117394 298732 117404 298788
rect 117460 298732 120120 298788
rect 373874 298508 373884 298564
rect 373940 298508 380072 298564
rect 439880 298508 442092 298564
rect 442148 298508 442158 298564
rect 199864 298284 202636 298340
rect 202692 298284 202702 298340
rect 57026 298172 57036 298228
rect 57092 298172 60088 298228
rect 109928 298172 117628 298228
rect 117684 298172 117694 298228
rect 369880 297948 375788 298004
rect 375844 297948 375854 298004
rect 595560 297892 597000 298088
rect 439880 297836 442764 297892
rect 442820 297836 442830 297892
rect 590146 297836 590156 297892
rect 590212 297864 597000 297892
rect 590212 297836 595672 297864
rect 200946 297724 200956 297780
rect 201012 297724 210056 297780
rect 112018 297612 112028 297668
rect 112084 297612 120120 297668
rect 3042 297500 3052 297556
rect 3108 297500 5096 297556
rect 56130 297500 56140 297556
rect 56196 297500 60088 297556
rect 109564 297332 109620 297528
rect 109554 297276 109564 297332
rect 109620 297276 109630 297332
rect 119970 297052 119980 297108
rect 120036 297052 120148 297108
rect 120092 296520 120148 297052
rect 199276 296772 199332 297192
rect 439880 297164 440636 297220
rect 440692 297164 440702 297220
rect 202626 297052 202636 297108
rect 202692 297052 210140 297108
rect 210196 297052 210206 297108
rect 369880 296828 372204 296884
rect 372260 296828 372270 296884
rect 199266 296716 199276 296772
rect 199332 296716 199342 296772
rect 439880 296492 440524 296548
rect 440580 296492 440590 296548
rect 563602 296492 563612 296548
rect 563668 296492 590156 296548
rect 590212 296492 590222 296548
rect 199266 296380 199276 296436
rect 199332 296380 199388 296436
rect 199444 296380 199454 296436
rect 109928 296156 115500 296212
rect 115556 296156 115566 296212
rect 199864 296044 201852 296100
rect 201908 296044 201918 296100
rect 439880 295820 441868 295876
rect 441924 295820 441934 295876
rect 369880 295708 373772 295764
rect 373828 295708 373838 295764
rect 112578 295596 112588 295652
rect 112644 295596 115276 295652
rect 115332 295596 115342 295652
rect 115826 295372 115836 295428
rect 115892 295372 120120 295428
rect 439880 295148 442316 295204
rect 442372 295148 442382 295204
rect 206322 295036 206332 295092
rect 206388 295036 210056 295092
rect 199864 294924 201740 294980
rect 201796 294924 201806 294980
rect 369880 294588 373772 294644
rect 373828 294588 373838 294644
rect 439880 294476 440188 294532
rect 440244 294476 440254 294532
rect 112018 294252 112028 294308
rect 112084 294252 120120 294308
rect 199864 293804 201740 293860
rect 201796 293804 201806 293860
rect 372866 293804 372876 293860
rect 372932 293804 380072 293860
rect 439880 293804 440524 293860
rect 440580 293804 440590 293860
rect 369880 293468 375452 293524
rect 375508 293468 375518 293524
rect 113586 293132 113596 293188
rect 113652 293132 120120 293188
rect 439880 293132 440300 293188
rect 440356 293132 440366 293188
rect 109928 292796 115388 292852
rect 115444 292796 115454 292852
rect 199864 292684 202524 292740
rect 202580 292684 202590 292740
rect 372642 292460 372652 292516
rect 372708 292460 380072 292516
rect 439880 292460 440188 292516
rect 440244 292460 440254 292516
rect 200834 292348 200844 292404
rect 200900 292348 210056 292404
rect 369880 292348 372092 292404
rect 372148 292348 372158 292404
rect 109928 292124 112700 292180
rect 112756 292124 112766 292180
rect 117170 292012 117180 292068
rect 117236 292012 120120 292068
rect 113474 291900 113484 291956
rect 113540 291900 114716 291956
rect 114772 291900 114782 291956
rect 439880 291788 441980 291844
rect 442036 291788 442046 291844
rect 199864 291564 201852 291620
rect 201908 291564 201918 291620
rect 109928 291452 112588 291508
rect 112644 291452 112654 291508
rect 113698 291340 113708 291396
rect 113764 291340 114268 291396
rect 114324 291340 114334 291396
rect 369880 291228 375676 291284
rect 375732 291228 375742 291284
rect 379362 291116 379372 291172
rect 379428 291116 380072 291172
rect 439880 291116 442428 291172
rect 442484 291116 442494 291172
rect -960 290836 480 291032
rect 113922 290892 113932 290948
rect 113988 290892 120120 290948
rect -960 290808 4732 290836
rect 392 290780 4732 290808
rect 4788 290780 4798 290836
rect 109928 290780 112812 290836
rect 112868 290780 112878 290836
rect 112690 290668 112700 290724
rect 112756 290668 119084 290724
rect 119140 290668 119150 290724
rect 199864 290444 200508 290500
rect 200564 290444 200574 290500
rect 377794 290444 377804 290500
rect 377860 290444 380072 290500
rect 439880 290444 440748 290500
rect 440804 290444 440814 290500
rect 369880 290108 373660 290164
rect 373716 290108 373726 290164
rect 114706 289772 114716 289828
rect 114772 289772 120120 289828
rect 376898 289772 376908 289828
rect 376964 289772 380072 289828
rect 439880 289772 442092 289828
rect 442148 289772 442158 289828
rect 204642 289660 204652 289716
rect 204708 289660 210056 289716
rect 54936 289436 58604 289492
rect 58660 289436 58670 289492
rect 109928 289436 114044 289492
rect 114100 289436 114110 289492
rect 199864 289324 201964 289380
rect 202020 289324 202030 289380
rect 380482 289100 380492 289156
rect 380548 289100 380558 289156
rect 369880 288988 372428 289044
rect 372484 288988 372494 289044
rect 54936 288764 59836 288820
rect 59892 288764 59902 288820
rect 109928 288764 112588 288820
rect 112644 288764 112654 288820
rect 114258 288652 114268 288708
rect 114324 288652 120120 288708
rect 379250 288428 379260 288484
rect 379316 288428 380072 288484
rect 54796 288316 59612 288372
rect 59668 288316 59678 288372
rect 54796 288120 54852 288316
rect 56130 288092 56140 288148
rect 56196 288092 60088 288148
rect 199276 287588 199332 288232
rect 369880 287868 373884 287924
rect 373940 287868 373950 287924
rect 379138 287756 379148 287812
rect 379204 287756 380072 287812
rect 113810 287532 113820 287588
rect 113876 287532 120120 287588
rect 199266 287532 199276 287588
rect 199332 287532 199342 287588
rect 54936 287420 58716 287476
rect 58772 287420 58782 287476
rect 199864 287084 201628 287140
rect 201684 287084 201694 287140
rect 378914 287084 378924 287140
rect 378980 287084 380072 287140
rect 209346 286972 209356 287028
rect 209412 286972 210056 287028
rect 369880 286748 372316 286804
rect 372372 286748 372382 286804
rect 117394 286412 117404 286468
rect 117460 286412 120120 286468
rect 380604 286132 380660 286440
rect 109928 286076 112700 286132
rect 112756 286076 112766 286132
rect 380594 286076 380604 286132
rect 380660 286076 380670 286132
rect 199864 285964 202076 286020
rect 202132 285964 202142 286020
rect 370626 285740 370636 285796
rect 370692 285740 380072 285796
rect 369880 285628 371980 285684
rect 372036 285628 372046 285684
rect 5170 285404 5180 285460
rect 5236 285404 5246 285460
rect 117170 285292 117180 285348
rect 117236 285292 120120 285348
rect 377234 285068 377244 285124
rect 377300 285068 380072 285124
rect 210018 284956 210028 285012
rect 210084 284956 210094 285012
rect 199864 284844 203644 284900
rect 203700 284844 203710 284900
rect 1474 284732 1484 284788
rect 1540 284732 5096 284788
rect 54936 284732 58716 284788
rect 58772 284732 58782 284788
rect 202402 284732 202412 284788
rect 202468 284732 207676 284788
rect 207732 284732 207742 284788
rect 111122 284508 111132 284564
rect 111188 284508 113372 284564
rect 113428 284508 113438 284564
rect 210028 284312 210084 284956
rect 595560 284676 597000 284872
rect 565282 284620 565292 284676
rect 565348 284648 597000 284676
rect 565348 284620 595672 284648
rect 369880 284508 373324 284564
rect 373380 284508 373390 284564
rect 379026 284396 379036 284452
rect 379092 284396 380072 284452
rect 115490 284172 115500 284228
rect 115556 284172 120120 284228
rect 5516 283892 5572 284088
rect 54936 284060 58716 284116
rect 58772 284060 58782 284116
rect 5506 283836 5516 283892
rect 5572 283836 5582 283892
rect 199864 283724 202188 283780
rect 202244 283724 202254 283780
rect 377906 283724 377916 283780
rect 377972 283724 380072 283780
rect 5282 283388 5292 283444
rect 5348 283388 5358 283444
rect 54936 283388 58716 283444
rect 58772 283388 58782 283444
rect 369880 283388 375564 283444
rect 375620 283388 375630 283444
rect 117506 283052 117516 283108
rect 117572 283052 120120 283108
rect 374434 283052 374444 283108
rect 374500 283052 380072 283108
rect 68786 282940 68796 282996
rect 68852 282940 119980 282996
rect 120036 282940 120046 282996
rect 87602 282828 87612 282884
rect 87668 282828 116956 282884
rect 117012 282828 117022 282884
rect 5740 282324 5796 282744
rect 199864 282604 200844 282660
rect 200900 282604 200910 282660
rect 5740 282268 7532 282324
rect 7588 282268 7598 282324
rect 115154 282268 115164 282324
rect 115220 282268 116004 282324
rect 369880 282268 373436 282324
rect 373492 282268 373502 282324
rect 115948 282212 116004 282268
rect 115948 282156 120148 282212
rect 109554 282044 109564 282100
rect 109620 282044 115164 282100
rect 115220 282044 115230 282100
rect 120092 281960 120148 282156
rect 53442 281820 53452 281876
rect 53508 281820 59612 281876
rect 59668 281820 59678 281876
rect 97346 281820 97356 281876
rect 97412 281820 119868 281876
rect 119924 281820 119934 281876
rect 40674 281708 40684 281764
rect 40740 281708 60060 281764
rect 60116 281708 60126 281764
rect 75506 281708 75516 281764
rect 75572 281708 117292 281764
rect 117348 281708 117358 281764
rect 25890 281596 25900 281652
rect 25956 281596 59836 281652
rect 59892 281596 59902 281652
rect 85586 281596 85596 281652
rect 85652 281596 117068 281652
rect 117124 281596 117134 281652
rect 204306 281596 204316 281652
rect 204372 281596 210056 281652
rect 26562 281484 26572 281540
rect 26628 281484 55132 281540
rect 55188 281484 55198 281540
rect 58146 281484 58156 281540
rect 58212 281484 119196 281540
rect 119252 281484 119262 281540
rect 2706 281372 2716 281428
rect 2772 281372 118860 281428
rect 118916 281372 118926 281428
rect 369880 281148 374892 281204
rect 374948 281148 374958 281204
rect 13132 280924 73948 280980
rect 85586 280924 85596 280980
rect 85652 280924 85662 280980
rect 97346 280924 97356 280980
rect 97412 280924 97422 280980
rect 13132 280644 13188 280924
rect 45378 280812 45388 280868
rect 45444 280812 54572 280868
rect 54628 280812 54638 280868
rect 73892 280756 73948 280924
rect 85596 280756 85652 280924
rect 97356 280756 97412 280924
rect 116834 280812 116844 280868
rect 116900 280812 120120 280868
rect 31892 280700 56924 280756
rect 56980 280700 56990 280756
rect 63746 280700 63756 280756
rect 63812 280700 70140 280756
rect 70196 280700 70206 280756
rect 73892 280700 74172 280756
rect 74228 280700 74238 280756
rect 74834 280700 74844 280756
rect 74900 280700 85652 280756
rect 87574 280700 87612 280756
rect 87668 280700 87678 280756
rect 89618 280700 89628 280756
rect 89684 280700 97412 280756
rect 121510 280700 121548 280756
rect 121604 280700 121614 280756
rect 199490 280700 199500 280756
rect 199556 280700 199948 280756
rect 200004 280700 200014 280756
rect 31892 280644 31948 280700
rect 13122 280588 13132 280644
rect 13188 280588 13198 280644
rect 23874 280588 23884 280644
rect 23940 280588 31948 280644
rect 40646 280588 40684 280644
rect 40740 280588 40750 280644
rect 44706 280588 44716 280644
rect 44772 280588 53452 280644
rect 53508 280588 53518 280644
rect 57810 280588 57820 280644
rect 57876 280588 141708 280644
rect 141764 280588 141774 280644
rect 157042 280588 157052 280644
rect 157108 280588 201628 280644
rect 201684 280588 201694 280644
rect 3154 280476 3164 280532
rect 3220 280476 5068 280532
rect 5124 280476 5134 280532
rect 25862 280476 25900 280532
rect 25956 280476 25966 280532
rect 26534 280476 26572 280532
rect 26628 280476 26638 280532
rect 45350 280476 45388 280532
rect 45444 280476 45454 280532
rect 58258 280476 58268 280532
rect 58324 280476 127484 280532
rect 127540 280476 127550 280532
rect 127670 280476 127708 280532
rect 127764 280476 127774 280532
rect 133606 280476 133644 280532
rect 133700 280476 133710 280532
rect 139654 280476 139692 280532
rect 139748 280476 139758 280532
rect 140998 280476 141036 280532
rect 141092 280476 141102 280532
rect 146374 280476 146412 280532
rect 146468 280476 146478 280532
rect 163622 280476 163660 280532
rect 163716 280476 163726 280532
rect 186386 280476 186396 280532
rect 186452 280476 194572 280532
rect 194628 280476 194638 280532
rect 198118 280476 198156 280532
rect 198212 280476 198222 280532
rect 44034 280364 44044 280420
rect 44100 280364 54684 280420
rect 54740 280364 54750 280420
rect 60386 280364 60396 280420
rect 60452 280364 151788 280420
rect 151844 280364 151854 280420
rect 186274 280364 186284 280420
rect 186340 280364 195020 280420
rect 195076 280364 195086 280420
rect 37986 280252 37996 280308
rect 38052 280252 49532 280308
rect 49588 280252 49598 280308
rect 54898 280252 54908 280308
rect 54964 280252 153132 280308
rect 153188 280252 153198 280308
rect 4610 280140 4620 280196
rect 4676 280140 166572 280196
rect 166628 280140 166638 280196
rect 23202 280028 23212 280084
rect 23268 280028 31948 280084
rect 74134 280028 74172 280084
rect 74228 280028 74238 280084
rect 75478 280028 75516 280084
rect 75572 280028 75582 280084
rect 77494 280028 77532 280084
rect 77588 280028 77598 280084
rect 119298 280028 119308 280084
rect 119364 280028 119374 280084
rect 121846 280028 121884 280084
rect 121940 280028 121950 280084
rect 122322 280028 122332 280084
rect 122388 280028 123004 280084
rect 123060 280028 123070 280084
rect 127474 280028 127484 280084
rect 127540 280028 137676 280084
rect 137732 280028 137742 280084
rect 149492 280028 159852 280084
rect 159908 280028 159918 280084
rect 194786 280028 194796 280084
rect 194852 280028 194862 280084
rect 369880 280028 374780 280084
rect 374836 280028 374846 280084
rect 31892 279972 31948 280028
rect 119308 279972 119364 280028
rect 149492 279972 149548 280028
rect 194796 279972 194852 280028
rect 31892 279916 81676 279972
rect 81732 279916 81742 279972
rect 119308 279916 123676 279972
rect 123732 279916 123742 279972
rect 125682 279916 125692 279972
rect 125748 279916 149548 279972
rect 194562 279916 194572 279972
rect 194628 279916 194852 279972
rect 27234 279804 27244 279860
rect 27300 279804 58044 279860
rect 58100 279804 58110 279860
rect 70802 279804 70812 279860
rect 70868 279804 111916 279860
rect 111972 279804 111982 279860
rect 119186 279804 119196 279860
rect 119252 279804 132300 279860
rect 132356 279804 132366 279860
rect 165666 279804 165676 279860
rect 165732 279804 206892 279860
rect 206948 279804 206958 279860
rect 76178 279692 76188 279748
rect 76244 279692 112700 279748
rect 112756 279692 112766 279748
rect 121426 279692 121436 279748
rect 121492 279692 125020 279748
rect 125076 279692 125086 279748
rect 137666 279692 137676 279748
rect 137732 279692 200732 279748
rect 200788 279692 200798 279748
rect 4722 279580 4732 279636
rect 4788 279580 167244 279636
rect 167300 279580 167310 279636
rect 115378 279468 115388 279524
rect 115444 279468 125692 279524
rect 125748 279468 125758 279524
rect 119970 279356 119980 279412
rect 120036 279356 134988 279412
rect 135044 279356 135054 279412
rect 105298 279020 105308 279076
rect 105364 279020 112588 279076
rect 112644 279020 114044 279076
rect 114100 279020 114110 279076
rect 111122 278908 111132 278964
rect 111188 278908 113484 278964
rect 113540 278908 113550 278964
rect 206210 278908 206220 278964
rect 206276 278908 210056 278964
rect 369880 278908 375004 278964
rect 375060 278908 375070 278964
rect 34626 278796 34636 278852
rect 34692 278796 52892 278852
rect 52948 278796 52958 278852
rect 72818 278796 72828 278852
rect 72884 278796 109228 278852
rect 109284 278796 109294 278852
rect 199154 278796 199164 278852
rect 199220 278796 200060 278852
rect 200116 278796 200126 278852
rect 54450 278684 54460 278740
rect 54516 278684 164556 278740
rect 164612 278684 164622 278740
rect 174598 278684 174636 278740
rect 174692 278684 174702 278740
rect 31266 278572 31276 278628
rect 31332 278572 54572 278628
rect 54628 278572 54638 278628
rect 58482 278572 58492 278628
rect 58548 278572 145068 278628
rect 145124 278572 145134 278628
rect 170482 278572 170492 278628
rect 170548 278572 193340 278628
rect 193396 278572 193406 278628
rect 36866 278460 36876 278516
rect 36932 278460 59724 278516
rect 59780 278460 59790 278516
rect 74134 278460 74172 278516
rect 74228 278460 74238 278516
rect 118850 278460 118860 278516
rect 118916 278460 173292 278516
rect 173348 278460 173358 278516
rect 187366 278460 187404 278516
rect 187460 278460 187470 278516
rect 12450 278348 12460 278404
rect 12516 278348 78204 278404
rect 78260 278348 78270 278404
rect 82226 278348 82236 278404
rect 82292 278348 109564 278404
rect 109620 278348 109630 278404
rect 111794 278348 111804 278404
rect 111860 278348 173964 278404
rect 174020 278348 174030 278404
rect 186162 278348 186172 278404
rect 186228 278348 196700 278404
rect 196756 278348 196766 278404
rect 42690 278236 42700 278292
rect 42756 278236 60620 278292
rect 60676 278236 60686 278292
rect 62066 278236 62076 278292
rect 62132 278236 113372 278292
rect 113428 278236 113438 278292
rect 136966 278236 137004 278292
rect 137060 278236 137070 278292
rect 168802 278236 168812 278292
rect 168868 278236 200620 278292
rect 200676 278236 200686 278292
rect 16818 278124 16828 278180
rect 16884 278124 56252 278180
rect 56308 278124 56318 278180
rect 60050 278124 60060 278180
rect 60116 278124 112700 278180
rect 112756 278124 112766 278180
rect 115014 278124 115052 278180
rect 115108 278124 115118 278180
rect 154466 278124 154476 278180
rect 154532 278124 197596 278180
rect 197652 278124 197662 278180
rect 26898 278012 26908 278068
rect 26964 278012 72828 278068
rect 72884 278012 72894 278068
rect 106866 278012 106876 278068
rect 106932 278012 201740 278068
rect 201796 278012 201806 278068
rect 530002 278012 530012 278068
rect 530068 278012 590492 278068
rect 590548 278012 590558 278068
rect 20514 277900 20524 277956
rect 20580 277900 60508 277956
rect 60564 277900 60574 277956
rect 62738 277900 62748 277956
rect 62804 277900 105308 277956
rect 105364 277900 105374 277956
rect 118626 277900 118636 277956
rect 118692 277900 184044 277956
rect 184100 277900 184110 277956
rect 5506 277788 5516 277844
rect 5572 277788 131628 277844
rect 131684 277788 131694 277844
rect 369880 277788 372092 277844
rect 372148 277788 372158 277844
rect 58706 277676 58716 277732
rect 58772 277676 126252 277732
rect 126308 277676 126318 277732
rect 7046 277116 7084 277172
rect 7140 277116 7150 277172
rect 7718 277116 7756 277172
rect 7812 277116 7822 277172
rect 35298 277116 35308 277172
rect 35364 277116 45276 277172
rect 45332 277116 45342 277172
rect 48710 277116 48748 277172
rect 48804 277116 48814 277172
rect 50082 277116 50092 277172
rect 50148 277116 56140 277172
rect 56196 277116 61404 277172
rect 61460 277116 61470 277172
rect 63858 277116 63868 277172
rect 63924 277116 65436 277172
rect 65492 277116 71932 277172
rect 71988 277116 71998 277172
rect 75618 277116 75628 277172
rect 75684 277116 76860 277172
rect 76916 277116 83580 277172
rect 83636 277116 83646 277172
rect 83804 277116 90300 277172
rect 90356 277116 90366 277172
rect 101042 277116 101052 277172
rect 101108 277116 110236 277172
rect 110292 277116 110302 277172
rect 119970 277116 119980 277172
rect 120036 277116 124348 277172
rect 124404 277116 124414 277172
rect 151078 277116 151116 277172
rect 151172 277116 151182 277172
rect 157938 277116 157948 277172
rect 158004 277116 159180 277172
rect 159236 277116 159246 277172
rect 159926 277116 159964 277172
rect 160020 277116 160030 277172
rect 165190 277116 165228 277172
rect 165284 277116 165294 277172
rect 165862 277116 165900 277172
rect 165956 277116 165966 277172
rect 175270 277116 175308 277172
rect 175364 277116 175374 277172
rect 178882 277116 178892 277172
rect 178948 277116 196588 277172
rect 196644 277116 196654 277172
rect 208292 277116 210364 277172
rect 210420 277116 210430 277172
rect 372082 277116 372092 277172
rect 372148 277116 441868 277172
rect 441924 277116 441934 277172
rect 83804 277060 83860 277116
rect 6402 277004 6412 277060
rect 6468 277004 16828 277060
rect 16884 277004 17612 277060
rect 17668 277004 17678 277060
rect 48066 277004 48076 277060
rect 48132 277004 57036 277060
rect 57092 277004 57102 277060
rect 63382 277004 63420 277060
rect 63476 277004 63486 277060
rect 81442 277004 81452 277060
rect 81508 277004 83860 277060
rect 84242 277004 84252 277060
rect 84308 277004 113596 277060
rect 113652 277004 113662 277060
rect 120530 277004 120540 277060
rect 120596 277004 149100 277060
rect 149156 277004 149166 277060
rect 166226 277004 166236 277060
rect 166292 277004 179340 277060
rect 179396 277004 179406 277060
rect 181346 277004 181356 277060
rect 181412 277004 195916 277060
rect 195972 277004 195982 277060
rect -960 276724 480 276920
rect 11106 276892 11116 276948
rect 11172 276892 60060 276948
rect 60116 276892 60126 276948
rect 62178 276892 62188 276948
rect 62244 276892 67452 276948
rect 67508 276892 80724 276948
rect 84802 276892 84812 276948
rect 84868 276892 84924 276948
rect 84980 276892 93660 276948
rect 93716 276892 93726 276948
rect 94322 276892 94332 276948
rect 94388 276892 110460 276948
rect 110516 276892 110526 276948
rect 120306 276892 120316 276948
rect 120372 276892 145740 276948
rect 145796 276892 145806 276948
rect 160402 276892 160412 276948
rect 160468 276892 167916 276948
rect 167972 276892 167982 276948
rect 5730 276780 5740 276836
rect 5796 276780 26908 276836
rect 26964 276780 26974 276836
rect 29250 276780 29260 276836
rect 29316 276780 76188 276836
rect 76244 276780 76254 276836
rect 80668 276724 80724 276892
rect 80882 276780 80892 276836
rect 80948 276780 82236 276836
rect 82292 276780 82302 276836
rect 97682 276780 97692 276836
rect 97748 276780 106764 276836
rect 106820 276780 106830 276836
rect 108322 276780 108332 276836
rect 108388 276780 120876 276836
rect 120932 276780 120942 276836
rect 147858 276780 147868 276836
rect 147924 276780 162540 276836
rect 162596 276780 162606 276836
rect 163762 276780 163772 276836
rect 163828 276780 190092 276836
rect 190148 276780 190158 276836
rect -960 276696 7980 276724
rect 392 276668 7980 276696
rect 8036 276668 8046 276724
rect 24546 276668 24556 276724
rect 24612 276668 62076 276724
rect 62132 276668 62142 276724
rect 64082 276668 64092 276724
rect 64148 276668 64204 276724
rect 64260 276668 64270 276724
rect 70354 276668 70364 276724
rect 70420 276668 79548 276724
rect 79604 276668 79614 276724
rect 80668 276668 82908 276724
rect 82964 276668 119196 276724
rect 119252 276668 119262 276724
rect 160514 276668 160524 276724
rect 160580 276668 192780 276724
rect 192836 276668 192846 276724
rect 208292 276612 208348 277116
rect 373314 277004 373324 277060
rect 373380 277004 440300 277060
rect 440356 277004 440366 277060
rect 373762 276892 373772 276948
rect 373828 276892 440636 276948
rect 440692 276892 440702 276948
rect 375442 276780 375452 276836
rect 375508 276780 442204 276836
rect 442260 276780 442270 276836
rect 369880 276668 373548 276724
rect 373604 276668 373614 276724
rect 375666 276668 375676 276724
rect 375732 276668 442428 276724
rect 442484 276668 442494 276724
rect 13794 276556 13804 276612
rect 13860 276556 26572 276612
rect 26628 276556 26638 276612
rect 29922 276556 29932 276612
rect 29988 276556 60396 276612
rect 60452 276556 60462 276612
rect 63410 276556 63420 276612
rect 63476 276556 69468 276612
rect 69524 276556 70252 276612
rect 70308 276556 70318 276612
rect 72146 276556 72156 276612
rect 72212 276556 88956 276612
rect 89012 276556 89022 276612
rect 114034 276556 114044 276612
rect 114100 276556 178892 276612
rect 178948 276556 178958 276612
rect 186386 276556 186396 276612
rect 186452 276556 208348 276612
rect 374770 276556 374780 276612
rect 374836 276556 442092 276612
rect 442148 276556 442158 276612
rect 10434 276444 10444 276500
rect 10500 276444 62748 276500
rect 62804 276444 62814 276500
rect 68114 276444 68124 276500
rect 68180 276444 68796 276500
rect 68852 276444 80892 276500
rect 80948 276444 80958 276500
rect 85652 276444 88284 276500
rect 88340 276444 189420 276500
rect 189476 276444 189486 276500
rect 9090 276332 9100 276388
rect 9156 276332 23436 276388
rect 23492 276332 23502 276388
rect 47394 276332 47404 276388
rect 47460 276332 56924 276388
rect 56980 276332 56990 276388
rect 63858 276332 63868 276388
rect 63924 276332 64764 276388
rect 64820 276332 73052 276388
rect 73108 276332 73118 276388
rect 78194 276332 78204 276388
rect 78260 276332 82236 276388
rect 82292 276332 82302 276388
rect 85652 276276 85708 276444
rect 97412 276332 188972 276388
rect 189028 276332 189532 276388
rect 189588 276332 189598 276388
rect 377906 276332 377916 276388
rect 377972 276332 440524 276388
rect 440580 276332 440590 276388
rect 97412 276276 97468 276332
rect 9762 276220 9772 276276
rect 9828 276220 60732 276276
rect 60788 276220 60798 276276
rect 73892 276220 85708 276276
rect 91532 276220 97468 276276
rect 118738 276220 118748 276276
rect 118804 276220 149772 276276
rect 149828 276220 149838 276276
rect 175942 276220 175980 276276
rect 176036 276220 176046 276276
rect 186694 276220 186732 276276
rect 186788 276220 186798 276276
rect 210690 276220 210700 276276
rect 210756 276220 210766 276276
rect 73892 276164 73948 276220
rect 38658 276108 38668 276164
rect 38724 276108 48636 276164
rect 48692 276108 48702 276164
rect 57026 276108 57036 276164
rect 57092 276108 73948 276164
rect 82226 276108 82236 276164
rect 82292 276108 90972 276164
rect 91028 276108 91038 276164
rect 91532 276052 91588 276220
rect 92978 276108 92988 276164
rect 93044 276108 118972 276164
rect 119028 276108 119038 276164
rect 197026 276108 197036 276164
rect 197092 276108 197484 276164
rect 197540 276108 197550 276164
rect 56914 275996 56924 276052
rect 56980 275996 80220 276052
rect 80276 275996 91588 276052
rect 94882 275996 94892 276052
rect 94948 275996 95676 276052
rect 95732 275996 95742 276052
rect 108658 275996 108668 276052
rect 108724 275996 122892 276052
rect 122948 275996 122958 276052
rect 188066 275884 188076 275940
rect 188132 275884 203420 275940
rect 203476 275884 203486 275940
rect 180002 275772 180012 275828
rect 180068 275772 181356 275828
rect 181412 275772 181422 275828
rect 184678 275772 184716 275828
rect 184772 275772 184782 275828
rect 199714 275772 199724 275828
rect 199780 275772 202412 275828
rect 202468 275772 202478 275828
rect 179778 275660 179788 275716
rect 179844 275660 180684 275716
rect 180740 275660 180750 275716
rect 183138 275660 183148 275716
rect 183204 275660 186060 275716
rect 186116 275660 186126 275716
rect 188066 275660 188076 275716
rect 188132 275660 194124 275716
rect 194180 275660 194190 275716
rect 372642 275660 372652 275716
rect 372708 275660 384748 275716
rect 384692 275604 384748 275660
rect 26002 275548 26012 275604
rect 26068 275548 26572 275604
rect 26628 275548 26638 275604
rect 36838 275548 36876 275604
rect 36932 275548 36942 275604
rect 41094 275548 41132 275604
rect 41188 275548 41198 275604
rect 61366 275548 61404 275604
rect 61460 275548 61470 275604
rect 64054 275548 64092 275604
rect 64148 275548 64158 275604
rect 65538 275548 65548 275604
rect 65604 275548 66780 275604
rect 66836 275548 72156 275604
rect 72212 275548 72222 275604
rect 100818 275548 100828 275604
rect 100884 275548 101724 275604
rect 101780 275548 103628 275604
rect 103684 275548 103694 275604
rect 168102 275548 168140 275604
rect 168196 275548 168206 275604
rect 169222 275548 169260 275604
rect 169316 275548 169326 275604
rect 169670 275548 169708 275604
rect 169764 275548 169774 275604
rect 176502 275548 176540 275604
rect 176596 275548 176606 275604
rect 177286 275548 177324 275604
rect 177380 275548 177390 275604
rect 178070 275548 178108 275604
rect 178164 275548 178174 275604
rect 179862 275548 179900 275604
rect 179956 275548 179966 275604
rect 181430 275548 181468 275604
rect 181524 275548 181534 275604
rect 184818 275548 184828 275604
rect 184884 275548 184922 275604
rect 188710 275548 188748 275604
rect 188804 275548 188814 275604
rect 189382 275548 189420 275604
rect 189476 275548 189486 275604
rect 190418 275548 190428 275604
rect 190484 275548 191436 275604
rect 191492 275548 191502 275604
rect 197698 275548 197708 275604
rect 197764 275548 201628 275604
rect 201684 275548 201694 275604
rect 369880 275548 375116 275604
rect 375172 275548 375182 275604
rect 384692 275548 442092 275604
rect 442148 275548 442158 275604
rect 15138 275436 15148 275492
rect 15204 275436 143052 275492
rect 143108 275436 143118 275492
rect 189074 275436 189084 275492
rect 189140 275436 199612 275492
rect 199668 275436 199678 275492
rect 373650 275436 373660 275492
rect 373716 275436 440748 275492
rect 440804 275436 440814 275492
rect 58370 275324 58380 275380
rect 58436 275324 161196 275380
rect 161252 275324 161262 275380
rect 374882 275324 374892 275380
rect 374948 275324 441980 275380
rect 442036 275324 442046 275380
rect 56690 275212 56700 275268
rect 56756 275212 158508 275268
rect 158564 275212 158574 275268
rect 375554 275212 375564 275268
rect 375620 275212 442316 275268
rect 442372 275212 442382 275268
rect 59490 275100 59500 275156
rect 59556 275100 157164 275156
rect 157220 275100 157230 275156
rect 373426 275100 373436 275156
rect 373492 275100 440188 275156
rect 440244 275100 440254 275156
rect 60274 274988 60284 275044
rect 60340 274988 152460 275044
rect 152516 274988 152526 275044
rect 46722 274876 46732 274932
rect 46788 274876 135660 274932
rect 135716 274876 135726 274932
rect 21858 274764 21868 274820
rect 21924 274764 84812 274820
rect 84868 274764 84878 274820
rect 86930 274764 86940 274820
rect 86996 274764 115164 274820
rect 115220 274764 115230 274820
rect 119186 274764 119196 274820
rect 119252 274764 199052 274820
rect 199108 274764 199118 274820
rect 375778 274764 375788 274820
rect 375844 274764 443660 274820
rect 443716 274764 443726 274820
rect 11778 274652 11788 274708
rect 11844 274652 65548 274708
rect 65604 274652 65614 274708
rect 68674 274652 68684 274708
rect 68740 274652 94892 274708
rect 94948 274652 94958 274708
rect 103394 274652 103404 274708
rect 103460 274652 202636 274708
rect 202692 274652 202702 274708
rect 371858 274652 371868 274708
rect 371924 274652 441980 274708
rect 442036 274652 442046 274708
rect 8418 274540 8428 274596
rect 8484 274540 68796 274596
rect 68852 274540 68862 274596
rect 72146 274540 72156 274596
rect 72212 274540 117068 274596
rect 117124 274540 117134 274596
rect 120194 274540 120204 274596
rect 120260 274540 150332 274596
rect 150388 274540 150398 274596
rect 369880 274428 375228 274484
rect 375284 274428 375294 274484
rect 25218 273756 25228 273812
rect 25284 273756 63868 273812
rect 63924 273756 63934 273812
rect 113362 273756 113372 273812
rect 113428 273756 196812 273812
rect 196868 273756 196878 273812
rect 372418 273756 372428 273812
rect 372484 273756 442764 273812
rect 442820 273756 442830 273812
rect 85586 273644 85596 273700
rect 85652 273644 115276 273700
rect 115332 273644 115342 273700
rect 118514 273644 118524 273700
rect 118580 273644 195468 273700
rect 195524 273644 195534 273700
rect 373874 273644 373884 273700
rect 373940 273644 440524 273700
rect 440580 273644 440590 273700
rect 56466 273532 56476 273588
rect 56532 273532 156492 273588
rect 156548 273532 156558 273588
rect 209234 273532 209244 273588
rect 209300 273532 210056 273588
rect 372194 273532 372204 273588
rect 372260 273532 413644 273588
rect 413700 273532 413710 273588
rect 58034 273420 58044 273476
rect 58100 273420 147868 273476
rect 147924 273420 147934 273476
rect 375778 273420 375788 273476
rect 375844 273420 408268 273476
rect 408324 273420 408334 273476
rect 31938 273308 31948 273364
rect 32004 273308 108332 273364
rect 108388 273308 108398 273364
rect 110002 273308 110012 273364
rect 110068 273308 194796 273364
rect 194852 273308 194862 273364
rect 369880 273308 373324 273364
rect 373380 273308 373390 273364
rect 375554 273308 375564 273364
rect 375620 273308 407596 273364
rect 407652 273308 407662 273364
rect 410274 273308 410284 273364
rect 410340 273308 422604 273364
rect 422660 273308 422670 273364
rect 60722 273196 60732 273252
rect 60788 273196 100828 273252
rect 100884 273196 100894 273252
rect 406466 273196 406476 273252
rect 406532 273196 423948 273252
rect 424004 273196 424014 273252
rect 19170 273084 19180 273140
rect 19236 273084 39676 273140
rect 39732 273084 66108 273140
rect 66164 273084 86268 273140
rect 86324 273084 86334 273140
rect 104962 273084 104972 273140
rect 105028 273084 202524 273140
rect 202580 273084 202590 273140
rect 374994 273084 375004 273140
rect 375060 273084 442092 273140
rect 442148 273084 442158 273140
rect 4162 272972 4172 273028
rect 4228 272972 166236 273028
rect 166292 272972 166302 273028
rect 370738 272972 370748 273028
rect 370804 272972 440188 273028
rect 440244 272972 440254 273028
rect 70354 272860 70364 272916
rect 70420 272860 79772 272916
rect 79828 272860 79838 272916
rect 21186 272748 21196 272804
rect 21252 272748 128940 272804
rect 128996 272748 129006 272804
rect 22530 272636 22540 272692
rect 22596 272636 126924 272692
rect 126980 272636 126990 272692
rect 369880 272188 404012 272244
rect 404068 272188 404078 272244
rect 111682 272076 111692 272132
rect 111748 272076 196140 272132
rect 196196 272076 196206 272132
rect 385382 272076 385420 272132
rect 385476 272076 385486 272132
rect 387202 272076 387212 272132
rect 387268 272076 390124 272132
rect 390180 272076 390190 272132
rect 27906 271964 27916 272020
rect 27972 271964 142380 272020
rect 142436 271964 142446 272020
rect 383842 271964 383852 272020
rect 383908 271964 406252 272020
rect 406308 271964 406318 272020
rect 419906 271964 419916 272020
rect 419972 271964 423388 272020
rect 423444 271964 423454 272020
rect 16482 271852 16492 271908
rect 16548 271852 130956 271908
rect 131012 271852 131022 271908
rect 387426 271852 387436 271908
rect 387492 271852 412972 271908
rect 413028 271852 413038 271908
rect 417452 271852 420028 271908
rect 417452 271796 417508 271852
rect 419972 271796 420028 271852
rect 35970 271740 35980 271796
rect 36036 271740 144396 271796
rect 144452 271740 144462 271796
rect 379922 271740 379932 271796
rect 379988 271740 417004 271796
rect 417060 271740 417070 271796
rect 417442 271740 417452 271796
rect 417508 271740 417518 271796
rect 419972 271740 431788 271796
rect 431844 271740 431854 271796
rect 51202 271628 51212 271684
rect 51268 271628 155820 271684
rect 155876 271628 155886 271684
rect 372418 271628 372428 271684
rect 372484 271628 409612 271684
rect 409668 271628 409678 271684
rect 416294 271628 416332 271684
rect 416388 271628 416398 271684
rect 419906 271628 419916 271684
rect 419972 271628 425068 271684
rect 425124 271628 425134 271684
rect 51426 271516 51436 271572
rect 51492 271516 155148 271572
rect 155204 271516 155214 271572
rect 373314 271516 373324 271572
rect 373380 271516 383404 271572
rect 383460 271516 383470 271572
rect 394146 271516 394156 271572
rect 394212 271516 431788 271572
rect 431844 271516 431854 271572
rect 595560 271460 597000 271656
rect 62962 271404 62972 271460
rect 63028 271404 163884 271460
rect 163940 271404 163950 271460
rect 374322 271404 374332 271460
rect 374388 271404 381388 271460
rect 381444 271404 381454 271460
rect 390114 271404 390124 271460
rect 390180 271404 430108 271460
rect 430164 271404 430174 271460
rect 550162 271404 550172 271460
rect 550228 271432 597000 271460
rect 550228 271404 595672 271432
rect 17154 271292 17164 271348
rect 17220 271292 28476 271348
rect 28532 271292 75628 271348
rect 75684 271292 75694 271348
rect 78866 271292 78876 271348
rect 78932 271292 116732 271348
rect 116788 271292 116798 271348
rect 167122 271292 167132 271348
rect 167188 271292 194348 271348
rect 194404 271292 194414 271348
rect 370962 271292 370972 271348
rect 371028 271292 384076 271348
rect 384132 271292 384142 271348
rect 387314 271292 387324 271348
rect 387380 271292 431900 271348
rect 431956 271292 431966 271348
rect 71922 271180 71932 271236
rect 71988 271180 100044 271236
rect 100100 271180 100110 271236
rect 118402 271180 118412 271236
rect 118468 271180 177996 271236
rect 178052 271180 178062 271236
rect 376226 271180 376236 271236
rect 376292 271180 380044 271236
rect 380100 271180 380110 271236
rect 409938 271180 409948 271236
rect 410004 271180 410956 271236
rect 411012 271180 411022 271236
rect 419972 271180 420140 271236
rect 420196 271180 420206 271236
rect 7522 271068 7532 271124
rect 7588 271068 132972 271124
rect 133028 271068 133038 271124
rect 369880 271068 381388 271124
rect 381444 271068 381454 271124
rect 388098 271068 388108 271124
rect 388164 271068 389452 271124
rect 389508 271068 389518 271124
rect 410022 271068 410060 271124
rect 410116 271068 410126 271124
rect 411618 271068 411628 271124
rect 411684 271068 412300 271124
rect 412356 271068 412366 271124
rect 413298 271068 413308 271124
rect 413364 271068 414316 271124
rect 414372 271068 414382 271124
rect 414978 271068 414988 271124
rect 415044 271068 415660 271124
rect 415716 271068 415726 271124
rect 418338 271068 418348 271124
rect 418404 271068 419692 271124
rect 419748 271068 419758 271124
rect 419972 271012 420028 271180
rect 373986 270956 373996 271012
rect 374052 270956 380716 271012
rect 380772 270956 380782 271012
rect 409826 270956 409836 271012
rect 409892 270956 420028 271012
rect 210242 270844 210252 270900
rect 210308 270844 210318 270900
rect 374994 270844 375004 270900
rect 375060 270844 382732 270900
rect 382788 270844 382798 270900
rect 374210 270732 374220 270788
rect 374276 270732 382060 270788
rect 382116 270732 382126 270788
rect 157042 270508 157052 270564
rect 157108 270508 176428 270564
rect 176484 270508 176494 270564
rect 7634 270396 7644 270452
rect 7700 270396 193452 270452
rect 193508 270396 193518 270452
rect 387986 270396 387996 270452
rect 388052 270396 441868 270452
rect 441924 270396 441934 270452
rect 18 270284 28 270340
rect 84 270284 172620 270340
rect 172676 270284 172686 270340
rect 371970 270284 371980 270340
rect 372036 270284 410788 270340
rect 410946 270284 410956 270340
rect 411012 270284 418460 270340
rect 418516 270284 418526 270340
rect 420354 270284 420364 270340
rect 420420 270284 422044 270340
rect 422100 270284 422110 270340
rect 410732 270228 410788 270284
rect 14466 270172 14476 270228
rect 14532 270172 127596 270228
rect 127652 270172 127662 270228
rect 372306 270172 372316 270228
rect 372372 270172 408940 270228
rect 408996 270172 409006 270228
rect 410732 270172 414988 270228
rect 415044 270172 415054 270228
rect 56242 270060 56252 270116
rect 56308 270060 154476 270116
rect 154532 270060 154542 270116
rect 194534 270060 194572 270116
rect 194628 270060 194638 270116
rect 375442 270060 375452 270116
rect 375508 270060 401548 270116
rect 401604 270060 401614 270116
rect 52994 269948 53004 270004
rect 53060 269948 150444 270004
rect 150500 269948 150510 270004
rect 172162 269948 172172 270004
rect 172228 269948 197372 270004
rect 197428 269948 197438 270004
rect 369880 269948 415660 270004
rect 415716 269948 415726 270004
rect 23426 269836 23436 269892
rect 23492 269836 68684 269892
rect 68740 269836 68750 269892
rect 105186 269836 105196 269892
rect 105252 269836 201852 269892
rect 201908 269836 201918 269892
rect 381378 269836 381388 269892
rect 381444 269836 404236 269892
rect 404292 269836 404302 269892
rect 405122 269836 405132 269892
rect 405188 269836 420028 269892
rect 420084 269836 420094 269892
rect 15810 269724 15820 269780
rect 15876 269724 21756 269780
rect 21812 269724 64092 269780
rect 64148 269724 64158 269780
rect 99922 269724 99932 269780
rect 99988 269724 201964 269780
rect 202020 269724 202030 269780
rect 377346 269724 377356 269780
rect 377412 269724 411628 269780
rect 411684 269724 411694 269780
rect 7522 269612 7532 269668
rect 7588 269612 190764 269668
rect 190820 269612 190830 269668
rect 372530 269612 372540 269668
rect 372596 269612 441084 269668
rect 441140 269612 441150 269668
rect 58594 269500 58604 269556
rect 58660 269500 134316 269556
rect 134372 269500 134382 269556
rect 370962 269500 370972 269556
rect 371028 269500 387436 269556
rect 387492 269500 387502 269556
rect 411730 268940 411740 268996
rect 411796 268940 418796 268996
rect 418852 268940 418862 268996
rect 369880 268828 440412 268884
rect 440468 268828 440478 268884
rect 4274 268716 4284 268772
rect 4340 268716 183372 268772
rect 183428 268716 183438 268772
rect 420018 268716 420028 268772
rect 420084 268716 421484 268772
rect 421540 268716 430444 268772
rect 430500 268716 430510 268772
rect 119074 268604 119084 268660
rect 119140 268604 185612 268660
rect 185668 268604 186396 268660
rect 186452 268604 186462 268660
rect 56354 268492 56364 268548
rect 56420 268492 157836 268548
rect 157892 268492 157902 268548
rect 375666 268492 375676 268548
rect 375732 268492 386764 268548
rect 386820 268492 386830 268548
rect 42018 268380 42028 268436
rect 42084 268380 139020 268436
rect 139076 268380 139086 268436
rect 139346 268380 139356 268436
rect 139412 268380 199836 268436
rect 199892 268380 199902 268436
rect 372754 268380 372764 268436
rect 372820 268380 384748 268436
rect 384804 268380 384814 268436
rect 49410 268268 49420 268324
rect 49476 268268 143724 268324
rect 143780 268268 143790 268324
rect 374546 268268 374556 268324
rect 374612 268268 388108 268324
rect 388164 268268 388174 268324
rect 56578 268156 56588 268212
rect 56644 268156 147756 268212
rect 147812 268156 147822 268212
rect 206098 268156 206108 268212
rect 206164 268156 210056 268212
rect 372418 268156 372428 268212
rect 372484 268156 386092 268212
rect 386148 268156 386158 268212
rect 82226 268044 82236 268100
rect 82292 268044 99932 268100
rect 99988 268044 99998 268100
rect 111682 268044 111692 268100
rect 111748 268044 192108 268100
rect 192164 268044 192174 268100
rect 381490 268044 381500 268100
rect 381556 268044 406924 268100
rect 406980 268044 406990 268100
rect 418338 268044 418348 268100
rect 418404 268044 426748 268100
rect 426804 268044 440188 268100
rect 440244 268044 440254 268100
rect 7746 267932 7756 267988
rect 7812 267932 171276 267988
rect 171332 267932 171342 267988
rect 380034 267932 380044 267988
rect 380100 267932 405580 267988
rect 405636 267932 405646 267988
rect 409602 267932 409612 267988
rect 409668 267932 419916 267988
rect 419972 267932 440412 267988
rect 440468 267932 440478 267988
rect 18498 267820 18508 267876
rect 18564 267820 129612 267876
rect 129668 267820 129678 267876
rect 424610 267820 424620 267876
rect 424676 267820 429772 267876
rect 429828 267820 429838 267876
rect 369880 267708 374668 267764
rect 374724 267708 374734 267764
rect 376002 267708 376012 267764
rect 376068 267708 408716 267764
rect 408772 267708 409836 267764
rect 409892 267708 409902 267764
rect 414978 267708 414988 267764
rect 415044 267708 426860 267764
rect 426916 267708 445228 267764
rect 445284 267708 445294 267764
rect 380146 267596 380156 267652
rect 380212 267596 417452 267652
rect 417508 267596 417518 267652
rect 403554 267484 403564 267540
rect 403620 267484 423052 267540
rect 423108 267484 423118 267540
rect 375218 267372 375228 267428
rect 375284 267372 405580 267428
rect 405636 267372 405646 267428
rect 423378 267372 423388 267428
rect 423444 267372 428428 267428
rect 428484 267372 428494 267428
rect 408930 267260 408940 267316
rect 408996 267260 419916 267316
rect 419972 267260 442316 267316
rect 442372 267260 442382 267316
rect 416322 267148 416332 267204
rect 416388 267148 418572 267204
rect 418628 267148 418638 267204
rect 420326 267148 420364 267204
rect 420420 267148 420430 267204
rect 7970 267036 7980 267092
rect 8036 267036 182700 267092
rect 182756 267036 182766 267092
rect 61282 266924 61292 266980
rect 61348 266924 153804 266980
rect 153860 266924 153870 266980
rect 380258 266924 380268 266980
rect 380324 266924 417676 266980
rect 417732 266924 417742 266980
rect 418572 266868 418628 267148
rect 46050 266812 46060 266868
rect 46116 266812 136332 266868
rect 136388 266812 136398 266868
rect 374658 266812 374668 266868
rect 374724 266812 412972 266868
rect 413028 266812 413038 266868
rect 418572 266812 443660 266868
rect 443716 266812 443726 266868
rect 60498 266700 60508 266756
rect 60564 266700 147084 266756
rect 147140 266700 147150 266756
rect 373538 266700 373548 266756
rect 373604 266700 440300 266756
rect 440356 266700 440366 266756
rect 59378 266588 59388 266644
rect 59444 266588 140364 266644
rect 140420 266588 140430 266644
rect 369880 266588 375676 266644
rect 375732 266588 375742 266644
rect 380034 266588 380044 266644
rect 380100 266588 420028 266644
rect 420084 266588 420094 266644
rect 122546 266476 122556 266532
rect 122612 266476 197484 266532
rect 197540 266476 197550 266532
rect 375106 266476 375116 266532
rect 375172 266476 441980 266532
rect 442036 266476 442046 266532
rect 17826 266364 17836 266420
rect 17892 266364 26796 266420
rect 26852 266364 81452 266420
rect 81508 266364 81518 266420
rect 83906 266364 83916 266420
rect 83972 266364 199612 266420
rect 199668 266364 199678 266420
rect 373314 266364 373324 266420
rect 373380 266364 440524 266420
rect 440580 266364 440590 266420
rect 7634 266252 7644 266308
rect 7700 266252 170604 266308
rect 170660 266252 170670 266308
rect 194226 266252 194236 266308
rect 194292 266252 202524 266308
rect 202580 266252 202590 266308
rect 370738 266252 370748 266308
rect 370804 266252 440972 266308
rect 441028 266252 441038 266308
rect 113698 266140 113708 266196
rect 113764 266140 181468 266196
rect 181524 266140 181534 266196
rect 209906 266028 209916 266084
rect 209972 266028 210084 266084
rect 185602 265468 185612 265524
rect 185668 265468 187404 265524
rect 187460 265468 187470 265524
rect 210028 265496 210084 266028
rect 403526 265692 403564 265748
rect 403620 265692 403630 265748
rect 410918 265692 410956 265748
rect 411012 265692 411022 265748
rect 375330 265580 375340 265636
rect 375396 265580 412300 265636
rect 412356 265580 412366 265636
rect 369880 265468 370076 265524
rect 370132 265468 370142 265524
rect 376114 265468 376124 265524
rect 376180 265468 414316 265524
rect 414372 265468 414382 265524
rect 115826 265356 115836 265412
rect 115892 265356 157052 265412
rect 157108 265356 157118 265412
rect 181458 265356 181468 265412
rect 181524 265356 183036 265412
rect 183092 265356 199276 265412
rect 199332 265356 199342 265412
rect 373202 265356 373212 265412
rect 373268 265356 407596 265412
rect 407652 265356 407662 265412
rect 410274 265356 410284 265412
rect 410340 265356 441980 265412
rect 442036 265356 442046 265412
rect 57922 265244 57932 265300
rect 57988 265244 161868 265300
rect 161924 265244 161934 265300
rect 375442 265244 375452 265300
rect 375508 265244 411628 265300
rect 411684 265244 411694 265300
rect 43362 265132 43372 265188
rect 43428 265132 138348 265188
rect 138404 265132 138414 265188
rect 373874 265132 373884 265188
rect 373940 265132 442428 265188
rect 442484 265132 442494 265188
rect 60162 265020 60172 265076
rect 60228 265020 148428 265076
rect 148484 265020 148494 265076
rect 373090 265020 373100 265076
rect 373156 265020 388780 265076
rect 388836 265020 388846 265076
rect 404002 265020 404012 265076
rect 404068 265020 442316 265076
rect 442372 265020 442382 265076
rect 119186 264908 119196 264964
rect 119252 264908 189084 264964
rect 189140 264908 189150 264964
rect 379250 264908 379260 264964
rect 379316 264908 442540 264964
rect 442596 264908 442606 264964
rect 19842 264796 19852 264852
rect 19908 264796 130284 264852
rect 130340 264796 130350 264852
rect 379138 264796 379148 264852
rect 379204 264796 442652 264852
rect 442708 264796 442718 264852
rect 73042 264684 73052 264740
rect 73108 264684 104972 264740
rect 105028 264684 105038 264740
rect 373874 264684 373884 264740
rect 373940 264684 439292 264740
rect 439348 264684 439358 264740
rect 6738 264572 6748 264628
rect 6804 264572 171948 264628
rect 172004 264572 172014 264628
rect 375218 264572 375228 264628
rect 375284 264572 442204 264628
rect 442260 264572 442270 264628
rect 379474 264460 379484 264516
rect 379540 264460 404908 264516
rect 404964 264460 404974 264516
rect 416994 264460 417004 264516
rect 417060 264460 423388 264516
rect 423444 264460 433468 264516
rect 433524 264460 433534 264516
rect 369880 264348 372204 264404
rect 372260 264348 372270 264404
rect 406242 264348 406252 264404
rect 406308 264348 406318 264404
rect 406252 264292 406308 264348
rect 403526 264236 403564 264292
rect 403620 264236 403630 264292
rect 406214 264236 406252 264292
rect 406308 264236 406318 264292
rect 406886 264236 406924 264292
rect 406980 264236 406990 264292
rect 410918 264236 410956 264292
rect 411012 264236 411022 264292
rect 413606 264236 413644 264292
rect 413700 264236 413710 264292
rect 189046 264124 189084 264180
rect 189140 264124 189150 264180
rect 373426 263900 373436 263956
rect 373492 263900 374444 263956
rect 374500 263900 374510 263956
rect 373650 263788 373660 263844
rect 373716 263788 374108 263844
rect 374164 263788 374174 263844
rect 380594 263676 380604 263732
rect 380660 263676 410956 263732
rect 411012 263676 411022 263732
rect 426178 263676 426188 263732
rect 426244 263676 434252 263732
rect 434308 263676 434318 263732
rect 379586 263564 379596 263620
rect 379652 263564 411628 263620
rect 411684 263564 411694 263620
rect 380146 263452 380156 263508
rect 380212 263452 414988 263508
rect 415044 263452 415054 263508
rect 379362 263340 379372 263396
rect 379428 263340 406252 263396
rect 406308 263340 406318 263396
rect 406914 263340 406924 263396
rect 406980 263340 411740 263396
rect 411796 263340 443548 263396
rect 443604 263340 443614 263396
rect 369880 263228 440972 263284
rect 441028 263228 441038 263284
rect 379810 263116 379820 263172
rect 379876 263116 413364 263172
rect 413634 263116 413644 263172
rect 413700 263116 431788 263172
rect 413308 263060 413364 263116
rect 431732 263060 431788 263116
rect 371186 263004 371196 263060
rect 371252 263004 410060 263060
rect 410116 263004 410126 263060
rect 413308 263004 418348 263060
rect 418404 263004 418414 263060
rect 431732 263004 433580 263060
rect 433636 263004 445340 263060
rect 445396 263004 445406 263060
rect 373762 262892 373772 262948
rect 373828 262892 440860 262948
rect 440916 262892 440926 262948
rect 392 262808 6748 262836
rect -960 262780 6748 262808
rect 6804 262780 6814 262836
rect 204418 262780 204428 262836
rect 204484 262780 210056 262836
rect -960 262584 480 262780
rect 369880 262108 370412 262164
rect 370468 262108 370478 262164
rect 375890 261660 375900 261716
rect 375956 261660 388108 261716
rect 388164 261660 388174 261716
rect 378802 261548 378812 261604
rect 378868 261548 409948 261604
rect 410004 261548 410014 261604
rect 369880 260988 373884 261044
rect 373940 260988 373950 261044
rect 210130 260092 210140 260148
rect 210196 260092 210206 260148
rect 369880 259868 375564 259924
rect 375620 259868 375630 259924
rect 369880 258748 372092 258804
rect 372148 258748 372158 258804
rect 595560 258244 597000 258440
rect 555202 258188 555212 258244
rect 555268 258216 597000 258244
rect 555268 258188 595672 258216
rect 369880 257628 372540 257684
rect 372596 257628 372606 257684
rect 210690 257404 210700 257460
rect 210756 257404 210766 257460
rect 369880 256508 375788 256564
rect 375844 256508 375854 256564
rect 372866 256060 372876 256116
rect 372932 256060 377580 256116
rect 377636 256060 380100 256116
rect 377122 255836 377132 255892
rect 377188 255836 377580 255892
rect 377636 255836 377646 255892
rect 369880 255388 375340 255444
rect 375396 255388 375406 255444
rect 380044 255416 380100 256060
rect 208002 254716 208012 254772
rect 208068 254716 210056 254772
rect 369880 254268 377132 254324
rect 377188 254268 377198 254324
rect 369880 253148 376124 253204
rect 376180 253148 376190 253204
rect 206098 252028 206108 252084
rect 206164 252028 207564 252084
rect 207620 252028 207630 252084
rect 207890 252028 207900 252084
rect 207956 252028 210056 252084
rect 369880 252028 376460 252084
rect 376516 252028 376526 252084
rect 369880 250908 373324 250964
rect 373380 250908 373390 250964
rect 375330 250012 375340 250068
rect 375396 250012 377580 250068
rect 377636 250012 380072 250068
rect 369880 249788 372988 249844
rect 373044 249788 373054 249844
rect 379922 249564 379932 249620
rect 379988 249564 380100 249620
rect 204306 249452 204316 249508
rect 204372 249452 208012 249508
rect 208068 249452 208078 249508
rect 207778 249340 207788 249396
rect 207844 249340 210056 249396
rect 380044 248948 380100 249564
rect 376114 248892 376124 248948
rect 376180 248892 380100 248948
rect 371074 248780 371084 248836
rect 371140 248780 373772 248836
rect 373828 248780 380100 248836
rect -960 248612 480 248696
rect 369880 248668 373212 248724
rect 373268 248668 373278 248724
rect 380044 248696 380100 248780
rect -960 248556 4956 248612
rect 5012 248556 5022 248612
rect -960 248472 480 248556
rect 376226 247996 376236 248052
rect 376292 247996 380072 248052
rect 369880 247548 375452 247604
rect 375508 247548 375518 247604
rect 376450 247324 376460 247380
rect 376516 247324 380072 247380
rect 373398 246876 373436 246932
rect 373492 246876 373502 246932
rect 375442 246876 375452 246932
rect 375508 246876 376236 246932
rect 376292 246876 376302 246932
rect 208114 246652 208124 246708
rect 208180 246652 210056 246708
rect 377458 246652 377468 246708
rect 377524 246652 379596 246708
rect 379652 246652 380072 246708
rect 369880 246428 376460 246484
rect 376516 246428 376526 246484
rect 370514 245980 370524 246036
rect 370580 245980 371196 246036
rect 371252 245980 380072 246036
rect 372932 245420 375228 245476
rect 375284 245420 375294 245476
rect 372932 245364 372988 245420
rect 369880 245308 372988 245364
rect 373762 245308 373772 245364
rect 373828 245308 380072 245364
rect 595560 245028 597000 245224
rect 587122 244972 587132 245028
rect 587188 245000 597000 245028
rect 587188 244972 595672 245000
rect 376450 244636 376460 244692
rect 376516 244636 380072 244692
rect 369880 244188 373884 244244
rect 373940 244188 373950 244244
rect 208226 243964 208236 244020
rect 208292 243964 210056 244020
rect 377570 243964 377580 244020
rect 377636 243964 379820 244020
rect 379876 243964 380072 244020
rect 377346 243292 377356 243348
rect 377412 243292 380072 243348
rect 380146 243180 380156 243236
rect 380212 243180 380222 243236
rect 369880 243068 376236 243124
rect 376292 243068 376302 243124
rect 373650 242732 373660 242788
rect 373716 242732 373884 242788
rect 373940 242732 373950 242788
rect 380156 242676 380212 243180
rect 378578 242620 378588 242676
rect 378644 242648 380212 242676
rect 378644 242620 380184 242648
rect 374546 242172 374556 242228
rect 374612 242172 380492 242228
rect 380548 242172 380558 242228
rect 371084 242060 373884 242116
rect 373940 242060 373950 242116
rect 371084 242004 371140 242060
rect 369880 241948 371140 242004
rect 372978 241948 372988 242004
rect 373044 241948 380072 242004
rect 439880 241948 440188 242004
rect 440244 241948 440254 242004
rect 380034 241724 380044 241780
rect 380100 241724 380110 241780
rect 380044 241332 380100 241724
rect 207666 241276 207676 241332
rect 207732 241276 210056 241332
rect 377234 241276 377244 241332
rect 377300 241304 380100 241332
rect 377300 241276 380072 241304
rect 379922 241164 379932 241220
rect 379988 241164 380100 241220
rect 369880 240828 373436 240884
rect 373492 240828 373502 240884
rect 380044 240660 380100 241164
rect 371970 240604 371980 240660
rect 372036 240632 380100 240660
rect 372036 240604 380072 240632
rect 439880 240604 440412 240660
rect 440468 240604 440478 240660
rect 373986 240380 373996 240436
rect 374052 240380 380604 240436
rect 380660 240380 380670 240436
rect 373622 240268 373660 240324
rect 373716 240268 373726 240324
rect 376226 240268 376236 240324
rect 376292 240268 379820 240324
rect 379876 240268 379886 240324
rect 372866 240156 372876 240212
rect 372932 240156 373772 240212
rect 373828 240156 373838 240212
rect 371074 240044 371084 240100
rect 371140 240044 372988 240100
rect 373044 240044 373054 240100
rect 369880 239708 370076 239764
rect 370132 239708 370142 239764
rect 380044 239540 380100 239960
rect 439852 239876 439908 239960
rect 439852 239820 439964 239876
rect 440020 239820 440030 239876
rect 372418 239484 372428 239540
rect 372484 239484 376684 239540
rect 376740 239484 376750 239540
rect 379652 239484 380100 239540
rect 379652 239428 379708 239484
rect 370850 239372 370860 239428
rect 370916 239372 378812 239428
rect 378868 239372 379708 239428
rect 376674 239260 376684 239316
rect 376740 239260 377132 239316
rect 377188 239260 380072 239316
rect 373538 238812 373548 238868
rect 373604 238812 373884 238868
rect 373940 238812 373950 238868
rect 372932 238700 375564 238756
rect 375620 238700 375630 238756
rect 372932 238644 372988 238700
rect 210018 238588 210028 238644
rect 210084 238588 210094 238644
rect 369880 238588 372988 238644
rect 373314 238588 373324 238644
rect 373380 238588 380072 238644
rect 380044 237860 380100 237944
rect 371186 237804 371196 237860
rect 371252 237804 379484 237860
rect 379540 237804 380100 237860
rect 375890 237692 375900 237748
rect 375956 237692 378924 237748
rect 378980 237692 378990 237748
rect 380258 237580 380268 237636
rect 380324 237580 380334 237636
rect 369880 237468 375900 237524
rect 375956 237468 375966 237524
rect 380268 236964 380324 237580
rect 439880 237244 442316 237300
rect 442372 237244 442382 237300
rect 379922 236908 379932 236964
rect 379988 236908 380324 236964
rect 372194 236796 372204 236852
rect 372260 236796 373660 236852
rect 373716 236796 373726 236852
rect 380034 236796 380044 236852
rect 380100 236796 380110 236852
rect 380044 236628 380100 236796
rect 377010 236572 377020 236628
rect 377076 236600 380100 236628
rect 377076 236572 380072 236600
rect 439880 236572 442092 236628
rect 442148 236572 442158 236628
rect 369880 236348 375116 236404
rect 375172 236348 375182 236404
rect 210690 235900 210700 235956
rect 210756 235900 210766 235956
rect 376226 235900 376236 235956
rect 376292 235900 380072 235956
rect 439880 235900 440300 235956
rect 440356 235900 440366 235956
rect 373650 235788 373660 235844
rect 373716 235788 380100 235844
rect 369880 235228 375228 235284
rect 375284 235228 375294 235284
rect 380044 235256 380100 235788
rect 375330 235116 375340 235172
rect 375396 235116 378028 235172
rect 378084 235116 378094 235172
rect 440962 235116 440972 235172
rect 441028 235116 441868 235172
rect 441924 235116 441934 235172
rect 371158 234780 371196 234836
rect 371252 234780 371262 234836
rect 392 234584 11004 234612
rect -960 234556 11004 234584
rect 11060 234556 11070 234612
rect 373762 234556 373772 234612
rect 373828 234556 380072 234612
rect -960 234360 480 234556
rect 370626 234332 370636 234388
rect 370692 234332 379708 234388
rect 379764 234332 379774 234388
rect 369880 234108 372316 234164
rect 372372 234108 372382 234164
rect 373874 233884 373884 233940
rect 373940 233884 380072 233940
rect 373398 233436 373436 233492
rect 373492 233436 373502 233492
rect 373986 233436 373996 233492
rect 374052 233436 375452 233492
rect 375508 233436 375518 233492
rect 207554 233212 207564 233268
rect 207620 233212 210056 233268
rect 371858 233212 371868 233268
rect 371924 233212 373884 233268
rect 373940 233212 380072 233268
rect 439880 233212 442204 233268
rect 442260 233212 442270 233268
rect 369880 232988 373660 233044
rect 373716 232988 373726 233044
rect 372306 232540 372316 232596
rect 372372 232540 372540 232596
rect 372596 232540 380072 232596
rect 439880 232540 441980 232596
rect 442036 232540 442046 232596
rect 595560 231924 597000 232008
rect 369880 231868 371868 231924
rect 371924 231868 371934 231924
rect 373986 231868 373996 231924
rect 374052 231868 380072 231924
rect 439880 231868 440524 231924
rect 440580 231868 440590 231924
rect 543554 231868 543564 231924
rect 543620 231868 597000 231924
rect 595560 231784 597000 231868
rect 370738 231196 370748 231252
rect 370804 231196 375340 231252
rect 375396 231196 380072 231252
rect 371746 230972 371756 231028
rect 371812 230972 379148 231028
rect 379204 230972 380100 231028
rect 369880 230748 370300 230804
rect 370356 230748 370366 230804
rect 209122 230524 209132 230580
rect 209188 230524 210056 230580
rect 380044 230552 380100 230972
rect 377122 229852 377132 229908
rect 377188 229852 380072 229908
rect 439880 229852 442428 229908
rect 442484 229852 442494 229908
rect 369880 229628 370132 229684
rect 370076 229012 370132 229628
rect 372642 229292 372652 229348
rect 372708 229292 378476 229348
rect 378532 229292 378542 229348
rect 371186 229180 371196 229236
rect 371252 229180 372652 229236
rect 372708 229180 380072 229236
rect 439880 229180 441868 229236
rect 441924 229180 441934 229236
rect 370076 228956 373436 229012
rect 373492 228956 373502 229012
rect 369880 228508 371644 228564
rect 371700 228508 371710 228564
rect 380370 228508 380380 228564
rect 380436 228508 380446 228564
rect 439880 228508 442204 228564
rect 442260 228508 442270 228564
rect 205986 227836 205996 227892
rect 206052 227836 210056 227892
rect 377682 227836 377692 227892
rect 377748 227836 378812 227892
rect 378868 227836 380072 227892
rect 369880 227388 370412 227444
rect 370468 227388 370478 227444
rect 375778 227164 375788 227220
rect 375844 227164 377580 227220
rect 377636 227164 380072 227220
rect 374882 226492 374892 226548
rect 374948 226492 379260 226548
rect 379316 226492 380072 226548
rect 439880 226492 442092 226548
rect 442148 226492 442158 226548
rect 369880 226268 370188 226324
rect 370244 226268 370254 226324
rect 372418 225932 372428 225988
rect 372484 225932 377468 225988
rect 377524 225932 380100 225988
rect 380044 225848 380100 225932
rect 376002 225260 376012 225316
rect 376068 225260 376236 225316
rect 376292 225260 376302 225316
rect 208292 225148 210056 225204
rect 369880 225148 375228 225204
rect 375284 225148 375294 225204
rect 376114 225148 376124 225204
rect 376180 225148 380072 225204
rect 208292 225092 208348 225148
rect 204978 225036 204988 225092
rect 205044 225036 208348 225092
rect 372978 225036 372988 225092
rect 373044 225036 373772 225092
rect 373828 225036 373838 225092
rect 376114 224476 376124 224532
rect 376180 224476 376796 224532
rect 376852 224476 380072 224532
rect 370626 224364 370636 224420
rect 370692 224364 372988 224420
rect 373044 224364 380100 224420
rect 369880 224028 370636 224084
rect 370692 224028 370702 224084
rect 380044 223832 380100 224364
rect 380258 223132 380268 223188
rect 380324 223132 380334 223188
rect 369880 222908 371980 222964
rect 372036 222908 372046 222964
rect 372642 222684 372652 222740
rect 372708 222684 378588 222740
rect 378644 222684 378654 222740
rect 370738 222572 370748 222628
rect 370804 222572 378700 222628
rect 378756 222572 380100 222628
rect 204978 222460 204988 222516
rect 205044 222460 210056 222516
rect 380044 222488 380100 222572
rect 369394 221788 369404 221844
rect 369460 221788 369470 221844
rect 378578 221788 378588 221844
rect 378644 221788 380072 221844
rect 379698 221676 379708 221732
rect 379764 221676 379932 221732
rect 379988 221676 379998 221732
rect 374658 221116 374668 221172
rect 374724 221116 377356 221172
rect 377412 221116 380072 221172
rect 369506 220668 369516 220724
rect 369572 220668 369582 220724
rect 392 220472 7756 220500
rect -960 220444 7756 220472
rect 7812 220444 7822 220500
rect 376226 220444 376236 220500
rect 376292 220444 380604 220500
rect 380660 220444 380670 220500
rect -960 220248 480 220444
rect 206658 219772 206668 219828
rect 206724 219772 210056 219828
rect 372082 219772 372092 219828
rect 372148 219772 380072 219828
rect 369880 219548 378700 219604
rect 378756 219548 378766 219604
rect 373538 219100 373548 219156
rect 373604 219100 376236 219156
rect 376292 219100 380072 219156
rect 372530 218652 372540 218708
rect 372596 218652 372764 218708
rect 372820 218652 380100 218708
rect 371746 218540 371756 218596
rect 371812 218540 374668 218596
rect 374724 218540 374734 218596
rect 369880 218428 373884 218484
rect 373940 218428 373950 218484
rect 380044 218456 380100 218652
rect 595560 218596 597000 218792
rect 543666 218540 543676 218596
rect 543732 218568 597000 218596
rect 543732 218540 595672 218568
rect 379922 218316 379932 218372
rect 379988 218316 380100 218372
rect 373090 217868 373100 217924
rect 373156 217868 379708 217924
rect 379764 217868 379774 217924
rect 380044 217812 380100 218316
rect 370738 217756 370748 217812
rect 370804 217784 380100 217812
rect 370804 217756 380072 217784
rect 369880 217308 379708 217364
rect 379764 217308 379774 217364
rect 206658 217084 206668 217140
rect 206724 217084 210056 217140
rect 374098 217084 374108 217140
rect 374164 217084 379484 217140
rect 379540 217084 380072 217140
rect 370626 216524 370636 216580
rect 370692 216524 373212 216580
rect 373268 216524 373278 216580
rect 380370 216412 380380 216468
rect 380436 216412 380446 216468
rect 369880 216188 373100 216244
rect 373156 216188 373166 216244
rect 375890 215740 375900 215796
rect 375956 215740 379484 215796
rect 379540 215740 380072 215796
rect 374210 215516 374220 215572
rect 374276 215516 379260 215572
rect 379316 215516 379326 215572
rect 374546 215404 374556 215460
rect 374612 215404 379484 215460
rect 379540 215404 379550 215460
rect 370188 215292 380380 215348
rect 380436 215292 380446 215348
rect 370188 215124 370244 215292
rect 370514 215180 370524 215236
rect 370580 215180 373548 215236
rect 373604 215180 380100 215236
rect 369880 215068 370244 215124
rect 373314 215068 373324 215124
rect 373380 215068 374556 215124
rect 374612 215068 374622 215124
rect 380044 215096 380100 215180
rect 373874 214508 373884 214564
rect 373940 214508 380324 214564
rect 206658 214396 206668 214452
rect 206724 214396 210056 214452
rect 369880 213948 373884 214004
rect 373940 213948 373950 214004
rect 380268 213668 380324 214508
rect 380258 213612 380268 213668
rect 380324 213612 380334 213668
rect 375414 213276 375452 213332
rect 375508 213276 375518 213332
rect 376114 213276 376124 213332
rect 376180 213276 376236 213332
rect 376292 213276 376302 213332
rect 373314 213164 373324 213220
rect 373380 213164 380268 213220
rect 380324 213164 380334 213220
rect 369880 212828 373884 212884
rect 373940 212828 373950 212884
rect 206658 211708 206668 211764
rect 206724 211708 210056 211764
rect 369880 211708 373884 211764
rect 373940 211708 373950 211764
rect 373398 211596 373436 211652
rect 373492 211596 373502 211652
rect 369880 210588 373660 210644
rect 373716 210588 373726 210644
rect 370710 209916 370748 209972
rect 370804 209916 370814 209972
rect 369880 209468 375452 209524
rect 375508 209468 375518 209524
rect 379698 209132 379708 209188
rect 379764 209132 380380 209188
rect 380436 209132 380446 209188
rect 206658 209020 206668 209076
rect 206724 209020 210056 209076
rect 372932 208460 375116 208516
rect 375172 208460 375182 208516
rect 372932 208404 372988 208460
rect 369880 208348 372988 208404
rect 378914 207340 378924 207396
rect 378980 207340 410956 207396
rect 411012 207340 411022 207396
rect 369880 207228 383068 207284
rect 383124 207228 383134 207284
rect 372082 207116 372092 207172
rect 372148 207116 399532 207172
rect 399588 207116 399598 207172
rect 370290 206668 370300 206724
rect 370356 206668 371756 206724
rect 371812 206668 371822 206724
rect 202374 206556 202412 206612
rect 202468 206556 208348 206612
rect 431778 206556 431788 206612
rect 431844 206556 442204 206612
rect 442260 206556 442270 206612
rect 208292 206388 208348 206556
rect 392 206360 4172 206388
rect -960 206332 4172 206360
rect 4228 206332 4238 206388
rect 208292 206332 210056 206388
rect 375218 206332 375228 206388
rect 375284 206332 385588 206388
rect -960 206136 480 206332
rect 385532 206276 385588 206332
rect 379362 206220 379372 206276
rect 379428 206220 385308 206276
rect 385364 206220 385374 206276
rect 385522 206220 385532 206276
rect 385588 206220 385598 206276
rect 369880 206108 403340 206164
rect 403396 206108 403406 206164
rect 375666 205996 375676 206052
rect 375732 205996 417004 206052
rect 417060 205996 417070 206052
rect 372306 205884 372316 205940
rect 372372 205884 396508 205940
rect 396452 205828 396508 205884
rect 380258 205772 380268 205828
rect 380324 205772 384804 205828
rect 396452 205772 407596 205828
rect 407652 205772 407662 205828
rect 384748 205716 384804 205772
rect 381798 205660 381836 205716
rect 381892 205660 381902 205716
rect 382050 205660 382060 205716
rect 382116 205660 382154 205716
rect 383366 205660 383404 205716
rect 383460 205660 383470 205716
rect 384738 205660 384748 205716
rect 384804 205660 384814 205716
rect 385522 205660 385532 205716
rect 385588 205660 442204 205716
rect 442260 205660 442270 205716
rect 373426 205548 373436 205604
rect 373492 205548 440636 205604
rect 440692 205548 440702 205604
rect 381154 205436 381164 205492
rect 381220 205436 383180 205492
rect 383236 205436 384076 205492
rect 384132 205436 384142 205492
rect 385298 205436 385308 205492
rect 385364 205436 414988 205492
rect 415044 205436 415054 205492
rect 416966 205436 417004 205492
rect 417060 205436 417070 205492
rect 595560 205380 597000 205576
rect 379138 205324 379148 205380
rect 379204 205324 419244 205380
rect 419300 205324 419310 205380
rect 560242 205324 560252 205380
rect 560308 205352 597000 205380
rect 560308 205324 595672 205352
rect 370850 205212 370860 205268
rect 370916 205212 385420 205268
rect 385476 205212 385486 205268
rect 386054 205212 386092 205268
rect 386148 205212 386158 205268
rect 386726 205212 386764 205268
rect 386820 205212 386830 205268
rect 389414 205212 389452 205268
rect 389508 205212 389518 205268
rect 395602 205212 395612 205268
rect 395668 205212 431788 205268
rect 431844 205212 431854 205268
rect 375228 205100 376516 205156
rect 399494 205100 399532 205156
rect 399588 205100 399598 205156
rect 403302 205100 403340 205156
rect 403396 205100 403406 205156
rect 410918 205100 410956 205156
rect 411012 205100 411022 205156
rect 413634 205100 413644 205156
rect 413700 205100 431900 205156
rect 431956 205100 431966 205156
rect 375228 205044 375284 205100
rect 376460 205044 376516 205100
rect 414764 205044 414820 205100
rect 369880 204988 375284 205044
rect 375442 204988 375452 205044
rect 375508 204988 376236 205044
rect 376292 204988 376302 205044
rect 376460 204988 391468 205044
rect 391524 204988 391534 205044
rect 407558 204988 407596 205044
rect 407652 204988 407662 205044
rect 414754 204988 414764 205044
rect 414820 204988 414830 205044
rect 414978 204988 414988 205044
rect 415044 204988 418572 205044
rect 418628 204988 418638 205044
rect 375554 204876 375564 204932
rect 375620 204876 408268 204932
rect 408324 204876 408334 204932
rect 372194 204764 372204 204820
rect 372260 204764 412300 204820
rect 412356 204764 412366 204820
rect 370402 204652 370412 204708
rect 370468 204652 410284 204708
rect 410340 204652 410350 204708
rect 379026 204540 379036 204596
rect 379092 204540 414316 204596
rect 414372 204540 414382 204596
rect 372530 204428 372540 204484
rect 372596 204428 406924 204484
rect 406980 204428 406990 204484
rect 375778 204316 375788 204372
rect 375844 204316 408940 204372
rect 408996 204316 409006 204372
rect 379250 204204 379260 204260
rect 379316 204204 416668 204260
rect 416724 204204 416734 204260
rect 419682 204204 419692 204260
rect 419748 204204 431788 204260
rect 431844 204204 431854 204260
rect 380482 204092 380492 204148
rect 380548 204092 418348 204148
rect 418404 204092 418414 204148
rect 370066 203980 370076 204036
rect 370132 203980 415660 204036
rect 415716 203980 415726 204036
rect 369880 203868 375900 203924
rect 375956 203868 375966 203924
rect 379250 203868 379260 203924
rect 379316 203868 380268 203924
rect 380324 203868 380334 203924
rect 402182 203868 402220 203924
rect 402276 203868 402286 203924
rect 204866 203644 204876 203700
rect 204932 203644 210056 203700
rect 382582 203196 382620 203252
rect 382676 203196 382686 203252
rect 383590 203196 383628 203252
rect 383684 203196 383694 203252
rect 388210 203196 388220 203252
rect 388276 203196 389452 203252
rect 389508 203196 389518 203252
rect 418338 203196 418348 203252
rect 418404 203196 427084 203252
rect 427140 203196 427150 203252
rect 370962 203084 370972 203140
rect 371028 203084 386428 203140
rect 386484 203084 387436 203140
rect 387492 203084 387502 203140
rect 418562 203084 418572 203140
rect 418628 203084 429772 203140
rect 429828 203084 429838 203140
rect 372754 202972 372764 203028
rect 372820 202972 377468 203028
rect 377524 202972 377534 203028
rect 381378 202972 381388 203028
rect 381444 202972 382396 203028
rect 382452 202972 382462 203028
rect 390572 202972 416332 203028
rect 416388 202972 416398 203028
rect 416658 202972 416668 203028
rect 416724 202972 423052 203028
rect 423108 202972 423118 203028
rect 390572 202916 390628 202972
rect 384412 202860 390628 202916
rect 390684 202860 412972 202916
rect 413028 202860 413038 202916
rect 414978 202860 414988 202916
rect 415044 202860 416556 202916
rect 416612 202860 440524 202916
rect 440580 202860 440590 202916
rect 369880 202748 384188 202804
rect 384244 202748 384254 202804
rect 384412 202692 384468 202860
rect 384626 202748 384636 202804
rect 384692 202748 390460 202804
rect 390516 202748 390526 202804
rect 390684 202692 390740 202860
rect 390898 202748 390908 202804
rect 390964 202748 400204 202804
rect 400260 202748 400270 202804
rect 376898 202636 376908 202692
rect 376964 202636 377916 202692
rect 377972 202636 377982 202692
rect 378476 202636 384468 202692
rect 384524 202636 390740 202692
rect 390796 202636 411628 202692
rect 411684 202636 411694 202692
rect 423042 202636 423052 202692
rect 423108 202636 433580 202692
rect 433636 202636 433646 202692
rect 378476 202580 378532 202636
rect 384524 202580 384580 202636
rect 372194 202524 372204 202580
rect 372260 202524 378476 202580
rect 378532 202524 378542 202580
rect 384300 202524 384580 202580
rect 384738 202524 384748 202580
rect 384804 202524 390572 202580
rect 390628 202524 390638 202580
rect 384300 202468 384356 202524
rect 390796 202468 390852 202636
rect 391010 202524 391020 202580
rect 391076 202524 417676 202580
rect 417732 202524 417742 202580
rect 427074 202524 427084 202580
rect 427140 202524 440524 202580
rect 440580 202524 440590 202580
rect 373202 202412 373212 202468
rect 373268 202412 374332 202468
rect 374388 202412 374398 202468
rect 377794 202412 377804 202468
rect 377860 202412 384356 202468
rect 384626 202412 384636 202468
rect 384692 202412 390852 202468
rect 414306 202412 414316 202468
rect 414372 202412 433692 202468
rect 433748 202412 433758 202468
rect 377458 202300 377468 202356
rect 377524 202300 418460 202356
rect 418516 202300 418526 202356
rect 370738 202188 370748 202244
rect 370804 202188 379708 202244
rect 379764 202188 419020 202244
rect 419076 202188 419086 202244
rect 377906 202076 377916 202132
rect 377972 202076 384636 202132
rect 384692 202076 384702 202132
rect 384066 201964 384076 202020
rect 384132 201964 384636 202020
rect 384692 201964 384702 202020
rect 397282 201852 397292 201908
rect 397348 201852 402220 201908
rect 402276 201852 402286 201908
rect 369880 201628 377468 201684
rect 377524 201628 377534 201684
rect 398178 201628 398188 201684
rect 398244 201628 404908 201684
rect 404964 201628 404974 201684
rect 429762 201628 429772 201684
rect 429828 201628 431900 201684
rect 431956 201628 431966 201684
rect 373538 201516 373548 201572
rect 373604 201516 374108 201572
rect 374164 201516 374174 201572
rect 374546 201516 374556 201572
rect 374612 201516 442092 201572
rect 442148 201516 442158 201572
rect 373314 201404 373324 201460
rect 373380 201404 373996 201460
rect 374052 201404 374062 201460
rect 380482 201404 380492 201460
rect 380548 201404 384748 201460
rect 384804 201404 388108 201460
rect 388164 201404 388174 201460
rect 404898 201404 404908 201460
rect 404964 201404 440300 201460
rect 440356 201404 440366 201460
rect 383842 201292 383852 201348
rect 383908 201292 388444 201348
rect 388500 201292 388780 201348
rect 388836 201292 388846 201348
rect 391458 201180 391468 201236
rect 391524 201180 411628 201236
rect 411684 201180 411694 201236
rect 392242 201068 392252 201124
rect 392308 201068 417676 201124
rect 417732 201068 417742 201124
rect 204978 200956 204988 201012
rect 205044 200956 210056 201012
rect 375890 200956 375900 201012
rect 375956 200956 413420 201012
rect 413476 200956 413486 201012
rect 373090 200844 373100 200900
rect 373156 200844 443772 200900
rect 443828 200844 443838 200900
rect 370290 200732 370300 200788
rect 370356 200732 441868 200788
rect 441924 200732 441934 200788
rect 369880 200508 445228 200564
rect 445284 200508 445294 200564
rect 384692 199668 384748 199892
rect 384804 199836 384814 199892
rect 381266 199612 381276 199668
rect 381332 199612 384748 199668
rect 416546 199612 416556 199668
rect 416612 199612 432012 199668
rect 432068 199612 432078 199668
rect 371858 199500 371868 199556
rect 371924 199500 408940 199556
rect 408996 199500 409006 199556
rect 414754 199500 414764 199556
rect 414820 199500 436828 199556
rect 436884 199500 436894 199556
rect 369880 199388 372092 199444
rect 372148 199388 372158 199444
rect 375218 199388 375228 199444
rect 375284 199388 410284 199444
rect 410340 199388 410350 199444
rect 410946 199388 410956 199444
rect 411012 199388 439404 199444
rect 439460 199388 439470 199444
rect 375890 199276 375900 199332
rect 375956 199276 417004 199332
rect 417060 199276 417070 199332
rect 371634 199164 371644 199220
rect 371700 199164 442316 199220
rect 442372 199164 442382 199220
rect 206658 199052 206668 199108
rect 206724 199052 208684 199108
rect 208740 199052 210084 199108
rect 370402 199052 370412 199108
rect 370468 199052 441980 199108
rect 442036 199052 442046 199108
rect 210028 198296 210084 199052
rect 379586 198492 379596 198548
rect 379652 198492 386092 198548
rect 386148 198492 386158 198548
rect 380258 198380 380268 198436
rect 380324 198380 384972 198436
rect 385028 198380 385038 198436
rect 369880 198268 375452 198324
rect 375508 198268 375518 198324
rect 380482 198268 380492 198324
rect 380548 198268 386764 198324
rect 386820 198268 386830 198324
rect 418310 198156 418348 198212
rect 418404 198156 418414 198212
rect 389750 198044 389788 198100
rect 389844 198044 389854 198100
rect 395714 197932 395724 197988
rect 395780 197932 412300 197988
rect 412356 197932 412366 197988
rect 383058 197820 383068 197876
rect 383124 197820 403564 197876
rect 403620 197820 403630 197876
rect 375106 197708 375116 197764
rect 375172 197708 405580 197764
rect 405636 197708 405646 197764
rect 375442 197596 375452 197652
rect 375508 197596 409612 197652
rect 409668 197596 409678 197652
rect 380370 197484 380380 197540
rect 380436 197484 416332 197540
rect 416388 197484 416398 197540
rect 379026 197372 379036 197428
rect 379092 197372 434252 197428
rect 434308 197372 434318 197428
rect 369880 197148 450268 197204
rect 450324 197148 450334 197204
rect 403330 197036 403340 197092
rect 403396 197036 410956 197092
rect 411012 197036 411022 197092
rect 373090 196700 373100 196756
rect 373156 196700 440300 196756
rect 440356 196700 440366 196756
rect 373202 196588 373212 196644
rect 373268 196588 448588 196644
rect 448644 196588 448654 196644
rect 382946 196364 382956 196420
rect 383012 196364 388444 196420
rect 388500 196364 388510 196420
rect 379138 196252 379148 196308
rect 379204 196252 388220 196308
rect 388276 196252 388286 196308
rect 379922 196140 379932 196196
rect 379988 196140 389788 196196
rect 389844 196140 389854 196196
rect 369880 196028 371420 196084
rect 371476 196028 371486 196084
rect 375890 196028 375900 196084
rect 375956 196028 386428 196084
rect 386484 196028 386494 196084
rect 373650 195916 373660 195972
rect 373716 195916 440300 195972
rect 440356 195916 440366 195972
rect 373874 195804 373884 195860
rect 373940 195804 443884 195860
rect 443940 195804 443950 195860
rect 371970 195692 371980 195748
rect 372036 195692 442876 195748
rect 442932 195692 442942 195748
rect 206882 195580 206892 195636
rect 206948 195580 207452 195636
rect 207508 195580 210056 195636
rect 375778 195132 375788 195188
rect 375844 195132 381724 195188
rect 381780 195132 381790 195188
rect 423332 195132 435148 195188
rect 423332 195076 423388 195132
rect 374434 195020 374444 195076
rect 374500 195020 423388 195076
rect 435092 195076 435148 195132
rect 435092 195020 446908 195076
rect 446964 195020 446974 195076
rect 369880 194908 373100 194964
rect 373156 194908 373166 194964
rect 373762 194908 373772 194964
rect 373828 194908 447020 194964
rect 447076 194908 447086 194964
rect 373986 194796 373996 194852
rect 374052 194796 423500 194852
rect 423556 194796 423566 194852
rect 423714 194796 423724 194852
rect 423780 194796 435148 194852
rect 435092 194740 435148 194796
rect 373874 194684 373884 194740
rect 373940 194684 423332 194740
rect 423388 194684 423398 194740
rect 435092 194684 443548 194740
rect 443604 194684 443614 194740
rect 378914 194572 378924 194628
rect 378980 194572 398188 194628
rect 398244 194572 398254 194628
rect 423490 194572 423500 194628
rect 423556 194572 445452 194628
rect 445508 194572 445518 194628
rect 374322 194460 374332 194516
rect 374388 194460 441868 194516
rect 441924 194460 441934 194516
rect 373650 194348 373660 194404
rect 373716 194348 442428 194404
rect 442484 194348 442494 194404
rect 3266 194012 3276 194068
rect 3332 194012 10892 194068
rect 10948 194012 10958 194068
rect 369880 193788 448588 193844
rect 448644 193788 448654 193844
rect 441970 193340 441980 193396
rect 442036 193340 442316 193396
rect 442372 193340 442382 193396
rect 373090 193228 373100 193284
rect 373156 193228 445564 193284
rect 445620 193228 445630 193284
rect 205202 192892 205212 192948
rect 205268 192892 210056 192948
rect 369880 192668 446908 192724
rect 446964 192668 446974 192724
rect 379138 192556 379148 192612
rect 379204 192556 397292 192612
rect 397348 192556 397358 192612
rect 375666 192444 375676 192500
rect 375732 192444 433468 192500
rect 433524 192444 433534 192500
rect 370178 192332 370188 192388
rect 370244 192332 442764 192388
rect 442820 192332 442830 192388
rect 392 192248 10892 192276
rect -960 192220 10892 192248
rect 10948 192220 10958 192276
rect -960 192024 480 192220
rect 595560 192164 597000 192360
rect 548482 192108 548492 192164
rect 548548 192136 597000 192164
rect 548548 192108 595672 192136
rect 373650 191772 373660 191828
rect 373716 191772 440188 191828
rect 440244 191772 440254 191828
rect 442166 191772 442204 191828
rect 442260 191772 442270 191828
rect 374098 191660 374108 191716
rect 374164 191660 443772 191716
rect 443828 191660 443838 191716
rect 369880 191548 445340 191604
rect 445396 191548 445406 191604
rect 369880 190428 373212 190484
rect 373268 190428 373278 190484
rect 204978 190204 204988 190260
rect 205044 190204 210056 190260
rect 375442 190092 375452 190148
rect 375508 190092 376236 190148
rect 376292 190092 380072 190148
rect 369880 189308 373772 189364
rect 373828 189308 373838 189364
rect 373062 188972 373100 189028
rect 373156 188972 373166 189028
rect 369880 188188 373884 188244
rect 373940 188188 373950 188244
rect 203410 187516 203420 187572
rect 203476 187516 204092 187572
rect 204148 187516 210056 187572
rect 369880 187068 371308 187124
rect 371364 187068 371374 187124
rect 375190 186508 375228 186564
rect 375284 186508 375294 186564
rect 369880 185948 373884 186004
rect 373940 185948 373950 186004
rect 204978 184940 204988 184996
rect 205044 184940 205884 184996
rect 205940 184940 208348 184996
rect 208292 184884 208348 184940
rect 208292 184828 210056 184884
rect 369880 184828 374444 184884
rect 374500 184828 374510 184884
rect 370066 184716 370076 184772
rect 370132 184716 380072 184772
rect 372754 184044 372764 184100
rect 372820 184044 375340 184100
rect 375396 184044 380072 184100
rect 369880 183708 373660 183764
rect 373716 183708 373726 183764
rect 371074 183372 371084 183428
rect 371140 183372 373884 183428
rect 373940 183372 380072 183428
rect 203410 182812 203420 182868
rect 203476 182812 204204 182868
rect 204260 182812 204270 182868
rect 370850 182700 370860 182756
rect 370916 182700 372204 182756
rect 372260 182700 380072 182756
rect 369880 182588 373100 182644
rect 373156 182588 373166 182644
rect 204194 182140 204204 182196
rect 204260 182140 210056 182196
rect 372866 182028 372876 182084
rect 372932 182028 379708 182084
rect 379764 182028 380072 182084
rect 369880 181468 374108 181524
rect 374164 181468 374174 181524
rect 371186 181356 371196 181412
rect 371252 181356 380072 181412
rect 374434 180684 374444 180740
rect 374500 180684 378700 180740
rect 378756 180684 380072 180740
rect 369880 180348 373660 180404
rect 373716 180348 373726 180404
rect 372530 180012 372540 180068
rect 372596 180012 373884 180068
rect 373940 180012 380072 180068
rect 204978 179452 204988 179508
rect 205044 179452 205772 179508
rect 205828 179452 210056 179508
rect 371074 179340 371084 179396
rect 371140 179340 373324 179396
rect 373380 179340 380072 179396
rect 439880 179340 442092 179396
rect 442148 179340 442158 179396
rect 369880 179228 373772 179284
rect 373828 179228 373838 179284
rect 595560 178948 597000 179144
rect 553522 178892 553532 178948
rect 553588 178920 597000 178948
rect 553588 178892 595672 178920
rect 377458 178668 377468 178724
rect 377524 178668 380072 178724
rect 439880 178668 441868 178724
rect 441924 178668 441934 178724
rect -960 178052 480 178136
rect 369880 178108 373996 178164
rect 374052 178108 374062 178164
rect -960 177996 7644 178052
rect 7700 177996 7710 178052
rect 375890 177996 375900 178052
rect 375956 177996 376236 178052
rect 376292 177996 380072 178052
rect 439880 177996 442428 178052
rect 442484 177996 442494 178052
rect -960 177912 480 177996
rect 372418 177324 372428 177380
rect 372484 177324 375788 177380
rect 375844 177324 380072 177380
rect 439880 177324 441868 177380
rect 441924 177324 441934 177380
rect 369880 176988 375900 177044
rect 375956 176988 375966 177044
rect 206658 176764 206668 176820
rect 206724 176764 208460 176820
rect 208516 176764 210056 176820
rect 370178 176652 370188 176708
rect 370244 176652 372316 176708
rect 372372 176652 380072 176708
rect 439880 176652 442540 176708
rect 442596 176652 442606 176708
rect 373650 176316 373660 176372
rect 373716 176316 374332 176372
rect 374388 176316 374398 176372
rect 379922 176316 379932 176372
rect 379988 176316 380100 176372
rect 380044 176036 380100 176316
rect 377458 175980 377468 176036
rect 377524 176008 380100 176036
rect 377524 175980 380072 176008
rect 439880 175980 442764 176036
rect 442820 175980 442830 176036
rect 369880 175868 373324 175924
rect 373380 175868 373390 175924
rect 377570 175308 377580 175364
rect 377636 175308 380072 175364
rect 439880 175308 442316 175364
rect 442372 175308 442382 175364
rect 372932 174860 373660 174916
rect 373716 174860 373726 174916
rect 372932 174804 372988 174860
rect 369880 174748 372988 174804
rect 371410 174636 371420 174692
rect 371476 174636 372316 174692
rect 372372 174636 372382 174692
rect 375554 174636 375564 174692
rect 375620 174636 380072 174692
rect 439880 174636 442652 174692
rect 442708 174636 442718 174692
rect 206882 174076 206892 174132
rect 206948 174076 208460 174132
rect 208516 174076 210056 174132
rect 373538 173964 373548 174020
rect 373604 173964 380072 174020
rect 439880 173964 440300 174020
rect 440356 173964 440366 174020
rect 369880 173628 371868 173684
rect 371924 173628 371934 173684
rect 370962 173292 370972 173348
rect 371028 173292 376012 173348
rect 376068 173292 380072 173348
rect 439880 173292 441980 173348
rect 442036 173292 442046 173348
rect 372642 173068 372652 173124
rect 372708 173068 373548 173124
rect 373604 173068 373614 173124
rect 379362 172620 379372 172676
rect 379428 172620 380072 172676
rect 439880 172620 442204 172676
rect 442260 172620 442270 172676
rect 369880 172508 375340 172564
rect 375396 172508 375406 172564
rect 376226 171948 376236 172004
rect 376292 171948 379484 172004
rect 379540 171948 380072 172004
rect 439880 171948 440636 172004
rect 440692 171948 440702 172004
rect 204978 171388 204988 171444
rect 205044 171388 210056 171444
rect 369880 171388 370076 171444
rect 370132 171388 370142 171444
rect 378914 171388 378924 171444
rect 378980 171388 379372 171444
rect 379428 171388 379438 171444
rect 374882 171276 374892 171332
rect 374948 171276 380072 171332
rect 439880 171276 443884 171332
rect 443940 171276 443950 171332
rect 370626 170604 370636 170660
rect 370692 170604 371756 170660
rect 371812 170604 380072 170660
rect 439880 170604 442092 170660
rect 442148 170604 442158 170660
rect 369880 170268 375564 170324
rect 375620 170268 375630 170324
rect 375106 169932 375116 169988
rect 375172 169932 380072 169988
rect 439880 169932 442876 169988
rect 442932 169932 442942 169988
rect 374882 169708 374892 169764
rect 374948 169708 376012 169764
rect 376068 169708 376078 169764
rect 439880 169260 443772 169316
rect 443828 169260 443838 169316
rect 369880 169148 370076 169204
rect 370132 169148 370142 169204
rect 201506 168700 201516 168756
rect 201572 168700 210056 168756
rect 199378 168028 199388 168084
rect 199444 168028 202300 168084
rect 202356 168028 202366 168084
rect 369880 168028 375564 168084
rect 375620 168028 375630 168084
rect 199154 167468 199164 167524
rect 199220 167468 202076 167524
rect 202132 167468 202142 167524
rect 377010 167244 377020 167300
rect 377076 167244 379708 167300
rect 379764 167244 380072 167300
rect 369880 166908 375676 166964
rect 375732 166908 375742 166964
rect 377122 166572 377132 166628
rect 377188 166572 380380 166628
rect 380436 166572 380446 166628
rect 20626 165676 20636 165732
rect 20692 165676 21756 165732
rect 21812 165676 21822 165732
rect 26674 165676 26684 165732
rect 26740 165676 26796 165732
rect 26852 165676 26862 165732
rect 28018 165676 28028 165732
rect 28084 165676 28476 165732
rect 28532 165676 28542 165732
rect 39638 165676 39676 165732
rect 39732 165676 39742 165732
rect 71698 165676 71708 165732
rect 71764 165676 72156 165732
rect 72212 165676 72222 165732
rect 82198 165676 82236 165732
rect 82292 165676 82302 165732
rect 84018 165676 84028 165732
rect 84084 165676 203308 165732
rect 203364 165676 203374 165732
rect 83794 165564 83804 165620
rect 83860 165564 84812 165620
rect 84868 165564 84878 165620
rect 120054 165564 120092 165620
rect 120148 165564 120158 165620
rect 122098 165564 122108 165620
rect 122164 165564 122556 165620
rect 122612 165564 122622 165620
rect 127558 165564 127596 165620
rect 127652 165564 127662 165620
rect 154018 165564 154028 165620
rect 154084 165564 154476 165620
rect 154532 165564 154542 165620
rect 182466 165564 182476 165620
rect 182532 165564 183036 165620
rect 183092 165564 183102 165620
rect 183810 165564 183820 165620
rect 183876 165564 184492 165620
rect 184548 165564 184558 165620
rect 184706 165564 184716 165620
rect 184772 165564 188972 165620
rect 189028 165564 189532 165620
rect 189588 165564 189598 165620
rect 192294 165564 192332 165620
rect 192388 165564 192398 165620
rect 183708 165452 200172 165508
rect 200228 165452 200238 165508
rect 183708 165396 183764 165452
rect 183698 165340 183708 165396
rect 183764 165340 183774 165396
rect 189522 164892 189532 164948
rect 189588 164892 196588 164948
rect 199266 164892 199276 164948
rect 199332 164892 202188 164948
rect 202244 164892 202254 164948
rect 196532 164724 196588 164892
rect 210028 164724 210084 166040
rect 377234 165900 377244 165956
rect 377300 165900 380072 165956
rect 369880 165788 375788 165844
rect 375844 165788 375854 165844
rect 595560 165732 597000 165928
rect 590482 165676 590492 165732
rect 590548 165704 597000 165732
rect 590548 165676 595672 165704
rect 370850 165228 370860 165284
rect 370916 165228 379820 165284
rect 379876 165228 380072 165284
rect 183250 164668 183260 164724
rect 183316 164668 184716 164724
rect 184772 164668 184782 164724
rect 196532 164668 210084 164724
rect 369880 164668 372204 164724
rect 372260 164668 372270 164724
rect 375330 164668 375340 164724
rect 375396 164668 377244 164724
rect 377300 164668 377310 164724
rect 92082 164556 92092 164612
rect 92148 164556 94892 164612
rect 94948 164556 94958 164612
rect 138786 164556 138796 164612
rect 138852 164556 160524 164612
rect 160580 164556 160590 164612
rect 171490 164556 171500 164612
rect 171556 164556 175532 164612
rect 175588 164556 175598 164612
rect 184034 164556 184044 164612
rect 184100 164556 199388 164612
rect 199444 164556 199454 164612
rect 374210 164556 374220 164612
rect 374276 164556 377356 164612
rect 377412 164556 380072 164612
rect 439880 164556 442652 164612
rect 442708 164556 442718 164612
rect 37874 164444 37884 164500
rect 37940 164444 172172 164500
rect 172228 164444 172238 164500
rect 189382 164444 189420 164500
rect 189476 164444 189486 164500
rect 191650 164444 191660 164500
rect 191716 164444 200844 164500
rect 200900 164444 200910 164500
rect 1474 164332 1484 164388
rect 1540 164332 46172 164388
rect 46228 164332 46238 164388
rect 179218 164332 179228 164388
rect 179284 164332 199164 164388
rect 199220 164332 199230 164388
rect 2930 164220 2940 164276
rect 2996 164220 45500 164276
rect 45556 164220 45566 164276
rect 128482 164220 128492 164276
rect 128548 164220 210476 164276
rect 210532 164220 210542 164276
rect 4834 164108 4844 164164
rect 4900 164108 44156 164164
rect 44212 164108 44222 164164
rect 120866 164108 120876 164164
rect 120932 164108 200508 164164
rect 200564 164108 200574 164164
rect -960 163828 480 164024
rect 38322 163996 38332 164052
rect 38388 163996 201852 164052
rect 201908 163996 201918 164052
rect 72370 163884 72380 163940
rect 72436 163884 165676 163940
rect 165732 163884 165742 163940
rect 181794 163884 181804 163940
rect 181860 163884 199276 163940
rect 199332 163884 199342 163940
rect 375666 163884 375676 163940
rect 375732 163884 378140 163940
rect 378196 163884 380072 163940
rect 439880 163884 442540 163940
rect 442596 163884 442606 163940
rect -960 163800 108332 163828
rect 392 163772 108332 163800
rect 108388 163772 108398 163828
rect 127138 163772 127148 163828
rect 127204 163772 201964 163828
rect 202020 163772 202030 163828
rect 45490 163548 45500 163604
rect 45556 163548 46396 163604
rect 46452 163548 46462 163604
rect 369880 163548 371980 163604
rect 372036 163548 372046 163604
rect 189410 163324 189420 163380
rect 189476 163324 210056 163380
rect 377458 163212 377468 163268
rect 377524 163212 377692 163268
rect 377748 163212 380072 163268
rect 439880 163212 440636 163268
rect 440692 163212 441980 163268
rect 442036 163212 442046 163268
rect 179218 163100 179228 163156
rect 179284 163100 179294 163156
rect 179228 163044 179284 163100
rect 44146 162988 44156 163044
rect 44212 162988 44940 163044
rect 44996 162988 45006 163044
rect 63970 162988 63980 163044
rect 64036 162988 144340 163044
rect 166114 162988 166124 163044
rect 166180 162988 179284 163044
rect 199266 162988 199276 163044
rect 199332 162988 204988 163044
rect 205044 162988 205054 163044
rect 371298 162988 371308 163044
rect 371364 162988 372092 163044
rect 372148 162988 372158 163044
rect 144284 162932 144340 162988
rect 20822 162876 20860 162932
rect 20916 162876 20926 162932
rect 27094 162876 27132 162932
rect 27188 162876 27198 162932
rect 91186 162876 91196 162932
rect 91252 162876 99932 162932
rect 99988 162876 99998 162932
rect 126214 162876 126252 162932
rect 126308 162876 126318 162932
rect 144284 162876 145180 162932
rect 145236 162876 146076 162932
rect 146132 162876 146142 162932
rect 165666 162876 165676 162932
rect 165732 162876 166236 162932
rect 166292 162876 170492 162932
rect 170548 162876 170558 162932
rect 191202 162876 191212 162932
rect 191268 162876 195804 162932
rect 195860 162876 195870 162932
rect 439852 162876 442316 162932
rect 442372 162876 442382 162932
rect 10882 162764 10892 162820
rect 10948 162764 45276 162820
rect 45332 162764 45342 162820
rect 91634 162764 91644 162820
rect 91700 162764 105196 162820
rect 105252 162764 105262 162820
rect 138338 162764 138348 162820
rect 138404 162764 157052 162820
rect 157108 162764 157118 162820
rect 183138 162764 183148 162820
rect 183204 162764 199276 162820
rect 199332 162764 199342 162820
rect 4498 162652 4508 162708
rect 4564 162652 26236 162708
rect 26292 162652 26302 162708
rect 82674 162652 82684 162708
rect 82740 162652 106652 162708
rect 106708 162652 106718 162708
rect 144452 162652 165228 162708
rect 165284 162652 203308 162708
rect 203364 162652 203374 162708
rect 1586 162540 1596 162596
rect 1652 162540 21308 162596
rect 21364 162540 21374 162596
rect 83122 162540 83132 162596
rect 83188 162540 104972 162596
rect 105028 162540 105038 162596
rect 2370 162428 2380 162484
rect 2436 162428 44380 162484
rect 44436 162428 47852 162484
rect 47908 162428 47918 162484
rect 71922 162428 71932 162484
rect 71988 162428 106876 162484
rect 106932 162428 106942 162484
rect 81778 162316 81788 162372
rect 81844 162316 108556 162372
rect 108612 162316 108622 162372
rect 64978 162204 64988 162260
rect 65044 162204 66108 162260
rect 66164 162204 143836 162260
rect 143892 162204 143902 162260
rect 144452 162148 144508 162652
rect 172386 162540 172396 162596
rect 172452 162540 206780 162596
rect 206836 162540 206846 162596
rect 373874 162540 373884 162596
rect 373940 162540 379820 162596
rect 379876 162540 380072 162596
rect 439852 162568 439908 162876
rect 171938 162428 171948 162484
rect 172004 162428 199164 162484
rect 199220 162428 199230 162484
rect 369880 162428 373548 162484
rect 373604 162428 373614 162484
rect 167906 162316 167916 162372
rect 167972 162316 208348 162372
rect 208404 162316 208414 162372
rect 182690 162204 182700 162260
rect 182756 162204 203644 162260
rect 203700 162204 203710 162260
rect 2258 162092 2268 162148
rect 2324 162092 44828 162148
rect 44884 162092 65212 162148
rect 65268 162092 144732 162148
rect 144788 162092 144798 162148
rect 146066 162092 146076 162148
rect 146132 162092 164780 162148
rect 164836 162092 199164 162148
rect 199220 162092 199230 162148
rect 137890 161980 137900 162036
rect 137956 161980 210140 162036
rect 210196 161980 210206 162036
rect 375666 161868 375676 161924
rect 375732 161868 380156 161924
rect 380212 161868 380222 161924
rect 439880 161868 440412 161924
rect 440468 161868 440478 161924
rect 143826 161532 143836 161588
rect 143892 161532 166124 161588
rect 166180 161532 166190 161588
rect 65650 161420 65660 161476
rect 65716 161420 144060 161476
rect 144116 161420 166236 161476
rect 166292 161420 166302 161476
rect 144274 161308 144284 161364
rect 144340 161308 166572 161364
rect 166628 161308 167916 161364
rect 167972 161308 167982 161364
rect 199238 161308 199276 161364
rect 199332 161308 199342 161364
rect 210578 161308 210588 161364
rect 210644 161308 210654 161364
rect 369880 161308 374612 161364
rect 17602 161196 17612 161252
rect 17668 161196 205100 161252
rect 205156 161196 205166 161252
rect 28466 161084 28476 161140
rect 28532 161084 210364 161140
rect 210420 161084 210430 161140
rect 210588 161028 210644 161308
rect 370188 161252 370244 161308
rect 374556 161252 374612 161308
rect 370178 161196 370188 161252
rect 370244 161196 370254 161252
rect 374556 161196 379036 161252
rect 379092 161196 380072 161252
rect 439880 161196 442204 161252
rect 442260 161196 442270 161252
rect 53666 160972 53676 161028
rect 53732 160972 210644 161028
rect 126914 160860 126924 160916
rect 126980 160860 177212 160916
rect 177268 160860 177278 160916
rect 128258 160748 128268 160804
rect 128324 160748 173852 160804
rect 173908 160748 173918 160804
rect 144834 160636 144844 160692
rect 144900 160636 146076 160692
rect 146132 160636 146142 160692
rect 181906 160636 181916 160692
rect 181972 160636 189084 160692
rect 189140 160636 189150 160692
rect 205090 160636 205100 160692
rect 205156 160636 210056 160692
rect 181458 160524 181468 160580
rect 181524 160524 205100 160580
rect 205156 160524 205166 160580
rect 377570 160524 377580 160580
rect 377636 160524 380072 160580
rect 439880 160524 442428 160580
rect 442484 160524 442494 160580
rect 65538 160412 65548 160468
rect 65604 160412 66332 160468
rect 66388 160412 143388 160468
rect 143444 160412 143454 160468
rect 156818 160412 156828 160468
rect 156884 160412 203532 160468
rect 203588 160412 203598 160468
rect 369880 160188 375228 160244
rect 375284 160188 376348 160244
rect 376404 160188 376414 160244
rect 377346 159852 377356 159908
rect 377412 159852 379596 159908
rect 379652 159852 380072 159908
rect 439880 159852 442092 159908
rect 442148 159852 442158 159908
rect 17602 159628 17612 159684
rect 17668 159628 17948 159684
rect 18004 159628 18014 159684
rect 143378 159628 143388 159684
rect 143444 159628 144284 159684
rect 144340 159628 144350 159684
rect 26002 159516 26012 159572
rect 26068 159516 181356 159572
rect 181412 159516 181422 159572
rect 377458 159516 377468 159572
rect 377524 159516 378812 159572
rect 378868 159516 378878 159572
rect 27794 159404 27804 159460
rect 27860 159404 167132 159460
rect 167188 159404 167198 159460
rect 171154 159180 171164 159236
rect 171220 159180 187292 159236
rect 187348 159180 187358 159236
rect 379474 159180 379484 159236
rect 379540 159180 380044 159236
rect 380100 159180 380110 159236
rect 439880 159180 442316 159236
rect 442372 159180 442382 159236
rect 182354 159068 182364 159124
rect 182420 159068 205212 159124
rect 205268 159068 205278 159124
rect 369880 159068 377468 159124
rect 377524 159068 377534 159124
rect 43474 158956 43484 159012
rect 43540 158956 65548 159012
rect 65604 158956 65614 159012
rect 127250 158956 127260 159012
rect 127316 158956 208796 159012
rect 208852 158956 208862 159012
rect 4274 158844 4284 158900
rect 4340 158844 160412 158900
rect 160468 158844 160478 158900
rect 172050 158844 172060 158900
rect 172116 158844 208572 158900
rect 208628 158844 208638 158900
rect 38098 158732 38108 158788
rect 38164 158732 200508 158788
rect 200564 158732 200574 158788
rect 439880 158508 441868 158564
rect 441924 158508 441934 158564
rect 379652 158060 380380 158116
rect 380436 158060 380446 158116
rect 379652 158004 379708 158060
rect 26002 157948 26012 158004
rect 26068 157948 26460 158004
rect 26516 157948 26526 158004
rect 181346 157948 181356 158004
rect 181412 157948 210056 158004
rect 369880 157948 379708 158004
rect 377010 157836 377020 157892
rect 377076 157836 377804 157892
rect 377860 157836 377870 157892
rect 372194 157724 372204 157780
rect 372260 157724 378252 157780
rect 378308 157724 378318 157780
rect 46610 157500 46620 157556
rect 46676 157500 63980 157556
rect 64036 157500 64046 157556
rect 118514 157500 118524 157556
rect 118580 157500 204204 157556
rect 204260 157500 204270 157556
rect 380044 157444 380100 157864
rect 439880 157836 441868 157892
rect 441924 157836 441934 157892
rect 43922 157388 43932 157444
rect 43988 157388 64988 157444
rect 65044 157388 65054 157444
rect 73042 157388 73052 157444
rect 73108 157388 89852 157444
rect 89908 157388 89918 157444
rect 116722 157388 116732 157444
rect 116788 157388 204540 157444
rect 204596 157388 204606 157444
rect 378242 157388 378252 157444
rect 378308 157388 380100 157444
rect 44930 157276 44940 157332
rect 44996 157276 66108 157332
rect 66164 157276 66174 157332
rect 82898 157276 82908 157332
rect 82964 157276 200172 157332
rect 200228 157276 200238 157332
rect 56914 157164 56924 157220
rect 56980 157164 206668 157220
rect 206724 157164 206734 157220
rect 377794 157164 377804 157220
rect 377860 157164 380072 157220
rect 27346 157052 27356 157108
rect 27412 157052 206668 157108
rect 206724 157052 206734 157108
rect 369880 156828 373996 156884
rect 374052 156828 374062 156884
rect 376338 156492 376348 156548
rect 376404 156492 379820 156548
rect 379876 156492 380072 156548
rect 145058 156268 145068 156324
rect 145124 156268 145740 156324
rect 145796 156268 145806 156324
rect 36866 156156 36876 156212
rect 36932 156156 191548 156212
rect 191604 156156 191614 156212
rect 377906 155820 377916 155876
rect 377972 155820 380072 155876
rect 369880 155708 379036 155764
rect 379092 155708 379102 155764
rect 45378 155596 45388 155652
rect 45444 155596 64876 155652
rect 64932 155596 64942 155652
rect 116834 155596 116844 155652
rect 116900 155596 207452 155652
rect 207508 155596 207518 155652
rect 27794 155484 27804 155540
rect 27860 155484 36876 155540
rect 36932 155484 36942 155540
rect 44370 155484 44380 155540
rect 44436 155484 65660 155540
rect 65716 155484 65726 155540
rect 89170 155484 89180 155540
rect 89236 155484 202300 155540
rect 202356 155484 202366 155540
rect 372194 155484 372204 155540
rect 372260 155484 379932 155540
rect 379988 155484 379998 155540
rect 18386 155372 18396 155428
rect 18452 155372 200396 155428
rect 200452 155372 200462 155428
rect 203298 155372 203308 155428
rect 203364 155372 207676 155428
rect 207732 155372 207742 155428
rect 373286 155372 373324 155428
rect 373380 155372 373390 155428
rect 375218 155372 375228 155428
rect 375284 155372 375788 155428
rect 375844 155372 375854 155428
rect 127698 155260 127708 155316
rect 127764 155260 129052 155316
rect 129108 155260 129118 155316
rect 191538 155260 191548 155316
rect 191604 155260 193004 155316
rect 193060 155260 210056 155316
rect 373426 155148 373436 155204
rect 373492 155148 377132 155204
rect 377188 155148 380072 155204
rect 372932 154700 380604 154756
rect 380660 154700 380670 154756
rect 372932 154644 372988 154700
rect 369880 154588 372988 154644
rect 377458 154476 377468 154532
rect 377524 154476 378700 154532
rect 378756 154476 380072 154532
rect 372754 153916 372764 153972
rect 372820 153916 376796 153972
rect 376852 153916 376862 153972
rect 120418 153804 120428 153860
rect 120484 153804 204092 153860
rect 204148 153804 204158 153860
rect 370738 153804 370748 153860
rect 370804 153804 377244 153860
rect 377300 153804 380072 153860
rect 118402 153692 118412 153748
rect 118468 153692 204428 153748
rect 204484 153692 204494 153748
rect 369880 153468 372988 153524
rect 372932 152852 372988 153468
rect 376786 153132 376796 153188
rect 376852 153132 377468 153188
rect 377524 153132 380072 153188
rect 38434 152796 38444 152852
rect 38500 152796 41132 152852
rect 41188 152796 193116 152852
rect 193172 152796 196588 152852
rect 372932 152796 379596 152852
rect 379652 152796 380100 152852
rect 196532 152628 196588 152796
rect 374546 152684 374556 152740
rect 374612 152684 376348 152740
rect 376404 152684 376414 152740
rect 377122 152684 377132 152740
rect 377188 152684 378924 152740
rect 378980 152684 378990 152740
rect 196532 152572 210056 152628
rect 380044 152488 380100 152796
rect 595560 152516 597000 152712
rect 543778 152460 543788 152516
rect 543844 152488 597000 152516
rect 543844 152460 595672 152488
rect 166226 152348 166236 152404
rect 166292 152348 202748 152404
rect 202804 152348 202814 152404
rect 369880 152348 377132 152404
rect 377188 152348 377198 152404
rect 128146 152236 128156 152292
rect 128212 152236 203420 152292
rect 203476 152236 203486 152292
rect 47842 152124 47852 152180
rect 47908 152124 65324 152180
rect 65380 152124 65390 152180
rect 74722 152124 74732 152180
rect 74788 152124 83468 152180
rect 83524 152124 83534 152180
rect 83682 152124 83692 152180
rect 83748 152124 108444 152180
rect 108500 152124 108510 152180
rect 116946 152124 116956 152180
rect 117012 152124 204652 152180
rect 204708 152124 204718 152180
rect 45042 152012 45052 152068
rect 45108 152012 67116 152068
rect 67172 152012 67182 152068
rect 71586 152012 71596 152068
rect 71652 152012 202524 152068
rect 202580 152012 202590 152068
rect 376338 151788 376348 151844
rect 376404 151788 380072 151844
rect 369880 151228 379148 151284
rect 379204 151228 379214 151284
rect 67106 151116 67116 151172
rect 67172 151116 142828 151172
rect 142884 151116 142894 151172
rect 374546 151116 374556 151172
rect 374612 151116 375452 151172
rect 375508 151116 375518 151172
rect 377234 151116 377244 151172
rect 377300 151116 379372 151172
rect 379428 151116 380072 151172
rect 380594 151004 380604 151060
rect 380660 151004 380670 151060
rect 182802 150780 182812 150836
rect 182868 150780 200284 150836
rect 200340 150780 200350 150836
rect 126802 150668 126812 150724
rect 126868 150668 202860 150724
rect 202916 150668 202926 150724
rect 69682 150556 69692 150612
rect 69748 150556 71148 150612
rect 71204 150556 208348 150612
rect 208404 150556 210084 150612
rect 26786 150444 26796 150500
rect 26852 150444 200284 150500
rect 200340 150444 200350 150500
rect 138646 150332 138684 150388
rect 138740 150332 138750 150388
rect 142818 150332 142828 150388
rect 142884 150332 144396 150388
rect 144452 150332 166236 150388
rect 166292 150332 166302 150388
rect 171602 150332 171612 150388
rect 171668 150332 200396 150388
rect 200452 150332 200462 150388
rect 210028 149912 210084 150556
rect 380604 150500 380660 151004
rect 379362 150444 379372 150500
rect 379428 150472 380660 150500
rect 379428 150444 380632 150472
rect 369880 150108 372988 150164
rect 373044 150108 373054 150164
rect -960 149716 480 149912
rect 380072 149800 380604 149828
rect 380044 149772 380604 149800
rect 380660 149772 380670 149828
rect -960 149688 103292 149716
rect 392 149660 103292 149688
rect 103348 149660 103358 149716
rect 380044 149604 380100 149772
rect 378700 149548 380100 149604
rect 83458 149436 83468 149492
rect 83524 149436 194460 149492
rect 194516 149436 194526 149492
rect 378700 149380 378756 149548
rect 89842 149324 89852 149380
rect 89908 149324 195692 149380
rect 195748 149324 206892 149380
rect 206948 149324 206958 149380
rect 378690 149324 378700 149380
rect 378756 149324 378766 149380
rect 64866 149212 64876 149268
rect 64932 149212 145740 149268
rect 145796 149212 164892 149268
rect 164948 149212 164958 149268
rect 65314 149100 65324 149156
rect 65380 149100 146076 149156
rect 146132 149100 146142 149156
rect 372978 149100 372988 149156
rect 373044 149100 379260 149156
rect 379316 149100 380072 149156
rect 66098 148988 66108 149044
rect 66164 148988 137452 149044
rect 137508 148988 137518 149044
rect 138002 148988 138012 149044
rect 138068 148988 139356 149044
rect 139412 148988 139422 149044
rect 142818 148988 142828 149044
rect 142884 148988 144172 149044
rect 144228 148988 165788 149044
rect 165844 148988 165854 149044
rect 369880 148988 378700 149044
rect 378756 148988 378766 149044
rect 2930 148876 2940 148932
rect 2996 148876 18732 148932
rect 18788 148876 18798 148932
rect 37538 148876 37548 148932
rect 37604 148876 54684 148932
rect 54740 148876 54750 148932
rect 65426 148876 65436 148932
rect 65492 148876 145628 148932
rect 145684 148876 145694 148932
rect 146066 148876 146076 148932
rect 146132 148876 165340 148932
rect 165396 148876 165406 148932
rect 189074 148876 189084 148932
rect 189140 148876 200732 148932
rect 200788 148876 200798 148932
rect 1586 148764 1596 148820
rect 1652 148764 25900 148820
rect 25956 148764 25966 148820
rect 46162 148764 46172 148820
rect 46228 148764 63980 148820
rect 64036 148764 145964 148820
rect 146020 148764 164556 148820
rect 164612 148764 164622 148820
rect 194450 148764 194460 148820
rect 194516 148764 206780 148820
rect 206836 148764 206846 148820
rect 2482 148652 2492 148708
rect 2548 148652 28140 148708
rect 28196 148652 28206 148708
rect 46386 148652 46396 148708
rect 46452 148652 64428 148708
rect 64484 148652 65436 148708
rect 65492 148652 65502 148708
rect 79762 148652 79772 148708
rect 79828 148652 81900 148708
rect 81956 148652 194236 148708
rect 194292 148652 206668 148708
rect 206724 148652 206734 148708
rect 88610 148540 88620 148596
rect 88676 148540 110236 148596
rect 110292 148540 110302 148596
rect 112354 148540 112364 148596
rect 112420 148540 125916 148596
rect 125972 148540 125982 148596
rect 137442 148540 137452 148596
rect 137508 148540 142828 148596
rect 142884 148540 142894 148596
rect 145618 148540 145628 148596
rect 145684 148540 149548 148596
rect 188626 148540 188636 148596
rect 188692 148540 199388 148596
rect 199444 148540 199454 148596
rect 137330 148428 137340 148484
rect 137396 148428 137676 148484
rect 137732 148428 137742 148484
rect 118710 148092 118748 148148
rect 118804 148092 118814 148148
rect 118290 147980 118300 148036
rect 118356 147980 119196 148036
rect 119252 147980 119262 148036
rect 149492 147924 149548 148540
rect 379138 148428 379148 148484
rect 379204 148428 379596 148484
rect 379652 148428 380072 148484
rect 164882 148204 164892 148260
rect 164948 148204 194908 148260
rect 194964 148204 194974 148260
rect 165330 148092 165340 148148
rect 165396 148092 199948 148148
rect 200004 148092 201180 148148
rect 201236 148092 201246 148148
rect 164546 147980 164556 148036
rect 164612 147980 200116 148036
rect 200060 147924 200116 147980
rect 45154 147868 45164 147924
rect 45220 147868 46620 147924
rect 46676 147868 46686 147924
rect 72006 147868 72044 147924
rect 72100 147868 72110 147924
rect 81414 147868 81452 147924
rect 81508 147868 81518 147924
rect 82338 147868 82348 147924
rect 82404 147868 83916 147924
rect 83972 147868 83982 147924
rect 117842 147868 117852 147924
rect 117908 147868 118636 147924
rect 118692 147868 118702 147924
rect 126354 147868 126364 147924
rect 126420 147868 126812 147924
rect 126868 147868 126878 147924
rect 149492 147868 164444 147924
rect 164500 147868 199892 147924
rect 200050 147868 200060 147924
rect 200116 147868 200956 147924
rect 201012 147868 201022 147924
rect 201180 147868 201628 147924
rect 201684 147868 202636 147924
rect 202692 147868 202702 147924
rect 369880 147868 370300 147924
rect 370356 147868 372820 147924
rect 376002 147868 376012 147924
rect 376068 147868 378924 147924
rect 378980 147868 378990 147924
rect 199836 147812 199892 147868
rect 201180 147812 201236 147868
rect 372764 147812 372820 147868
rect 199836 147756 201236 147812
rect 372754 147756 372764 147812
rect 372820 147756 380072 147812
rect 194898 147420 194908 147476
rect 194964 147420 199724 147476
rect 199780 147420 199790 147476
rect 155362 147308 155372 147364
rect 155428 147308 207788 147364
rect 207844 147308 207854 147364
rect 165778 147196 165788 147252
rect 165844 147196 199052 147252
rect 199108 147196 199118 147252
rect 206658 147196 206668 147252
rect 206724 147196 210056 147252
rect 150322 147084 150332 147140
rect 150388 147084 208124 147140
rect 208180 147084 208190 147140
rect 375218 147084 375228 147140
rect 375284 147084 380072 147140
rect 120306 146972 120316 147028
rect 120372 146972 204316 147028
rect 204372 146972 204382 147028
rect 369880 146748 372428 146804
rect 372484 146748 380212 146804
rect 380156 146244 380212 146748
rect 380146 146188 380156 146244
rect 380212 146188 380222 146244
rect 377122 145740 377132 145796
rect 377188 145740 380044 145796
rect 380100 145740 380110 145796
rect 369880 145628 375228 145684
rect 375284 145628 375452 145684
rect 375508 145628 375518 145684
rect 167906 145516 167916 145572
rect 167972 145516 200844 145572
rect 200900 145516 200910 145572
rect 121650 145404 121660 145460
rect 121716 145404 207900 145460
rect 207956 145404 207966 145460
rect 121762 145292 121772 145348
rect 121828 145292 208236 145348
rect 208292 145292 208302 145348
rect 378802 145068 378812 145124
rect 378868 145068 380604 145124
rect 380660 145068 380670 145124
rect 166226 144620 166236 144676
rect 166292 144620 166302 144676
rect 166236 144564 166292 144620
rect 166226 144508 166236 144564
rect 166292 144508 199052 144564
rect 199108 144508 199118 144564
rect 206770 144508 206780 144564
rect 206836 144508 210056 144564
rect 369880 144508 378812 144564
rect 378868 144508 378878 144564
rect 369880 143388 377244 143444
rect 377300 143388 379708 143444
rect 379764 143388 379774 143444
rect 369880 142268 376348 142324
rect 376404 142268 378812 142324
rect 378868 142268 378878 142324
rect 206882 141820 206892 141876
rect 206948 141820 210056 141876
rect 369880 141148 377468 141204
rect 377524 141148 380604 141204
rect 380660 141148 380670 141204
rect 377234 141036 377244 141092
rect 377300 141036 378812 141092
rect 378868 141036 378878 141092
rect 369880 140028 377244 140084
rect 377300 140028 377310 140084
rect 378242 139356 378252 139412
rect 378308 139356 378924 139412
rect 378980 139356 378990 139412
rect 595560 139300 597000 139496
rect 543890 139244 543900 139300
rect 543956 139272 597000 139300
rect 543956 139244 595672 139272
rect 204194 139132 204204 139188
rect 204260 139132 210056 139188
rect 369880 138908 377132 138964
rect 377188 138908 380492 138964
rect 380548 138908 380558 138964
rect 382498 137900 382508 137956
rect 382564 137900 383068 137956
rect 383124 137900 383134 137956
rect 369880 137788 378924 137844
rect 378980 137788 378990 137844
rect 372194 137452 372204 137508
rect 372260 137452 380044 137508
rect 380100 137452 380110 137508
rect 379026 137340 379036 137396
rect 379092 137340 396844 137396
rect 396900 137340 396910 137396
rect 442082 137340 442092 137396
rect 442148 137340 442652 137396
rect 442708 137340 442718 137396
rect 373986 137228 373996 137284
rect 374052 137228 397516 137284
rect 397572 137228 397582 137284
rect 408034 137228 408044 137284
rect 408100 137228 443660 137284
rect 443716 137228 443726 137284
rect 375442 137116 375452 137172
rect 375508 137116 393932 137172
rect 393988 137116 393998 137172
rect 408146 137116 408156 137172
rect 408212 137116 445340 137172
rect 445396 137116 445406 137172
rect 379586 137004 379596 137060
rect 379652 137004 442092 137060
rect 442148 137004 442158 137060
rect 374322 136892 374332 136948
rect 374388 136892 440412 136948
rect 440468 136892 440478 136948
rect 369880 136668 377916 136724
rect 377972 136668 379708 136724
rect 380370 136668 380380 136724
rect 380436 136668 385420 136724
rect 385476 136668 385486 136724
rect 379652 136612 379708 136668
rect 379652 136556 387212 136612
rect 387268 136556 387278 136612
rect 205986 136444 205996 136500
rect 206052 136444 210056 136500
rect 397506 136220 397516 136276
rect 397572 136220 408044 136276
rect 408100 136220 408110 136276
rect 396806 136108 396844 136164
rect 396900 136108 408156 136164
rect 408212 136108 408222 136164
rect 381378 135996 381388 136052
rect 381444 135996 382396 136052
rect 382452 135996 382462 136052
rect 377346 135884 377356 135940
rect 377412 135884 395724 135940
rect 395780 135884 395790 135940
rect 392 135800 7644 135828
rect -960 135772 7644 135800
rect 7700 135772 7710 135828
rect 373762 135772 373772 135828
rect 373828 135772 379708 135828
rect 382946 135772 382956 135828
rect 383012 135772 388108 135828
rect 388164 135772 388836 135828
rect -960 135576 480 135772
rect 379652 135604 379708 135772
rect 388780 135716 388836 135772
rect 396844 135716 396900 136108
rect 380706 135660 380716 135716
rect 380772 135660 380940 135716
rect 380996 135660 381006 135716
rect 382050 135660 382060 135716
rect 382116 135660 382172 135716
rect 382228 135660 382238 135716
rect 383590 135660 383628 135716
rect 383684 135660 383694 135716
rect 385382 135660 385420 135716
rect 385476 135660 385486 135716
rect 388770 135660 388780 135716
rect 388836 135660 388846 135716
rect 396834 135660 396844 135716
rect 396900 135660 396910 135716
rect 397478 135660 397516 135716
rect 397572 135660 397582 135716
rect 369880 135548 377020 135604
rect 377076 135548 377086 135604
rect 379652 135548 385532 135604
rect 385588 135548 385598 135604
rect 385746 135548 385756 135604
rect 385812 135548 442876 135604
rect 442932 135548 442942 135604
rect 378690 135436 378700 135492
rect 378756 135436 441980 135492
rect 442036 135436 442046 135492
rect 377906 135324 377916 135380
rect 377972 135324 442428 135380
rect 442484 135324 442494 135380
rect 379250 135212 379260 135268
rect 379316 135212 384748 135268
rect 384804 135212 384814 135268
rect 385522 135212 385532 135268
rect 385588 135212 440300 135268
rect 440356 135212 440366 135268
rect 380034 135100 380044 135156
rect 380100 135100 385756 135156
rect 385812 135100 385822 135156
rect 398178 135100 398188 135156
rect 398244 135100 445228 135156
rect 445284 135100 445294 135156
rect 379652 134988 441868 135044
rect 441924 134988 441934 135044
rect 379652 134820 379708 134988
rect 380370 134876 380380 134932
rect 380436 134876 398188 134932
rect 398244 134876 398254 134932
rect 377346 134764 377356 134820
rect 377412 134764 379708 134820
rect 381602 134764 381612 134820
rect 381668 134764 382732 134820
rect 382788 134764 382798 134820
rect 377010 134652 377020 134708
rect 377076 134652 385532 134708
rect 385588 134652 385598 134708
rect 374322 134540 374332 134596
rect 374388 134540 377356 134596
rect 377412 134540 377422 134596
rect 369880 134428 377356 134484
rect 377412 134428 377422 134484
rect 372306 134316 372316 134372
rect 372372 134316 372540 134372
rect 372596 134316 377916 134372
rect 377972 134316 377982 134372
rect 381266 134316 381276 134372
rect 381332 134316 388108 134372
rect 388164 134316 388174 134372
rect 396452 134316 442204 134372
rect 442260 134316 442270 134372
rect 379586 134204 379596 134260
rect 379652 134204 385644 134260
rect 385700 134204 386092 134260
rect 386148 134204 386158 134260
rect 379138 134092 379148 134148
rect 379204 134092 379708 134148
rect 380482 134092 380492 134148
rect 380548 134092 386428 134148
rect 386484 134092 386764 134148
rect 386820 134092 386830 134148
rect 379652 134036 379708 134092
rect 379652 133980 389452 134036
rect 389508 133980 389518 134036
rect 375890 133868 375900 133924
rect 375956 133868 386540 133924
rect 386596 133868 387436 133924
rect 387492 133868 387502 133924
rect 396452 133812 396508 134316
rect 419010 134204 419020 134260
rect 419076 134204 440524 134260
rect 440580 134204 440590 134260
rect 209682 133756 209692 133812
rect 209748 133756 210056 133812
rect 380258 133756 380268 133812
rect 380324 133756 396508 133812
rect 379250 133644 379260 133700
rect 379316 133644 442764 133700
rect 442820 133644 442830 133700
rect 373650 133532 373660 133588
rect 373716 133532 443772 133588
rect 443828 133532 443838 133588
rect 372932 133420 377580 133476
rect 377636 133420 394044 133476
rect 394100 133420 394110 133476
rect 372932 133364 372988 133420
rect 369880 133308 372988 133364
rect 390562 132748 390572 132804
rect 390628 132748 399868 132804
rect 372642 132636 372652 132692
rect 372708 132636 373100 132692
rect 373156 132636 376908 132692
rect 376964 132636 376974 132692
rect 381350 132636 381388 132692
rect 381444 132636 381454 132692
rect 381798 132636 381836 132692
rect 381892 132636 381902 132692
rect 383394 132636 383404 132692
rect 383460 132636 384524 132692
rect 384580 132636 384590 132692
rect 385868 132636 388108 132692
rect 383170 132524 383180 132580
rect 383236 132524 384076 132580
rect 384132 132524 384142 132580
rect 384300 132524 384748 132580
rect 384934 132524 384972 132580
rect 385028 132524 385038 132580
rect 385606 132524 385644 132580
rect 385700 132524 385710 132580
rect 384300 132468 384356 132524
rect 380034 132412 380044 132468
rect 380100 132412 381500 132468
rect 381556 132412 381566 132468
rect 381714 132412 381724 132468
rect 381780 132412 384356 132468
rect 384692 132468 384748 132524
rect 385868 132468 385924 132636
rect 386502 132524 386540 132580
rect 386596 132524 386606 132580
rect 384692 132412 385924 132468
rect 388052 132468 388108 132636
rect 399812 132580 399868 132748
rect 414866 132636 414876 132692
rect 414932 132636 418348 132692
rect 418404 132636 433692 132692
rect 433748 132636 433758 132692
rect 399812 132524 414316 132580
rect 414372 132524 414382 132580
rect 415650 132524 415660 132580
rect 415716 132524 439404 132580
rect 439460 132524 439470 132580
rect 388052 132412 412300 132468
rect 412356 132412 412366 132468
rect 414978 132412 414988 132468
rect 415044 132412 436828 132468
rect 436884 132412 436894 132468
rect 379026 132300 379036 132356
rect 379092 132300 379932 132356
rect 379988 132300 390572 132356
rect 390628 132300 390638 132356
rect 390786 132300 390796 132356
rect 390852 132300 412972 132356
rect 413028 132300 413038 132356
rect 417442 132300 417452 132356
rect 417508 132300 433580 132356
rect 433636 132300 433646 132356
rect 369880 132188 372988 132244
rect 376114 132188 376124 132244
rect 376180 132188 384356 132244
rect 384514 132188 384524 132244
rect 384580 132188 410956 132244
rect 411012 132188 411022 132244
rect 416322 132188 416332 132244
rect 416388 132188 432012 132244
rect 432068 132188 432078 132244
rect 372932 131572 372988 132188
rect 384300 132132 384356 132188
rect 377458 132076 377468 132132
rect 377524 132076 378028 132132
rect 378084 132076 381724 132132
rect 381780 132076 381790 132132
rect 384300 132076 410284 132132
rect 410340 132076 410350 132132
rect 416994 132076 417004 132132
rect 417060 132076 417900 132132
rect 417956 132076 431788 132132
rect 431844 132076 431854 132132
rect 377794 131964 377804 132020
rect 377860 131964 411628 132020
rect 411684 131964 411694 132020
rect 419234 131964 419244 132020
rect 419300 131964 431900 132020
rect 431956 131964 431966 132020
rect 377906 131852 377916 131908
rect 377972 131852 413644 131908
rect 413700 131852 413710 131908
rect 378578 131740 378588 131796
rect 378644 131740 379372 131796
rect 379428 131740 390796 131796
rect 390852 131740 390862 131796
rect 404226 131740 404236 131796
rect 404292 131740 440188 131796
rect 440244 131740 440254 131796
rect 377570 131628 377580 131684
rect 377636 131628 384524 131684
rect 384580 131628 384590 131684
rect 386390 131628 386428 131684
rect 386484 131628 386494 131684
rect 411506 131628 411516 131684
rect 411572 131628 415660 131684
rect 415716 131628 415726 131684
rect 372932 131516 377692 131572
rect 377748 131516 392252 131572
rect 392308 131516 392318 131572
rect 388210 131404 388220 131460
rect 388276 131404 389452 131460
rect 389508 131404 389518 131460
rect 414082 131180 414092 131236
rect 414148 131180 414988 131236
rect 415044 131180 415054 131236
rect 208002 131068 208012 131124
rect 208068 131068 210056 131124
rect 369880 131068 374220 131124
rect 374276 131068 377300 131124
rect 398150 131068 398188 131124
rect 398244 131068 398254 131124
rect 377244 131012 377300 131068
rect 371074 130956 371084 131012
rect 371140 130956 375228 131012
rect 375284 130956 375294 131012
rect 377244 130956 395836 131012
rect 395892 130956 395902 131012
rect 373762 130844 373772 130900
rect 373828 130844 374108 130900
rect 374164 130844 377580 130900
rect 377636 130844 377646 130900
rect 370514 130732 370524 130788
rect 370580 130732 376348 130788
rect 376404 130732 377804 130788
rect 377860 130732 377870 130788
rect 371970 130620 371980 130676
rect 372036 130620 372204 130676
rect 372260 130620 377916 130676
rect 377972 130620 377982 130676
rect 383058 130284 383068 130340
rect 383124 130284 429212 130340
rect 429268 130284 429278 130340
rect 376114 130172 376124 130228
rect 376180 130172 442316 130228
rect 442372 130172 442382 130228
rect 369880 129948 374332 130004
rect 374388 129948 374398 130004
rect 199042 129276 199052 129332
rect 199108 129276 200732 129332
rect 200788 129276 200798 129332
rect 375190 129276 375228 129332
rect 375284 129276 409612 129332
rect 409668 129276 409678 129332
rect 375330 129164 375340 129220
rect 375396 129164 376124 129220
rect 376180 129164 376190 129220
rect 388098 129164 388108 129220
rect 388164 129164 389788 129220
rect 389844 129164 389854 129220
rect 382162 129052 382172 129108
rect 382228 129052 404236 129108
rect 404292 129052 404302 129108
rect 384738 128940 384748 128996
rect 384804 128940 390012 128996
rect 390068 128940 390078 128996
rect 392466 128940 392476 128996
rect 392532 128940 414876 128996
rect 414932 128940 414942 128996
rect 369880 128828 375340 128884
rect 375396 128828 377132 128884
rect 377188 128828 377198 128884
rect 381378 128828 381388 128884
rect 381444 128828 388332 128884
rect 388388 128828 388398 128884
rect 408146 128828 408156 128884
rect 408212 128828 433468 128884
rect 433524 128828 433534 128884
rect 377906 128716 377916 128772
rect 377972 128716 442988 128772
rect 443044 128716 443054 128772
rect 377234 128604 377244 128660
rect 377300 128604 442652 128660
rect 442708 128604 442718 128660
rect 373314 128492 373324 128548
rect 373380 128492 443660 128548
rect 443716 128492 443726 128548
rect 209458 128380 209468 128436
rect 209524 128380 210056 128436
rect 374322 127932 374332 127988
rect 374388 127932 378028 127988
rect 378084 127932 381724 127988
rect 381780 127932 381790 127988
rect 369880 127708 374332 127764
rect 374388 127708 374398 127764
rect 370514 127596 370524 127652
rect 370580 127596 377916 127652
rect 377972 127596 377982 127652
rect 374322 127484 374332 127540
rect 374388 127484 377804 127540
rect 377860 127484 379708 127540
rect 379764 127484 379774 127540
rect 370738 127148 370748 127204
rect 370804 127148 373996 127204
rect 374052 127148 377244 127204
rect 377300 127148 377310 127204
rect 380370 127148 380380 127204
rect 380436 127148 411516 127204
rect 411572 127148 411582 127204
rect 408034 127036 408044 127092
rect 408100 127036 431788 127092
rect 431844 127036 431854 127092
rect 375890 126924 375900 126980
rect 375956 126924 441868 126980
rect 441924 126924 441934 126980
rect 373538 126812 373548 126868
rect 373604 126812 440412 126868
rect 440468 126812 440478 126868
rect 369880 126588 372988 126644
rect 373044 126588 373054 126644
rect 595560 126084 597000 126280
rect 572002 126028 572012 126084
rect 572068 126056 597000 126084
rect 572068 126028 595672 126056
rect 381938 125916 381948 125972
rect 382004 125916 442540 125972
rect 442596 125916 442606 125972
rect 204082 125692 204092 125748
rect 204148 125692 210056 125748
rect 369880 125468 370412 125524
rect 370468 125468 379484 125524
rect 379540 125468 379550 125524
rect 384514 125468 384524 125524
rect 384580 125468 393148 125524
rect 393204 125468 393214 125524
rect 392354 125356 392364 125412
rect 392420 125356 417900 125412
rect 417956 125356 417966 125412
rect 378690 125244 378700 125300
rect 378756 125244 419244 125300
rect 419300 125244 419310 125300
rect 372306 125132 372316 125188
rect 372372 125132 442316 125188
rect 442372 125132 442382 125188
rect 372978 124572 372988 124628
rect 373044 124572 377692 124628
rect 377748 124572 377758 124628
rect 373762 124460 373772 124516
rect 373828 124460 381948 124516
rect 382004 124460 382014 124516
rect 369880 124348 373212 124404
rect 373268 124348 373884 124404
rect 373940 124348 373950 124404
rect 377682 124348 377692 124404
rect 377748 124348 379820 124404
rect 379876 124348 379886 124404
rect 429202 124236 429212 124292
rect 429268 124236 443548 124292
rect 443604 124236 443614 124292
rect 382274 124012 382284 124068
rect 382340 124012 390572 124068
rect 390628 124012 390638 124068
rect 379138 123900 379148 123956
rect 379204 123900 414092 123956
rect 414148 123900 414158 123956
rect 379474 123788 379484 123844
rect 379540 123788 417452 123844
rect 417508 123788 417518 123844
rect 380258 123676 380268 123732
rect 380324 123676 419132 123732
rect 419188 123676 419198 123732
rect 371858 123564 371868 123620
rect 371924 123564 442204 123620
rect 442260 123564 442270 123620
rect 372082 123452 372092 123508
rect 372148 123452 442428 123508
rect 442484 123452 442494 123508
rect 369880 123228 375788 123284
rect 375844 123228 375854 123284
rect 209234 123004 209244 123060
rect 209300 123004 210056 123060
rect 372642 122220 372652 122276
rect 372708 122220 382172 122276
rect 382228 122220 382238 122276
rect 369880 122108 378140 122164
rect 378196 122108 378206 122164
rect 379250 121996 379260 122052
rect 379316 121996 416332 122052
rect 416388 121996 416398 122052
rect 392 121688 7532 121716
rect -960 121660 7532 121688
rect 7588 121660 7598 121716
rect -960 121464 480 121660
rect 369880 120988 372652 121044
rect 372708 120988 372718 121044
rect 378130 120988 378140 121044
rect 378196 120988 379596 121044
rect 379652 120988 379662 121044
rect 205874 120316 205884 120372
rect 205940 120316 210056 120372
rect 369880 119868 370300 119924
rect 370356 119868 373884 119924
rect 373940 119868 373950 119924
rect 369880 118748 374220 118804
rect 374276 118748 374286 118804
rect 204642 117628 204652 117684
rect 204708 117628 210056 117684
rect 369880 117628 380156 117684
rect 380212 117628 380222 117684
rect 369880 116508 372540 116564
rect 372596 116508 373772 116564
rect 373828 116508 373838 116564
rect 374210 116284 374220 116340
rect 374276 116284 379596 116340
rect 379652 116284 379662 116340
rect 374546 115612 374556 115668
rect 374612 115612 380072 115668
rect 369880 115388 370300 115444
rect 370356 115388 370366 115444
rect 207442 114940 207452 114996
rect 207508 114940 210056 114996
rect 373538 114940 373548 114996
rect 373604 114940 380380 114996
rect 380436 114940 380446 114996
rect 369880 114268 373548 114324
rect 373604 114268 373614 114324
rect 369880 113148 372316 113204
rect 372372 113148 372382 113204
rect 595560 112868 597000 113064
rect 546802 112812 546812 112868
rect 546868 112840 597000 112868
rect 546868 112812 595672 112840
rect 204530 112252 204540 112308
rect 204596 112252 210056 112308
rect 369880 112028 375340 112084
rect 375396 112028 375406 112084
rect 375330 111020 375340 111076
rect 375396 111020 375900 111076
rect 375956 111020 375966 111076
rect 369880 110908 373996 110964
rect 374052 110908 375676 110964
rect 375732 110908 375742 110964
rect 369880 109788 372428 109844
rect 372484 109788 374332 109844
rect 374388 109788 374398 109844
rect 204194 109564 204204 109620
rect 204260 109564 210056 109620
rect 369880 108668 373100 108724
rect 373156 108668 373166 108724
rect 372932 108164 372988 108668
rect 372932 108108 373884 108164
rect 373940 108108 373950 108164
rect -960 107492 480 107576
rect 369880 107548 374556 107604
rect 374612 107548 378700 107604
rect 378756 107548 378766 107604
rect -960 107436 7532 107492
rect 7588 107436 7598 107492
rect -960 107352 480 107436
rect 204418 106876 204428 106932
rect 204484 106876 210056 106932
rect 369880 106428 375900 106484
rect 375956 106428 380268 106484
rect 380324 106428 380334 106484
rect 369880 105308 374220 105364
rect 374276 105308 379484 105364
rect 379540 105308 379550 105364
rect 209122 104188 209132 104244
rect 209188 104188 210056 104244
rect 369880 104188 375452 104244
rect 375508 104188 376124 104244
rect 376180 104188 376190 104244
rect 200722 104076 200732 104132
rect 200788 104076 203196 104132
rect 203252 104076 203262 104132
rect 374322 104076 374332 104132
rect 374388 104076 379260 104132
rect 379316 104076 379326 104132
rect 369880 103068 374332 103124
rect 374388 103068 374398 103124
rect 369880 101948 377580 102004
rect 377636 101948 377646 102004
rect 204082 101500 204092 101556
rect 204148 101500 210056 101556
rect 369880 100828 377580 100884
rect 377636 100828 380380 100884
rect 380436 100828 380446 100884
rect 369880 99708 377356 99764
rect 377412 99708 377422 99764
rect 595560 99652 597000 99848
rect 590146 99596 590156 99652
rect 590212 99624 597000 99652
rect 590212 99596 595672 99624
rect 377346 99148 377356 99204
rect 377412 99148 379148 99204
rect 379204 99148 379214 99204
rect 370626 99036 370636 99092
rect 370692 99036 373100 99092
rect 373156 99036 373166 99092
rect 204306 98812 204316 98868
rect 204372 98812 210056 98868
rect 372082 98812 372092 98868
rect 372148 98812 376236 98868
rect 376292 98812 380072 98868
rect 369880 98588 374108 98644
rect 374164 98588 377020 98644
rect 377076 98588 377086 98644
rect 551842 98252 551852 98308
rect 551908 98252 590156 98308
rect 590212 98252 590222 98308
rect 373762 98140 373772 98196
rect 373828 98140 380072 98196
rect 372932 97692 376124 97748
rect 376180 97692 380380 97748
rect 380436 97692 380446 97748
rect 372932 97524 372988 97692
rect 203410 97468 203420 97524
rect 203476 97468 205044 97524
rect 369880 97468 372988 97524
rect 373090 97468 373100 97524
rect 373156 97468 380072 97524
rect 204988 97412 205044 97468
rect 204988 97356 207452 97412
rect 207508 97356 207518 97412
rect 380044 96628 380100 96824
rect 372530 96572 372540 96628
rect 372596 96572 376460 96628
rect 376516 96572 380100 96628
rect 369880 96348 377468 96404
rect 377524 96348 379260 96404
rect 379316 96348 379326 96404
rect 208226 96124 208236 96180
rect 208292 96124 210056 96180
rect 372418 96124 372428 96180
rect 372484 96124 380072 96180
rect 372530 95676 372540 95732
rect 372596 95676 373212 95732
rect 373268 95676 373278 95732
rect 373538 95676 373548 95732
rect 373604 95676 374108 95732
rect 374164 95676 374174 95732
rect 370850 95452 370860 95508
rect 370916 95452 372988 95508
rect 373044 95452 380072 95508
rect 369880 95228 376348 95284
rect 376404 95228 379484 95284
rect 379540 95228 379550 95284
rect 372194 95004 372204 95060
rect 372260 95004 379148 95060
rect 379204 95004 379214 95060
rect 376002 94780 376012 94836
rect 376068 94780 380072 94836
rect 372838 94444 372876 94500
rect 372932 94444 372942 94500
rect 370188 94220 372204 94276
rect 372260 94220 372270 94276
rect 372978 94220 372988 94276
rect 373044 94220 374948 94276
rect 370188 94164 370244 94220
rect 374892 94164 374948 94220
rect 369880 94108 370244 94164
rect 370402 94108 370412 94164
rect 370468 94108 373772 94164
rect 373828 94108 373838 94164
rect 374892 94108 380072 94164
rect 372838 93772 372876 93828
rect 372932 93772 372942 93828
rect 392 93464 4284 93492
rect -960 93436 4284 93464
rect 4340 93436 4350 93492
rect 207890 93436 207900 93492
rect 207956 93436 210056 93492
rect 371970 93436 371980 93492
rect 372036 93436 380072 93492
rect -960 93240 480 93436
rect 369880 92988 379036 93044
rect 379092 92988 379102 93044
rect 372194 92764 372204 92820
rect 372260 92764 380072 92820
rect 375778 92092 375788 92148
rect 375844 92092 380072 92148
rect 369880 91868 379372 91924
rect 379428 91868 379438 91924
rect 376002 91420 376012 91476
rect 376068 91420 380072 91476
rect 439880 91420 443772 91476
rect 443828 91420 443838 91476
rect 370962 90860 370972 90916
rect 371028 90860 373212 90916
rect 373268 90860 376404 90916
rect 376348 90804 376404 90860
rect 208114 90748 208124 90804
rect 208180 90748 210056 90804
rect 369880 90748 375228 90804
rect 375284 90748 376124 90804
rect 376180 90748 376190 90804
rect 376348 90748 380072 90804
rect 439880 90748 443660 90804
rect 443716 90748 443726 90804
rect 373762 90636 373772 90692
rect 373828 90636 376012 90692
rect 376068 90636 376078 90692
rect 370402 90076 370412 90132
rect 370468 90076 380072 90132
rect 439880 90076 447020 90132
rect 447076 90076 447086 90132
rect 369880 89628 373100 89684
rect 373156 89628 373166 89684
rect 370178 89404 370188 89460
rect 370244 89404 380072 89460
rect 439880 89404 442428 89460
rect 442484 89404 442494 89460
rect 369880 88508 376012 88564
rect 376068 88508 376078 88564
rect 380044 88340 380100 88760
rect 439880 88732 443548 88788
rect 443604 88732 443614 88788
rect 370178 88284 370188 88340
rect 370244 88284 370860 88340
rect 370916 88284 380100 88340
rect 207778 88060 207788 88116
rect 207844 88060 210056 88116
rect 375666 88060 375676 88116
rect 375732 88060 380072 88116
rect 439880 88060 445340 88116
rect 445396 88060 445406 88116
rect 369880 87388 370860 87444
rect 370916 87388 370926 87444
rect 372866 87388 372876 87444
rect 372932 87388 374780 87444
rect 374836 87388 380072 87444
rect 439880 87388 442316 87444
rect 442372 87388 442382 87444
rect 374434 87276 374444 87332
rect 374500 87276 374510 87332
rect 374444 87220 374500 87276
rect 374444 87164 376460 87220
rect 376516 87164 380100 87220
rect 380044 86744 380100 87164
rect 439880 86716 450268 86772
rect 450324 86716 450334 86772
rect 595560 86436 597000 86632
rect 556882 86380 556892 86436
rect 556948 86408 597000 86436
rect 556948 86380 595672 86408
rect 369880 86268 373772 86324
rect 373828 86268 373838 86324
rect 371074 86044 371084 86100
rect 371140 86044 371308 86100
rect 371364 86044 380072 86100
rect 439880 86044 446908 86100
rect 446964 86044 446974 86100
rect 372642 85596 372652 85652
rect 372708 85596 374444 85652
rect 374500 85596 374510 85652
rect 205762 85372 205772 85428
rect 205828 85372 210056 85428
rect 371186 85372 371196 85428
rect 371252 85372 373100 85428
rect 373156 85372 380072 85428
rect 439880 85372 448588 85428
rect 448644 85372 448654 85428
rect 369880 85148 372988 85204
rect 373044 85148 373054 85204
rect 377234 84700 377244 84756
rect 377300 84700 377356 84756
rect 377412 84700 380072 84756
rect 439880 84700 448588 84756
rect 448644 84700 448654 84756
rect 369880 84028 372988 84084
rect 373044 84028 373054 84084
rect 373314 84028 373324 84084
rect 373380 84028 374444 84084
rect 374500 84028 380072 84084
rect 439880 84028 441980 84084
rect 442036 84028 442046 84084
rect 372082 83356 372092 83412
rect 372148 83356 380072 83412
rect 439880 83356 440300 83412
rect 440356 83356 440366 83412
rect 369880 82908 376460 82964
rect 376516 82908 376526 82964
rect 199042 82684 199052 82740
rect 199108 82684 210056 82740
rect 375778 82684 375788 82740
rect 375844 82684 380072 82740
rect 439880 82684 440300 82740
rect 440356 82684 440366 82740
rect 379586 82012 379596 82068
rect 379652 82012 380072 82068
rect 439880 82012 440188 82068
rect 440244 82012 440254 82068
rect 369880 81788 378812 81844
rect 378868 81788 378878 81844
rect 375442 81340 375452 81396
rect 375508 81340 380072 81396
rect 439880 81340 440412 81396
rect 440468 81340 440478 81396
rect 371084 80780 378812 80836
rect 378868 80780 378878 80836
rect 371084 80724 371140 80780
rect 369880 80668 371140 80724
rect 372642 80668 372652 80724
rect 372708 80668 380072 80724
rect 439880 80668 442204 80724
rect 442260 80668 442270 80724
rect 201170 79996 201180 80052
rect 201236 79996 210056 80052
rect 372530 79996 372540 80052
rect 372596 79996 380072 80052
rect 439880 79996 445228 80052
rect 445284 79996 445294 80052
rect 369880 79548 378812 79604
rect 378868 79548 378878 79604
rect 392 79352 4172 79380
rect -960 79324 4172 79352
rect 4228 79324 4238 79380
rect 377570 79324 377580 79380
rect 377636 79324 380072 79380
rect 439880 79324 440412 79380
rect 440468 79324 440478 79380
rect -960 79128 480 79324
rect 370066 78652 370076 78708
rect 370132 78652 380072 78708
rect 439880 78652 446908 78708
rect 446964 78652 446974 78708
rect 369880 78428 378812 78484
rect 378868 78428 378878 78484
rect 370290 77980 370300 78036
rect 370356 77980 380072 78036
rect 439880 77980 445564 78036
rect 445620 77980 445630 78036
rect 207666 77308 207676 77364
rect 207732 77308 210056 77364
rect 369880 77308 378812 77364
rect 378868 77308 378878 77364
rect 379474 77308 379484 77364
rect 379540 77308 380072 77364
rect 439880 77308 445452 77364
rect 445508 77308 445518 77364
rect 375554 76636 375564 76692
rect 375620 76636 380072 76692
rect 439880 76636 441868 76692
rect 441924 76636 441934 76692
rect 369880 76188 379596 76244
rect 379652 76188 379662 76244
rect 376226 75964 376236 76020
rect 376292 75964 380072 76020
rect 439880 75964 443772 76020
rect 443828 75964 443838 76020
rect 380146 75292 380156 75348
rect 380212 75292 380222 75348
rect 439880 75292 443660 75348
rect 443716 75292 443726 75348
rect 369880 75068 379596 75124
rect 379652 75068 379662 75124
rect 202738 74620 202748 74676
rect 202804 74620 210056 74676
rect 372530 74620 372540 74676
rect 372596 74620 380072 74676
rect 372932 74060 378588 74116
rect 378644 74060 378654 74116
rect 372932 74004 372988 74060
rect 369880 73948 372988 74004
rect 377682 73948 377692 74004
rect 377748 73948 380072 74004
rect 377794 73276 377804 73332
rect 377860 73276 380072 73332
rect 595560 73220 597000 73416
rect 545122 73164 545132 73220
rect 545188 73192 597000 73220
rect 545188 73164 595672 73192
rect 369880 72828 378812 72884
rect 378868 72828 378878 72884
rect 370290 72604 370300 72660
rect 370356 72604 380072 72660
rect 374434 72156 374444 72212
rect 374500 72156 376460 72212
rect 376516 72156 376526 72212
rect 199266 71932 199276 71988
rect 199332 71932 210056 71988
rect 377122 71932 377132 71988
rect 377188 71932 380072 71988
rect 369880 71708 377580 71764
rect 377636 71708 377646 71764
rect 374098 71260 374108 71316
rect 374164 71260 380072 71316
rect 372932 70700 373212 70756
rect 373268 70700 373278 70756
rect 372932 70644 372988 70700
rect 369880 70588 372988 70644
rect 377906 70588 377916 70644
rect 377972 70588 380072 70644
rect 509880 70588 513212 70644
rect 513268 70588 513278 70644
rect 376226 70476 376236 70532
rect 376292 70476 377244 70532
rect 377300 70476 377310 70532
rect 372306 69916 372316 69972
rect 372372 69916 380072 69972
rect 439880 69916 442876 69972
rect 442932 69916 442942 69972
rect 457762 69916 457772 69972
rect 457828 69916 460040 69972
rect 509880 69916 512428 69972
rect 512484 69916 512494 69972
rect 369880 69468 373772 69524
rect 373828 69468 373838 69524
rect 200834 69244 200844 69300
rect 200900 69244 210056 69300
rect 375890 69244 375900 69300
rect 375956 69244 380072 69300
rect 439880 69244 441980 69300
rect 442036 69244 442046 69300
rect 509880 69244 512540 69300
rect 512596 69244 512606 69300
rect 375666 68572 375676 68628
rect 375732 68572 380072 68628
rect 439880 68572 442764 68628
rect 442820 68572 442830 68628
rect 509880 68572 530012 68628
rect 530068 68572 530078 68628
rect 369880 68348 372092 68404
rect 372148 68348 372158 68404
rect 372418 67900 372428 67956
rect 372484 67900 380072 67956
rect 372932 67452 380604 67508
rect 380660 67452 380670 67508
rect 372932 67284 372988 67452
rect 369880 67228 372988 67284
rect 373874 67228 373884 67284
rect 373940 67228 380072 67284
rect 199714 66556 199724 66612
rect 199780 66556 210056 66612
rect 377346 66556 377356 66612
rect 377412 66556 380072 66612
rect 439880 66556 441868 66612
rect 441924 66556 441934 66612
rect 369880 66108 379932 66164
rect 379988 66108 379998 66164
rect 377010 65884 377020 65940
rect 377076 65884 380072 65940
rect 379810 65548 379820 65604
rect 379876 65548 379932 65604
rect 379988 65548 379998 65604
rect 392 65240 4172 65268
rect -960 65212 4172 65240
rect 4228 65212 4238 65268
rect 377570 65212 377580 65268
rect 377636 65212 380072 65268
rect -960 65016 480 65212
rect 369880 64988 377580 65044
rect 377636 64988 377646 65044
rect 374546 64540 374556 64596
rect 374612 64540 380072 64596
rect 202626 63868 202636 63924
rect 202692 63868 210056 63924
rect 369880 63868 377580 63924
rect 377636 63868 377646 63924
rect 375890 63196 375900 63252
rect 375956 63196 380072 63252
rect 369880 62748 377580 62804
rect 377636 62748 377646 62804
rect 374210 62524 374220 62580
rect 374276 62524 380072 62580
rect 375442 61852 375452 61908
rect 375508 61852 380072 61908
rect 369880 61628 372428 61684
rect 372484 61628 372494 61684
rect 200946 61180 200956 61236
rect 201012 61180 210056 61236
rect 374322 61180 374332 61236
rect 374388 61180 380072 61236
rect 369880 60508 373100 60564
rect 373156 60508 373166 60564
rect 595560 60004 597000 60200
rect 544002 59948 544012 60004
rect 544068 59976 597000 60004
rect 544068 59948 595672 59976
rect 369880 59388 374444 59444
rect 374500 59388 374510 59444
rect 207666 58492 207676 58548
rect 207732 58492 210056 58548
rect 369880 58268 373324 58324
rect 373380 58268 373390 58324
rect 207442 57820 207452 57876
rect 207508 57820 209916 57876
rect 209972 57820 209982 57876
rect 369880 57148 374780 57204
rect 374836 57148 374846 57204
rect 369880 56028 371308 56084
rect 371364 56028 371374 56084
rect 202514 55804 202524 55860
rect 202580 55804 210056 55860
rect 369880 54908 376348 54964
rect 376404 54908 376414 54964
rect 369880 53788 377132 53844
rect 377188 53788 377198 53844
rect 207442 53116 207452 53172
rect 207508 53116 210056 53172
rect 369880 52668 374556 52724
rect 374612 52668 376236 52724
rect 376292 52668 376302 52724
rect 372932 52108 376236 52164
rect 376292 52108 376302 52164
rect 372932 51604 372988 52108
rect 369880 51548 370412 51604
rect 370468 51548 372988 51604
rect 130 51212 140 51268
rect 196 51212 532 51268
rect 476 51156 532 51212
rect 392 51128 532 51156
rect -960 51100 532 51128
rect -960 50904 480 51100
rect 207554 50428 207564 50484
rect 207620 50428 210056 50484
rect 394034 47964 394044 48020
rect 394100 47964 403564 48020
rect 403620 47964 403630 48020
rect 379362 47852 379372 47908
rect 379428 47852 417676 47908
rect 417732 47852 417742 47908
rect 208114 47740 208124 47796
rect 208180 47740 210056 47796
rect 394818 46956 394828 47012
rect 394884 46956 457772 47012
rect 457828 46956 457838 47012
rect 595560 46788 597000 46984
rect 590594 46732 590604 46788
rect 590660 46760 597000 46788
rect 590660 46732 595672 46760
rect 379250 46284 379260 46340
rect 379316 46284 396844 46340
rect 396900 46284 396910 46340
rect 379474 46172 379484 46228
rect 379540 46172 398188 46228
rect 398244 46172 398254 46228
rect 380482 45948 380492 46004
rect 380548 45948 393820 46004
rect 393876 45948 393886 46004
rect 385522 45836 385532 45892
rect 385588 45836 393652 45892
rect 381350 45724 381388 45780
rect 381444 45724 381454 45780
rect 381602 45724 381612 45780
rect 381668 45724 382060 45780
rect 382116 45724 382126 45780
rect 383058 45724 383068 45780
rect 383124 45724 384076 45780
rect 384132 45724 384142 45780
rect 384738 45724 384748 45780
rect 384804 45724 385644 45780
rect 385700 45724 385710 45780
rect 388098 45724 388108 45780
rect 388164 45724 389788 45780
rect 389844 45724 389854 45780
rect 379652 45612 390460 45668
rect 390516 45612 390526 45668
rect 379652 45556 379708 45612
rect 378802 45500 378812 45556
rect 378868 45500 379708 45556
rect 381490 45500 381500 45556
rect 381556 45500 382732 45556
rect 382788 45500 382798 45556
rect 383814 45500 383852 45556
rect 383908 45500 383918 45556
rect 384934 45500 384972 45556
rect 385028 45500 385038 45556
rect 386390 45500 386428 45556
rect 386484 45500 386494 45556
rect 386950 45500 386988 45556
rect 387044 45500 387054 45556
rect 388322 45500 388332 45556
rect 388388 45500 389004 45556
rect 389060 45500 389070 45556
rect 391458 45500 391468 45556
rect 391524 45500 391916 45556
rect 391972 45500 391982 45556
rect 393596 45444 393652 45836
rect 396806 45724 396844 45780
rect 396900 45724 396910 45780
rect 398150 45724 398188 45780
rect 398244 45724 398254 45780
rect 403526 45724 403564 45780
rect 403620 45724 403630 45780
rect 417638 45724 417676 45780
rect 417732 45724 417742 45780
rect 397842 45612 397852 45668
rect 397908 45612 418348 45668
rect 418404 45612 418414 45668
rect 393810 45500 393820 45556
rect 393876 45500 412972 45556
rect 413028 45500 413038 45556
rect 388098 45388 388108 45444
rect 388164 45388 388332 45444
rect 388388 45388 388398 45444
rect 393596 45388 407596 45444
rect 407652 45388 407662 45444
rect 199154 45276 199164 45332
rect 199220 45276 512540 45332
rect 512596 45276 512606 45332
rect 386082 45164 386092 45220
rect 386148 45164 389900 45220
rect 389956 45164 389966 45220
rect 392242 45164 392252 45220
rect 392308 45164 392318 45220
rect 395714 45164 395724 45220
rect 395780 45164 405580 45220
rect 405636 45164 405646 45220
rect 392252 45108 392308 45164
rect 392252 45052 402892 45108
rect 402948 45052 402958 45108
rect 408212 45052 416332 45108
rect 416388 45052 416398 45108
rect 485538 45052 485548 45108
rect 485604 45052 573692 45108
rect 573748 45052 573758 45108
rect 408212 44996 408268 45052
rect 380594 44940 380604 44996
rect 380660 44940 408268 44996
rect 378914 44828 378924 44884
rect 378980 44828 410956 44884
rect 411012 44828 411022 44884
rect 375554 44716 375564 44772
rect 375620 44716 406252 44772
rect 406308 44716 406318 44772
rect 380258 44604 380268 44660
rect 380324 44604 423052 44660
rect 423108 44604 423118 44660
rect 370066 44380 370076 44436
rect 370132 44380 376348 44436
rect 385746 44380 385756 44436
rect 385812 44380 406924 44436
rect 406980 44380 406990 44436
rect 376292 44212 376348 44380
rect 379138 44268 379148 44324
rect 379204 44268 398860 44324
rect 398916 44268 398926 44324
rect 376292 44156 385756 44212
rect 385812 44156 385822 44212
rect 395826 43596 395836 43652
rect 395892 43596 400876 43652
rect 400932 43596 400942 43652
rect 419654 43596 419692 43652
rect 419748 43596 419758 43652
rect 420354 43596 420364 43652
rect 420420 43596 429212 43652
rect 429268 43596 429278 43652
rect 484866 43596 484876 43652
rect 484932 43596 540092 43652
rect 540148 43596 540158 43652
rect 394146 43484 394156 43540
rect 394212 43484 404236 43540
rect 404292 43484 404302 43540
rect 415650 43484 415660 43540
rect 415716 43484 431788 43540
rect 431844 43484 431854 43540
rect 484194 43484 484204 43540
rect 484260 43484 511532 43540
rect 511588 43484 511598 43540
rect 390562 43372 390572 43428
rect 390628 43372 421036 43428
rect 421092 43372 421102 43428
rect 393922 43260 393932 43316
rect 393988 43260 422380 43316
rect 422436 43260 422446 43316
rect 379362 43148 379372 43204
rect 379428 43148 400204 43204
rect 400260 43148 400270 43204
rect 416994 43148 417004 43204
rect 417060 43148 433468 43204
rect 433524 43148 433534 43204
rect 378802 43036 378812 43092
rect 378868 43036 414316 43092
rect 414372 43036 414382 43092
rect 380370 42924 380380 42980
rect 380436 42924 396172 42980
rect 396228 42924 396238 42980
rect 396386 42924 396396 42980
rect 396452 42924 413644 42980
rect 413700 42924 413710 42980
rect 378690 42812 378700 42868
rect 378756 42812 410284 42868
rect 410340 42812 410350 42868
rect 379026 42700 379036 42756
rect 379092 42700 399532 42756
rect 399588 42700 399598 42756
rect 374546 41916 374556 41972
rect 374612 41916 512428 41972
rect 512484 41916 512494 41972
rect 372754 41804 372764 41860
rect 372820 41804 423724 41860
rect 423780 41804 423790 41860
rect 387202 41692 387212 41748
rect 387268 41692 409612 41748
rect 409668 41692 409678 41748
rect 379810 40236 379820 40292
rect 379876 40236 408940 40292
rect 408996 40236 409006 40292
rect -960 36820 480 37016
rect -960 36792 110012 36820
rect 392 36764 110012 36792
rect 110068 36764 110078 36820
rect 595560 33684 597000 33768
rect 550274 33628 550284 33684
rect 550340 33628 597000 33684
rect 595560 33544 597000 33628
rect 539896 32844 543452 32900
rect 543508 32844 543518 32900
rect 539896 31724 563612 31780
rect 563668 31724 563678 31780
rect 539896 30604 565292 30660
rect 565348 30604 565358 30660
rect 539896 29484 550172 29540
rect 550228 29484 550238 29540
rect 544226 29372 544236 29428
rect 544292 29372 587132 29428
rect 587188 29372 587198 29428
rect 539896 28364 555212 28420
rect 555268 28364 555278 28420
rect 539896 27244 544236 27300
rect 544292 27244 544302 27300
rect 539896 26124 543564 26180
rect 543620 26124 543630 26180
rect 539896 25004 543676 25060
rect 543732 25004 543742 25060
rect 544338 24332 544348 24388
rect 544404 24332 590492 24388
rect 590548 24332 590558 24388
rect 539896 23884 560252 23940
rect 560308 23884 560318 23940
rect 18 22988 28 23044
rect 84 22988 532 23044
rect 476 22932 532 22988
rect 392 22904 532 22932
rect -960 22876 532 22904
rect -960 22680 480 22876
rect 539896 22764 548492 22820
rect 548548 22764 548558 22820
rect 539896 21644 553532 21700
rect 553588 21644 553598 21700
rect 539896 20524 544348 20580
rect 544404 20524 544414 20580
rect 595560 20356 597000 20552
rect 591266 20300 591276 20356
rect 591332 20328 597000 20356
rect 591332 20300 595672 20328
rect 539896 19404 543788 19460
rect 543844 19404 543854 19460
rect 548482 19292 548492 19348
rect 548548 19292 591276 19348
rect 591332 19292 591342 19348
rect 539896 18284 543900 18340
rect 543956 18284 543966 18340
rect 539896 17164 572012 17220
rect 572068 17164 572078 17220
rect 539896 16044 546812 16100
rect 546868 16044 546878 16100
rect 539896 14924 551852 14980
rect 551908 14924 551918 14980
rect 539896 13804 556892 13860
rect 556948 13804 556958 13860
rect 539896 12684 545132 12740
rect 545188 12684 545198 12740
rect 544338 12572 544348 12628
rect 544404 12572 590604 12628
rect 590660 12572 590670 12628
rect 539896 11564 544012 11620
rect 544068 11564 544078 11620
rect 539896 10444 544348 10500
rect 544404 10444 544414 10500
rect 539896 9324 550284 9380
rect 550340 9324 550350 9380
rect 392 8792 4284 8820
rect -960 8764 4284 8792
rect 4340 8764 4350 8820
rect -960 8568 480 8764
rect 539896 8204 548492 8260
rect 548548 8204 548558 8260
rect 595560 7140 597000 7336
rect 539896 7112 597000 7140
rect 539896 7084 595672 7112
rect 396386 5516 396396 5572
rect 396452 5516 437612 5572
rect 437668 5516 437678 5572
rect 483074 5516 483084 5572
rect 483140 5516 523516 5572
rect 523572 5516 523582 5572
rect 401314 5404 401324 5460
rect 401380 5404 443548 5460
rect 443604 5404 443614 5460
rect 462466 5404 462476 5460
rect 462532 5404 506380 5460
rect 506436 5404 506446 5460
rect 382498 5292 382508 5348
rect 382564 5292 408268 5348
rect 420130 5292 420140 5348
rect 420196 5292 465724 5348
rect 465780 5292 465790 5348
rect 474338 5292 474348 5348
rect 474404 5292 533036 5348
rect 533092 5292 533102 5348
rect 353602 5180 353612 5236
rect 353668 5180 386652 5236
rect 386708 5180 386718 5236
rect 408212 5124 408268 5292
rect 429538 5180 429548 5236
rect 429604 5180 478156 5236
rect 478212 5180 478222 5236
rect 493154 5180 493164 5236
rect 493220 5180 555884 5236
rect 555940 5180 555950 5236
rect 15362 5068 15372 5124
rect 15428 5068 47852 5124
rect 47908 5068 47918 5124
rect 68684 5068 91756 5124
rect 91812 5068 91822 5124
rect 333218 5068 333228 5124
rect 333284 5068 361676 5124
rect 361732 5068 361742 5124
rect 367714 5068 367724 5124
rect 367780 5068 403116 5124
rect 403172 5068 403182 5124
rect 408212 5068 420364 5124
rect 420420 5068 420430 5124
rect 434242 5068 434252 5124
rect 434308 5068 442820 5124
rect 442950 5068 442988 5124
rect 443044 5068 443054 5124
rect 443212 5068 482860 5124
rect 482916 5068 482926 5124
rect 495394 5068 495404 5124
rect 495460 5068 498988 5124
rect 499044 5068 499054 5124
rect 507266 5068 507276 5124
rect 507332 5068 573020 5124
rect 573076 5068 573086 5124
rect 68684 5012 68740 5068
rect 442764 5012 442820 5068
rect 443212 5012 443268 5068
rect 28690 4956 28700 5012
rect 28756 4956 58940 5012
rect 58996 4956 59006 5012
rect 68674 4956 68684 5012
rect 68740 4956 68750 5012
rect 73042 4956 73052 5012
rect 73108 4956 84812 5012
rect 84868 4956 84878 5012
rect 85810 4956 85820 5012
rect 85876 4956 105980 5012
rect 106036 4956 106046 5012
rect 106754 4956 106764 5012
rect 106820 4956 122668 5012
rect 122724 4956 122734 5012
rect 123890 4956 123900 5012
rect 123956 4956 136556 5012
rect 136612 4956 136622 5012
rect 139122 4956 139132 5012
rect 139188 4956 149548 5012
rect 149604 4956 149614 5012
rect 160066 4956 160076 5012
rect 160132 4956 166348 5012
rect 166404 4956 166414 5012
rect 294690 4956 294700 5012
rect 294756 4956 314188 5012
rect 314244 4956 314254 5012
rect 316642 4956 316652 5012
rect 316708 4956 340732 5012
rect 340788 4956 340798 5012
rect 341730 4956 341740 5012
rect 341796 4956 371308 5012
rect 371364 4956 371374 5012
rect 393026 4956 393036 5012
rect 393092 4956 434364 5012
rect 434420 4956 434430 5012
rect 442764 4956 443268 5012
rect 454626 4956 454636 5012
rect 454692 4956 508284 5012
rect 508340 4956 508350 5012
rect 515666 4956 515676 5012
rect 515732 4956 584444 5012
rect 584500 4956 584510 5012
rect 30594 4844 30604 4900
rect 30660 4844 60396 4900
rect 60452 4844 60462 4900
rect 64866 4844 64876 4900
rect 64932 4844 88620 4900
rect 88676 4844 88686 4900
rect 89618 4844 89628 4900
rect 89684 4844 109004 4900
rect 109060 4844 109070 4900
rect 110562 4844 110572 4900
rect 110628 4844 126252 4900
rect 126308 4844 126318 4900
rect 127586 4844 127596 4900
rect 127652 4844 140364 4900
rect 140420 4844 140430 4900
rect 141026 4844 141036 4900
rect 141092 4844 151340 4900
rect 151396 4844 151406 4900
rect 284610 4844 284620 4900
rect 284676 4844 302652 4900
rect 302708 4844 302718 4900
rect 304994 4844 305004 4900
rect 305060 4844 327404 4900
rect 327460 4844 327470 4900
rect 337922 4844 337932 4900
rect 337988 4844 367388 4900
rect 367444 4844 367454 4900
rect 425730 4844 425740 4900
rect 425796 4844 474012 4900
rect 474068 4844 474078 4900
rect 496290 4844 496300 4900
rect 496356 4844 559692 4900
rect 559748 4844 559758 4900
rect 40114 4732 40124 4788
rect 40180 4732 68236 4788
rect 68292 4732 68302 4788
rect 70466 4732 70476 4788
rect 70532 4732 93324 4788
rect 93380 4732 93390 4788
rect 95330 4732 95340 4788
rect 95396 4732 113708 4788
rect 113764 4732 113774 4788
rect 120082 4732 120092 4788
rect 120148 4732 134092 4788
rect 134148 4732 134158 4788
rect 142930 4732 142940 4788
rect 142996 4732 152908 4788
rect 152964 4732 152974 4788
rect 283042 4732 283052 4788
rect 283108 4732 300748 4788
rect 300804 4732 300814 4788
rect 301858 4732 301868 4788
rect 301924 4732 323596 4788
rect 323652 4732 323662 4788
rect 336354 4732 336364 4788
rect 336420 4732 365484 4788
rect 365540 4732 365550 4788
rect 486882 4732 486892 4788
rect 486948 4732 548268 4788
rect 548324 4732 548334 4788
rect 43922 4620 43932 4676
rect 43988 4620 71372 4676
rect 71428 4620 71438 4676
rect 72482 4620 72492 4676
rect 72548 4620 94892 4676
rect 94948 4620 94958 4676
rect 99026 4620 99036 4676
rect 99092 4620 116844 4676
rect 116900 4620 116910 4676
rect 125794 4620 125804 4676
rect 125860 4620 138796 4676
rect 138852 4620 138862 4676
rect 144834 4620 144844 4676
rect 144900 4620 154476 4676
rect 154532 4620 154542 4676
rect 158162 4620 158172 4676
rect 158228 4620 165452 4676
rect 165508 4620 165518 4676
rect 242274 4620 242284 4676
rect 242340 4620 251244 4676
rect 251300 4620 251310 4676
rect 298722 4620 298732 4676
rect 298788 4620 319788 4676
rect 319844 4620 319854 4676
rect 328514 4620 328524 4676
rect 328580 4620 355964 4676
rect 356020 4620 356030 4676
rect 477474 4620 477484 4676
rect 477540 4620 536844 4676
rect 536900 4620 536910 4676
rect 45826 4508 45836 4564
rect 45892 4508 72940 4564
rect 72996 4508 73006 4564
rect 74386 4508 74396 4564
rect 74452 4508 96460 4564
rect 96516 4508 96526 4564
rect 101042 4508 101052 4564
rect 101108 4508 118412 4564
rect 118468 4508 118478 4564
rect 129602 4508 129612 4564
rect 129668 4508 141932 4564
rect 141988 4508 141998 4564
rect 146738 4508 146748 4564
rect 146804 4508 156044 4564
rect 156100 4508 156110 4564
rect 240706 4508 240716 4564
rect 240772 4508 249340 4564
rect 249396 4508 249406 4564
rect 297154 4508 297164 4564
rect 297220 4508 317884 4564
rect 317940 4508 317950 4564
rect 326946 4508 326956 4564
rect 327012 4508 354060 4564
rect 354116 4508 354126 4564
rect 468066 4508 468076 4564
rect 468132 4508 525420 4564
rect 525476 4508 525486 4564
rect 47730 4396 47740 4452
rect 47796 4396 74508 4452
rect 74564 4396 74574 4452
rect 76290 4396 76300 4452
rect 76356 4396 98028 4452
rect 98084 4396 98094 4452
rect 102946 4396 102956 4452
rect 103012 4396 119980 4452
rect 120036 4396 120046 4452
rect 131506 4396 131516 4452
rect 131572 4396 143500 4452
rect 143556 4396 143566 4452
rect 148642 4396 148652 4452
rect 148708 4396 157612 4452
rect 157668 4396 157678 4452
rect 239138 4396 239148 4452
rect 239204 4396 247436 4452
rect 247492 4396 247502 4452
rect 295586 4396 295596 4452
rect 295652 4396 315980 4452
rect 316036 4396 316046 4452
rect 322242 4396 322252 4452
rect 322308 4396 348348 4452
rect 348404 4396 348414 4452
rect 463362 4396 463372 4452
rect 463428 4396 519708 4452
rect 519764 4396 519774 4452
rect 51538 4284 51548 4340
rect 51604 4284 77644 4340
rect 77700 4284 77710 4340
rect 78194 4284 78204 4340
rect 78260 4284 99596 4340
rect 99652 4284 99662 4340
rect 104850 4284 104860 4340
rect 104916 4284 121548 4340
rect 121604 4284 121614 4340
rect 290882 4284 290892 4340
rect 290948 4284 310268 4340
rect 310324 4284 310334 4340
rect 320674 4284 320684 4340
rect 320740 4284 346444 4340
rect 346500 4284 346510 4340
rect 444546 4284 444556 4340
rect 444612 4284 496860 4340
rect 496916 4284 496926 4340
rect 53442 4172 53452 4228
rect 53508 4172 79212 4228
rect 79268 4172 79278 4228
rect 82002 4172 82012 4228
rect 82068 4172 102732 4228
rect 102788 4172 102798 4228
rect 108658 4172 108668 4228
rect 108724 4172 124684 4228
rect 124740 4172 124750 4228
rect 289314 4172 289324 4228
rect 289380 4172 308364 4228
rect 308420 4172 308430 4228
rect 319106 4172 319116 4228
rect 319172 4172 344540 4228
rect 344596 4172 344606 4228
rect 411506 4172 411516 4228
rect 411572 4172 430220 4228
rect 430276 4172 430286 4228
rect 57362 4060 57372 4116
rect 57428 4060 82348 4116
rect 82404 4060 82414 4116
rect 83906 4060 83916 4116
rect 83972 4060 104300 4116
rect 104356 4060 104366 4116
rect 112466 4060 112476 4116
rect 112532 4060 127820 4116
rect 127876 4060 127886 4116
rect 287746 4060 287756 4116
rect 287812 4060 306460 4116
rect 306516 4060 306526 4116
rect 317538 4060 317548 4116
rect 317604 4060 342748 4116
rect 342804 4060 342814 4116
rect 401426 4060 401436 4116
rect 401492 4060 416892 4116
rect 416948 4060 416958 4116
rect 61058 3948 61068 4004
rect 61124 3948 73052 4004
rect 73108 3948 73118 4004
rect 281474 3948 281484 4004
rect 281540 3948 298844 4004
rect 298900 3948 298910 4004
rect 314402 3948 314412 4004
rect 314468 3948 338828 4004
rect 338884 3948 338894 4004
rect 389554 3948 389564 4004
rect 389620 3948 399868 4004
rect 399924 3948 399934 4004
rect 412290 3948 412300 4004
rect 412356 3948 456988 4004
rect 457044 3948 457054 4004
rect 161970 3836 161980 3892
rect 162036 3836 168588 3892
rect 168644 3836 168654 3892
rect 351026 3836 351036 3892
rect 351092 3836 382620 3892
rect 382676 3836 382686 3892
rect 387986 3836 387996 3892
rect 388052 3836 422604 3892
rect 422660 3836 422670 3892
rect 428418 3836 428428 3892
rect 428484 3836 439740 3892
rect 439796 3836 439806 3892
rect 150546 3724 150556 3780
rect 150612 3724 159180 3780
rect 159236 3724 159246 3780
rect 164098 3724 164108 3780
rect 164164 3724 170156 3780
rect 170212 3724 170222 3780
rect 245410 3724 245420 3780
rect 245476 3724 255052 3780
rect 255108 3724 255118 3780
rect 381378 3724 381388 3780
rect 381444 3724 409276 3780
rect 409332 3724 409342 3780
rect 416658 3724 416668 3780
rect 416724 3724 428540 3780
rect 428596 3724 428606 3780
rect 435810 3724 435820 3780
rect 435876 3724 485548 3780
rect 485604 3724 485614 3780
rect 503794 3724 503804 3780
rect 503860 3724 514108 3780
rect 514164 3724 514174 3780
rect 152450 3612 152460 3668
rect 152516 3612 160748 3668
rect 160804 3612 160814 3668
rect 165778 3612 165788 3668
rect 165844 3612 171724 3668
rect 171780 3612 171790 3668
rect 218754 3612 218764 3668
rect 218820 3612 222684 3668
rect 222740 3612 222750 3668
rect 223458 3612 223468 3668
rect 223524 3612 228508 3668
rect 228564 3612 228574 3668
rect 243842 3612 243852 3668
rect 243908 3612 253148 3668
rect 253204 3612 253214 3668
rect 366146 3612 366156 3668
rect 366212 3612 394044 3668
rect 394100 3612 394110 3668
rect 407586 3612 407596 3668
rect 407652 3612 449652 3668
rect 450258 3612 450268 3668
rect 450324 3612 462588 3668
rect 462644 3612 462654 3668
rect 480386 3612 480396 3668
rect 480452 3612 491148 3668
rect 491204 3612 491214 3668
rect 512418 3612 512428 3668
rect 512484 3612 580636 3668
rect 580692 3612 580702 3668
rect 449596 3556 449652 3612
rect 154354 3500 154364 3556
rect 154420 3500 162316 3556
rect 162372 3500 162382 3556
rect 167682 3500 167692 3556
rect 167748 3500 173292 3556
rect 173348 3500 173358 3556
rect 186722 3500 186732 3556
rect 186788 3500 188972 3556
rect 189028 3500 189038 3556
rect 210914 3500 210924 3556
rect 210980 3500 213164 3556
rect 213220 3500 213230 3556
rect 214050 3500 214060 3556
rect 214116 3500 216972 3556
rect 217028 3500 217038 3556
rect 217186 3500 217196 3556
rect 217252 3500 220780 3556
rect 220836 3500 220846 3556
rect 221890 3500 221900 3556
rect 221956 3500 226492 3556
rect 226548 3500 226558 3556
rect 237570 3500 237580 3556
rect 237636 3500 245532 3556
rect 245588 3500 245598 3556
rect 359538 3500 359548 3556
rect 359604 3500 376908 3556
rect 376964 3500 376974 3556
rect 377906 3500 377916 3556
rect 377972 3500 411180 3556
rect 411236 3500 411246 3556
rect 440178 3500 440188 3556
rect 440244 3500 449372 3556
rect 449428 3500 449438 3556
rect 449596 3500 451164 3556
rect 451220 3500 451230 3556
rect 456866 3500 456876 3556
rect 456932 3500 468300 3556
rect 468356 3500 468366 3556
rect 492146 3500 492156 3556
rect 492212 3500 502572 3556
rect 502628 3500 502638 3556
rect 524178 3500 524188 3556
rect 524244 3500 531132 3556
rect 531188 3500 531198 3556
rect 21074 3388 21084 3444
rect 21140 3388 51996 3444
rect 52052 3388 52062 3444
rect 156146 3388 156156 3444
rect 156212 3388 163884 3444
rect 163940 3388 163950 3444
rect 169586 3388 169596 3444
rect 169652 3388 174860 3444
rect 174916 3388 174926 3444
rect 188626 3388 188636 3444
rect 188692 3388 190540 3444
rect 190596 3388 190606 3444
rect 209346 3388 209356 3444
rect 209412 3388 211260 3444
rect 211316 3388 211326 3444
rect 212482 3388 212492 3444
rect 212548 3388 215068 3444
rect 215124 3388 215134 3444
rect 215618 3388 215628 3444
rect 215684 3388 218876 3444
rect 218932 3388 218942 3444
rect 220322 3388 220332 3444
rect 220388 3388 224588 3444
rect 224644 3388 224654 3444
rect 236002 3388 236012 3444
rect 236068 3388 243628 3444
rect 243684 3388 243694 3444
rect 246978 3388 246988 3444
rect 247044 3388 257068 3444
rect 257124 3388 257134 3444
rect 372932 3388 388332 3444
rect 388388 3388 388398 3444
rect 435026 3388 435036 3444
rect 435092 3388 445452 3444
rect 445508 3388 445518 3444
rect 449260 3388 454972 3444
rect 455028 3388 455038 3444
rect 471986 3388 471996 3444
rect 472052 3388 479724 3444
rect 479780 3388 479790 3444
rect 484652 3388 493052 3444
rect 493108 3388 493118 3444
rect 494918 3388 494956 3444
rect 495012 3388 495022 3444
rect 498978 3388 498988 3444
rect 499044 3388 500668 3444
rect 500724 3388 500734 3444
rect 503906 3388 503916 3444
rect 503972 3388 510188 3444
rect 510244 3388 510254 3444
rect 510514 3388 510524 3444
rect 510580 3388 515900 3444
rect 515956 3388 515966 3444
rect 529190 3388 529228 3444
rect 529284 3388 529294 3444
rect 557750 3388 557788 3444
rect 557844 3388 557854 3444
rect 565366 3388 565404 3444
rect 565460 3388 565470 3444
rect 372932 3332 372988 3388
rect 253250 3276 253260 3332
rect 253316 3276 264572 3332
rect 264628 3276 264638 3332
rect 268930 3276 268940 3332
rect 268996 3276 283612 3332
rect 283668 3276 283678 3332
rect 323810 3276 323820 3332
rect 323876 3276 350252 3332
rect 350308 3276 350318 3332
rect 359874 3276 359884 3332
rect 359940 3276 366156 3332
rect 366212 3276 366222 3332
rect 367052 3276 372988 3332
rect 373986 3276 373996 3332
rect 374052 3276 377916 3332
rect 377972 3276 377982 3332
rect 383394 3276 383404 3332
rect 383460 3276 387996 3332
rect 388052 3276 388062 3332
rect 447654 3276 447692 3332
rect 447748 3276 447758 3332
rect 367052 3220 367108 3276
rect 449260 3220 449316 3388
rect 471202 3276 471212 3332
rect 471268 3276 475468 3332
rect 475524 3276 475534 3332
rect 36306 3164 36316 3220
rect 36372 3164 65100 3220
rect 65156 3164 65166 3220
rect 254818 3164 254828 3220
rect 254884 3164 266476 3220
rect 266532 3164 266542 3220
rect 272066 3164 272076 3220
rect 272132 3164 287420 3220
rect 287476 3164 287486 3220
rect 300290 3164 300300 3220
rect 300356 3164 321692 3220
rect 321748 3164 321758 3220
rect 325378 3164 325388 3220
rect 325444 3164 352156 3220
rect 352212 3164 352222 3220
rect 355170 3164 355180 3220
rect 355236 3164 367108 3220
rect 372418 3164 372428 3220
rect 372484 3164 381388 3220
rect 381444 3164 381454 3220
rect 410050 3164 410060 3220
rect 410116 3164 449316 3220
rect 452386 3164 452396 3220
rect 452452 3164 462476 3220
rect 462532 3164 462542 3220
rect 466498 3164 466508 3220
rect 466564 3164 483084 3220
rect 483140 3164 483150 3220
rect 484652 3108 484708 3388
rect 499398 3276 499436 3332
rect 499492 3276 499502 3332
rect 500994 3276 501004 3332
rect 501060 3276 501676 3332
rect 501732 3276 501742 3332
rect 34402 3052 34412 3108
rect 34468 3052 63532 3108
rect 63588 3052 63598 3108
rect 256386 3052 256396 3108
rect 256452 3052 268380 3108
rect 268436 3052 268446 3108
rect 273634 3052 273644 3108
rect 273700 3052 289324 3108
rect 289380 3052 289390 3108
rect 303426 3052 303436 3108
rect 303492 3052 325500 3108
rect 325556 3052 325566 3108
rect 330082 3052 330092 3108
rect 330148 3052 357868 3108
rect 357924 3052 357934 3108
rect 386530 3052 386540 3108
rect 386596 3052 426412 3108
rect 426468 3052 426478 3108
rect 441410 3052 441420 3108
rect 441476 3052 484708 3108
rect 485314 3052 485324 3108
rect 485380 3052 546364 3108
rect 546420 3052 546430 3108
rect 32498 2940 32508 2996
rect 32564 2940 61964 2996
rect 62020 2940 62030 2996
rect 80098 2940 80108 2996
rect 80164 2940 101164 2996
rect 101220 2940 101230 2996
rect 259522 2940 259532 2996
rect 259588 2940 272188 2996
rect 272244 2940 272254 2996
rect 276770 2940 276780 2996
rect 276836 2940 293132 2996
rect 293188 2940 293198 2996
rect 306562 2940 306572 2996
rect 306628 2940 329308 2996
rect 329364 2940 329374 2996
rect 334786 2940 334796 2996
rect 334852 2940 363580 2996
rect 363636 2940 363646 2996
rect 378690 2940 378700 2996
rect 378756 2940 401436 2996
rect 401492 2940 401502 2996
rect 405346 2940 405356 2996
rect 405412 2940 440188 2996
rect 440244 2940 440254 2996
rect 457062 2940 457100 2996
rect 457156 2940 457166 2996
rect 490018 2940 490028 2996
rect 490084 2940 552076 2996
rect 552132 2940 552142 2996
rect 26786 2828 26796 2884
rect 26852 2828 57260 2884
rect 57316 2828 57326 2884
rect 66770 2828 66780 2884
rect 66836 2828 90188 2884
rect 90244 2828 90254 2884
rect 97234 2828 97244 2884
rect 97300 2828 115276 2884
rect 115332 2828 115342 2884
rect 121986 2828 121996 2884
rect 122052 2828 135660 2884
rect 135716 2828 135726 2884
rect 229730 2828 229740 2884
rect 229796 2828 236012 2884
rect 236068 2828 236078 2884
rect 262658 2828 262668 2884
rect 262724 2828 275996 2884
rect 276052 2828 276062 2884
rect 278338 2828 278348 2884
rect 278404 2828 295036 2884
rect 295092 2828 295102 2884
rect 309698 2828 309708 2884
rect 309764 2828 333116 2884
rect 333172 2828 333182 2884
rect 339490 2828 339500 2884
rect 339556 2828 369292 2884
rect 369348 2828 369358 2884
rect 402210 2828 402220 2884
rect 402276 2828 435036 2884
rect 435092 2828 435102 2884
rect 439842 2828 439852 2884
rect 439908 2828 480396 2884
rect 480452 2828 480462 2884
rect 491586 2828 491596 2884
rect 491652 2828 553980 2884
rect 554036 2828 554046 2884
rect 24882 2716 24892 2772
rect 24948 2716 55692 2772
rect 55748 2716 55758 2772
rect 62962 2716 62972 2772
rect 63028 2716 87052 2772
rect 87108 2716 87118 2772
rect 93426 2716 93436 2772
rect 93492 2716 112140 2772
rect 112196 2716 112206 2772
rect 118178 2716 118188 2772
rect 118244 2716 132524 2772
rect 132580 2716 132590 2772
rect 137218 2716 137228 2772
rect 137284 2716 148204 2772
rect 148260 2716 148270 2772
rect 175298 2716 175308 2772
rect 175364 2716 179564 2772
rect 179620 2716 179630 2772
rect 231298 2716 231308 2772
rect 231364 2716 237916 2772
rect 237972 2716 237982 2772
rect 248546 2716 248556 2772
rect 248612 2716 258860 2772
rect 258916 2716 258926 2772
rect 264226 2716 264236 2772
rect 264292 2716 277900 2772
rect 277956 2716 277966 2772
rect 279906 2716 279916 2772
rect 279972 2716 296940 2772
rect 296996 2716 297006 2772
rect 311266 2716 311276 2772
rect 311332 2716 335020 2772
rect 335076 2716 335086 2772
rect 348898 2716 348908 2772
rect 348964 2716 380716 2772
rect 380772 2716 380782 2772
rect 389666 2716 389676 2772
rect 389732 2716 411516 2772
rect 411572 2716 411582 2772
rect 414754 2716 414764 2772
rect 414820 2716 460684 2772
rect 460740 2716 460750 2772
rect 508834 2716 508844 2772
rect 508900 2716 574924 2772
rect 574980 2716 574990 2772
rect 19170 2604 19180 2660
rect 19236 2604 50988 2660
rect 51044 2604 51054 2660
rect 59154 2604 59164 2660
rect 59220 2604 83244 2660
rect 83300 2604 83310 2660
rect 91522 2604 91532 2660
rect 91588 2604 109900 2660
rect 109956 2604 109966 2660
rect 116274 2604 116284 2660
rect 116340 2604 130956 2660
rect 131012 2604 131022 2660
rect 135314 2604 135324 2660
rect 135380 2604 146636 2660
rect 146692 2604 146702 2660
rect 173394 2604 173404 2660
rect 173460 2604 177996 2660
rect 178052 2604 178062 2660
rect 179106 2604 179116 2660
rect 179172 2604 182700 2660
rect 182756 2604 182766 2660
rect 182914 2604 182924 2660
rect 182980 2604 185836 2660
rect 185892 2604 185902 2660
rect 226594 2604 226604 2660
rect 226660 2604 232204 2660
rect 232260 2604 232270 2660
rect 234434 2604 234444 2660
rect 234500 2604 241724 2660
rect 241780 2604 241790 2660
rect 257954 2604 257964 2660
rect 258020 2604 270284 2660
rect 270340 2604 270350 2660
rect 270498 2604 270508 2660
rect 270564 2604 285628 2660
rect 285684 2604 285694 2660
rect 286178 2604 286188 2660
rect 286244 2604 304556 2660
rect 304612 2604 304622 2660
rect 308130 2604 308140 2660
rect 308196 2604 331212 2660
rect 331268 2604 331278 2660
rect 331650 2604 331660 2660
rect 331716 2604 359772 2660
rect 359828 2604 359838 2660
rect 363010 2604 363020 2660
rect 363076 2604 397852 2660
rect 397908 2604 397918 2660
rect 424162 2604 424172 2660
rect 424228 2604 472108 2660
rect 472164 2604 472174 2660
rect 475906 2604 475916 2660
rect 475972 2604 507276 2660
rect 507332 2604 507342 2660
rect 510402 2604 510412 2660
rect 510468 2604 576828 2660
rect 576884 2604 576894 2660
rect 17266 2492 17276 2548
rect 17332 2492 49420 2548
rect 49476 2492 49486 2548
rect 55346 2492 55356 2548
rect 55412 2492 80780 2548
rect 80836 2492 80846 2548
rect 87714 2492 87724 2548
rect 87780 2492 107436 2548
rect 107492 2492 107502 2548
rect 114370 2492 114380 2548
rect 114436 2492 129388 2548
rect 129444 2492 129454 2548
rect 133410 2492 133420 2548
rect 133476 2492 145068 2548
rect 145124 2492 145134 2548
rect 171490 2492 171500 2548
rect 171556 2492 176428 2548
rect 176484 2492 176494 2548
rect 181010 2492 181020 2548
rect 181076 2492 184268 2548
rect 184324 2492 184334 2548
rect 184706 2492 184716 2548
rect 184772 2492 187404 2548
rect 187460 2492 187470 2548
rect 225026 2492 225036 2548
rect 225092 2492 230300 2548
rect 230356 2492 230366 2548
rect 232866 2492 232876 2548
rect 232932 2492 239820 2548
rect 239876 2492 239886 2548
rect 250114 2492 250124 2548
rect 250180 2492 260764 2548
rect 260820 2492 260830 2548
rect 261090 2492 261100 2548
rect 261156 2492 274092 2548
rect 274148 2492 274158 2548
rect 275202 2492 275212 2548
rect 275268 2492 291228 2548
rect 291284 2492 291294 2548
rect 292450 2492 292460 2548
rect 292516 2492 312172 2548
rect 312228 2492 312238 2548
rect 312834 2492 312844 2548
rect 312900 2492 336924 2548
rect 336980 2492 336990 2548
rect 344194 2492 344204 2548
rect 344260 2492 375004 2548
rect 375060 2492 375070 2548
rect 377122 2492 377132 2548
rect 377188 2492 414988 2548
rect 415044 2492 415054 2548
rect 438274 2492 438284 2548
rect 438340 2492 489244 2548
rect 489300 2492 489310 2548
rect 504102 2492 504140 2548
rect 504196 2492 504206 2548
rect 505698 2492 505708 2548
rect 505764 2492 510748 2548
rect 510804 2492 510814 2548
rect 513538 2492 513548 2548
rect 513604 2492 582540 2548
rect 582596 2492 582606 2548
rect 41906 2380 41916 2436
rect 41972 2380 69804 2436
rect 69860 2380 69870 2436
rect 177202 2380 177212 2436
rect 177268 2380 181132 2436
rect 181188 2380 181198 2436
rect 228162 2380 228172 2436
rect 228228 2380 234108 2436
rect 234164 2380 234174 2436
rect 251682 2380 251692 2436
rect 251748 2380 262668 2436
rect 262724 2380 262734 2436
rect 267362 2380 267372 2436
rect 267428 2380 281708 2436
rect 281764 2380 281774 2436
rect 358306 2380 358316 2436
rect 358372 2380 392140 2436
rect 392196 2380 392206 2436
rect 408212 2380 432124 2436
rect 432180 2380 432190 2436
rect 472770 2380 472780 2436
rect 472836 2380 524188 2436
rect 524244 2380 524254 2436
rect 49634 2268 49644 2324
rect 49700 2268 76076 2324
rect 76132 2268 76142 2324
rect 265794 2268 265804 2324
rect 265860 2268 279804 2324
rect 279860 2268 279870 2324
rect 345762 2268 345772 2324
rect 345828 2268 359548 2324
rect 359604 2268 359614 2324
rect 369506 2268 369516 2324
rect 369572 2268 405468 2324
rect 405524 2268 405534 2324
rect 408212 2212 408268 2380
rect 421026 2268 421036 2324
rect 421092 2268 456876 2324
rect 456932 2268 456942 2324
rect 480610 2268 480620 2324
rect 480676 2268 509068 2324
rect 509124 2268 509134 2324
rect 38210 2156 38220 2212
rect 38276 2156 66668 2212
rect 66724 2156 66734 2212
rect 364578 2156 364588 2212
rect 364644 2156 389564 2212
rect 389620 2156 389630 2212
rect 391234 2156 391244 2212
rect 391300 2156 408268 2212
rect 416322 2156 416332 2212
rect 416388 2156 450268 2212
rect 450324 2156 450334 2212
rect 458658 2156 458668 2212
rect 458724 2156 503804 2212
rect 503860 2156 503870 2212
rect 397506 2044 397516 2100
rect 397572 2044 428428 2100
rect 428484 2044 428494 2100
rect 461794 2044 461804 2100
rect 461860 2044 517804 2100
rect 517860 2044 517870 2100
rect 388098 1932 388108 1988
rect 388164 1932 416668 1988
rect 416724 1932 416734 1988
rect 430434 1932 430444 1988
rect 430500 1932 471996 1988
rect 472052 1932 472062 1988
rect 482178 1932 482188 1988
rect 482244 1932 525868 1988
rect 361442 1820 361452 1876
rect 361508 1820 364476 1876
rect 364532 1820 364542 1876
rect 436706 1820 436716 1876
rect 436772 1820 436828 1876
rect 436884 1820 436894 1876
rect 449250 1820 449260 1876
rect 449316 1820 492156 1876
rect 492212 1820 492222 1876
rect 525812 1764 525868 1932
rect 525812 1708 542556 1764
rect 542612 1708 542622 1764
rect 563462 1708 563500 1764
rect 563556 1708 563566 1764
rect 394370 1596 394380 1652
rect 394436 1596 435932 1652
rect 435988 1596 435998 1652
rect 497858 1596 497868 1652
rect 497924 1596 561596 1652
rect 561652 1596 561662 1652
rect 384962 1484 384972 1540
rect 385028 1484 424508 1540
rect 424564 1484 424574 1540
rect 460226 1484 460236 1540
rect 460292 1484 510524 1540
rect 510580 1484 510590 1540
rect 423266 1372 423276 1428
rect 423332 1372 470204 1428
rect 470260 1372 470270 1428
rect 455522 1260 455532 1316
rect 455588 1260 503916 1316
rect 503972 1260 503982 1316
rect 413186 1148 413196 1204
rect 413252 1148 420028 1204
rect 483746 1148 483756 1204
rect 483812 1148 487676 1204
rect 487732 1148 487742 1204
rect 419972 980 420028 1148
rect 419972 924 458780 980
rect 458836 924 458846 980
rect 507266 924 507276 980
rect 507332 924 514108 980
rect 514052 868 514108 924
rect 352034 812 352044 868
rect 352100 812 384524 868
rect 384580 812 384590 868
rect 403778 812 403788 868
rect 403844 812 447356 868
rect 447412 812 447422 868
rect 450818 812 450828 868
rect 450884 812 504476 868
rect 504532 812 504542 868
rect 509058 812 509068 868
rect 509124 812 512372 868
rect 514052 812 534940 868
rect 534996 812 535006 868
rect 512316 756 512372 812
rect 347778 700 347788 756
rect 347844 700 378812 756
rect 378868 700 378878 756
rect 399074 700 399084 756
rect 399140 700 441644 756
rect 441700 700 441710 756
rect 446114 700 446124 756
rect 446180 700 498764 756
rect 498820 700 498830 756
rect 512054 700 512092 756
rect 512148 700 512158 756
rect 512316 700 540652 756
rect 540708 700 540718 756
rect 364466 588 364476 644
rect 364532 588 395948 644
rect 396004 588 396014 644
rect 396452 588 401660 644
rect 401716 588 401726 644
rect 408482 588 408492 644
rect 408548 588 453068 644
rect 453124 588 453134 644
rect 464930 588 464940 644
rect 464996 588 521612 644
rect 521668 588 521678 644
rect 537572 588 538748 644
rect 538804 588 538814 644
rect 569174 588 569212 644
rect 569268 588 569278 644
rect 571190 588 571228 644
rect 571284 588 571294 644
rect 342514 476 342524 532
rect 342580 476 349468 532
rect 356738 476 356748 532
rect 356804 476 390124 532
rect 390180 476 390190 532
rect 23090 252 23100 308
rect 23156 252 54124 308
rect 54180 252 54190 308
rect 349412 196 349468 476
rect 396452 420 396508 588
rect 417890 476 417900 532
rect 417956 476 464380 532
rect 464436 476 464446 532
rect 469634 476 469644 532
rect 469700 476 527212 532
rect 527268 476 527278 532
rect 537572 420 537628 588
rect 366370 364 366380 420
rect 366436 364 396508 420
rect 427298 364 427308 420
rect 427364 364 475804 420
rect 475860 364 475870 420
rect 487452 364 537628 420
rect 370850 252 370860 308
rect 370916 252 407260 308
rect 407316 252 407326 308
rect 433010 252 433020 308
rect 433076 252 481516 308
rect 481572 252 481582 308
rect 13570 140 13580 196
rect 13636 140 46284 196
rect 46340 140 46350 196
rect 349412 140 372988 196
rect 373044 140 373054 196
rect 376226 140 376236 196
rect 376292 140 412972 196
rect 413028 140 413038 196
rect 436818 140 436828 196
rect 436884 140 487228 196
rect 487284 140 487294 196
rect 487452 84 487508 364
rect 487666 252 487676 308
rect 487732 252 544348 308
rect 544404 252 544414 308
rect 488450 140 488460 196
rect 488516 140 550060 196
rect 550116 140 550126 196
rect 11666 28 11676 84
rect 11732 28 44716 84
rect 44772 28 44782 84
rect 380034 28 380044 84
rect 380100 28 418684 84
rect 418740 28 418750 84
rect 479042 28 479052 84
rect 479108 28 487508 84
rect 503458 28 503468 84
rect 503524 28 567196 84
rect 567252 28 567262 84
<< via3 >>
rect 111692 590940 111748 590996
rect 120092 590716 120148 590772
rect 199948 590716 200004 590772
rect 106652 590604 106708 590660
rect 52892 590492 52948 590548
rect 584668 590156 584724 590212
rect 590492 588588 590548 588644
rect 199836 587132 199892 587188
rect 54572 575372 54628 575428
rect 120204 573020 120260 573076
rect 590604 562156 590660 562212
rect 111804 558908 111860 558964
rect 108332 544796 108388 544852
rect 59836 535724 59892 535780
rect 2492 530684 2548 530740
rect 54460 523292 54516 523348
rect 590604 523292 590660 523348
rect 28 516460 84 516516
rect 200060 511532 200116 511588
rect 49532 496076 49588 496132
rect 4172 488348 4228 488404
rect 59612 482972 59668 483028
rect 590492 482972 590548 483028
rect 62972 482860 63028 482916
rect 114268 474236 114324 474292
rect 1484 469644 1540 469700
rect 60620 456428 60676 456484
rect 4396 446012 4452 446068
rect 60508 437612 60564 437668
rect 110012 431900 110068 431956
rect 57932 430108 57988 430164
rect 140 403564 196 403620
rect 3164 403564 3220 403620
rect 203420 390572 203476 390628
rect 513212 390348 513268 390404
rect 387212 374668 387268 374724
rect 212156 373324 212212 373380
rect 211932 373212 211988 373268
rect 54684 373100 54740 373156
rect 197708 371756 197764 371812
rect 211708 371644 211764 371700
rect 210252 371420 210308 371476
rect 210140 370300 210196 370356
rect 196588 370188 196644 370244
rect 194908 370076 194964 370132
rect 199500 368620 199556 368676
rect 213388 367948 213444 368004
rect 204204 366828 204260 366884
rect 210028 366604 210084 366660
rect 195020 366380 195076 366436
rect 112476 365484 112532 365540
rect 209692 365372 209748 365428
rect 209244 365260 209300 365316
rect 209468 365148 209524 365204
rect 213500 364812 213556 364868
rect 199724 364588 199780 364644
rect 590492 363916 590548 363972
rect 171276 363692 171332 363748
rect 204316 363468 204372 363524
rect 114156 363356 114212 363412
rect 196700 363356 196756 363412
rect 160748 363020 160804 363076
rect 164668 363020 164724 363076
rect 194572 363020 194628 363076
rect 151340 362908 151396 362964
rect 152012 362908 152068 362964
rect 156156 362908 156212 362964
rect 157836 362908 157892 362964
rect 163436 362124 163492 362180
rect 193340 362124 193396 362180
rect 199948 362124 200004 362180
rect 200284 362124 200340 362180
rect 155372 361900 155428 361956
rect 205996 361900 206052 361956
rect 207564 361788 207620 361844
rect 150668 361564 150724 361620
rect 155372 361564 155428 361620
rect 211820 361564 211876 361620
rect 161420 361116 161476 361172
rect 197372 360556 197428 360612
rect 194684 360108 194740 360164
rect 166124 359548 166180 359604
rect 173516 359548 173572 359604
rect 190764 359548 190820 359604
rect 190988 359548 191044 359604
rect 192556 359548 192612 359604
rect 194236 359548 194292 359604
rect 195692 359548 195748 359604
rect 197372 359548 197428 359604
rect 182252 359436 182308 359492
rect 186956 359436 187012 359492
rect 189532 359436 189588 359492
rect 193004 359436 193060 359492
rect 194348 359436 194404 359492
rect 200060 358652 200116 358708
rect 200396 358652 200452 358708
rect 63756 358092 63812 358148
rect 199276 357644 199332 357700
rect 199276 357084 199332 357140
rect 199388 355964 199444 356020
rect 117404 355852 117460 355908
rect 58268 354732 58324 354788
rect 202076 354284 202132 354340
rect 58604 353612 58660 353668
rect 117180 352492 117236 352548
rect 91532 351372 91588 351428
rect 116620 350252 116676 350308
rect 201852 349804 201908 349860
rect 61292 348012 61348 348068
rect 112588 346892 112644 346948
rect 107436 345772 107492 345828
rect 64652 344652 64708 344708
rect 200620 344204 200676 344260
rect 58492 343532 58548 343588
rect 57820 342412 57876 342468
rect 202188 341964 202244 342020
rect 56588 340284 56644 340340
rect 107436 340284 107492 340340
rect 116732 340172 116788 340228
rect 117068 340172 117124 340228
rect 201964 339724 202020 339780
rect 108668 339388 108724 339444
rect 118636 339276 118692 339332
rect 60060 338828 60116 338884
rect 116620 338828 116676 338884
rect 56812 338716 56868 338772
rect 112588 338716 112644 338772
rect 116844 338604 116900 338660
rect 119196 337484 119252 337540
rect 210364 337484 210420 337540
rect 58716 337260 58772 337316
rect 117180 337260 117236 337316
rect 109116 337148 109172 337204
rect 119196 336924 119252 336980
rect 199276 336364 199332 336420
rect 109116 336028 109172 336084
rect 116956 336028 117012 336084
rect 206892 335244 206948 335300
rect 7532 335132 7588 335188
rect 118748 334796 118804 334852
rect 120540 334460 120596 334516
rect 56924 334348 56980 334404
rect 64652 334348 64708 334404
rect 202076 334124 202132 334180
rect 51212 333452 51268 333508
rect 63532 333452 63588 333508
rect 51436 333340 51492 333396
rect 4284 333116 4340 333172
rect 60396 333004 60452 333060
rect 203308 333004 203364 333060
rect 53004 332892 53060 332948
rect 63644 332668 63700 332724
rect 56700 331772 56756 331828
rect 91532 331772 91588 331828
rect 201964 331884 202020 331940
rect 119196 331660 119252 331716
rect 119868 331548 119924 331604
rect 114156 330988 114212 331044
rect 57708 330876 57764 330932
rect 62972 330876 63028 330932
rect 56476 330764 56532 330820
rect 61292 330764 61348 330820
rect 58044 330204 58100 330260
rect 199276 330204 199332 330260
rect 119644 329980 119700 330036
rect 115052 329756 115108 329812
rect 120316 329308 120372 329364
rect 200060 329252 200116 329308
rect 200284 329196 200340 329252
rect 118860 329084 118916 329140
rect 115948 328972 116004 329028
rect 210476 328524 210532 328580
rect 111916 328412 111972 328468
rect 423948 328076 424004 328132
rect 431788 327964 431844 328020
rect 112252 327852 112308 327908
rect 420140 327852 420196 327908
rect 112588 327740 112644 327796
rect 380268 327740 380324 327796
rect 420028 327740 420084 327796
rect 426860 327740 426916 327796
rect 370636 327628 370692 327684
rect 426748 327628 426804 327684
rect 428428 326172 428484 326228
rect 433468 326060 433524 326116
rect 379708 325948 379764 326004
rect 57932 325724 57988 325780
rect 113484 325724 113540 325780
rect 115276 325612 115332 325668
rect 199276 325164 199332 325220
rect 5292 324828 5348 324884
rect 4956 324604 5012 324660
rect 57036 325052 57092 325108
rect 113820 325052 113876 325108
rect 208124 325052 208180 325108
rect 212268 325052 212324 325108
rect 410732 324940 410788 324996
rect 423388 324940 423444 324996
rect 377580 324828 377636 324884
rect 442092 324828 442148 324884
rect 376124 324716 376180 324772
rect 441868 324716 441924 324772
rect 58380 324604 58436 324660
rect 373884 324604 373940 324660
rect 440300 324604 440356 324660
rect 115500 324492 115556 324548
rect 380380 324492 380436 324548
rect 432124 324492 432180 324548
rect 112028 324380 112084 324436
rect 410732 324380 410788 324436
rect 411404 324380 411460 324436
rect 418348 324380 418404 324436
rect 418796 324380 418852 324436
rect 421260 324380 421316 324436
rect 422044 324380 422100 324436
rect 422604 324380 422660 324436
rect 424172 324380 424228 324436
rect 425068 324380 425124 324436
rect 426188 324380 426244 324436
rect 426412 324380 426468 324436
rect 114268 324156 114324 324212
rect 199388 324044 199444 324100
rect 57932 323708 57988 323764
rect 113708 323708 113764 323764
rect 113260 323372 113316 323428
rect 426412 323372 426468 323428
rect 436828 323372 436884 323428
rect 58156 323036 58212 323092
rect 113036 323036 113092 323092
rect 379036 323036 379092 323092
rect 442316 323036 442372 323092
rect 201852 322924 201908 322980
rect 378812 322924 378868 322980
rect 442204 322924 442260 322980
rect 375452 322812 375508 322868
rect 441980 322812 442036 322868
rect 373660 322700 373716 322756
rect 440412 322700 440468 322756
rect 373772 322588 373828 322644
rect 440188 322588 440244 322644
rect 58604 322364 58660 322420
rect 113596 322364 113652 322420
rect 115612 322252 115668 322308
rect 206668 321804 206724 321860
rect 58716 321692 58772 321748
rect 113372 321692 113428 321748
rect 114828 321132 114884 321188
rect 56140 321020 56196 321076
rect 57820 321020 57876 321076
rect 60172 321020 60228 321076
rect 117404 321020 117460 321076
rect 57148 320908 57204 320964
rect 56700 320348 56756 320404
rect 117292 320348 117348 320404
rect 115388 320012 115444 320068
rect 210588 320012 210644 320068
rect 60060 319676 60116 319732
rect 113148 319676 113204 319732
rect 116620 319004 116676 319060
rect 5068 318332 5124 318388
rect 117180 318332 117236 318388
rect 373884 318108 373940 318164
rect 199276 317772 199332 317828
rect 115164 317660 115220 317716
rect 58268 317436 58324 317492
rect 112588 317436 112644 317492
rect 202300 317324 202356 317380
rect 115948 316988 116004 317044
rect 115836 316652 115892 316708
rect 376012 316652 376068 316708
rect 56476 316316 56532 316372
rect 113932 316316 113988 316372
rect 200172 316204 200228 316260
rect 377468 315980 377524 316036
rect 377580 315868 377636 315924
rect 115724 315644 115780 315700
rect 117180 315532 117236 315588
rect 376796 315308 376852 315364
rect 199612 315084 199668 315140
rect 117180 314972 117236 315028
rect 373772 314748 373828 314804
rect 117292 314412 117348 314468
rect 58268 314300 58324 314356
rect 115836 314300 115892 314356
rect 56252 314188 56308 314244
rect 116956 313964 117012 314020
rect 120428 313964 120484 314020
rect 202524 313964 202580 314020
rect 56812 313628 56868 313684
rect 379036 313628 379092 313684
rect 116620 313292 116676 313348
rect 200508 312844 200564 312900
rect 443548 312620 443604 312676
rect 114044 312508 114100 312564
rect 373772 312508 373828 312564
rect 113148 312172 113204 312228
rect 441868 311948 441924 312004
rect 378812 311388 378868 311444
rect 445228 311276 445284 311332
rect 113372 311052 113428 311108
rect 543452 311052 543508 311108
rect 3052 310940 3108 310996
rect 114268 310940 114324 310996
rect 116956 310716 117012 310772
rect 200284 310604 200340 310660
rect 377356 310604 377412 310660
rect 115948 309932 116004 309988
rect 200396 309484 200452 309540
rect 57036 309148 57092 309204
rect 58492 309148 58548 309204
rect 375452 309148 375508 309204
rect 58716 308924 58772 308980
rect 5292 308700 5348 308756
rect 445340 308588 445396 308644
rect 118524 308364 118580 308420
rect 373884 308028 373940 308084
rect 442540 307916 442596 307972
rect 373660 306908 373716 306964
rect 117292 306572 117348 306628
rect 443660 306572 443716 306628
rect 114828 306236 114884 306292
rect 115052 305452 115108 305508
rect 440860 305228 440916 305284
rect 118412 305004 118468 305060
rect 57708 304892 57764 304948
rect 57148 304668 57204 304724
rect 442652 304556 442708 304612
rect 115724 304332 115780 304388
rect 56588 304220 56644 304276
rect 199836 303884 199892 303940
rect 442204 303884 442260 303940
rect 58492 303548 58548 303604
rect 118860 303212 118916 303268
rect 376236 303212 376292 303268
rect 441980 303212 442036 303268
rect 56364 302876 56420 302932
rect 115612 302876 115668 302932
rect 441084 302540 441140 302596
rect 377244 302428 377300 302484
rect 376460 301868 376516 301924
rect 440972 301868 441028 301924
rect 54460 301532 54516 301588
rect 56924 301532 56980 301588
rect 199276 301196 199332 301252
rect 440300 301196 440356 301252
rect 59724 300860 59780 300916
rect 110908 300860 110964 300916
rect 206780 300748 206836 300804
rect 113820 300524 113876 300580
rect 115836 300524 115892 300580
rect 199276 300524 199332 300580
rect 56476 300188 56532 300244
rect 113260 300188 113316 300244
rect 376460 300188 376516 300244
rect 442204 300524 442260 300580
rect 111916 299964 111972 300020
rect 202188 299404 202244 299460
rect 377244 299852 377300 299908
rect 440412 299852 440468 299908
rect 373660 299180 373716 299236
rect 442316 299180 442372 299236
rect 112252 299068 112308 299124
rect 112700 299068 112756 299124
rect 117404 298732 117460 298788
rect 373884 298508 373940 298564
rect 442092 298508 442148 298564
rect 202636 298284 202692 298340
rect 57036 298172 57092 298228
rect 117628 298172 117684 298228
rect 442764 297836 442820 297892
rect 590156 297836 590212 297892
rect 112028 297612 112084 297668
rect 3052 297500 3108 297556
rect 56140 297500 56196 297556
rect 440636 297164 440692 297220
rect 199276 296716 199332 296772
rect 440524 296492 440580 296548
rect 563612 296492 563668 296548
rect 590156 296492 590212 296548
rect 199276 296380 199332 296436
rect 115500 296156 115556 296212
rect 201852 296044 201908 296100
rect 441868 295820 441924 295876
rect 373772 295708 373828 295764
rect 112588 295596 112644 295652
rect 115276 295596 115332 295652
rect 115836 295372 115892 295428
rect 442316 295148 442372 295204
rect 373772 294588 373828 294644
rect 440188 294476 440244 294532
rect 201740 293804 201796 293860
rect 372876 293804 372932 293860
rect 440524 293804 440580 293860
rect 375452 293468 375508 293524
rect 113596 293132 113652 293188
rect 440300 293132 440356 293188
rect 115388 292796 115444 292852
rect 440188 292460 440244 292516
rect 372092 292348 372148 292404
rect 117180 292012 117236 292068
rect 113484 291900 113540 291956
rect 114716 291900 114772 291956
rect 441980 291788 442036 291844
rect 112588 291452 112644 291508
rect 113708 291340 113764 291396
rect 114268 291340 114324 291396
rect 375676 291228 375732 291284
rect 379372 291116 379428 291172
rect 442428 291116 442484 291172
rect 113932 290892 113988 290948
rect 4732 290780 4788 290836
rect 112812 290780 112868 290836
rect 440748 290444 440804 290500
rect 373660 290108 373716 290164
rect 114716 289772 114772 289828
rect 442092 289772 442148 289828
rect 114044 289436 114100 289492
rect 380492 289100 380548 289156
rect 372428 288988 372484 289044
rect 114268 288652 114324 288708
rect 59612 288316 59668 288372
rect 373884 287868 373940 287924
rect 199276 287532 199332 287588
rect 58716 287420 58772 287476
rect 112700 286076 112756 286132
rect 380604 286076 380660 286132
rect 5180 285404 5236 285460
rect 377244 285068 377300 285124
rect 1484 284732 1540 284788
rect 202412 284732 202468 284788
rect 207676 284732 207732 284788
rect 113372 284508 113428 284564
rect 565292 284620 565348 284676
rect 373324 284508 373380 284564
rect 58716 284060 58772 284116
rect 5292 283388 5348 283444
rect 58716 283388 58772 283444
rect 375564 283388 375620 283444
rect 68796 282940 68852 282996
rect 87612 282828 87668 282884
rect 7532 282268 7588 282324
rect 115164 282268 115220 282324
rect 373436 282268 373492 282324
rect 115164 282044 115220 282100
rect 97356 281820 97412 281876
rect 40684 281708 40740 281764
rect 75516 281708 75572 281764
rect 25900 281596 25956 281652
rect 59836 281596 59892 281652
rect 85596 281596 85652 281652
rect 26572 281484 26628 281540
rect 118860 281372 118916 281428
rect 374892 281148 374948 281204
rect 85596 280924 85652 280980
rect 97356 280924 97412 280980
rect 45388 280812 45444 280868
rect 63756 280700 63812 280756
rect 74172 280700 74228 280756
rect 87612 280700 87668 280756
rect 121548 280700 121604 280756
rect 199948 280700 200004 280756
rect 40684 280588 40740 280644
rect 157052 280588 157108 280644
rect 3164 280476 3220 280532
rect 25900 280476 25956 280532
rect 26572 280476 26628 280532
rect 45388 280476 45444 280532
rect 127484 280476 127540 280532
rect 127708 280476 127764 280532
rect 133644 280476 133700 280532
rect 139692 280476 139748 280532
rect 141036 280476 141092 280532
rect 146412 280476 146468 280532
rect 163660 280476 163716 280532
rect 186396 280476 186452 280532
rect 194572 280476 194628 280532
rect 198156 280476 198212 280532
rect 186284 280364 186340 280420
rect 195020 280364 195076 280420
rect 49532 280252 49588 280308
rect 74172 280028 74228 280084
rect 75516 280028 75572 280084
rect 77532 280028 77588 280084
rect 119308 280028 119364 280084
rect 121884 280028 121940 280084
rect 122332 280028 122388 280084
rect 127484 280028 127540 280084
rect 194796 280028 194852 280084
rect 374780 280028 374836 280084
rect 58044 279804 58100 279860
rect 165676 279804 165732 279860
rect 206892 279804 206948 279860
rect 121436 279692 121492 279748
rect 137676 279692 137732 279748
rect 200732 279692 200788 279748
rect 105308 279020 105364 279076
rect 111132 278908 111188 278964
rect 375004 278908 375060 278964
rect 52892 278796 52948 278852
rect 200060 278796 200116 278852
rect 174636 278684 174692 278740
rect 54572 278572 54628 278628
rect 170492 278572 170548 278628
rect 193340 278572 193396 278628
rect 74172 278460 74228 278516
rect 187404 278460 187460 278516
rect 186172 278348 186228 278404
rect 196700 278348 196756 278404
rect 60620 278236 60676 278292
rect 113372 278236 113428 278292
rect 137004 278236 137060 278292
rect 168812 278236 168868 278292
rect 56252 278124 56308 278180
rect 112700 278124 112756 278180
rect 115052 278124 115108 278180
rect 154476 278124 154532 278180
rect 197596 278124 197652 278180
rect 530012 278012 530068 278068
rect 590492 278012 590548 278068
rect 60508 277900 60564 277956
rect 105308 277900 105364 277956
rect 7084 277116 7140 277172
rect 7756 277116 7812 277172
rect 45276 277116 45332 277172
rect 48748 277116 48804 277172
rect 63868 277116 63924 277172
rect 119980 277116 120036 277172
rect 151116 277116 151172 277172
rect 157948 277116 158004 277172
rect 159964 277116 160020 277172
rect 165228 277116 165284 277172
rect 165900 277116 165956 277172
rect 175308 277116 175364 277172
rect 178892 277116 178948 277172
rect 196588 277116 196644 277172
rect 372092 277116 372148 277172
rect 441868 277116 441924 277172
rect 17612 277004 17668 277060
rect 63420 277004 63476 277060
rect 181356 277004 181412 277060
rect 195916 277004 195972 277060
rect 62188 276892 62244 276948
rect 84812 276892 84868 276948
rect 160412 276892 160468 276948
rect 106764 276780 106820 276836
rect 163772 276780 163828 276836
rect 64204 276668 64260 276724
rect 70364 276668 70420 276724
rect 160524 276668 160580 276724
rect 373324 277004 373380 277060
rect 440300 277004 440356 277060
rect 373772 276892 373828 276948
rect 440636 276892 440692 276948
rect 375452 276780 375508 276836
rect 442204 276780 442260 276836
rect 373548 276668 373604 276724
rect 375676 276668 375732 276724
rect 442428 276668 442484 276724
rect 60396 276556 60452 276612
rect 63420 276556 63476 276612
rect 70252 276556 70308 276612
rect 72156 276556 72212 276612
rect 178892 276556 178948 276612
rect 374780 276556 374836 276612
rect 442092 276556 442148 276612
rect 189420 276444 189476 276500
rect 82236 276332 82292 276388
rect 188972 276332 189028 276388
rect 189532 276332 189588 276388
rect 175980 276220 176036 276276
rect 186732 276220 186788 276276
rect 210700 276220 210756 276276
rect 48636 276108 48692 276164
rect 82236 276108 82292 276164
rect 197036 276108 197092 276164
rect 94892 275996 94948 276052
rect 108668 275996 108724 276052
rect 203420 275884 203476 275940
rect 180012 275772 180068 275828
rect 184716 275772 184772 275828
rect 199724 275772 199780 275828
rect 179788 275660 179844 275716
rect 183148 275660 183204 275716
rect 188076 275660 188132 275716
rect 372652 275660 372708 275716
rect 26012 275548 26068 275604
rect 36876 275548 36932 275604
rect 41132 275548 41188 275604
rect 61404 275548 61460 275604
rect 64092 275548 64148 275604
rect 72156 275548 72212 275604
rect 103628 275548 103684 275604
rect 168140 275548 168196 275604
rect 169260 275548 169316 275604
rect 169708 275548 169764 275604
rect 176540 275548 176596 275604
rect 177324 275548 177380 275604
rect 178108 275548 178164 275604
rect 179900 275548 179956 275604
rect 181468 275548 181524 275604
rect 184828 275548 184884 275604
rect 188748 275548 188804 275604
rect 189420 275548 189476 275604
rect 190428 275548 190484 275604
rect 197708 275548 197764 275604
rect 375116 275548 375172 275604
rect 373660 275436 373716 275492
rect 440748 275436 440804 275492
rect 374892 275324 374948 275380
rect 441980 275324 442036 275380
rect 375564 275212 375620 275268
rect 442316 275212 442372 275268
rect 373436 275100 373492 275156
rect 440188 275100 440244 275156
rect 84812 274764 84868 274820
rect 119196 274764 119252 274820
rect 199052 274764 199108 274820
rect 375788 274764 375844 274820
rect 443660 274764 443716 274820
rect 94892 274652 94948 274708
rect 103404 274652 103460 274708
rect 202636 274652 202692 274708
rect 117068 274540 117124 274596
rect 150332 274540 150388 274596
rect 375228 274428 375284 274484
rect 372428 273756 372484 273812
rect 442764 273756 442820 273812
rect 373884 273644 373940 273700
rect 440524 273644 440580 273700
rect 373324 273308 373380 273364
rect 422604 273308 422660 273364
rect 423948 273196 424004 273252
rect 39676 273084 39732 273140
rect 375004 273084 375060 273140
rect 442092 273084 442148 273140
rect 70364 272860 70420 272916
rect 79772 272860 79828 272916
rect 404012 272188 404068 272244
rect 385420 272076 385476 272132
rect 387212 272076 387268 272132
rect 383852 271964 383908 272020
rect 419916 271964 419972 272020
rect 423388 271964 423444 272020
rect 387436 271852 387492 271908
rect 431788 271740 431844 271796
rect 51212 271628 51268 271684
rect 416332 271628 416388 271684
rect 425068 271628 425124 271684
rect 51436 271516 51492 271572
rect 431788 271516 431844 271572
rect 62972 271404 63028 271460
rect 430108 271404 430164 271460
rect 550172 271404 550228 271460
rect 28476 271292 28532 271348
rect 167132 271292 167188 271348
rect 194348 271292 194404 271348
rect 370972 271292 371028 271348
rect 387324 271292 387380 271348
rect 431900 271292 431956 271348
rect 100044 271180 100100 271236
rect 409948 271180 410004 271236
rect 420140 271180 420196 271236
rect 7532 271068 7588 271124
rect 388108 271068 388164 271124
rect 410060 271068 410116 271124
rect 411628 271068 411684 271124
rect 413308 271068 413364 271124
rect 414988 271068 415044 271124
rect 418348 271068 418404 271124
rect 210252 270844 210308 270900
rect 375004 270844 375060 270900
rect 176428 270508 176484 270564
rect 7644 270396 7700 270452
rect 387996 270396 388052 270452
rect 418460 270284 418516 270340
rect 422044 270284 422100 270340
rect 194572 270060 194628 270116
rect 53004 269948 53060 270004
rect 172172 269948 172228 270004
rect 197372 269948 197428 270004
rect 420028 269836 420084 269892
rect 21756 269724 21812 269780
rect 64092 269724 64148 269780
rect 201964 269724 202020 269780
rect 372540 269612 372596 269668
rect 441084 269612 441140 269668
rect 411740 268940 411796 268996
rect 418796 268940 418852 268996
rect 440412 268828 440468 268884
rect 421484 268716 421540 268772
rect 375676 268492 375732 268548
rect 139356 268380 139412 268436
rect 199836 268380 199892 268436
rect 372764 268380 372820 268436
rect 372428 268156 372484 268212
rect 99932 268044 99988 268100
rect 111692 268044 111748 268100
rect 381500 268044 381556 268100
rect 426748 268044 426804 268100
rect 424620 267820 424676 267876
rect 426860 267708 426916 267764
rect 380156 267596 380212 267652
rect 428428 267372 428484 267428
rect 419916 267260 419972 267316
rect 418572 267148 418628 267204
rect 420364 267148 420420 267204
rect 61292 266924 61348 266980
rect 373548 266700 373604 266756
rect 440300 266700 440356 266756
rect 380044 266588 380100 266644
rect 122556 266476 122612 266532
rect 197484 266476 197540 266532
rect 375116 266476 375172 266532
rect 441980 266476 442036 266532
rect 26796 266364 26852 266420
rect 83916 266364 83972 266420
rect 199612 266364 199668 266420
rect 373324 266364 373380 266420
rect 440524 266364 440580 266420
rect 370748 266252 370804 266308
rect 440972 266252 441028 266308
rect 187404 265468 187460 265524
rect 403564 265692 403620 265748
rect 410956 265692 411012 265748
rect 183036 265356 183092 265412
rect 373884 265132 373940 265188
rect 442428 265132 442484 265188
rect 404012 265020 404068 265076
rect 442316 265020 442372 265076
rect 379260 264908 379316 264964
rect 442540 264908 442596 264964
rect 379148 264796 379204 264852
rect 442652 264796 442708 264852
rect 104972 264684 105028 264740
rect 375228 264572 375284 264628
rect 442204 264572 442260 264628
rect 433468 264460 433524 264516
rect 403564 264236 403620 264292
rect 406252 264236 406308 264292
rect 406924 264236 406980 264292
rect 410956 264236 411012 264292
rect 413644 264236 413700 264292
rect 189084 264124 189140 264180
rect 373436 263900 373492 263956
rect 373660 263788 373716 263844
rect 380604 263676 380660 263732
rect 410956 263676 411012 263732
rect 426188 263676 426244 263732
rect 434252 263676 434308 263732
rect 411628 263564 411684 263620
rect 414988 263452 415044 263508
rect 406252 263340 406308 263396
rect 406924 263340 406980 263396
rect 411740 263340 411796 263396
rect 440972 263228 441028 263284
rect 413644 263116 413700 263172
rect 410060 263004 410116 263060
rect 418348 263004 418404 263060
rect 433580 263004 433636 263060
rect 373772 262892 373828 262948
rect 440860 262892 440916 262948
rect 388108 261660 388164 261716
rect 409948 261548 410004 261604
rect 373884 260988 373940 261044
rect 210140 260092 210196 260148
rect 372092 258748 372148 258804
rect 555212 258188 555268 258244
rect 210700 257404 210756 257460
rect 377580 256060 377636 256116
rect 377132 255836 377188 255892
rect 377580 255836 377636 255892
rect 377132 254268 377188 254324
rect 206108 252028 206164 252084
rect 376460 252028 376516 252084
rect 373324 250908 373380 250964
rect 377580 250012 377636 250068
rect 372988 249788 373044 249844
rect 379932 249564 379988 249620
rect 204316 249452 204372 249508
rect 371084 248780 371140 248836
rect 373772 248780 373828 248836
rect 4956 248556 5012 248612
rect 376236 247996 376292 248052
rect 376460 247324 376516 247380
rect 373436 246876 373492 246932
rect 376236 246876 376292 246932
rect 376460 246428 376516 246484
rect 373772 245308 373828 245364
rect 587132 244972 587188 245028
rect 376460 244636 376516 244692
rect 373884 244188 373940 244244
rect 376236 243068 376292 243124
rect 373660 242732 373716 242788
rect 378588 242620 378644 242676
rect 373884 242060 373940 242116
rect 372988 241948 373044 242004
rect 440188 241948 440244 242004
rect 380044 241724 380100 241780
rect 373436 240828 373492 240884
rect 440412 240604 440468 240660
rect 373660 240268 373716 240324
rect 370076 239708 370132 239764
rect 439964 239820 440020 239876
rect 373548 238812 373604 238868
rect 375564 238700 375620 238756
rect 210028 238588 210084 238644
rect 373324 238588 373380 238644
rect 371196 237804 371252 237860
rect 379484 237804 379540 237860
rect 378924 237692 378980 237748
rect 442316 237244 442372 237300
rect 379932 236908 379988 236964
rect 372204 236796 372260 236852
rect 373660 236796 373716 236852
rect 442092 236572 442148 236628
rect 375116 236348 375172 236404
rect 210700 235900 210756 235956
rect 376236 235900 376292 235956
rect 440300 235900 440356 235956
rect 373660 235788 373716 235844
rect 440972 235116 441028 235172
rect 441868 235116 441924 235172
rect 371196 234780 371252 234836
rect 11004 234556 11060 234612
rect 373772 234556 373828 234612
rect 373884 233884 373940 233940
rect 373436 233436 373492 233492
rect 375452 233436 375508 233492
rect 207564 233212 207620 233268
rect 442204 233212 442260 233268
rect 373660 232988 373716 233044
rect 372316 232540 372372 232596
rect 372540 232540 372596 232596
rect 441980 232540 442036 232596
rect 440524 231868 440580 231924
rect 543564 231868 543620 231924
rect 370748 231196 370804 231252
rect 375340 231196 375396 231252
rect 371756 230972 371812 231028
rect 379148 230972 379204 231028
rect 370300 230748 370356 230804
rect 377132 229852 377188 229908
rect 442428 229852 442484 229908
rect 378476 229292 378532 229348
rect 371196 229180 371252 229236
rect 372652 229180 372708 229236
rect 441868 229180 441924 229236
rect 373436 228956 373492 229012
rect 371644 228508 371700 228564
rect 380380 228508 380436 228564
rect 370412 227388 370468 227444
rect 375788 227164 375844 227220
rect 377580 227164 377636 227220
rect 374892 226492 374948 226548
rect 379260 226492 379316 226548
rect 370188 226268 370244 226324
rect 377468 225932 377524 225988
rect 376012 225260 376068 225316
rect 375228 225148 375284 225204
rect 376124 225148 376180 225204
rect 204988 225036 205044 225092
rect 373772 225036 373828 225092
rect 376124 224476 376180 224532
rect 376796 224476 376852 224532
rect 370636 224364 370692 224420
rect 370636 224028 370692 224084
rect 380268 223132 380324 223188
rect 371980 222908 372036 222964
rect 204988 222460 205044 222516
rect 369404 221788 369460 221844
rect 379708 221676 379764 221732
rect 377356 221116 377412 221172
rect 369516 220668 369572 220724
rect 380604 220444 380660 220500
rect 206668 219772 206724 219828
rect 372092 219772 372148 219828
rect 378700 219548 378756 219604
rect 372540 218652 372596 218708
rect 373884 218428 373940 218484
rect 543676 218540 543732 218596
rect 379708 217868 379764 217924
rect 379708 217308 379764 217364
rect 206668 217084 206724 217140
rect 379484 217084 379540 217140
rect 370636 216524 370692 216580
rect 373212 216524 373268 216580
rect 380380 216412 380436 216468
rect 373100 216188 373156 216244
rect 375900 215740 375956 215796
rect 379484 215740 379540 215796
rect 379260 215516 379316 215572
rect 379484 215404 379540 215460
rect 370524 215180 370580 215236
rect 373548 215180 373604 215236
rect 373324 215068 373380 215124
rect 373884 214508 373940 214564
rect 206668 214396 206724 214452
rect 373884 213948 373940 214004
rect 380268 213612 380324 213668
rect 375452 213276 375508 213332
rect 376124 213276 376180 213332
rect 380268 213164 380324 213220
rect 373884 212828 373940 212884
rect 206668 211708 206724 211764
rect 373884 211708 373940 211764
rect 373436 211596 373492 211652
rect 373660 210588 373716 210644
rect 370748 209916 370804 209972
rect 379708 209132 379764 209188
rect 380380 209132 380436 209188
rect 206668 209020 206724 209076
rect 410956 207340 411012 207396
rect 383068 207228 383124 207284
rect 399532 207116 399588 207172
rect 202412 206556 202468 206612
rect 431788 206556 431844 206612
rect 4172 206332 4228 206388
rect 375228 206332 375284 206388
rect 379372 206220 379428 206276
rect 385308 206220 385364 206276
rect 385532 206220 385588 206276
rect 403340 206108 403396 206164
rect 417004 205996 417060 206052
rect 380268 205772 380324 205828
rect 407596 205772 407652 205828
rect 381836 205660 381892 205716
rect 382060 205660 382116 205716
rect 383404 205660 383460 205716
rect 385532 205660 385588 205716
rect 442204 205660 442260 205716
rect 381164 205436 381220 205492
rect 383180 205436 383236 205492
rect 385308 205436 385364 205492
rect 414988 205436 415044 205492
rect 417004 205436 417060 205492
rect 560252 205324 560308 205380
rect 370860 205212 370916 205268
rect 386092 205212 386148 205268
rect 386764 205212 386820 205268
rect 389452 205212 389508 205268
rect 395612 205212 395668 205268
rect 431788 205212 431844 205268
rect 399532 205100 399588 205156
rect 403340 205100 403396 205156
rect 410956 205100 411012 205156
rect 431900 205100 431956 205156
rect 375452 204988 375508 205044
rect 407596 204988 407652 205044
rect 414988 204988 415044 205044
rect 431788 204204 431844 204260
rect 380492 204092 380548 204148
rect 380268 203868 380324 203924
rect 402220 203868 402276 203924
rect 204876 203644 204932 203700
rect 382620 203196 382676 203252
rect 383628 203196 383684 203252
rect 377468 202972 377524 203028
rect 382396 202972 382452 203028
rect 433580 202636 433636 202692
rect 378476 202524 378532 202580
rect 384748 202524 384804 202580
rect 390572 202524 390628 202580
rect 391020 202524 391076 202580
rect 373212 202412 373268 202468
rect 433692 202412 433748 202468
rect 377468 202300 377524 202356
rect 384076 201964 384132 202020
rect 384636 201964 384692 202020
rect 397292 201852 397348 201908
rect 377468 201628 377524 201684
rect 431900 201628 431956 201684
rect 373548 201516 373604 201572
rect 373324 201404 373380 201460
rect 384748 201404 384804 201460
rect 383852 201292 383908 201348
rect 392252 201068 392308 201124
rect 204988 200956 205044 201012
rect 373100 200844 373156 200900
rect 443772 200844 443828 200900
rect 370300 200732 370356 200788
rect 441868 200732 441924 200788
rect 445228 200508 445284 200564
rect 384748 199836 384804 199892
rect 381276 199612 381332 199668
rect 432012 199612 432068 199668
rect 436828 199500 436884 199556
rect 372092 199388 372148 199444
rect 371644 199164 371700 199220
rect 442316 199164 442372 199220
rect 206668 199052 206724 199108
rect 370412 199052 370468 199108
rect 441980 199052 442036 199108
rect 375452 198268 375508 198324
rect 380492 198268 380548 198324
rect 418348 198156 418404 198212
rect 389788 198044 389844 198100
rect 395724 197932 395780 197988
rect 383068 197820 383124 197876
rect 434252 197372 434308 197428
rect 450268 197148 450324 197204
rect 382956 196364 383012 196420
rect 371420 196028 371476 196084
rect 373660 195916 373716 195972
rect 440300 195916 440356 195972
rect 373884 195804 373940 195860
rect 443884 195804 443940 195860
rect 371980 195692 372036 195748
rect 442876 195692 442932 195748
rect 206892 195580 206948 195636
rect 381724 195132 381780 195188
rect 373772 194908 373828 194964
rect 447020 194908 447076 194964
rect 423724 194796 423780 194852
rect 373884 194684 373940 194740
rect 423332 194684 423388 194740
rect 443548 194684 443604 194740
rect 378924 194572 378980 194628
rect 373660 194348 373716 194404
rect 442428 194348 442484 194404
rect 448588 193788 448644 193844
rect 441980 193340 442036 193396
rect 205212 192892 205268 192948
rect 446908 192668 446964 192724
rect 379148 192556 379204 192612
rect 397292 192556 397348 192612
rect 433468 192444 433524 192500
rect 370188 192332 370244 192388
rect 442764 192332 442820 192388
rect 10892 192220 10948 192276
rect 548492 192108 548548 192164
rect 373660 191772 373716 191828
rect 440188 191772 440244 191828
rect 442204 191772 442260 191828
rect 445340 191548 445396 191604
rect 204988 190204 205044 190260
rect 373772 189308 373828 189364
rect 373100 188972 373156 189028
rect 373884 188188 373940 188244
rect 203420 187516 203476 187572
rect 371308 187068 371364 187124
rect 375228 186508 375284 186564
rect 373884 185948 373940 186004
rect 204988 184940 205044 184996
rect 370076 184716 370132 184772
rect 372764 184044 372820 184100
rect 375340 184044 375396 184100
rect 373660 183708 373716 183764
rect 371084 183372 371140 183428
rect 373884 183372 373940 183428
rect 203420 182812 203476 182868
rect 370860 182700 370916 182756
rect 372204 182700 372260 182756
rect 373100 182588 373156 182644
rect 372876 182028 372932 182084
rect 379708 182028 379764 182084
rect 371196 181356 371252 181412
rect 373660 180348 373716 180404
rect 204988 179452 205044 179508
rect 371084 179340 371140 179396
rect 373324 179340 373380 179396
rect 442092 179340 442148 179396
rect 373772 179228 373828 179284
rect 553532 178892 553588 178948
rect 377468 178668 377524 178724
rect 441868 178668 441924 178724
rect 375900 177996 375956 178052
rect 376236 177996 376292 178052
rect 442428 177996 442484 178052
rect 372428 177324 372484 177380
rect 375788 177324 375844 177380
rect 375900 176988 375956 177044
rect 206668 176764 206724 176820
rect 370188 176652 370244 176708
rect 372316 176652 372372 176708
rect 442540 176652 442596 176708
rect 373660 176316 373716 176372
rect 377468 175980 377524 176036
rect 442764 175980 442820 176036
rect 377580 175308 377636 175364
rect 442316 175308 442372 175364
rect 373660 174860 373716 174916
rect 371420 174636 371476 174692
rect 375564 174636 375620 174692
rect 442652 174636 442708 174692
rect 206892 174076 206948 174132
rect 208460 174076 208516 174132
rect 373548 173964 373604 174020
rect 440300 173964 440356 174020
rect 371868 173628 371924 173684
rect 441980 173292 442036 173348
rect 372652 173068 372708 173124
rect 373548 173068 373604 173124
rect 375340 172508 375396 172564
rect 204988 171388 205044 171444
rect 374892 171276 374948 171332
rect 443884 171276 443940 171332
rect 370636 170604 370692 170660
rect 371756 170604 371812 170660
rect 375116 169932 375172 169988
rect 442876 169932 442932 169988
rect 374892 169708 374948 169764
rect 376012 169708 376068 169764
rect 443772 169260 443828 169316
rect 370076 169148 370132 169204
rect 201516 168700 201572 168756
rect 375564 168028 375620 168084
rect 375676 166908 375732 166964
rect 380380 166572 380436 166628
rect 21756 165676 21812 165732
rect 26796 165676 26852 165732
rect 28476 165676 28532 165732
rect 39676 165676 39732 165732
rect 72156 165676 72212 165732
rect 82236 165676 82292 165732
rect 203308 165676 203364 165732
rect 84812 165564 84868 165620
rect 120092 165564 120148 165620
rect 122556 165564 122612 165620
rect 127596 165564 127652 165620
rect 154476 165564 154532 165620
rect 183036 165564 183092 165620
rect 184492 165564 184548 165620
rect 188972 165564 189028 165620
rect 189532 165564 189588 165620
rect 192332 165564 192388 165620
rect 189532 164892 189588 164948
rect 375788 165788 375844 165844
rect 590492 165676 590548 165732
rect 372204 164668 372260 164724
rect 94892 164556 94948 164612
rect 160524 164556 160580 164612
rect 175532 164556 175588 164612
rect 199388 164556 199444 164612
rect 172172 164444 172228 164500
rect 189420 164444 189476 164500
rect 179228 164332 179284 164388
rect 199164 164332 199220 164388
rect 210476 164220 210532 164276
rect 201852 163996 201908 164052
rect 165676 163884 165732 163940
rect 199276 163884 199332 163940
rect 108332 163772 108388 163828
rect 371980 163548 372036 163604
rect 440636 163212 440692 163268
rect 179228 163100 179284 163156
rect 199276 162988 199332 163044
rect 371308 162988 371364 163044
rect 20860 162876 20916 162932
rect 27132 162876 27188 162932
rect 126252 162876 126308 162932
rect 170492 162876 170548 162932
rect 195804 162876 195860 162932
rect 442316 162876 442372 162932
rect 157052 162764 157108 162820
rect 106652 162652 106708 162708
rect 1596 162540 1652 162596
rect 108556 162316 108612 162372
rect 379820 162540 379876 162596
rect 373548 162428 373604 162484
rect 380156 161868 380212 161924
rect 440412 161868 440468 161924
rect 199276 161308 199332 161364
rect 210588 161308 210644 161364
rect 17612 161196 17668 161252
rect 205100 161196 205156 161252
rect 210364 161084 210420 161140
rect 177212 160860 177268 160916
rect 173852 160748 173908 160804
rect 189084 160636 189140 160692
rect 205100 160636 205156 160692
rect 379596 159852 379652 159908
rect 17612 159628 17668 159684
rect 26012 159516 26068 159572
rect 181356 159516 181412 159572
rect 378812 159516 378868 159572
rect 167132 159404 167188 159460
rect 187292 159180 187348 159236
rect 380044 159180 380100 159236
rect 160412 158844 160468 158900
rect 200508 158732 200564 158788
rect 441868 158508 441924 158564
rect 380380 158060 380436 158116
rect 26012 157948 26068 158004
rect 181356 157948 181412 158004
rect 118524 157500 118580 157556
rect 73052 157388 73108 157444
rect 116732 157388 116788 157444
rect 200172 157276 200228 157332
rect 206668 157164 206724 157220
rect 379820 156492 379876 156548
rect 36876 156156 36932 156212
rect 191548 156156 191604 156212
rect 379036 155708 379092 155764
rect 116844 155596 116900 155652
rect 36876 155484 36932 155540
rect 202300 155484 202356 155540
rect 200396 155372 200452 155428
rect 373324 155372 373380 155428
rect 129052 155260 129108 155316
rect 191548 155260 191604 155316
rect 193004 155260 193060 155316
rect 373436 155148 373492 155204
rect 380604 154700 380660 154756
rect 378700 154476 378756 154532
rect 120428 153804 120484 153860
rect 118412 153692 118468 153748
rect 41132 152796 41188 152852
rect 193116 152796 193172 152852
rect 379596 152796 379652 152852
rect 376348 152684 376404 152740
rect 377132 152684 377188 152740
rect 378924 152684 378980 152740
rect 543788 152460 543844 152516
rect 377132 152348 377188 152404
rect 74732 152124 74788 152180
rect 108444 152124 108500 152180
rect 116956 152124 117012 152180
rect 202524 152012 202580 152068
rect 376348 151788 376404 151844
rect 379148 151228 379204 151284
rect 377244 151116 377300 151172
rect 379372 151116 379428 151172
rect 380604 151004 380660 151060
rect 69692 150556 69748 150612
rect 208348 150556 208404 150612
rect 200284 150444 200340 150500
rect 138684 150332 138740 150388
rect 379372 150444 379428 150500
rect 380604 149772 380660 149828
rect 103292 149660 103348 149716
rect 194460 149436 194516 149492
rect 195692 149324 195748 149380
rect 379260 149100 379316 149156
rect 137452 148988 137508 149044
rect 139356 148988 139412 149044
rect 2940 148876 2996 148932
rect 54684 148876 54740 148932
rect 194460 148764 194516 148820
rect 79772 148652 79828 148708
rect 194236 148652 194292 148708
rect 110236 148540 110292 148596
rect 112364 148540 112420 148596
rect 137452 148540 137508 148596
rect 137676 148428 137732 148484
rect 118748 148092 118804 148148
rect 119196 147980 119252 148036
rect 379148 148428 379204 148484
rect 379596 148428 379652 148484
rect 194908 148204 194964 148260
rect 72044 147868 72100 147924
rect 81452 147868 81508 147924
rect 83916 147868 83972 147924
rect 118636 147868 118692 147924
rect 126812 147868 126868 147924
rect 194908 147420 194964 147476
rect 155372 147308 155428 147364
rect 199052 147196 199108 147252
rect 150332 147084 150388 147140
rect 120316 146972 120372 147028
rect 377132 145740 377188 145796
rect 380044 145740 380100 145796
rect 121660 145404 121716 145460
rect 121772 145292 121828 145348
rect 380604 145068 380660 145124
rect 377244 143388 377300 143444
rect 379708 143388 379764 143444
rect 376348 142268 376404 142324
rect 378812 142268 378868 142324
rect 380604 141148 380660 141204
rect 543900 139244 543956 139300
rect 204204 139132 204260 139188
rect 382508 137900 382564 137956
rect 383068 137900 383124 137956
rect 379036 137340 379092 137396
rect 396844 137340 396900 137396
rect 397516 137228 397572 137284
rect 408044 137228 408100 137284
rect 393932 137116 393988 137172
rect 408156 137116 408212 137172
rect 379596 137004 379652 137060
rect 385420 136668 385476 136724
rect 387212 136556 387268 136612
rect 205996 136444 206052 136500
rect 397516 136220 397572 136276
rect 408044 136220 408100 136276
rect 396844 136108 396900 136164
rect 408156 136108 408212 136164
rect 382396 135996 382452 136052
rect 395724 135884 395780 135940
rect 7644 135772 7700 135828
rect 373772 135772 373828 135828
rect 382956 135772 383012 135828
rect 388108 135772 388164 135828
rect 382172 135660 382228 135716
rect 383628 135660 383684 135716
rect 385420 135660 385476 135716
rect 397516 135660 397572 135716
rect 385532 135548 385588 135604
rect 385756 135548 385812 135604
rect 384748 135212 384804 135268
rect 385532 135212 385588 135268
rect 440300 135212 440356 135268
rect 380044 135100 380100 135156
rect 385756 135100 385812 135156
rect 380380 134876 380436 134932
rect 377356 134764 377412 134820
rect 381612 134764 381668 134820
rect 382732 134764 382788 134820
rect 385532 134652 385588 134708
rect 377356 134540 377412 134596
rect 372316 134316 372372 134372
rect 372540 134316 372596 134372
rect 381276 134316 381332 134372
rect 380492 134092 380548 134148
rect 209692 133756 209748 133812
rect 380268 133756 380324 133812
rect 379260 133644 379316 133700
rect 373660 133532 373716 133588
rect 443772 133532 443828 133588
rect 394044 133420 394100 133476
rect 390572 132748 390628 132804
rect 376908 132636 376964 132692
rect 381388 132636 381444 132692
rect 381836 132636 381892 132692
rect 384524 132636 384580 132692
rect 383180 132524 383236 132580
rect 384972 132524 385028 132580
rect 385644 132524 385700 132580
rect 381500 132412 381556 132468
rect 386540 132524 386596 132580
rect 433692 132636 433748 132692
rect 436828 132412 436884 132468
rect 379932 132300 379988 132356
rect 390572 132300 390628 132356
rect 390796 132300 390852 132356
rect 433580 132300 433636 132356
rect 432012 132188 432068 132244
rect 431788 132076 431844 132132
rect 431900 131964 431956 132020
rect 378588 131740 378644 131796
rect 390796 131740 390852 131796
rect 386428 131628 386484 131684
rect 392252 131516 392308 131572
rect 388220 131404 388276 131460
rect 398188 131068 398244 131124
rect 395836 130956 395892 131012
rect 383068 130284 383124 130340
rect 429212 130284 429268 130340
rect 376124 130172 376180 130228
rect 375228 129276 375284 129332
rect 375340 129164 375396 129220
rect 376124 129164 376180 129220
rect 389788 129164 389844 129220
rect 384748 128940 384804 128996
rect 390012 128940 390068 128996
rect 392476 128940 392532 128996
rect 381388 128828 381444 128884
rect 388332 128828 388388 128884
rect 408156 128828 408212 128884
rect 433468 128828 433524 128884
rect 373324 128492 373380 128548
rect 209468 128380 209524 128436
rect 381724 127932 381780 127988
rect 370524 127596 370580 127652
rect 370748 127148 370804 127204
rect 408044 127036 408100 127092
rect 431788 127036 431844 127092
rect 375900 126924 375956 126980
rect 441868 126924 441924 126980
rect 373548 126812 373604 126868
rect 440412 126812 440468 126868
rect 572012 126028 572068 126084
rect 381948 125916 382004 125972
rect 204092 125692 204148 125748
rect 384524 125468 384580 125524
rect 393148 125468 393204 125524
rect 392364 125356 392420 125412
rect 381948 124460 382004 124516
rect 429212 124236 429268 124292
rect 382284 124012 382340 124068
rect 390572 124012 390628 124068
rect 371868 123564 371924 123620
rect 442204 123564 442260 123620
rect 209244 123004 209300 123060
rect 205884 120316 205940 120372
rect 373884 119868 373940 119924
rect 380156 117628 380212 117684
rect 372540 116508 372596 116564
rect 379596 116284 379652 116340
rect 370300 115388 370356 115444
rect 373548 114940 373604 114996
rect 380380 114940 380436 114996
rect 373548 114268 373604 114324
rect 372316 113148 372372 113204
rect 546812 112812 546868 112868
rect 375340 112028 375396 112084
rect 375340 111020 375396 111076
rect 375900 111020 375956 111076
rect 7532 107436 7588 107492
rect 209132 104188 209188 104244
rect 376124 104188 376180 104244
rect 377580 101948 377636 102004
rect 590156 99596 590212 99652
rect 370636 99036 370692 99092
rect 373100 99036 373156 99092
rect 551852 98252 551908 98308
rect 590156 98252 590212 98308
rect 373772 98140 373828 98196
rect 373100 97468 373156 97524
rect 372428 96124 372484 96180
rect 373548 95676 373604 95732
rect 370860 95452 370916 95508
rect 376012 94780 376068 94836
rect 372876 94444 372932 94500
rect 372988 94220 373044 94276
rect 370412 94108 370468 94164
rect 372876 93772 372932 93828
rect 4284 93436 4340 93492
rect 371980 93436 372036 93492
rect 372204 92764 372260 92820
rect 375788 92092 375844 92148
rect 443772 91420 443828 91476
rect 375228 90748 375284 90804
rect 376124 90748 376180 90804
rect 443660 90748 443716 90804
rect 447020 90076 447076 90132
rect 373100 89628 373156 89684
rect 376012 88508 376068 88564
rect 443548 88732 443604 88788
rect 370188 88284 370244 88340
rect 370860 88284 370916 88340
rect 375676 88060 375732 88116
rect 445340 88060 445396 88116
rect 370860 87388 370916 87444
rect 372876 87388 372932 87444
rect 374780 87388 374836 87444
rect 376460 87164 376516 87220
rect 450268 86716 450324 86772
rect 556892 86380 556948 86436
rect 373772 86268 373828 86324
rect 371084 86044 371140 86100
rect 371308 86044 371364 86100
rect 446908 86044 446964 86100
rect 372652 85596 372708 85652
rect 205772 85372 205828 85428
rect 371196 85372 371252 85428
rect 448588 85372 448644 85428
rect 372988 85148 373044 85204
rect 377356 84700 377412 84756
rect 441980 84028 442036 84084
rect 372092 83356 372148 83412
rect 199052 82684 199108 82740
rect 440300 82684 440356 82740
rect 440188 82012 440244 82068
rect 378812 81788 378868 81844
rect 375452 81340 375508 81396
rect 378812 80780 378868 80836
rect 442204 80668 442260 80724
rect 445228 79996 445284 80052
rect 378812 79548 378868 79604
rect 4172 79324 4228 79380
rect 377580 79324 377636 79380
rect 440412 79324 440468 79380
rect 370076 78652 370132 78708
rect 378812 78428 378868 78484
rect 378812 77308 378868 77364
rect 379484 77308 379540 77364
rect 375564 76636 375620 76692
rect 441868 76636 441924 76692
rect 379596 76188 379652 76244
rect 376236 75964 376292 76020
rect 380156 75292 380212 75348
rect 379596 75068 379652 75124
rect 372540 74620 372596 74676
rect 378588 74060 378644 74116
rect 545132 73164 545188 73220
rect 378812 72828 378868 72884
rect 370300 72604 370356 72660
rect 376460 72156 376516 72212
rect 377580 71708 377636 71764
rect 513212 70588 513268 70644
rect 372316 69916 372372 69972
rect 375900 69244 375956 69300
rect 530012 68572 530068 68628
rect 379932 66108 379988 66164
rect 379932 65548 379988 65604
rect 377580 64988 377636 65044
rect 377580 63868 377636 63924
rect 377580 62748 377636 62804
rect 372428 61628 372484 61684
rect 544012 59948 544068 60004
rect 207676 58492 207732 58548
rect 209916 57820 209972 57876
rect 374780 57148 374836 57204
rect 371308 56028 371364 56084
rect 376348 54908 376404 54964
rect 377132 53788 377188 53844
rect 207452 53116 207508 53172
rect 376236 52108 376292 52164
rect 370412 51548 370468 51604
rect 140 51212 196 51268
rect 394044 47964 394100 48020
rect 403564 47964 403620 48020
rect 379372 47852 379428 47908
rect 417676 47852 417732 47908
rect 208124 47740 208180 47796
rect 394828 46956 394884 47012
rect 590604 46732 590660 46788
rect 396844 46284 396900 46340
rect 398188 46172 398244 46228
rect 393820 45948 393876 46004
rect 385532 45836 385588 45892
rect 381388 45724 381444 45780
rect 381612 45724 381668 45780
rect 383068 45724 383124 45780
rect 385644 45724 385700 45780
rect 389788 45724 389844 45780
rect 378812 45500 378868 45556
rect 381500 45500 381556 45556
rect 383852 45500 383908 45556
rect 384972 45500 385028 45556
rect 386428 45500 386484 45556
rect 386988 45500 387044 45556
rect 388332 45500 388388 45556
rect 391468 45500 391524 45556
rect 396844 45724 396900 45780
rect 398188 45724 398244 45780
rect 403564 45724 403620 45780
rect 417676 45724 417732 45780
rect 393820 45500 393876 45556
rect 388108 45388 388164 45444
rect 389900 45164 389956 45220
rect 392252 45164 392308 45220
rect 395724 45164 395780 45220
rect 380604 44940 380660 44996
rect 385756 44380 385812 44436
rect 385756 44156 385812 44212
rect 395836 43596 395892 43652
rect 419692 43596 419748 43652
rect 429212 43596 429268 43652
rect 394156 43484 394212 43540
rect 431788 43484 431844 43540
rect 390572 43372 390628 43428
rect 393932 43260 393988 43316
rect 433468 43148 433524 43204
rect 396396 42924 396452 42980
rect 378700 42812 378756 42868
rect 387212 41692 387268 41748
rect 379820 40236 379876 40292
rect 110012 36764 110068 36820
rect 550284 33628 550340 33684
rect 543452 32844 543508 32900
rect 563612 31724 563668 31780
rect 565292 30604 565348 30660
rect 550172 29484 550228 29540
rect 544236 29372 544292 29428
rect 587132 29372 587188 29428
rect 555212 28364 555268 28420
rect 544236 27244 544292 27300
rect 543564 26124 543620 26180
rect 543676 25004 543732 25060
rect 544348 24332 544404 24388
rect 590492 24332 590548 24388
rect 560252 23884 560308 23940
rect 28 22988 84 23044
rect 548492 22764 548548 22820
rect 553532 21644 553588 21700
rect 544348 20524 544404 20580
rect 591276 20300 591332 20356
rect 543788 19404 543844 19460
rect 548492 19292 548548 19348
rect 591276 19292 591332 19348
rect 543900 18284 543956 18340
rect 572012 17164 572068 17220
rect 546812 16044 546868 16100
rect 551852 14924 551908 14980
rect 556892 13804 556948 13860
rect 545132 12684 545188 12740
rect 544348 12572 544404 12628
rect 590604 12572 590660 12628
rect 544012 11564 544068 11620
rect 544348 10444 544404 10500
rect 550284 9324 550340 9380
rect 548492 8204 548548 8260
rect 442988 5068 443044 5124
rect 498988 5068 499044 5124
rect 494956 3388 495012 3444
rect 498988 3388 499044 3444
rect 529228 3388 529284 3444
rect 557788 3388 557844 3444
rect 565404 3388 565460 3444
rect 447692 3276 447748 3332
rect 475468 3276 475524 3332
rect 499436 3276 499492 3332
rect 501676 3276 501732 3332
rect 457100 2940 457156 2996
rect 504140 2492 504196 2548
rect 510748 2492 510804 2548
rect 436828 1820 436884 1876
rect 563500 1708 563556 1764
rect 487676 1148 487732 1204
rect 512092 700 512148 756
rect 569212 588 569268 644
rect 571228 588 571284 644
rect 436828 140 436884 196
rect 487676 252 487732 308
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect 5418 597212 6038 598268
rect 5418 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 6038 597212
rect 5418 597088 6038 597156
rect 5418 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 6038 597088
rect 5418 596964 6038 597032
rect 5418 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 6038 596964
rect 5418 596840 6038 596908
rect 5418 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 6038 596840
rect 5418 580350 6038 596784
rect 5418 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 6038 580350
rect 5418 580226 6038 580294
rect 5418 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 6038 580226
rect 5418 580102 6038 580170
rect 5418 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 6038 580102
rect 5418 579978 6038 580046
rect 5418 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 6038 579978
rect 5418 562350 6038 579922
rect 5418 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 6038 562350
rect 5418 562226 6038 562294
rect 5418 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 6038 562226
rect 5418 562102 6038 562170
rect 5418 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 6038 562102
rect 5418 561978 6038 562046
rect 5418 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 6038 561978
rect 5418 544350 6038 561922
rect 5418 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 6038 544350
rect 5418 544226 6038 544294
rect 5418 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 6038 544226
rect 5418 544102 6038 544170
rect 5418 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 6038 544102
rect 5418 543978 6038 544046
rect 5418 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 6038 543978
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect 2492 530740 2548 530750
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect 28 516516 84 516526
rect 28 273538 84 516460
rect 1484 469700 1540 469710
rect 28 273472 84 273482
rect 140 403620 196 403630
rect 140 271918 196 403564
rect 1484 284788 1540 469644
rect 1484 284722 1540 284732
rect 1596 361378 1652 361388
rect 140 271852 196 271862
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect 28 267958 84 267968
rect 28 23044 84 267902
rect 140 266518 196 266528
rect 140 51268 196 266462
rect 1596 162596 1652 361322
rect 2492 273718 2548 530684
rect 5418 526350 6038 543922
rect 5418 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 6038 526350
rect 5418 526226 6038 526294
rect 5418 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 6038 526226
rect 5418 526102 6038 526170
rect 5418 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 6038 526102
rect 5418 525978 6038 526046
rect 5418 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 6038 525978
rect 5418 508350 6038 525922
rect 5418 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 6038 508350
rect 5418 508226 6038 508294
rect 5418 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 6038 508226
rect 5418 508102 6038 508170
rect 5418 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 6038 508102
rect 5418 507978 6038 508046
rect 5418 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 6038 507978
rect 5418 490350 6038 507922
rect 5418 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 6038 490350
rect 5418 490226 6038 490294
rect 5418 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 6038 490226
rect 5418 490102 6038 490170
rect 5418 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 6038 490102
rect 5418 489978 6038 490046
rect 5418 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 6038 489978
rect 4172 488404 4228 488414
rect 3164 403620 3220 403630
rect 2492 273652 2548 273662
rect 2940 366418 2996 366428
rect 1596 162530 1652 162540
rect 2940 148932 2996 366362
rect 3052 332038 3108 332048
rect 3052 310996 3108 331982
rect 3052 310930 3108 310940
rect 3052 297556 3108 297566
rect 3052 281638 3108 297500
rect 3052 281572 3108 281582
rect 3164 280532 3220 403564
rect 3164 280466 3220 280476
rect 4172 270298 4228 488348
rect 5418 472350 6038 489922
rect 5418 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 6038 472350
rect 5418 472226 6038 472294
rect 5418 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 6038 472226
rect 5418 472102 6038 472170
rect 5418 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 6038 472102
rect 5418 471978 6038 472046
rect 5418 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 6038 471978
rect 5418 454350 6038 471922
rect 5418 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 6038 454350
rect 5418 454226 6038 454294
rect 5418 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 6038 454226
rect 5418 454102 6038 454170
rect 5418 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 6038 454102
rect 5418 453978 6038 454046
rect 5418 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 6038 453978
rect 4396 446068 4452 446078
rect 4284 333172 4340 333182
rect 4284 272098 4340 333116
rect 4284 272032 4340 272042
rect 4396 270478 4452 446012
rect 5418 436350 6038 453922
rect 5418 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 6038 436350
rect 5418 436226 6038 436294
rect 5418 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 6038 436226
rect 5418 436102 6038 436170
rect 5418 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 6038 436102
rect 5418 435978 6038 436046
rect 5418 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 6038 435978
rect 5418 418350 6038 435922
rect 5418 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 6038 418350
rect 5418 418226 6038 418294
rect 5418 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 6038 418226
rect 5418 418102 6038 418170
rect 5418 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 6038 418102
rect 5418 417978 6038 418046
rect 5418 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 6038 417978
rect 5418 400350 6038 417922
rect 5418 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 6038 400350
rect 5418 400226 6038 400294
rect 5418 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 6038 400226
rect 5418 400102 6038 400170
rect 5418 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 6038 400102
rect 5418 399978 6038 400046
rect 5418 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 6038 399978
rect 5418 382350 6038 399922
rect 5418 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 6038 382350
rect 5418 382226 6038 382294
rect 5418 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 6038 382226
rect 5418 382102 6038 382170
rect 5418 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 6038 382102
rect 5418 381978 6038 382046
rect 5418 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 6038 381978
rect 5418 364350 6038 381922
rect 5418 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 6038 364350
rect 5418 364226 6038 364294
rect 5418 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 6038 364226
rect 5418 364102 6038 364170
rect 5418 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 6038 364102
rect 5418 363978 6038 364046
rect 5418 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 6038 363978
rect 5418 346350 6038 363922
rect 5418 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 6038 346350
rect 5418 346226 6038 346294
rect 5418 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 6038 346226
rect 5418 346102 6038 346170
rect 5418 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 6038 346102
rect 5418 345978 6038 346046
rect 5418 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 6038 345978
rect 5068 331858 5124 331868
rect 4956 324660 5012 324670
rect 4732 290836 4788 290846
rect 4732 290742 4788 290762
rect 4956 278038 5012 324604
rect 5068 318388 5124 331802
rect 5418 328350 6038 345922
rect 9138 598172 9758 598268
rect 9138 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 9758 598172
rect 9138 598048 9758 598116
rect 9138 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 9758 598048
rect 9138 597924 9758 597992
rect 9138 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 9758 597924
rect 9138 597800 9758 597868
rect 9138 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 9758 597800
rect 9138 586350 9758 597744
rect 9138 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 9758 586350
rect 9138 586226 9758 586294
rect 9138 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 9758 586226
rect 9138 586102 9758 586170
rect 9138 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 9758 586102
rect 9138 585978 9758 586046
rect 9138 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 9758 585978
rect 9138 568350 9758 585922
rect 9138 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 9758 568350
rect 9138 568226 9758 568294
rect 9138 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 9758 568226
rect 9138 568102 9758 568170
rect 9138 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 9758 568102
rect 9138 567978 9758 568046
rect 9138 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 9758 567978
rect 9138 550350 9758 567922
rect 9138 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 9758 550350
rect 9138 550226 9758 550294
rect 9138 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 9758 550226
rect 9138 550102 9758 550170
rect 9138 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 9758 550102
rect 9138 549978 9758 550046
rect 9138 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 9758 549978
rect 9138 532350 9758 549922
rect 9138 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 9758 532350
rect 9138 532226 9758 532294
rect 9138 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 9758 532226
rect 9138 532102 9758 532170
rect 9138 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 9758 532102
rect 9138 531978 9758 532046
rect 9138 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 9758 531978
rect 9138 514350 9758 531922
rect 9138 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 9758 514350
rect 9138 514226 9758 514294
rect 9138 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 9758 514226
rect 9138 514102 9758 514170
rect 9138 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 9758 514102
rect 9138 513978 9758 514046
rect 9138 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 9758 513978
rect 9138 496350 9758 513922
rect 9138 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 9758 496350
rect 9138 496226 9758 496294
rect 9138 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 9758 496226
rect 9138 496102 9758 496170
rect 9138 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 9758 496102
rect 9138 495978 9758 496046
rect 9138 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 9758 495978
rect 9138 478350 9758 495922
rect 9138 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 9758 478350
rect 9138 478226 9758 478294
rect 9138 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 9758 478226
rect 9138 478102 9758 478170
rect 9138 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 9758 478102
rect 9138 477978 9758 478046
rect 9138 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 9758 477978
rect 9138 460350 9758 477922
rect 9138 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 9758 460350
rect 9138 460226 9758 460294
rect 9138 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 9758 460226
rect 9138 460102 9758 460170
rect 9138 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 9758 460102
rect 9138 459978 9758 460046
rect 9138 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 9758 459978
rect 9138 442350 9758 459922
rect 9138 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 9758 442350
rect 9138 442226 9758 442294
rect 9138 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 9758 442226
rect 9138 442102 9758 442170
rect 9138 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 9758 442102
rect 9138 441978 9758 442046
rect 9138 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 9758 441978
rect 9138 424350 9758 441922
rect 9138 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 9758 424350
rect 9138 424226 9758 424294
rect 9138 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 9758 424226
rect 9138 424102 9758 424170
rect 9138 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 9758 424102
rect 9138 423978 9758 424046
rect 9138 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 9758 423978
rect 9138 406350 9758 423922
rect 9138 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 9758 406350
rect 9138 406226 9758 406294
rect 9138 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 9758 406226
rect 9138 406102 9758 406170
rect 9138 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 9758 406102
rect 9138 405978 9758 406046
rect 9138 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 9758 405978
rect 9138 388350 9758 405922
rect 9138 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 9758 388350
rect 9138 388226 9758 388294
rect 9138 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 9758 388226
rect 9138 388102 9758 388170
rect 9138 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 9758 388102
rect 9138 387978 9758 388046
rect 9138 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 9758 387978
rect 9138 370350 9758 387922
rect 9138 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 9758 370350
rect 9138 370226 9758 370294
rect 9138 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 9758 370226
rect 9138 370102 9758 370170
rect 9138 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 9758 370102
rect 9138 369978 9758 370046
rect 9138 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 9758 369978
rect 9138 352350 9758 369922
rect 9138 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 9758 352350
rect 9138 352226 9758 352294
rect 9138 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 9758 352226
rect 9138 352102 9758 352170
rect 9138 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 9758 352102
rect 9138 351978 9758 352046
rect 9138 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 9758 351978
rect 5418 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 6038 328350
rect 5418 328226 6038 328294
rect 5418 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 6038 328226
rect 5418 328102 6038 328170
rect 5418 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 6038 328102
rect 5418 327978 6038 328046
rect 5418 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 6038 327978
rect 5292 325018 5348 325028
rect 5292 324884 5348 324962
rect 5292 324818 5348 324828
rect 5068 318322 5124 318332
rect 5418 310350 6038 327922
rect 5418 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 6038 310350
rect 5418 310226 6038 310294
rect 5418 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 6038 310226
rect 5418 310102 6038 310170
rect 5418 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 6038 310102
rect 5418 309978 6038 310046
rect 5418 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 6038 309978
rect 5292 308998 5348 309008
rect 5292 308756 5348 308942
rect 5292 308690 5348 308700
rect 5418 292350 6038 309922
rect 7532 335188 7588 335198
rect 7532 308998 7588 335132
rect 9138 334350 9758 351922
rect 9138 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 9758 334350
rect 9138 334226 9758 334294
rect 9138 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 9758 334226
rect 9138 334102 9758 334170
rect 9138 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 9758 334102
rect 9138 333978 9758 334046
rect 9138 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 9758 333978
rect 9138 328428 9758 333922
rect 36138 597212 36758 598268
rect 36138 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 36758 597212
rect 36138 597088 36758 597156
rect 36138 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 36758 597088
rect 36138 596964 36758 597032
rect 36138 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 36758 596964
rect 36138 596840 36758 596908
rect 36138 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 36758 596840
rect 36138 580350 36758 596784
rect 36138 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 36758 580350
rect 36138 580226 36758 580294
rect 36138 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 36758 580226
rect 36138 580102 36758 580170
rect 36138 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 36758 580102
rect 36138 579978 36758 580046
rect 36138 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 36758 579978
rect 36138 562350 36758 579922
rect 36138 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 36758 562350
rect 36138 562226 36758 562294
rect 36138 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 36758 562226
rect 36138 562102 36758 562170
rect 36138 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 36758 562102
rect 36138 561978 36758 562046
rect 36138 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 36758 561978
rect 36138 544350 36758 561922
rect 36138 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 36758 544350
rect 36138 544226 36758 544294
rect 36138 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 36758 544226
rect 36138 544102 36758 544170
rect 36138 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 36758 544102
rect 36138 543978 36758 544046
rect 36138 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 36758 543978
rect 36138 526350 36758 543922
rect 36138 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 36758 526350
rect 36138 526226 36758 526294
rect 36138 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 36758 526226
rect 36138 526102 36758 526170
rect 36138 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 36758 526102
rect 36138 525978 36758 526046
rect 36138 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 36758 525978
rect 36138 508350 36758 525922
rect 36138 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 36758 508350
rect 36138 508226 36758 508294
rect 36138 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 36758 508226
rect 36138 508102 36758 508170
rect 36138 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 36758 508102
rect 36138 507978 36758 508046
rect 36138 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 36758 507978
rect 36138 490350 36758 507922
rect 36138 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 36758 490350
rect 36138 490226 36758 490294
rect 36138 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 36758 490226
rect 36138 490102 36758 490170
rect 36138 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 36758 490102
rect 36138 489978 36758 490046
rect 36138 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 36758 489978
rect 36138 472350 36758 489922
rect 36138 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 36758 472350
rect 36138 472226 36758 472294
rect 36138 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 36758 472226
rect 36138 472102 36758 472170
rect 36138 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 36758 472102
rect 36138 471978 36758 472046
rect 36138 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 36758 471978
rect 36138 454350 36758 471922
rect 36138 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 36758 454350
rect 36138 454226 36758 454294
rect 36138 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 36758 454226
rect 36138 454102 36758 454170
rect 36138 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 36758 454102
rect 36138 453978 36758 454046
rect 36138 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 36758 453978
rect 36138 436350 36758 453922
rect 36138 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 36758 436350
rect 36138 436226 36758 436294
rect 36138 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 36758 436226
rect 36138 436102 36758 436170
rect 36138 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 36758 436102
rect 36138 435978 36758 436046
rect 36138 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 36758 435978
rect 36138 418350 36758 435922
rect 36138 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 36758 418350
rect 36138 418226 36758 418294
rect 36138 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 36758 418226
rect 36138 418102 36758 418170
rect 36138 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 36758 418102
rect 36138 417978 36758 418046
rect 36138 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 36758 417978
rect 36138 400350 36758 417922
rect 36138 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 36758 400350
rect 36138 400226 36758 400294
rect 36138 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 36758 400226
rect 36138 400102 36758 400170
rect 36138 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 36758 400102
rect 36138 399978 36758 400046
rect 36138 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 36758 399978
rect 36138 382350 36758 399922
rect 36138 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 36758 382350
rect 36138 382226 36758 382294
rect 36138 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 36758 382226
rect 36138 382102 36758 382170
rect 36138 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 36758 382102
rect 36138 381978 36758 382046
rect 36138 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 36758 381978
rect 36138 364350 36758 381922
rect 36138 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 36758 364350
rect 36138 364226 36758 364294
rect 36138 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 36758 364226
rect 36138 364102 36758 364170
rect 36138 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 36758 364102
rect 36138 363978 36758 364046
rect 36138 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 36758 363978
rect 36138 346350 36758 363922
rect 36138 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 36758 346350
rect 36138 346226 36758 346294
rect 36138 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 36758 346226
rect 36138 346102 36758 346170
rect 36138 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 36758 346102
rect 36138 345978 36758 346046
rect 36138 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 36758 345978
rect 36138 328350 36758 345922
rect 39858 598172 40478 598268
rect 39858 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 40478 598172
rect 39858 598048 40478 598116
rect 39858 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 40478 598048
rect 39858 597924 40478 597992
rect 39858 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 40478 597924
rect 39858 597800 40478 597868
rect 39858 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 40478 597800
rect 39858 586350 40478 597744
rect 66858 597212 67478 598268
rect 66858 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 67478 597212
rect 66858 597088 67478 597156
rect 66858 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 67478 597088
rect 66858 596964 67478 597032
rect 66858 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 67478 596964
rect 66858 596840 67478 596908
rect 66858 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 67478 596840
rect 39858 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 40478 586350
rect 39858 586226 40478 586294
rect 39858 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 40478 586226
rect 39858 586102 40478 586170
rect 39858 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 40478 586102
rect 39858 585978 40478 586046
rect 39858 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 40478 585978
rect 39858 568350 40478 585922
rect 39858 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 40478 568350
rect 39858 568226 40478 568294
rect 39858 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 40478 568226
rect 39858 568102 40478 568170
rect 39858 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 40478 568102
rect 39858 567978 40478 568046
rect 39858 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 40478 567978
rect 39858 550350 40478 567922
rect 39858 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 40478 550350
rect 39858 550226 40478 550294
rect 39858 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 40478 550226
rect 39858 550102 40478 550170
rect 39858 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 40478 550102
rect 39858 549978 40478 550046
rect 39858 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 40478 549978
rect 39858 532350 40478 549922
rect 39858 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532294 40478 532350
rect 39858 532226 40478 532294
rect 39858 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 40478 532226
rect 39858 532102 40478 532170
rect 39858 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 40478 532102
rect 39858 531978 40478 532046
rect 39858 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531922 40478 531978
rect 39858 514350 40478 531922
rect 39858 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 40478 514350
rect 39858 514226 40478 514294
rect 39858 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 40478 514226
rect 39858 514102 40478 514170
rect 39858 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 40478 514102
rect 39858 513978 40478 514046
rect 39858 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 40478 513978
rect 39858 496350 40478 513922
rect 39858 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 40478 496350
rect 39858 496226 40478 496294
rect 39858 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 40478 496226
rect 39858 496102 40478 496170
rect 52892 590548 52948 590558
rect 39858 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496046 40478 496102
rect 39858 495978 40478 496046
rect 39858 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495922 40478 495978
rect 39858 478350 40478 495922
rect 39858 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 40478 478350
rect 39858 478226 40478 478294
rect 39858 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 40478 478226
rect 39858 478102 40478 478170
rect 39858 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 40478 478102
rect 39858 477978 40478 478046
rect 39858 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 40478 477978
rect 39858 460350 40478 477922
rect 39858 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 40478 460350
rect 39858 460226 40478 460294
rect 39858 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 40478 460226
rect 39858 460102 40478 460170
rect 39858 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 40478 460102
rect 39858 459978 40478 460046
rect 39858 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 40478 459978
rect 39858 442350 40478 459922
rect 39858 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 40478 442350
rect 39858 442226 40478 442294
rect 39858 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 40478 442226
rect 39858 442102 40478 442170
rect 39858 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 40478 442102
rect 39858 441978 40478 442046
rect 39858 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 40478 441978
rect 39858 424350 40478 441922
rect 39858 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 40478 424350
rect 39858 424226 40478 424294
rect 39858 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 40478 424226
rect 39858 424102 40478 424170
rect 39858 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 40478 424102
rect 39858 423978 40478 424046
rect 39858 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 40478 423978
rect 39858 406350 40478 423922
rect 39858 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 40478 406350
rect 39858 406226 40478 406294
rect 39858 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 40478 406226
rect 39858 406102 40478 406170
rect 39858 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 40478 406102
rect 39858 405978 40478 406046
rect 39858 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 40478 405978
rect 39858 388350 40478 405922
rect 39858 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 40478 388350
rect 39858 388226 40478 388294
rect 39858 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 40478 388226
rect 39858 388102 40478 388170
rect 39858 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 40478 388102
rect 39858 387978 40478 388046
rect 39858 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 40478 387978
rect 39858 370350 40478 387922
rect 39858 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 40478 370350
rect 39858 370226 40478 370294
rect 39858 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 40478 370226
rect 39858 370102 40478 370170
rect 39858 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 40478 370102
rect 39858 369978 40478 370046
rect 39858 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 40478 369978
rect 39858 352350 40478 369922
rect 39858 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 40478 352350
rect 39858 352226 40478 352294
rect 39858 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 40478 352226
rect 39858 352102 40478 352170
rect 39858 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 40478 352102
rect 39858 351978 40478 352046
rect 39858 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 40478 351978
rect 39858 334350 40478 351922
rect 39858 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 40478 334350
rect 39858 334226 40478 334294
rect 39858 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 40478 334226
rect 39858 334102 40478 334170
rect 39858 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 40478 334102
rect 39858 333978 40478 334046
rect 39858 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 40478 333978
rect 39858 328428 40478 333922
rect 49532 496132 49588 496142
rect 36138 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 36758 328350
rect 36138 328226 36758 328294
rect 36138 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 36758 328226
rect 36138 328102 36758 328170
rect 36138 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 36758 328102
rect 36138 327978 36758 328046
rect 36138 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 36758 327978
rect 36138 326670 36758 327922
rect 24808 316350 25128 316384
rect 24808 316294 24878 316350
rect 24934 316294 25002 316350
rect 25058 316294 25128 316350
rect 24808 316226 25128 316294
rect 24808 316170 24878 316226
rect 24934 316170 25002 316226
rect 25058 316170 25128 316226
rect 24808 316102 25128 316170
rect 24808 316046 24878 316102
rect 24934 316046 25002 316102
rect 25058 316046 25128 316102
rect 24808 315978 25128 316046
rect 24808 315922 24878 315978
rect 24934 315922 25002 315978
rect 25058 315922 25128 315978
rect 24808 315888 25128 315922
rect 9448 310350 9768 310384
rect 9448 310294 9518 310350
rect 9574 310294 9642 310350
rect 9698 310294 9768 310350
rect 9448 310226 9768 310294
rect 9448 310170 9518 310226
rect 9574 310170 9642 310226
rect 9698 310170 9768 310226
rect 9448 310102 9768 310170
rect 9448 310046 9518 310102
rect 9574 310046 9642 310102
rect 9698 310046 9768 310102
rect 9448 309978 9768 310046
rect 9448 309922 9518 309978
rect 9574 309922 9642 309978
rect 9698 309922 9768 309978
rect 9448 309888 9768 309922
rect 40168 310350 40488 310384
rect 40168 310294 40238 310350
rect 40294 310294 40362 310350
rect 40418 310294 40488 310350
rect 40168 310226 40488 310294
rect 40168 310170 40238 310226
rect 40294 310170 40362 310226
rect 40418 310170 40488 310226
rect 40168 310102 40488 310170
rect 40168 310046 40238 310102
rect 40294 310046 40362 310102
rect 40418 310046 40488 310102
rect 40168 309978 40488 310046
rect 40168 309922 40238 309978
rect 40294 309922 40362 309978
rect 40418 309922 40488 309978
rect 40168 309888 40488 309922
rect 7532 308932 7588 308942
rect 24808 298350 25128 298384
rect 24808 298294 24878 298350
rect 24934 298294 25002 298350
rect 25058 298294 25128 298350
rect 24808 298226 25128 298294
rect 24808 298170 24878 298226
rect 24934 298170 25002 298226
rect 25058 298170 25128 298226
rect 24808 298102 25128 298170
rect 24808 298046 24878 298102
rect 24934 298046 25002 298102
rect 25058 298046 25128 298102
rect 24808 297978 25128 298046
rect 24808 297922 24878 297978
rect 24934 297922 25002 297978
rect 25058 297922 25128 297978
rect 24808 297888 25128 297922
rect 5418 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 6038 292350
rect 5418 292226 6038 292294
rect 5418 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 6038 292226
rect 5418 292102 6038 292170
rect 5418 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 6038 292102
rect 5418 291978 6038 292046
rect 5418 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 6038 291978
rect 5180 285460 5236 285470
rect 5180 281458 5236 285404
rect 5292 283444 5348 283454
rect 5292 281818 5348 283388
rect 5292 281752 5348 281762
rect 5292 281458 5348 281468
rect 5180 281402 5292 281458
rect 5292 281392 5348 281402
rect 4956 277972 5012 277982
rect 4396 270412 4452 270422
rect 5418 274350 6038 291922
rect 9448 292350 9768 292384
rect 9448 292294 9518 292350
rect 9574 292294 9642 292350
rect 9698 292294 9768 292350
rect 9448 292226 9768 292294
rect 9448 292170 9518 292226
rect 9574 292170 9642 292226
rect 9698 292170 9768 292226
rect 9448 292102 9768 292170
rect 9448 292046 9518 292102
rect 9574 292046 9642 292102
rect 9698 292046 9768 292102
rect 9448 291978 9768 292046
rect 9448 291922 9518 291978
rect 9574 291922 9642 291978
rect 9698 291922 9768 291978
rect 9448 291888 9768 291922
rect 40168 292350 40488 292384
rect 40168 292294 40238 292350
rect 40294 292294 40362 292350
rect 40418 292294 40488 292350
rect 40168 292226 40488 292294
rect 40168 292170 40238 292226
rect 40294 292170 40362 292226
rect 40418 292170 40488 292226
rect 40168 292102 40488 292170
rect 40168 292046 40238 292102
rect 40294 292046 40362 292102
rect 40418 292046 40488 292102
rect 40168 291978 40488 292046
rect 40168 291922 40238 291978
rect 40294 291922 40362 291978
rect 40418 291922 40488 291978
rect 40168 291888 40488 291922
rect 7644 290818 7700 290828
rect 7532 282324 7588 282334
rect 7084 277172 7140 277182
rect 7084 275518 7140 277116
rect 7084 275452 7140 275462
rect 5418 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 6038 274350
rect 5418 274226 6038 274294
rect 5418 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 6038 274226
rect 5418 274102 6038 274170
rect 5418 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 6038 274102
rect 5418 273978 6038 274046
rect 5418 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 6038 273978
rect 4172 270232 4228 270242
rect 4284 268318 4340 268328
rect 4172 266698 4228 266708
rect 4172 208348 4228 266642
rect 4060 208292 4228 208348
rect 4060 196588 4116 208292
rect 4172 206578 4228 206588
rect 4172 206388 4228 206522
rect 4172 206322 4228 206332
rect 4060 196532 4228 196588
rect 2940 148866 2996 148876
rect 4172 79380 4228 196532
rect 4284 93492 4340 268262
rect 4956 257878 5012 257888
rect 4956 248612 5012 257822
rect 4956 248546 5012 248556
rect 5418 256350 6038 273922
rect 7532 271124 7588 282268
rect 7532 271058 7588 271068
rect 7644 270452 7700 290762
rect 40684 281764 40740 281774
rect 25900 281652 25956 281662
rect 9138 280350 9758 280964
rect 25900 280532 25956 281596
rect 25900 280466 25956 280476
rect 26572 281540 26628 281550
rect 26572 280532 26628 281484
rect 26572 280466 26628 280476
rect 9138 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 9758 280350
rect 9138 280226 9758 280294
rect 9138 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 9758 280226
rect 9138 280102 9758 280170
rect 9138 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 9758 280102
rect 9138 279978 9758 280046
rect 9138 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 9758 279978
rect 7756 277318 7812 277328
rect 7756 277172 7812 277262
rect 7756 277106 7812 277116
rect 7644 270386 7700 270396
rect 5418 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 6038 256350
rect 5418 256226 6038 256294
rect 5418 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 6038 256226
rect 5418 256102 6038 256170
rect 5418 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 6038 256102
rect 5418 255978 6038 256046
rect 5418 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 6038 255978
rect 4284 93426 4340 93436
rect 5418 238350 6038 255922
rect 5418 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 6038 238350
rect 5418 238226 6038 238294
rect 5418 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 6038 238226
rect 5418 238102 6038 238170
rect 5418 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 6038 238102
rect 5418 237978 6038 238046
rect 5418 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 6038 237978
rect 5418 220350 6038 237922
rect 5418 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 6038 220350
rect 5418 220226 6038 220294
rect 5418 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 6038 220226
rect 5418 220102 6038 220170
rect 5418 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 6038 220102
rect 5418 219978 6038 220046
rect 5418 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 6038 219978
rect 5418 202350 6038 219922
rect 5418 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 6038 202350
rect 5418 202226 6038 202294
rect 5418 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 6038 202226
rect 5418 202102 6038 202170
rect 5418 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 6038 202102
rect 5418 201978 6038 202046
rect 5418 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 6038 201978
rect 5418 184350 6038 201922
rect 5418 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 6038 184350
rect 5418 184226 6038 184294
rect 5418 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 6038 184226
rect 5418 184102 6038 184170
rect 5418 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 6038 184102
rect 5418 183978 6038 184046
rect 5418 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 6038 183978
rect 5418 166350 6038 183922
rect 5418 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 6038 166350
rect 5418 166226 6038 166294
rect 5418 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 6038 166226
rect 5418 166102 6038 166170
rect 5418 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 6038 166102
rect 5418 165978 6038 166046
rect 5418 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 6038 165978
rect 5418 148350 6038 165922
rect 5418 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 6038 148350
rect 5418 148226 6038 148294
rect 5418 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 6038 148226
rect 5418 148102 6038 148170
rect 5418 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 6038 148102
rect 5418 147978 6038 148046
rect 5418 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 6038 147978
rect 5418 130350 6038 147922
rect 5418 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 6038 130350
rect 5418 130226 6038 130294
rect 5418 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 6038 130226
rect 5418 130102 6038 130170
rect 5418 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 6038 130102
rect 5418 129978 6038 130046
rect 5418 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 6038 129978
rect 5418 112350 6038 129922
rect 5418 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 6038 112350
rect 5418 112226 6038 112294
rect 5418 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 6038 112226
rect 5418 112102 6038 112170
rect 5418 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 6038 112102
rect 5418 111978 6038 112046
rect 5418 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 6038 111978
rect 5418 94350 6038 111922
rect 7532 266338 7588 266348
rect 7532 107492 7588 266282
rect 7644 264718 7700 264728
rect 7644 135828 7700 264662
rect 7644 135762 7700 135772
rect 9138 262350 9758 279922
rect 17612 277060 17668 277070
rect 9138 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 9758 262350
rect 9138 262226 9758 262294
rect 9138 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 9758 262226
rect 9138 262102 9758 262170
rect 9138 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 9758 262102
rect 9138 261978 9758 262046
rect 9138 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 9758 261978
rect 9138 244350 9758 261922
rect 9138 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 9758 244350
rect 9138 244226 9758 244294
rect 9138 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 9758 244226
rect 9138 244102 9758 244170
rect 9138 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 9758 244102
rect 9138 243978 9758 244046
rect 9138 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 9758 243978
rect 9138 226350 9758 243922
rect 9138 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 9758 226350
rect 9138 226226 9758 226294
rect 9138 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 9758 226226
rect 9138 226102 9758 226170
rect 9138 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 9758 226102
rect 9138 225978 9758 226046
rect 9138 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 9758 225978
rect 9138 208350 9758 225922
rect 9138 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 9758 208350
rect 9138 208226 9758 208294
rect 9138 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 9758 208226
rect 9138 208102 9758 208170
rect 9138 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 9758 208102
rect 9138 207978 9758 208046
rect 9138 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 9758 207978
rect 9138 190350 9758 207922
rect 10892 268138 10948 268148
rect 10892 192276 10948 268082
rect 11004 264538 11060 264548
rect 11004 234612 11060 264482
rect 13736 256350 14212 256384
rect 13736 256294 13760 256350
rect 13816 256294 13884 256350
rect 13940 256294 14008 256350
rect 14064 256294 14132 256350
rect 14188 256294 14212 256350
rect 13736 256226 14212 256294
rect 13736 256170 13760 256226
rect 13816 256170 13884 256226
rect 13940 256170 14008 256226
rect 14064 256170 14132 256226
rect 14188 256170 14212 256226
rect 13736 256102 14212 256170
rect 13736 256046 13760 256102
rect 13816 256046 13884 256102
rect 13940 256046 14008 256102
rect 14064 256046 14132 256102
rect 14188 256046 14212 256102
rect 13736 255978 14212 256046
rect 13736 255922 13760 255978
rect 13816 255922 13884 255978
rect 13940 255922 14008 255978
rect 14064 255922 14132 255978
rect 14188 255922 14212 255978
rect 13736 255888 14212 255922
rect 12936 244350 13412 244384
rect 12936 244294 12960 244350
rect 13016 244294 13084 244350
rect 13140 244294 13208 244350
rect 13264 244294 13332 244350
rect 13388 244294 13412 244350
rect 12936 244226 13412 244294
rect 12936 244170 12960 244226
rect 13016 244170 13084 244226
rect 13140 244170 13208 244226
rect 13264 244170 13332 244226
rect 13388 244170 13412 244226
rect 12936 244102 13412 244170
rect 12936 244046 12960 244102
rect 13016 244046 13084 244102
rect 13140 244046 13208 244102
rect 13264 244046 13332 244102
rect 13388 244046 13412 244102
rect 12936 243978 13412 244046
rect 12936 243922 12960 243978
rect 13016 243922 13084 243978
rect 13140 243922 13208 243978
rect 13264 243922 13332 243978
rect 13388 243922 13412 243978
rect 12936 243888 13412 243922
rect 13736 238350 14212 238384
rect 13736 238294 13760 238350
rect 13816 238294 13884 238350
rect 13940 238294 14008 238350
rect 14064 238294 14132 238350
rect 14188 238294 14212 238350
rect 13736 238226 14212 238294
rect 13736 238170 13760 238226
rect 13816 238170 13884 238226
rect 13940 238170 14008 238226
rect 14064 238170 14132 238226
rect 14188 238170 14212 238226
rect 13736 238102 14212 238170
rect 13736 238046 13760 238102
rect 13816 238046 13884 238102
rect 13940 238046 14008 238102
rect 14064 238046 14132 238102
rect 14188 238046 14212 238102
rect 13736 237978 14212 238046
rect 13736 237922 13760 237978
rect 13816 237922 13884 237978
rect 13940 237922 14008 237978
rect 14064 237922 14132 237978
rect 14188 237922 14212 237978
rect 13736 237888 14212 237922
rect 11004 234546 11060 234556
rect 12936 226350 13412 226384
rect 12936 226294 12960 226350
rect 13016 226294 13084 226350
rect 13140 226294 13208 226350
rect 13264 226294 13332 226350
rect 13388 226294 13412 226350
rect 12936 226226 13412 226294
rect 12936 226170 12960 226226
rect 13016 226170 13084 226226
rect 13140 226170 13208 226226
rect 13264 226170 13332 226226
rect 13388 226170 13412 226226
rect 12936 226102 13412 226170
rect 12936 226046 12960 226102
rect 13016 226046 13084 226102
rect 13140 226046 13208 226102
rect 13264 226046 13332 226102
rect 13388 226046 13412 226102
rect 12936 225978 13412 226046
rect 12936 225922 12960 225978
rect 13016 225922 13084 225978
rect 13140 225922 13208 225978
rect 13264 225922 13332 225978
rect 13388 225922 13412 225978
rect 12936 225888 13412 225922
rect 13736 220350 14212 220384
rect 13736 220294 13760 220350
rect 13816 220294 13884 220350
rect 13940 220294 14008 220350
rect 14064 220294 14132 220350
rect 14188 220294 14212 220350
rect 13736 220226 14212 220294
rect 13736 220170 13760 220226
rect 13816 220170 13884 220226
rect 13940 220170 14008 220226
rect 14064 220170 14132 220226
rect 14188 220170 14212 220226
rect 13736 220102 14212 220170
rect 13736 220046 13760 220102
rect 13816 220046 13884 220102
rect 13940 220046 14008 220102
rect 14064 220046 14132 220102
rect 14188 220046 14212 220102
rect 13736 219978 14212 220046
rect 13736 219922 13760 219978
rect 13816 219922 13884 219978
rect 13940 219922 14008 219978
rect 14064 219922 14132 219978
rect 14188 219922 14212 219978
rect 13736 219888 14212 219922
rect 12936 208350 13412 208384
rect 12936 208294 12960 208350
rect 13016 208294 13084 208350
rect 13140 208294 13208 208350
rect 13264 208294 13332 208350
rect 13388 208294 13412 208350
rect 12936 208226 13412 208294
rect 12936 208170 12960 208226
rect 13016 208170 13084 208226
rect 13140 208170 13208 208226
rect 13264 208170 13332 208226
rect 13388 208170 13412 208226
rect 12936 208102 13412 208170
rect 12936 208046 12960 208102
rect 13016 208046 13084 208102
rect 13140 208046 13208 208102
rect 13264 208046 13332 208102
rect 13388 208046 13412 208102
rect 12936 207978 13412 208046
rect 12936 207922 12960 207978
rect 13016 207922 13084 207978
rect 13140 207922 13208 207978
rect 13264 207922 13332 207978
rect 13388 207922 13412 207978
rect 12936 207888 13412 207922
rect 13736 202350 14212 202384
rect 13736 202294 13760 202350
rect 13816 202294 13884 202350
rect 13940 202294 14008 202350
rect 14064 202294 14132 202350
rect 14188 202294 14212 202350
rect 13736 202226 14212 202294
rect 13736 202170 13760 202226
rect 13816 202170 13884 202226
rect 13940 202170 14008 202226
rect 14064 202170 14132 202226
rect 14188 202170 14212 202226
rect 13736 202102 14212 202170
rect 13736 202046 13760 202102
rect 13816 202046 13884 202102
rect 13940 202046 14008 202102
rect 14064 202046 14132 202102
rect 14188 202046 14212 202102
rect 13736 201978 14212 202046
rect 13736 201922 13760 201978
rect 13816 201922 13884 201978
rect 13940 201922 14008 201978
rect 14064 201922 14132 201978
rect 14188 201922 14212 201978
rect 13736 201888 14212 201922
rect 10892 192210 10948 192220
rect 9138 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 9758 190350
rect 9138 190226 9758 190294
rect 9138 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 9758 190226
rect 9138 190102 9758 190170
rect 9138 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 9758 190102
rect 9138 189978 9758 190046
rect 9138 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 9758 189978
rect 9138 172350 9758 189922
rect 12936 190350 13412 190384
rect 12936 190294 12960 190350
rect 13016 190294 13084 190350
rect 13140 190294 13208 190350
rect 13264 190294 13332 190350
rect 13388 190294 13412 190350
rect 12936 190226 13412 190294
rect 12936 190170 12960 190226
rect 13016 190170 13084 190226
rect 13140 190170 13208 190226
rect 13264 190170 13332 190226
rect 13388 190170 13412 190226
rect 12936 190102 13412 190170
rect 12936 190046 12960 190102
rect 13016 190046 13084 190102
rect 13140 190046 13208 190102
rect 13264 190046 13332 190102
rect 13388 190046 13412 190102
rect 12936 189978 13412 190046
rect 12936 189922 12960 189978
rect 13016 189922 13084 189978
rect 13140 189922 13208 189978
rect 13264 189922 13332 189978
rect 13388 189922 13412 189978
rect 12936 189888 13412 189922
rect 13736 184350 14212 184384
rect 13736 184294 13760 184350
rect 13816 184294 13884 184350
rect 13940 184294 14008 184350
rect 14064 184294 14132 184350
rect 14188 184294 14212 184350
rect 13736 184226 14212 184294
rect 13736 184170 13760 184226
rect 13816 184170 13884 184226
rect 13940 184170 14008 184226
rect 14064 184170 14132 184226
rect 14188 184170 14212 184226
rect 13736 184102 14212 184170
rect 13736 184046 13760 184102
rect 13816 184046 13884 184102
rect 13940 184046 14008 184102
rect 14064 184046 14132 184102
rect 14188 184046 14212 184102
rect 13736 183978 14212 184046
rect 13736 183922 13760 183978
rect 13816 183922 13884 183978
rect 13940 183922 14008 183978
rect 14064 183922 14132 183978
rect 14188 183922 14212 183978
rect 13736 183888 14212 183922
rect 9138 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 9758 172350
rect 9138 172226 9758 172294
rect 9138 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 9758 172226
rect 9138 172102 9758 172170
rect 9138 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 9758 172102
rect 9138 171978 9758 172046
rect 9138 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 9758 171978
rect 9138 154350 9758 171922
rect 12936 172350 13412 172384
rect 12936 172294 12960 172350
rect 13016 172294 13084 172350
rect 13140 172294 13208 172350
rect 13264 172294 13332 172350
rect 13388 172294 13412 172350
rect 12936 172226 13412 172294
rect 12936 172170 12960 172226
rect 13016 172170 13084 172226
rect 13140 172170 13208 172226
rect 13264 172170 13332 172226
rect 13388 172170 13412 172226
rect 12936 172102 13412 172170
rect 12936 172046 12960 172102
rect 13016 172046 13084 172102
rect 13140 172046 13208 172102
rect 13264 172046 13332 172102
rect 13388 172046 13412 172102
rect 12936 171978 13412 172046
rect 12936 171922 12960 171978
rect 13016 171922 13084 171978
rect 13140 171922 13208 171978
rect 13264 171922 13332 171978
rect 13388 171922 13412 171978
rect 12936 171888 13412 171922
rect 17612 161252 17668 277004
rect 26012 275604 26068 275614
rect 21756 269780 21812 269790
rect 21756 185698 21812 269724
rect 21756 165732 21812 185642
rect 21756 165666 21812 165676
rect 20860 162932 20916 162942
rect 20860 162838 20916 162876
rect 20860 162772 20916 162782
rect 17612 159684 17668 161196
rect 17612 159618 17668 159628
rect 26012 159572 26068 275548
rect 36138 274350 36758 281266
rect 39858 280350 40478 280964
rect 40684 280644 40740 281708
rect 40684 280578 40740 280588
rect 45388 280868 45444 280878
rect 45388 280532 45444 280812
rect 45388 280466 45444 280476
rect 39858 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 40478 280350
rect 39858 280226 40478 280294
rect 49532 280308 49588 496076
rect 49532 280242 49588 280252
rect 51212 333508 51268 333518
rect 39858 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 40478 280226
rect 39858 280102 40478 280170
rect 39858 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 40478 280102
rect 39858 279978 40478 280046
rect 39858 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 40478 279978
rect 36138 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 36758 274350
rect 36138 274226 36758 274294
rect 36138 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 36758 274226
rect 36138 274102 36758 274170
rect 36138 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 36758 274102
rect 36138 273978 36758 274046
rect 36138 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 36758 273978
rect 28476 271348 28532 271358
rect 26796 266420 26852 266430
rect 26796 187318 26852 266364
rect 26796 165732 26852 187262
rect 26796 165666 26852 165676
rect 28476 191458 28532 271292
rect 28476 165732 28532 191402
rect 28476 165666 28532 165676
rect 36138 256350 36758 273922
rect 36138 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 36758 256350
rect 36138 256226 36758 256294
rect 36138 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 36758 256226
rect 36138 256102 36758 256170
rect 36138 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 36758 256102
rect 36138 255978 36758 256046
rect 36138 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 36758 255978
rect 36138 238350 36758 255922
rect 36138 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 36758 238350
rect 36138 238226 36758 238294
rect 36138 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 36758 238226
rect 36138 238102 36758 238170
rect 36138 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 36758 238102
rect 36138 237978 36758 238046
rect 36138 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 36758 237978
rect 36138 220350 36758 237922
rect 36138 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 36758 220350
rect 36138 220226 36758 220294
rect 36138 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 36758 220226
rect 36138 220102 36758 220170
rect 36138 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 36758 220102
rect 36138 219978 36758 220046
rect 36138 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 36758 219978
rect 36138 202350 36758 219922
rect 36138 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 36758 202350
rect 36138 202226 36758 202294
rect 36138 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 36758 202226
rect 36138 202102 36758 202170
rect 36138 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 36758 202102
rect 36138 201978 36758 202046
rect 36138 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 36758 201978
rect 36138 184350 36758 201922
rect 36138 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 36758 184350
rect 36138 184226 36758 184294
rect 36138 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 36758 184226
rect 36138 184102 36758 184170
rect 36138 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 36758 184102
rect 36138 183978 36758 184046
rect 36138 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 36758 183978
rect 36138 166350 36758 183922
rect 36138 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 36758 166350
rect 36138 166226 36758 166294
rect 36138 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 36758 166226
rect 36138 166102 36758 166170
rect 36138 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 36758 166102
rect 36138 165978 36758 166046
rect 36138 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 36758 165978
rect 27132 162932 27188 162942
rect 27132 162658 27188 162876
rect 27132 162592 27188 162602
rect 26012 158004 26068 159516
rect 26012 157938 26068 157948
rect 9138 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 9758 154350
rect 9138 154226 9758 154294
rect 9138 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 9758 154226
rect 9138 154102 9758 154170
rect 9138 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 9758 154102
rect 9138 153978 9758 154046
rect 9138 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 9758 153978
rect 9138 136350 9758 153922
rect 36138 148350 36758 165922
rect 36876 275604 36932 275614
rect 36876 156212 36932 275548
rect 39676 273140 39732 273150
rect 39676 193078 39732 273084
rect 39676 165732 39732 193022
rect 39676 165666 39732 165676
rect 39858 262350 40478 279922
rect 45276 277172 45332 277182
rect 45276 277072 45332 277082
rect 48748 277172 48804 277182
rect 48636 276958 48692 276968
rect 48636 276164 48692 276902
rect 48748 276598 48804 277116
rect 48748 276532 48804 276542
rect 48636 276098 48692 276108
rect 39858 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 40478 262350
rect 39858 262226 40478 262294
rect 39858 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 40478 262226
rect 39858 262102 40478 262170
rect 39858 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 40478 262102
rect 39858 261978 40478 262046
rect 39858 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 40478 261978
rect 39858 244350 40478 261922
rect 39858 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 40478 244350
rect 39858 244226 40478 244294
rect 39858 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 40478 244226
rect 39858 244102 40478 244170
rect 39858 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 40478 244102
rect 39858 243978 40478 244046
rect 39858 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 40478 243978
rect 39858 226350 40478 243922
rect 39858 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 40478 226350
rect 39858 226226 40478 226294
rect 39858 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 40478 226226
rect 39858 226102 40478 226170
rect 39858 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 40478 226102
rect 39858 225978 40478 226046
rect 39858 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 40478 225978
rect 39858 208350 40478 225922
rect 39858 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 40478 208350
rect 39858 208226 40478 208294
rect 39858 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 40478 208226
rect 39858 208102 40478 208170
rect 39858 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 40478 208102
rect 39858 207978 40478 208046
rect 39858 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 40478 207978
rect 39858 190350 40478 207922
rect 39858 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 40478 190350
rect 39858 190226 40478 190294
rect 39858 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 40478 190226
rect 39858 190102 40478 190170
rect 39858 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 40478 190102
rect 39858 189978 40478 190046
rect 39858 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 40478 189978
rect 39858 172350 40478 189922
rect 39858 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 40478 172350
rect 39858 172226 40478 172294
rect 39858 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 40478 172226
rect 39858 172102 40478 172170
rect 39858 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 40478 172102
rect 39858 171978 40478 172046
rect 39858 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 40478 171978
rect 36876 155540 36932 156156
rect 36876 155474 36932 155484
rect 36138 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 36758 148350
rect 36138 148226 36758 148294
rect 36138 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 36758 148226
rect 36138 148102 36758 148170
rect 36138 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 36758 148102
rect 36138 147978 36758 148046
rect 36138 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 36758 147978
rect 9138 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 9758 136350
rect 9138 136226 9758 136294
rect 9138 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 9758 136226
rect 9138 136102 9758 136170
rect 9138 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 9758 136102
rect 9138 135978 9758 136046
rect 9138 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 9758 135978
rect 7532 107426 7588 107436
rect 9138 118350 9758 135922
rect 11906 136350 12382 136384
rect 11906 136294 11930 136350
rect 11986 136294 12054 136350
rect 12110 136294 12178 136350
rect 12234 136294 12302 136350
rect 12358 136294 12382 136350
rect 11906 136226 12382 136294
rect 11906 136170 11930 136226
rect 11986 136170 12054 136226
rect 12110 136170 12178 136226
rect 12234 136170 12302 136226
rect 12358 136170 12382 136226
rect 11906 136102 12382 136170
rect 11906 136046 11930 136102
rect 11986 136046 12054 136102
rect 12110 136046 12178 136102
rect 12234 136046 12302 136102
rect 12358 136046 12382 136102
rect 11906 135978 12382 136046
rect 11906 135922 11930 135978
rect 11986 135922 12054 135978
rect 12110 135922 12178 135978
rect 12234 135922 12302 135978
rect 12358 135922 12382 135978
rect 11906 135888 12382 135922
rect 11106 130350 11582 130384
rect 11106 130294 11130 130350
rect 11186 130294 11254 130350
rect 11310 130294 11378 130350
rect 11434 130294 11502 130350
rect 11558 130294 11582 130350
rect 11106 130226 11582 130294
rect 11106 130170 11130 130226
rect 11186 130170 11254 130226
rect 11310 130170 11378 130226
rect 11434 130170 11502 130226
rect 11558 130170 11582 130226
rect 11106 130102 11582 130170
rect 11106 130046 11130 130102
rect 11186 130046 11254 130102
rect 11310 130046 11378 130102
rect 11434 130046 11502 130102
rect 11558 130046 11582 130102
rect 11106 129978 11582 130046
rect 11106 129922 11130 129978
rect 11186 129922 11254 129978
rect 11310 129922 11378 129978
rect 11434 129922 11502 129978
rect 11558 129922 11582 129978
rect 11106 129888 11582 129922
rect 36138 130350 36758 147922
rect 36138 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 36758 130350
rect 36138 130226 36758 130294
rect 36138 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 36758 130226
rect 36138 130102 36758 130170
rect 36138 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 36758 130102
rect 36138 129978 36758 130046
rect 36138 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 36758 129978
rect 9138 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 9758 118350
rect 9138 118226 9758 118294
rect 9138 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 9758 118226
rect 9138 118102 9758 118170
rect 9138 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 9758 118102
rect 9138 117978 9758 118046
rect 9138 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 9758 117978
rect 5418 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 6038 94350
rect 5418 94226 6038 94294
rect 5418 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 6038 94226
rect 5418 94102 6038 94170
rect 5418 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 6038 94102
rect 5418 93978 6038 94046
rect 5418 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 6038 93978
rect 4172 79314 4228 79324
rect 140 51202 196 51212
rect 5418 76350 6038 93922
rect 5418 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 6038 76350
rect 5418 76226 6038 76294
rect 5418 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 6038 76226
rect 5418 76102 6038 76170
rect 5418 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 6038 76102
rect 5418 75978 6038 76046
rect 5418 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 6038 75978
rect 5418 58350 6038 75922
rect 5418 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 6038 58350
rect 5418 58226 6038 58294
rect 5418 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 6038 58226
rect 5418 58102 6038 58170
rect 5418 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 6038 58102
rect 5418 57978 6038 58046
rect 5418 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 6038 57978
rect 28 22978 84 22988
rect 5418 40350 6038 57922
rect 5418 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 6038 40350
rect 5418 40226 6038 40294
rect 5418 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 6038 40226
rect 5418 40102 6038 40170
rect 5418 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 6038 40102
rect 5418 39978 6038 40046
rect 5418 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 6038 39978
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 5418 22350 6038 39922
rect 5418 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 6038 22350
rect 5418 22226 6038 22294
rect 5418 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 6038 22226
rect 5418 22102 6038 22170
rect 5418 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 6038 22102
rect 5418 21978 6038 22046
rect 5418 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 6038 21978
rect 5418 4350 6038 21922
rect 5418 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 6038 4350
rect 5418 4226 6038 4294
rect 5418 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 6038 4226
rect 5418 4102 6038 4170
rect 5418 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 6038 4102
rect 5418 3978 6038 4046
rect 5418 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 6038 3978
rect 5418 -160 6038 3922
rect 5418 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 6038 -160
rect 5418 -284 6038 -216
rect 5418 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 6038 -284
rect 5418 -408 6038 -340
rect 5418 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 6038 -408
rect 5418 -532 6038 -464
rect 5418 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 6038 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 5418 -1644 6038 -588
rect 9138 100350 9758 117922
rect 11906 118350 12382 118384
rect 11906 118294 11930 118350
rect 11986 118294 12054 118350
rect 12110 118294 12178 118350
rect 12234 118294 12302 118350
rect 12358 118294 12382 118350
rect 11906 118226 12382 118294
rect 11906 118170 11930 118226
rect 11986 118170 12054 118226
rect 12110 118170 12178 118226
rect 12234 118170 12302 118226
rect 12358 118170 12382 118226
rect 11906 118102 12382 118170
rect 11906 118046 11930 118102
rect 11986 118046 12054 118102
rect 12110 118046 12178 118102
rect 12234 118046 12302 118102
rect 12358 118046 12382 118102
rect 11906 117978 12382 118046
rect 11906 117922 11930 117978
rect 11986 117922 12054 117978
rect 12110 117922 12178 117978
rect 12234 117922 12302 117978
rect 12358 117922 12382 117978
rect 11906 117888 12382 117922
rect 11106 112350 11582 112384
rect 11106 112294 11130 112350
rect 11186 112294 11254 112350
rect 11310 112294 11378 112350
rect 11434 112294 11502 112350
rect 11558 112294 11582 112350
rect 11106 112226 11582 112294
rect 11106 112170 11130 112226
rect 11186 112170 11254 112226
rect 11310 112170 11378 112226
rect 11434 112170 11502 112226
rect 11558 112170 11582 112226
rect 11106 112102 11582 112170
rect 11106 112046 11130 112102
rect 11186 112046 11254 112102
rect 11310 112046 11378 112102
rect 11434 112046 11502 112102
rect 11558 112046 11582 112102
rect 11106 111978 11582 112046
rect 11106 111922 11130 111978
rect 11186 111922 11254 111978
rect 11310 111922 11378 111978
rect 11434 111922 11502 111978
rect 11558 111922 11582 111978
rect 11106 111888 11582 111922
rect 36138 112350 36758 129922
rect 36138 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 36758 112350
rect 36138 112226 36758 112294
rect 36138 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 36758 112226
rect 36138 112102 36758 112170
rect 36138 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 36758 112102
rect 36138 111978 36758 112046
rect 36138 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 36758 111978
rect 9138 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 9758 100350
rect 9138 100226 9758 100294
rect 9138 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 9758 100226
rect 9138 100102 9758 100170
rect 9138 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 9758 100102
rect 9138 99978 9758 100046
rect 9138 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 9758 99978
rect 9138 82350 9758 99922
rect 11906 100350 12382 100384
rect 11906 100294 11930 100350
rect 11986 100294 12054 100350
rect 12110 100294 12178 100350
rect 12234 100294 12302 100350
rect 12358 100294 12382 100350
rect 11906 100226 12382 100294
rect 11906 100170 11930 100226
rect 11986 100170 12054 100226
rect 12110 100170 12178 100226
rect 12234 100170 12302 100226
rect 12358 100170 12382 100226
rect 11906 100102 12382 100170
rect 11906 100046 11930 100102
rect 11986 100046 12054 100102
rect 12110 100046 12178 100102
rect 12234 100046 12302 100102
rect 12358 100046 12382 100102
rect 11906 99978 12382 100046
rect 11906 99922 11930 99978
rect 11986 99922 12054 99978
rect 12110 99922 12178 99978
rect 12234 99922 12302 99978
rect 12358 99922 12382 99978
rect 11906 99888 12382 99922
rect 11106 94350 11582 94384
rect 11106 94294 11130 94350
rect 11186 94294 11254 94350
rect 11310 94294 11378 94350
rect 11434 94294 11502 94350
rect 11558 94294 11582 94350
rect 11106 94226 11582 94294
rect 11106 94170 11130 94226
rect 11186 94170 11254 94226
rect 11310 94170 11378 94226
rect 11434 94170 11502 94226
rect 11558 94170 11582 94226
rect 11106 94102 11582 94170
rect 11106 94046 11130 94102
rect 11186 94046 11254 94102
rect 11310 94046 11378 94102
rect 11434 94046 11502 94102
rect 11558 94046 11582 94102
rect 11106 93978 11582 94046
rect 11106 93922 11130 93978
rect 11186 93922 11254 93978
rect 11310 93922 11378 93978
rect 11434 93922 11502 93978
rect 11558 93922 11582 93978
rect 11106 93888 11582 93922
rect 36138 94350 36758 111922
rect 36138 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 36758 94350
rect 36138 94226 36758 94294
rect 36138 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 36758 94226
rect 36138 94102 36758 94170
rect 36138 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 36758 94102
rect 36138 93978 36758 94046
rect 36138 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 36758 93978
rect 9138 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 9758 82350
rect 9138 82226 9758 82294
rect 9138 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 9758 82226
rect 9138 82102 9758 82170
rect 9138 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 9758 82102
rect 9138 81978 9758 82046
rect 9138 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 9758 81978
rect 9138 64350 9758 81922
rect 11906 82350 12382 82384
rect 11906 82294 11930 82350
rect 11986 82294 12054 82350
rect 12110 82294 12178 82350
rect 12234 82294 12302 82350
rect 12358 82294 12382 82350
rect 11906 82226 12382 82294
rect 11906 82170 11930 82226
rect 11986 82170 12054 82226
rect 12110 82170 12178 82226
rect 12234 82170 12302 82226
rect 12358 82170 12382 82226
rect 11906 82102 12382 82170
rect 11906 82046 11930 82102
rect 11986 82046 12054 82102
rect 12110 82046 12178 82102
rect 12234 82046 12302 82102
rect 12358 82046 12382 82102
rect 11906 81978 12382 82046
rect 11906 81922 11930 81978
rect 11986 81922 12054 81978
rect 12110 81922 12178 81978
rect 12234 81922 12302 81978
rect 12358 81922 12382 81978
rect 11906 81888 12382 81922
rect 11106 76350 11582 76384
rect 11106 76294 11130 76350
rect 11186 76294 11254 76350
rect 11310 76294 11378 76350
rect 11434 76294 11502 76350
rect 11558 76294 11582 76350
rect 11106 76226 11582 76294
rect 11106 76170 11130 76226
rect 11186 76170 11254 76226
rect 11310 76170 11378 76226
rect 11434 76170 11502 76226
rect 11558 76170 11582 76226
rect 11106 76102 11582 76170
rect 11106 76046 11130 76102
rect 11186 76046 11254 76102
rect 11310 76046 11378 76102
rect 11434 76046 11502 76102
rect 11558 76046 11582 76102
rect 11106 75978 11582 76046
rect 11106 75922 11130 75978
rect 11186 75922 11254 75978
rect 11310 75922 11378 75978
rect 11434 75922 11502 75978
rect 11558 75922 11582 75978
rect 11106 75888 11582 75922
rect 36138 76350 36758 93922
rect 36138 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 36758 76350
rect 36138 76226 36758 76294
rect 36138 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 36758 76226
rect 36138 76102 36758 76170
rect 36138 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 36758 76102
rect 36138 75978 36758 76046
rect 36138 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 36758 75978
rect 9138 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 9758 64350
rect 9138 64226 9758 64294
rect 9138 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 9758 64226
rect 9138 64102 9758 64170
rect 9138 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 9758 64102
rect 9138 63978 9758 64046
rect 9138 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 9758 63978
rect 9138 46350 9758 63922
rect 11906 64350 12382 64384
rect 11906 64294 11930 64350
rect 11986 64294 12054 64350
rect 12110 64294 12178 64350
rect 12234 64294 12302 64350
rect 12358 64294 12382 64350
rect 11906 64226 12382 64294
rect 11906 64170 11930 64226
rect 11986 64170 12054 64226
rect 12110 64170 12178 64226
rect 12234 64170 12302 64226
rect 12358 64170 12382 64226
rect 11906 64102 12382 64170
rect 11906 64046 11930 64102
rect 11986 64046 12054 64102
rect 12110 64046 12178 64102
rect 12234 64046 12302 64102
rect 12358 64046 12382 64102
rect 11906 63978 12382 64046
rect 11906 63922 11930 63978
rect 11986 63922 12054 63978
rect 12110 63922 12178 63978
rect 12234 63922 12302 63978
rect 12358 63922 12382 63978
rect 11906 63888 12382 63922
rect 11106 58350 11582 58384
rect 11106 58294 11130 58350
rect 11186 58294 11254 58350
rect 11310 58294 11378 58350
rect 11434 58294 11502 58350
rect 11558 58294 11582 58350
rect 11106 58226 11582 58294
rect 11106 58170 11130 58226
rect 11186 58170 11254 58226
rect 11310 58170 11378 58226
rect 11434 58170 11502 58226
rect 11558 58170 11582 58226
rect 11106 58102 11582 58170
rect 11106 58046 11130 58102
rect 11186 58046 11254 58102
rect 11310 58046 11378 58102
rect 11434 58046 11502 58102
rect 11558 58046 11582 58102
rect 11106 57978 11582 58046
rect 11106 57922 11130 57978
rect 11186 57922 11254 57978
rect 11310 57922 11378 57978
rect 11434 57922 11502 57978
rect 11558 57922 11582 57978
rect 11106 57888 11582 57922
rect 36138 58350 36758 75922
rect 36138 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 36758 58350
rect 36138 58226 36758 58294
rect 36138 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 36758 58226
rect 36138 58102 36758 58170
rect 36138 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 36758 58102
rect 36138 57978 36758 58046
rect 36138 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 36758 57978
rect 9138 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 9758 46350
rect 9138 46226 9758 46294
rect 9138 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 9758 46226
rect 9138 46102 9758 46170
rect 9138 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 9758 46102
rect 9138 45978 9758 46046
rect 9138 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 9758 45978
rect 9138 28350 9758 45922
rect 9138 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 9758 28350
rect 9138 28226 9758 28294
rect 9138 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 9758 28226
rect 9138 28102 9758 28170
rect 9138 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 9758 28102
rect 9138 27978 9758 28046
rect 9138 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 9758 27978
rect 9138 10350 9758 27922
rect 9138 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 9758 10350
rect 9138 10226 9758 10294
rect 9138 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 9758 10226
rect 9138 10102 9758 10170
rect 9138 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 9758 10102
rect 9138 9978 9758 10046
rect 9138 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 9758 9978
rect 9138 -1120 9758 9922
rect 9138 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 9758 -1120
rect 9138 -1244 9758 -1176
rect 9138 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 9758 -1244
rect 9138 -1368 9758 -1300
rect 9138 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 9758 -1368
rect 9138 -1492 9758 -1424
rect 9138 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 9758 -1492
rect 9138 -1644 9758 -1548
rect 36138 40350 36758 57922
rect 36138 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 36758 40350
rect 36138 40226 36758 40294
rect 36138 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 36758 40226
rect 36138 40102 36758 40170
rect 36138 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 36758 40102
rect 36138 39978 36758 40046
rect 36138 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 36758 39978
rect 36138 22350 36758 39922
rect 36138 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 36758 22350
rect 36138 22226 36758 22294
rect 36138 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 36758 22226
rect 36138 22102 36758 22170
rect 36138 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 36758 22102
rect 36138 21978 36758 22046
rect 36138 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 36758 21978
rect 36138 4350 36758 21922
rect 36138 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 36758 4350
rect 36138 4226 36758 4294
rect 36138 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 36758 4226
rect 36138 4102 36758 4170
rect 36138 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 36758 4102
rect 36138 3978 36758 4046
rect 36138 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 36758 3978
rect 36138 -160 36758 3922
rect 36138 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 36758 -160
rect 36138 -284 36758 -216
rect 36138 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 36758 -284
rect 36138 -408 36758 -340
rect 36138 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 36758 -408
rect 36138 -532 36758 -464
rect 36138 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 36758 -532
rect 36138 -1644 36758 -588
rect 39858 154350 40478 171922
rect 39858 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 40478 154350
rect 39858 154226 40478 154294
rect 39858 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 40478 154226
rect 39858 154102 40478 154170
rect 39858 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 40478 154102
rect 39858 153978 40478 154046
rect 39858 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 40478 153978
rect 39858 136350 40478 153922
rect 41132 275604 41188 275614
rect 41132 152852 41188 275548
rect 51212 271684 51268 333452
rect 51212 271618 51268 271628
rect 51436 333396 51492 333406
rect 51436 271572 51492 333340
rect 52892 278852 52948 590492
rect 66858 580350 67478 596784
rect 66858 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 67478 580350
rect 66858 580226 67478 580294
rect 66858 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 67478 580226
rect 66858 580102 67478 580170
rect 66858 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 67478 580102
rect 66858 579978 67478 580046
rect 66858 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 67478 579978
rect 54572 575428 54628 575438
rect 54460 523348 54516 523358
rect 52892 278786 52948 278796
rect 53004 332948 53060 332958
rect 51436 271506 51492 271516
rect 53004 270004 53060 332892
rect 54460 301588 54516 523292
rect 54460 301522 54516 301532
rect 54572 278628 54628 575372
rect 66858 562350 67478 579922
rect 66858 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 67478 562350
rect 66858 562226 67478 562294
rect 66858 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 67478 562226
rect 66858 562102 67478 562170
rect 66858 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 67478 562102
rect 66858 561978 67478 562046
rect 66858 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 67478 561978
rect 66858 544350 67478 561922
rect 66858 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 67478 544350
rect 66858 544226 67478 544294
rect 66858 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 67478 544226
rect 66858 544102 67478 544170
rect 66858 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 67478 544102
rect 66858 543978 67478 544046
rect 66858 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 67478 543978
rect 59836 535780 59892 535790
rect 59612 483028 59668 483038
rect 57932 430164 57988 430174
rect 54572 278562 54628 278572
rect 54684 373156 54740 373166
rect 53004 269938 53060 269948
rect 41132 152786 41188 152796
rect 54684 148932 54740 373100
rect 57820 342468 57876 342478
rect 56588 340340 56644 340350
rect 56476 330820 56532 330830
rect 56140 321076 56196 321086
rect 56140 297556 56196 321020
rect 56476 316372 56532 330764
rect 56476 316306 56532 316316
rect 56140 297490 56196 297500
rect 56252 314244 56308 314254
rect 56252 278180 56308 314188
rect 56588 304276 56644 340284
rect 56812 338772 56868 338782
rect 56700 331828 56756 331838
rect 56700 320404 56756 331772
rect 56700 320338 56756 320348
rect 56812 313684 56868 338716
rect 56812 313618 56868 313628
rect 56924 334404 56980 334414
rect 56588 304210 56644 304220
rect 56364 302932 56420 302942
rect 56364 281998 56420 302876
rect 56924 301588 56980 334348
rect 57708 330932 57764 330942
rect 57036 325108 57092 325118
rect 57036 325018 57092 325052
rect 57036 324952 57092 324962
rect 57148 320964 57204 320974
rect 56924 301522 56980 301532
rect 57036 309204 57092 309214
rect 56476 300244 56532 300254
rect 56476 283078 56532 300188
rect 57036 298228 57092 309148
rect 57148 304724 57204 320908
rect 57708 304948 57764 330876
rect 57820 321076 57876 342412
rect 57932 325780 57988 430108
rect 58268 354788 58324 354798
rect 57932 325714 57988 325724
rect 58044 330260 58100 330270
rect 57820 321010 57876 321020
rect 57932 323764 57988 323774
rect 57708 304882 57764 304892
rect 57148 304658 57204 304668
rect 57036 298162 57092 298172
rect 57932 283438 57988 323708
rect 57932 283372 57988 283382
rect 56476 283012 56532 283022
rect 56364 281932 56420 281942
rect 56252 278114 56308 278124
rect 58044 279860 58100 330204
rect 58156 323092 58212 323102
rect 58156 284698 58212 323036
rect 58268 317492 58324 354732
rect 58604 353668 58660 353678
rect 58492 343588 58548 343598
rect 58268 317426 58324 317436
rect 58380 324660 58436 324670
rect 58156 284632 58212 284642
rect 58268 314356 58324 314366
rect 58268 282178 58324 314300
rect 58380 286498 58436 324604
rect 58492 309204 58548 343532
rect 58604 322420 58660 353612
rect 58604 322354 58660 322364
rect 58716 337316 58772 337326
rect 58716 321748 58772 337260
rect 58716 321682 58772 321692
rect 58492 309138 58548 309148
rect 58716 308980 58772 308990
rect 58716 307558 58772 308924
rect 58716 307492 58772 307502
rect 58380 286432 58436 286442
rect 58492 303604 58548 303614
rect 58492 283258 58548 303548
rect 59612 288372 59668 482972
rect 59724 368758 59780 368768
rect 59724 300916 59780 368702
rect 59724 300850 59780 300860
rect 59612 288306 59668 288316
rect 58716 287476 58772 287486
rect 58716 287398 58772 287420
rect 58716 287332 58772 287342
rect 58716 284116 58772 284126
rect 58716 283978 58772 284060
rect 58716 283912 58772 283922
rect 58492 283192 58548 283202
rect 58716 283444 58772 283454
rect 58716 282358 58772 283388
rect 58716 282292 58772 282302
rect 58268 282112 58324 282122
rect 59836 281652 59892 535724
rect 66858 526350 67478 543922
rect 66858 526294 66954 526350
rect 67010 526294 67078 526350
rect 67134 526294 67202 526350
rect 67258 526294 67326 526350
rect 67382 526294 67478 526350
rect 66858 526226 67478 526294
rect 66858 526170 66954 526226
rect 67010 526170 67078 526226
rect 67134 526170 67202 526226
rect 67258 526170 67326 526226
rect 67382 526170 67478 526226
rect 66858 526102 67478 526170
rect 66858 526046 66954 526102
rect 67010 526046 67078 526102
rect 67134 526046 67202 526102
rect 67258 526046 67326 526102
rect 67382 526046 67478 526102
rect 66858 525978 67478 526046
rect 66858 525922 66954 525978
rect 67010 525922 67078 525978
rect 67134 525922 67202 525978
rect 67258 525922 67326 525978
rect 67382 525922 67478 525978
rect 66858 508350 67478 525922
rect 66858 508294 66954 508350
rect 67010 508294 67078 508350
rect 67134 508294 67202 508350
rect 67258 508294 67326 508350
rect 67382 508294 67478 508350
rect 66858 508226 67478 508294
rect 66858 508170 66954 508226
rect 67010 508170 67078 508226
rect 67134 508170 67202 508226
rect 67258 508170 67326 508226
rect 67382 508170 67478 508226
rect 66858 508102 67478 508170
rect 66858 508046 66954 508102
rect 67010 508046 67078 508102
rect 67134 508046 67202 508102
rect 67258 508046 67326 508102
rect 67382 508046 67478 508102
rect 66858 507978 67478 508046
rect 66858 507922 66954 507978
rect 67010 507922 67078 507978
rect 67134 507922 67202 507978
rect 67258 507922 67326 507978
rect 67382 507922 67478 507978
rect 66858 490350 67478 507922
rect 66858 490294 66954 490350
rect 67010 490294 67078 490350
rect 67134 490294 67202 490350
rect 67258 490294 67326 490350
rect 67382 490294 67478 490350
rect 66858 490226 67478 490294
rect 66858 490170 66954 490226
rect 67010 490170 67078 490226
rect 67134 490170 67202 490226
rect 67258 490170 67326 490226
rect 67382 490170 67478 490226
rect 66858 490102 67478 490170
rect 66858 490046 66954 490102
rect 67010 490046 67078 490102
rect 67134 490046 67202 490102
rect 67258 490046 67326 490102
rect 67382 490046 67478 490102
rect 66858 489978 67478 490046
rect 66858 489922 66954 489978
rect 67010 489922 67078 489978
rect 67134 489922 67202 489978
rect 67258 489922 67326 489978
rect 67382 489922 67478 489978
rect 62972 482916 63028 482926
rect 60620 456484 60676 456494
rect 60508 437668 60564 437678
rect 60060 338884 60116 338894
rect 60060 319732 60116 338828
rect 60396 333060 60452 333070
rect 60172 321076 60228 321096
rect 60172 320992 60228 321002
rect 60060 319666 60116 319676
rect 59836 281586 59892 281596
rect 58044 276418 58100 279804
rect 58044 276352 58100 276362
rect 60396 276612 60452 333004
rect 60508 277956 60564 437612
rect 60620 278292 60676 456428
rect 61292 348068 61348 348078
rect 61292 330820 61348 348012
rect 62972 330932 63028 482860
rect 66858 472350 67478 489922
rect 66858 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 67478 472350
rect 66858 472226 67478 472294
rect 66858 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 67478 472226
rect 66858 472102 67478 472170
rect 66858 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 67478 472102
rect 66858 471978 67478 472046
rect 66858 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 67478 471978
rect 66858 454350 67478 471922
rect 66858 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 67478 454350
rect 66858 454226 67478 454294
rect 66858 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 67478 454226
rect 66858 454102 67478 454170
rect 66858 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 67478 454102
rect 66858 453978 67478 454046
rect 66858 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 67478 453978
rect 66858 436350 67478 453922
rect 66858 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 67478 436350
rect 66858 436226 67478 436294
rect 66858 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 67478 436226
rect 66858 436102 67478 436170
rect 66858 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 67478 436102
rect 66858 435978 67478 436046
rect 66858 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 67478 435978
rect 66858 418350 67478 435922
rect 66858 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 67478 418350
rect 66858 418226 67478 418294
rect 66858 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 67478 418226
rect 66858 418102 67478 418170
rect 66858 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 67478 418102
rect 66858 417978 67478 418046
rect 66858 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 67478 417978
rect 66858 400350 67478 417922
rect 66858 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 67478 400350
rect 66858 400226 67478 400294
rect 66858 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 67478 400226
rect 66858 400102 67478 400170
rect 66858 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 67478 400102
rect 66858 399978 67478 400046
rect 66858 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 67478 399978
rect 66858 382350 67478 399922
rect 66858 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 67478 382350
rect 66858 382226 67478 382294
rect 66858 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 67478 382226
rect 66858 382102 67478 382170
rect 66858 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 67478 382102
rect 66858 381978 67478 382046
rect 66858 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 67478 381978
rect 66858 364350 67478 381922
rect 66858 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 67478 364350
rect 66858 364226 67478 364294
rect 66858 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 67478 364226
rect 66858 364102 67478 364170
rect 66858 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 67478 364102
rect 66858 363978 67478 364046
rect 66858 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 67478 363978
rect 63756 358148 63812 358158
rect 62972 330866 63028 330876
rect 63532 333508 63588 333518
rect 61292 330754 61348 330764
rect 60620 278226 60676 278236
rect 61292 321058 61348 321068
rect 60508 277890 60564 277900
rect 60396 276058 60452 276556
rect 60396 275992 60452 276002
rect 61292 266980 61348 321002
rect 62972 307558 63028 307568
rect 62188 276948 62244 276958
rect 62188 276598 62244 276892
rect 62188 276532 62244 276542
rect 61292 266914 61348 266924
rect 61404 275604 61460 275614
rect 61404 260398 61460 275548
rect 62972 271460 63028 307502
rect 63420 277060 63476 277070
rect 63420 276612 63476 277004
rect 63532 276958 63588 333452
rect 63532 276892 63588 276902
rect 63644 332724 63700 332734
rect 63644 277138 63700 332668
rect 63756 280756 63812 358092
rect 66858 346350 67478 363922
rect 66858 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 67478 346350
rect 66858 346226 67478 346294
rect 66858 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 67478 346226
rect 66858 346102 67478 346170
rect 66858 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 67478 346102
rect 66858 345978 67478 346046
rect 66858 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 67478 345978
rect 64652 344708 64708 344718
rect 64652 334404 64708 344652
rect 64652 334338 64708 334348
rect 66858 330590 67478 345922
rect 70578 598172 71198 598268
rect 70578 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 71198 598172
rect 70578 598048 71198 598116
rect 70578 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 71198 598048
rect 70578 597924 71198 597992
rect 70578 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 71198 597924
rect 70578 597800 71198 597868
rect 70578 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 71198 597800
rect 70578 586350 71198 597744
rect 70578 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 71198 586350
rect 70578 586226 71198 586294
rect 70578 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 71198 586226
rect 70578 586102 71198 586170
rect 70578 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 71198 586102
rect 70578 585978 71198 586046
rect 70578 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 71198 585978
rect 70578 568350 71198 585922
rect 70578 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 71198 568350
rect 70578 568226 71198 568294
rect 70578 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 71198 568226
rect 70578 568102 71198 568170
rect 70578 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 71198 568102
rect 70578 567978 71198 568046
rect 70578 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 71198 567978
rect 70578 550350 71198 567922
rect 70578 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 71198 550350
rect 70578 550226 71198 550294
rect 70578 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 71198 550226
rect 70578 550102 71198 550170
rect 70578 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 71198 550102
rect 70578 549978 71198 550046
rect 70578 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 71198 549978
rect 70578 532350 71198 549922
rect 70578 532294 70674 532350
rect 70730 532294 70798 532350
rect 70854 532294 70922 532350
rect 70978 532294 71046 532350
rect 71102 532294 71198 532350
rect 70578 532226 71198 532294
rect 70578 532170 70674 532226
rect 70730 532170 70798 532226
rect 70854 532170 70922 532226
rect 70978 532170 71046 532226
rect 71102 532170 71198 532226
rect 70578 532102 71198 532170
rect 70578 532046 70674 532102
rect 70730 532046 70798 532102
rect 70854 532046 70922 532102
rect 70978 532046 71046 532102
rect 71102 532046 71198 532102
rect 70578 531978 71198 532046
rect 70578 531922 70674 531978
rect 70730 531922 70798 531978
rect 70854 531922 70922 531978
rect 70978 531922 71046 531978
rect 71102 531922 71198 531978
rect 70578 514350 71198 531922
rect 70578 514294 70674 514350
rect 70730 514294 70798 514350
rect 70854 514294 70922 514350
rect 70978 514294 71046 514350
rect 71102 514294 71198 514350
rect 70578 514226 71198 514294
rect 70578 514170 70674 514226
rect 70730 514170 70798 514226
rect 70854 514170 70922 514226
rect 70978 514170 71046 514226
rect 71102 514170 71198 514226
rect 70578 514102 71198 514170
rect 70578 514046 70674 514102
rect 70730 514046 70798 514102
rect 70854 514046 70922 514102
rect 70978 514046 71046 514102
rect 71102 514046 71198 514102
rect 70578 513978 71198 514046
rect 70578 513922 70674 513978
rect 70730 513922 70798 513978
rect 70854 513922 70922 513978
rect 70978 513922 71046 513978
rect 71102 513922 71198 513978
rect 70578 496350 71198 513922
rect 70578 496294 70674 496350
rect 70730 496294 70798 496350
rect 70854 496294 70922 496350
rect 70978 496294 71046 496350
rect 71102 496294 71198 496350
rect 70578 496226 71198 496294
rect 70578 496170 70674 496226
rect 70730 496170 70798 496226
rect 70854 496170 70922 496226
rect 70978 496170 71046 496226
rect 71102 496170 71198 496226
rect 70578 496102 71198 496170
rect 70578 496046 70674 496102
rect 70730 496046 70798 496102
rect 70854 496046 70922 496102
rect 70978 496046 71046 496102
rect 71102 496046 71198 496102
rect 70578 495978 71198 496046
rect 70578 495922 70674 495978
rect 70730 495922 70798 495978
rect 70854 495922 70922 495978
rect 70978 495922 71046 495978
rect 71102 495922 71198 495978
rect 70578 478350 71198 495922
rect 70578 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 71198 478350
rect 70578 478226 71198 478294
rect 70578 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 71198 478226
rect 70578 478102 71198 478170
rect 70578 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 71198 478102
rect 70578 477978 71198 478046
rect 70578 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 71198 477978
rect 70578 460350 71198 477922
rect 70578 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 71198 460350
rect 70578 460226 71198 460294
rect 70578 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 71198 460226
rect 70578 460102 71198 460170
rect 70578 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 71198 460102
rect 70578 459978 71198 460046
rect 70578 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 71198 459978
rect 70578 442350 71198 459922
rect 70578 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 71198 442350
rect 70578 442226 71198 442294
rect 70578 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 71198 442226
rect 70578 442102 71198 442170
rect 70578 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 71198 442102
rect 70578 441978 71198 442046
rect 70578 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 71198 441978
rect 70578 424350 71198 441922
rect 70578 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 71198 424350
rect 70578 424226 71198 424294
rect 70578 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 71198 424226
rect 70578 424102 71198 424170
rect 70578 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 71198 424102
rect 70578 423978 71198 424046
rect 70578 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 71198 423978
rect 70578 406350 71198 423922
rect 70578 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 71198 406350
rect 70578 406226 71198 406294
rect 70578 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 71198 406226
rect 70578 406102 71198 406170
rect 70578 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 71198 406102
rect 70578 405978 71198 406046
rect 70578 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 71198 405978
rect 70578 388350 71198 405922
rect 70578 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 71198 388350
rect 70578 388226 71198 388294
rect 70578 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 71198 388226
rect 70578 388102 71198 388170
rect 70578 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 71198 388102
rect 70578 387978 71198 388046
rect 70578 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 71198 387978
rect 70578 370350 71198 387922
rect 70578 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 71198 370350
rect 70578 370226 71198 370294
rect 70578 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 71198 370226
rect 70578 370102 71198 370170
rect 70578 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 71198 370102
rect 70578 369978 71198 370046
rect 70578 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 71198 369978
rect 70578 352350 71198 369922
rect 70578 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 71198 352350
rect 70578 352226 71198 352294
rect 70578 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 71198 352226
rect 70578 352102 71198 352170
rect 70578 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 71198 352102
rect 70578 351978 71198 352046
rect 70578 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 71198 351978
rect 70578 334350 71198 351922
rect 97578 597212 98198 598268
rect 97578 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 98198 597212
rect 97578 597088 98198 597156
rect 97578 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 98198 597088
rect 97578 596964 98198 597032
rect 97578 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 98198 596964
rect 97578 596840 98198 596908
rect 97578 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 98198 596840
rect 97578 580350 98198 596784
rect 97578 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 98198 580350
rect 97578 580226 98198 580294
rect 97578 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 98198 580226
rect 97578 580102 98198 580170
rect 97578 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 98198 580102
rect 97578 579978 98198 580046
rect 97578 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 98198 579978
rect 97578 562350 98198 579922
rect 97578 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 98198 562350
rect 97578 562226 98198 562294
rect 97578 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 98198 562226
rect 97578 562102 98198 562170
rect 97578 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 98198 562102
rect 97578 561978 98198 562046
rect 97578 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 98198 561978
rect 97578 544350 98198 561922
rect 97578 544294 97674 544350
rect 97730 544294 97798 544350
rect 97854 544294 97922 544350
rect 97978 544294 98046 544350
rect 98102 544294 98198 544350
rect 97578 544226 98198 544294
rect 97578 544170 97674 544226
rect 97730 544170 97798 544226
rect 97854 544170 97922 544226
rect 97978 544170 98046 544226
rect 98102 544170 98198 544226
rect 97578 544102 98198 544170
rect 97578 544046 97674 544102
rect 97730 544046 97798 544102
rect 97854 544046 97922 544102
rect 97978 544046 98046 544102
rect 98102 544046 98198 544102
rect 97578 543978 98198 544046
rect 97578 543922 97674 543978
rect 97730 543922 97798 543978
rect 97854 543922 97922 543978
rect 97978 543922 98046 543978
rect 98102 543922 98198 543978
rect 97578 526350 98198 543922
rect 97578 526294 97674 526350
rect 97730 526294 97798 526350
rect 97854 526294 97922 526350
rect 97978 526294 98046 526350
rect 98102 526294 98198 526350
rect 97578 526226 98198 526294
rect 97578 526170 97674 526226
rect 97730 526170 97798 526226
rect 97854 526170 97922 526226
rect 97978 526170 98046 526226
rect 98102 526170 98198 526226
rect 97578 526102 98198 526170
rect 97578 526046 97674 526102
rect 97730 526046 97798 526102
rect 97854 526046 97922 526102
rect 97978 526046 98046 526102
rect 98102 526046 98198 526102
rect 97578 525978 98198 526046
rect 97578 525922 97674 525978
rect 97730 525922 97798 525978
rect 97854 525922 97922 525978
rect 97978 525922 98046 525978
rect 98102 525922 98198 525978
rect 97578 508350 98198 525922
rect 97578 508294 97674 508350
rect 97730 508294 97798 508350
rect 97854 508294 97922 508350
rect 97978 508294 98046 508350
rect 98102 508294 98198 508350
rect 97578 508226 98198 508294
rect 97578 508170 97674 508226
rect 97730 508170 97798 508226
rect 97854 508170 97922 508226
rect 97978 508170 98046 508226
rect 98102 508170 98198 508226
rect 97578 508102 98198 508170
rect 97578 508046 97674 508102
rect 97730 508046 97798 508102
rect 97854 508046 97922 508102
rect 97978 508046 98046 508102
rect 98102 508046 98198 508102
rect 97578 507978 98198 508046
rect 97578 507922 97674 507978
rect 97730 507922 97798 507978
rect 97854 507922 97922 507978
rect 97978 507922 98046 507978
rect 98102 507922 98198 507978
rect 97578 490350 98198 507922
rect 97578 490294 97674 490350
rect 97730 490294 97798 490350
rect 97854 490294 97922 490350
rect 97978 490294 98046 490350
rect 98102 490294 98198 490350
rect 97578 490226 98198 490294
rect 97578 490170 97674 490226
rect 97730 490170 97798 490226
rect 97854 490170 97922 490226
rect 97978 490170 98046 490226
rect 98102 490170 98198 490226
rect 97578 490102 98198 490170
rect 97578 490046 97674 490102
rect 97730 490046 97798 490102
rect 97854 490046 97922 490102
rect 97978 490046 98046 490102
rect 98102 490046 98198 490102
rect 97578 489978 98198 490046
rect 97578 489922 97674 489978
rect 97730 489922 97798 489978
rect 97854 489922 97922 489978
rect 97978 489922 98046 489978
rect 98102 489922 98198 489978
rect 97578 472350 98198 489922
rect 97578 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 98198 472350
rect 97578 472226 98198 472294
rect 97578 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 98198 472226
rect 97578 472102 98198 472170
rect 97578 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 98198 472102
rect 97578 471978 98198 472046
rect 97578 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 98198 471978
rect 97578 454350 98198 471922
rect 97578 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 98198 454350
rect 97578 454226 98198 454294
rect 97578 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 98198 454226
rect 97578 454102 98198 454170
rect 97578 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 98198 454102
rect 97578 453978 98198 454046
rect 97578 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 98198 453978
rect 97578 436350 98198 453922
rect 97578 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 98198 436350
rect 97578 436226 98198 436294
rect 97578 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 98198 436226
rect 97578 436102 98198 436170
rect 97578 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 98198 436102
rect 97578 435978 98198 436046
rect 97578 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 98198 435978
rect 97578 418350 98198 435922
rect 97578 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 98198 418350
rect 97578 418226 98198 418294
rect 97578 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 98198 418226
rect 97578 418102 98198 418170
rect 97578 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 98198 418102
rect 97578 417978 98198 418046
rect 97578 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 98198 417978
rect 97578 400350 98198 417922
rect 97578 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 98198 400350
rect 97578 400226 98198 400294
rect 97578 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 98198 400226
rect 97578 400102 98198 400170
rect 97578 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 98198 400102
rect 97578 399978 98198 400046
rect 97578 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 98198 399978
rect 97578 382350 98198 399922
rect 97578 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 98198 382350
rect 97578 382226 98198 382294
rect 97578 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 98198 382226
rect 97578 382102 98198 382170
rect 97578 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 98198 382102
rect 97578 381978 98198 382046
rect 97578 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 98198 381978
rect 97578 364350 98198 381922
rect 97578 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 98198 364350
rect 97578 364226 98198 364294
rect 97578 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 98198 364226
rect 97578 364102 98198 364170
rect 97578 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 98198 364102
rect 97578 363978 98198 364046
rect 97578 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 98198 363978
rect 70578 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 71198 334350
rect 70578 334226 71198 334294
rect 70578 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 71198 334226
rect 70578 334102 71198 334170
rect 70578 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 71198 334102
rect 70578 333978 71198 334046
rect 70578 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 71198 333978
rect 70578 330590 71198 333922
rect 91532 351428 91588 351438
rect 91532 331828 91588 351372
rect 91532 331762 91588 331772
rect 97578 346350 98198 363922
rect 97578 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 98198 346350
rect 97578 346226 98198 346294
rect 97578 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 98198 346226
rect 97578 346102 98198 346170
rect 97578 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 98198 346102
rect 97578 345978 98198 346046
rect 97578 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 98198 345978
rect 97578 330590 98198 345922
rect 101298 598172 101918 598268
rect 101298 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 101918 598172
rect 101298 598048 101918 598116
rect 101298 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 101918 598048
rect 101298 597924 101918 597992
rect 101298 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 101918 597924
rect 101298 597800 101918 597868
rect 101298 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 101918 597800
rect 101298 586350 101918 597744
rect 128298 597212 128918 598268
rect 128298 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 128918 597212
rect 128298 597088 128918 597156
rect 128298 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 128918 597088
rect 128298 596964 128918 597032
rect 128298 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 128918 596964
rect 128298 596840 128918 596908
rect 128298 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 128918 596840
rect 111692 590996 111748 591006
rect 101298 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 101918 586350
rect 101298 586226 101918 586294
rect 101298 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 101918 586226
rect 101298 586102 101918 586170
rect 101298 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 101918 586102
rect 101298 585978 101918 586046
rect 101298 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 101918 585978
rect 101298 568350 101918 585922
rect 101298 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 101918 568350
rect 101298 568226 101918 568294
rect 101298 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 101918 568226
rect 101298 568102 101918 568170
rect 101298 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 101918 568102
rect 101298 567978 101918 568046
rect 101298 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 101918 567978
rect 101298 550350 101918 567922
rect 101298 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 101918 550350
rect 101298 550226 101918 550294
rect 101298 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 101918 550226
rect 101298 550102 101918 550170
rect 101298 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 101918 550102
rect 101298 549978 101918 550046
rect 101298 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 101918 549978
rect 101298 532350 101918 549922
rect 101298 532294 101394 532350
rect 101450 532294 101518 532350
rect 101574 532294 101642 532350
rect 101698 532294 101766 532350
rect 101822 532294 101918 532350
rect 101298 532226 101918 532294
rect 101298 532170 101394 532226
rect 101450 532170 101518 532226
rect 101574 532170 101642 532226
rect 101698 532170 101766 532226
rect 101822 532170 101918 532226
rect 101298 532102 101918 532170
rect 101298 532046 101394 532102
rect 101450 532046 101518 532102
rect 101574 532046 101642 532102
rect 101698 532046 101766 532102
rect 101822 532046 101918 532102
rect 101298 531978 101918 532046
rect 101298 531922 101394 531978
rect 101450 531922 101518 531978
rect 101574 531922 101642 531978
rect 101698 531922 101766 531978
rect 101822 531922 101918 531978
rect 101298 514350 101918 531922
rect 101298 514294 101394 514350
rect 101450 514294 101518 514350
rect 101574 514294 101642 514350
rect 101698 514294 101766 514350
rect 101822 514294 101918 514350
rect 101298 514226 101918 514294
rect 101298 514170 101394 514226
rect 101450 514170 101518 514226
rect 101574 514170 101642 514226
rect 101698 514170 101766 514226
rect 101822 514170 101918 514226
rect 101298 514102 101918 514170
rect 101298 514046 101394 514102
rect 101450 514046 101518 514102
rect 101574 514046 101642 514102
rect 101698 514046 101766 514102
rect 101822 514046 101918 514102
rect 101298 513978 101918 514046
rect 101298 513922 101394 513978
rect 101450 513922 101518 513978
rect 101574 513922 101642 513978
rect 101698 513922 101766 513978
rect 101822 513922 101918 513978
rect 101298 496350 101918 513922
rect 101298 496294 101394 496350
rect 101450 496294 101518 496350
rect 101574 496294 101642 496350
rect 101698 496294 101766 496350
rect 101822 496294 101918 496350
rect 101298 496226 101918 496294
rect 101298 496170 101394 496226
rect 101450 496170 101518 496226
rect 101574 496170 101642 496226
rect 101698 496170 101766 496226
rect 101822 496170 101918 496226
rect 101298 496102 101918 496170
rect 101298 496046 101394 496102
rect 101450 496046 101518 496102
rect 101574 496046 101642 496102
rect 101698 496046 101766 496102
rect 101822 496046 101918 496102
rect 101298 495978 101918 496046
rect 101298 495922 101394 495978
rect 101450 495922 101518 495978
rect 101574 495922 101642 495978
rect 101698 495922 101766 495978
rect 101822 495922 101918 495978
rect 101298 478350 101918 495922
rect 101298 478294 101394 478350
rect 101450 478294 101518 478350
rect 101574 478294 101642 478350
rect 101698 478294 101766 478350
rect 101822 478294 101918 478350
rect 101298 478226 101918 478294
rect 101298 478170 101394 478226
rect 101450 478170 101518 478226
rect 101574 478170 101642 478226
rect 101698 478170 101766 478226
rect 101822 478170 101918 478226
rect 101298 478102 101918 478170
rect 101298 478046 101394 478102
rect 101450 478046 101518 478102
rect 101574 478046 101642 478102
rect 101698 478046 101766 478102
rect 101822 478046 101918 478102
rect 101298 477978 101918 478046
rect 101298 477922 101394 477978
rect 101450 477922 101518 477978
rect 101574 477922 101642 477978
rect 101698 477922 101766 477978
rect 101822 477922 101918 477978
rect 101298 460350 101918 477922
rect 101298 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 101918 460350
rect 101298 460226 101918 460294
rect 101298 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 101918 460226
rect 101298 460102 101918 460170
rect 101298 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 101918 460102
rect 101298 459978 101918 460046
rect 101298 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 101918 459978
rect 101298 442350 101918 459922
rect 101298 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 101918 442350
rect 101298 442226 101918 442294
rect 101298 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 101918 442226
rect 101298 442102 101918 442170
rect 101298 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 101918 442102
rect 101298 441978 101918 442046
rect 101298 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 101918 441978
rect 101298 424350 101918 441922
rect 101298 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 101918 424350
rect 101298 424226 101918 424294
rect 101298 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 101918 424226
rect 101298 424102 101918 424170
rect 101298 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 101918 424102
rect 101298 423978 101918 424046
rect 101298 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 101918 423978
rect 101298 406350 101918 423922
rect 101298 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 101918 406350
rect 101298 406226 101918 406294
rect 101298 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 101918 406226
rect 101298 406102 101918 406170
rect 101298 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 101918 406102
rect 101298 405978 101918 406046
rect 101298 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 101918 405978
rect 101298 388350 101918 405922
rect 101298 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 101918 388350
rect 101298 388226 101918 388294
rect 101298 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 101918 388226
rect 101298 388102 101918 388170
rect 101298 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 101918 388102
rect 101298 387978 101918 388046
rect 101298 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 101918 387978
rect 101298 370350 101918 387922
rect 101298 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 101918 370350
rect 101298 370226 101918 370294
rect 101298 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 101918 370226
rect 101298 370102 101918 370170
rect 101298 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 101918 370102
rect 101298 369978 101918 370046
rect 101298 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 101918 369978
rect 101298 352350 101918 369922
rect 101298 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 101918 352350
rect 101298 352226 101918 352294
rect 101298 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 101918 352226
rect 101298 352102 101918 352170
rect 101298 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 101918 352102
rect 101298 351978 101918 352046
rect 101298 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 101918 351978
rect 101298 334350 101918 351922
rect 101298 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 101918 334350
rect 101298 334226 101918 334294
rect 101298 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 101918 334226
rect 101298 334102 101918 334170
rect 101298 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 101918 334102
rect 101298 333978 101918 334046
rect 101298 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 101918 333978
rect 101298 330590 101918 333922
rect 106652 590660 106708 590670
rect 79808 316350 80128 316384
rect 79808 316294 79878 316350
rect 79934 316294 80002 316350
rect 80058 316294 80128 316350
rect 79808 316226 80128 316294
rect 79808 316170 79878 316226
rect 79934 316170 80002 316226
rect 80058 316170 80128 316226
rect 79808 316102 80128 316170
rect 79808 316046 79878 316102
rect 79934 316046 80002 316102
rect 80058 316046 80128 316102
rect 79808 315978 80128 316046
rect 79808 315922 79878 315978
rect 79934 315922 80002 315978
rect 80058 315922 80128 315978
rect 79808 315888 80128 315922
rect 64448 310350 64768 310384
rect 64448 310294 64518 310350
rect 64574 310294 64642 310350
rect 64698 310294 64768 310350
rect 64448 310226 64768 310294
rect 64448 310170 64518 310226
rect 64574 310170 64642 310226
rect 64698 310170 64768 310226
rect 64448 310102 64768 310170
rect 64448 310046 64518 310102
rect 64574 310046 64642 310102
rect 64698 310046 64768 310102
rect 64448 309978 64768 310046
rect 64448 309922 64518 309978
rect 64574 309922 64642 309978
rect 64698 309922 64768 309978
rect 64448 309888 64768 309922
rect 95168 310350 95488 310384
rect 95168 310294 95238 310350
rect 95294 310294 95362 310350
rect 95418 310294 95488 310350
rect 95168 310226 95488 310294
rect 95168 310170 95238 310226
rect 95294 310170 95362 310226
rect 95418 310170 95488 310226
rect 95168 310102 95488 310170
rect 95168 310046 95238 310102
rect 95294 310046 95362 310102
rect 95418 310046 95488 310102
rect 95168 309978 95488 310046
rect 95168 309922 95238 309978
rect 95294 309922 95362 309978
rect 95418 309922 95488 309978
rect 95168 309888 95488 309922
rect 79808 298350 80128 298384
rect 79808 298294 79878 298350
rect 79934 298294 80002 298350
rect 80058 298294 80128 298350
rect 79808 298226 80128 298294
rect 79808 298170 79878 298226
rect 79934 298170 80002 298226
rect 80058 298170 80128 298226
rect 79808 298102 80128 298170
rect 79808 298046 79878 298102
rect 79934 298046 80002 298102
rect 80058 298046 80128 298102
rect 79808 297978 80128 298046
rect 79808 297922 79878 297978
rect 79934 297922 80002 297978
rect 80058 297922 80128 297978
rect 79808 297888 80128 297922
rect 64448 292350 64768 292384
rect 64448 292294 64518 292350
rect 64574 292294 64642 292350
rect 64698 292294 64768 292350
rect 64448 292226 64768 292294
rect 64448 292170 64518 292226
rect 64574 292170 64642 292226
rect 64698 292170 64768 292226
rect 64448 292102 64768 292170
rect 64448 292046 64518 292102
rect 64574 292046 64642 292102
rect 64698 292046 64768 292102
rect 64448 291978 64768 292046
rect 64448 291922 64518 291978
rect 64574 291922 64642 291978
rect 64698 291922 64768 291978
rect 64448 291888 64768 291922
rect 95168 292350 95488 292384
rect 95168 292294 95238 292350
rect 95294 292294 95362 292350
rect 95418 292294 95488 292350
rect 95168 292226 95488 292294
rect 95168 292170 95238 292226
rect 95294 292170 95362 292226
rect 95418 292170 95488 292226
rect 95168 292102 95488 292170
rect 95168 292046 95238 292102
rect 95294 292046 95362 292102
rect 95418 292046 95488 292102
rect 95168 291978 95488 292046
rect 95168 291922 95238 291978
rect 95294 291922 95362 291978
rect 95418 291922 95488 291978
rect 95168 291888 95488 291922
rect 68796 287398 68852 287408
rect 63756 280690 63812 280700
rect 63868 277318 63924 277328
rect 63868 277172 63924 277262
rect 63868 277106 63924 277116
rect 63420 275518 63476 276556
rect 63644 276238 63700 277082
rect 64204 276778 64260 276788
rect 64204 276658 64260 276668
rect 63644 276172 63700 276182
rect 63420 275452 63476 275462
rect 64092 275604 64148 275614
rect 62972 271394 63028 271404
rect 64092 269780 64148 275548
rect 64092 269714 64148 269724
rect 66858 274350 67478 286194
rect 68796 282996 68852 287342
rect 77532 286678 77588 286688
rect 68796 282930 68852 282940
rect 70578 280350 71198 286194
rect 75516 281764 75572 281774
rect 70578 280294 70674 280350
rect 70730 280294 70798 280350
rect 70854 280294 70922 280350
rect 70978 280294 71046 280350
rect 71102 280294 71198 280350
rect 70578 280226 71198 280294
rect 70578 280170 70674 280226
rect 70730 280170 70798 280226
rect 70854 280170 70922 280226
rect 70978 280170 71046 280226
rect 71102 280170 71198 280226
rect 70578 280102 71198 280170
rect 70578 280046 70674 280102
rect 70730 280046 70798 280102
rect 70854 280046 70922 280102
rect 70978 280046 71046 280102
rect 71102 280046 71198 280102
rect 70578 279978 71198 280046
rect 74172 280756 74228 280766
rect 74172 280084 74228 280700
rect 74172 280018 74228 280028
rect 75516 280084 75572 281708
rect 75516 280018 75572 280028
rect 77532 280084 77588 286622
rect 106652 286678 106708 590604
rect 108332 544852 108388 544862
rect 107436 345828 107492 345838
rect 107436 340340 107492 345772
rect 107436 340274 107492 340284
rect 106652 286612 106708 286622
rect 106764 326098 106820 326108
rect 87612 282884 87668 282894
rect 85596 281652 85652 281662
rect 85596 280980 85652 281596
rect 85596 280914 85652 280924
rect 87612 280756 87668 282828
rect 97356 281876 97412 281886
rect 97356 280980 97412 281820
rect 97356 280914 97412 280924
rect 87612 280690 87668 280700
rect 77532 280018 77588 280028
rect 101298 280350 101918 286194
rect 101298 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 101918 280350
rect 101298 280226 101918 280294
rect 101298 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 101918 280226
rect 101298 280102 101918 280170
rect 101298 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 101918 280102
rect 70578 279922 70674 279978
rect 70730 279922 70798 279978
rect 70854 279922 70922 279978
rect 70978 279922 71046 279978
rect 71102 279922 71198 279978
rect 70364 276778 70420 276788
rect 70364 276658 70420 276668
rect 70252 276612 70308 276622
rect 66858 274294 66954 274350
rect 67010 274294 67078 274350
rect 67134 274294 67202 274350
rect 67258 274294 67326 274350
rect 67382 274294 67478 274350
rect 66858 274226 67478 274294
rect 66858 274170 66954 274226
rect 67010 274170 67078 274226
rect 67134 274170 67202 274226
rect 67258 274170 67326 274226
rect 67382 274170 67478 274226
rect 66858 274102 67478 274170
rect 66858 274046 66954 274102
rect 67010 274046 67078 274102
rect 67134 274046 67202 274102
rect 67258 274046 67326 274102
rect 67382 274046 67478 274102
rect 66858 273978 67478 274046
rect 66858 273922 66954 273978
rect 67010 273922 67078 273978
rect 67134 273922 67202 273978
rect 67258 273922 67326 273978
rect 67382 273922 67478 273978
rect 61404 260332 61460 260342
rect 54684 148866 54740 148876
rect 66858 256350 67478 273922
rect 66858 256294 66954 256350
rect 67010 256294 67078 256350
rect 67134 256294 67202 256350
rect 67258 256294 67326 256350
rect 67382 256294 67478 256350
rect 66858 256226 67478 256294
rect 66858 256170 66954 256226
rect 67010 256170 67078 256226
rect 67134 256170 67202 256226
rect 67258 256170 67326 256226
rect 67382 256170 67478 256226
rect 66858 256102 67478 256170
rect 66858 256046 66954 256102
rect 67010 256046 67078 256102
rect 67134 256046 67202 256102
rect 67258 256046 67326 256102
rect 67382 256046 67478 256102
rect 66858 255978 67478 256046
rect 66858 255922 66954 255978
rect 67010 255922 67078 255978
rect 67134 255922 67202 255978
rect 67258 255922 67326 255978
rect 67382 255922 67478 255978
rect 66858 238350 67478 255922
rect 66858 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 67478 238350
rect 66858 238226 67478 238294
rect 66858 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 67478 238226
rect 66858 238102 67478 238170
rect 66858 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 67478 238102
rect 66858 237978 67478 238046
rect 66858 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 67478 237978
rect 66858 220350 67478 237922
rect 66858 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 67478 220350
rect 66858 220226 67478 220294
rect 66858 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 67478 220226
rect 66858 220102 67478 220170
rect 66858 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 67478 220102
rect 66858 219978 67478 220046
rect 66858 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 67478 219978
rect 66858 202350 67478 219922
rect 66858 202294 66954 202350
rect 67010 202294 67078 202350
rect 67134 202294 67202 202350
rect 67258 202294 67326 202350
rect 67382 202294 67478 202350
rect 66858 202226 67478 202294
rect 66858 202170 66954 202226
rect 67010 202170 67078 202226
rect 67134 202170 67202 202226
rect 67258 202170 67326 202226
rect 67382 202170 67478 202226
rect 66858 202102 67478 202170
rect 66858 202046 66954 202102
rect 67010 202046 67078 202102
rect 67134 202046 67202 202102
rect 67258 202046 67326 202102
rect 67382 202046 67478 202102
rect 66858 201978 67478 202046
rect 66858 201922 66954 201978
rect 67010 201922 67078 201978
rect 67134 201922 67202 201978
rect 67258 201922 67326 201978
rect 67382 201922 67478 201978
rect 66858 184350 67478 201922
rect 66858 184294 66954 184350
rect 67010 184294 67078 184350
rect 67134 184294 67202 184350
rect 67258 184294 67326 184350
rect 67382 184294 67478 184350
rect 66858 184226 67478 184294
rect 66858 184170 66954 184226
rect 67010 184170 67078 184226
rect 67134 184170 67202 184226
rect 67258 184170 67326 184226
rect 67382 184170 67478 184226
rect 66858 184102 67478 184170
rect 66858 184046 66954 184102
rect 67010 184046 67078 184102
rect 67134 184046 67202 184102
rect 67258 184046 67326 184102
rect 67382 184046 67478 184102
rect 66858 183978 67478 184046
rect 66858 183922 66954 183978
rect 67010 183922 67078 183978
rect 67134 183922 67202 183978
rect 67258 183922 67326 183978
rect 67382 183922 67478 183978
rect 66858 166350 67478 183922
rect 66858 166294 66954 166350
rect 67010 166294 67078 166350
rect 67134 166294 67202 166350
rect 67258 166294 67326 166350
rect 67382 166294 67478 166350
rect 66858 166226 67478 166294
rect 66858 166170 66954 166226
rect 67010 166170 67078 166226
rect 67134 166170 67202 166226
rect 67258 166170 67326 166226
rect 67382 166170 67478 166226
rect 66858 166102 67478 166170
rect 66858 166046 66954 166102
rect 67010 166046 67078 166102
rect 67134 166046 67202 166102
rect 67258 166046 67326 166102
rect 67382 166046 67478 166102
rect 66858 165978 67478 166046
rect 66858 165922 66954 165978
rect 67010 165922 67078 165978
rect 67134 165922 67202 165978
rect 67258 165922 67326 165978
rect 67382 165922 67478 165978
rect 39858 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 40478 136350
rect 39858 136226 40478 136294
rect 39858 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 40478 136226
rect 39858 136102 40478 136170
rect 39858 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 40478 136102
rect 39858 135978 40478 136046
rect 39858 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 40478 135978
rect 39858 118350 40478 135922
rect 39858 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 40478 118350
rect 39858 118226 40478 118294
rect 39858 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 40478 118226
rect 39858 118102 40478 118170
rect 39858 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 40478 118102
rect 39858 117978 40478 118046
rect 39858 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 40478 117978
rect 39858 100350 40478 117922
rect 39858 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 40478 100350
rect 39858 100226 40478 100294
rect 39858 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 40478 100226
rect 39858 100102 40478 100170
rect 39858 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 40478 100102
rect 39858 99978 40478 100046
rect 39858 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 40478 99978
rect 39858 82350 40478 99922
rect 39858 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 40478 82350
rect 39858 82226 40478 82294
rect 39858 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 40478 82226
rect 39858 82102 40478 82170
rect 39858 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 40478 82102
rect 39858 81978 40478 82046
rect 39858 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 40478 81978
rect 39858 64350 40478 81922
rect 39858 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 40478 64350
rect 39858 64226 40478 64294
rect 39858 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 40478 64226
rect 39858 64102 40478 64170
rect 39858 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 40478 64102
rect 39858 63978 40478 64046
rect 39858 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 40478 63978
rect 39858 46350 40478 63922
rect 39858 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 40478 46350
rect 39858 46226 40478 46294
rect 39858 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 40478 46226
rect 39858 46102 40478 46170
rect 39858 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 40478 46102
rect 39858 45978 40478 46046
rect 39858 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 40478 45978
rect 39858 28350 40478 45922
rect 39858 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 40478 28350
rect 39858 28226 40478 28294
rect 39858 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 40478 28226
rect 39858 28102 40478 28170
rect 39858 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 40478 28102
rect 39858 27978 40478 28046
rect 39858 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 40478 27978
rect 39858 10350 40478 27922
rect 39858 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 40478 10350
rect 39858 10226 40478 10294
rect 39858 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 40478 10226
rect 39858 10102 40478 10170
rect 39858 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 40478 10102
rect 39858 9978 40478 10046
rect 39858 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 40478 9978
rect 39858 -1120 40478 9922
rect 39858 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 40478 -1120
rect 39858 -1244 40478 -1176
rect 39858 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 40478 -1244
rect 39858 -1368 40478 -1300
rect 39858 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 40478 -1368
rect 39858 -1492 40478 -1424
rect 39858 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 40478 -1492
rect 39858 -1644 40478 -1548
rect 66858 148350 67478 165922
rect 69692 276238 69748 276248
rect 69692 150612 69748 276182
rect 70252 271378 70308 276556
rect 70364 276058 70420 276068
rect 70364 272916 70420 276002
rect 70364 272850 70420 272860
rect 70364 271378 70420 271388
rect 70252 271322 70364 271378
rect 70364 271312 70420 271322
rect 69692 150546 69748 150556
rect 70578 262350 71198 279922
rect 101298 279978 101918 280046
rect 101298 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 101918 279978
rect 74172 278516 74228 278526
rect 74172 278218 74228 278460
rect 74172 278152 74228 278162
rect 73052 276958 73108 276968
rect 70578 262294 70674 262350
rect 70730 262294 70798 262350
rect 70854 262294 70922 262350
rect 70978 262294 71046 262350
rect 71102 262294 71198 262350
rect 70578 262226 71198 262294
rect 70578 262170 70674 262226
rect 70730 262170 70798 262226
rect 70854 262170 70922 262226
rect 70978 262170 71046 262226
rect 71102 262170 71198 262226
rect 70578 262102 71198 262170
rect 70578 262046 70674 262102
rect 70730 262046 70798 262102
rect 70854 262046 70922 262102
rect 70978 262046 71046 262102
rect 71102 262046 71198 262102
rect 70578 261978 71198 262046
rect 70578 261922 70674 261978
rect 70730 261922 70798 261978
rect 70854 261922 70922 261978
rect 70978 261922 71046 261978
rect 71102 261922 71198 261978
rect 70578 244350 71198 261922
rect 70578 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 71198 244350
rect 70578 244226 71198 244294
rect 70578 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 71198 244226
rect 70578 244102 71198 244170
rect 70578 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 71198 244102
rect 70578 243978 71198 244046
rect 70578 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 71198 243978
rect 70578 226350 71198 243922
rect 70578 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 71198 226350
rect 70578 226226 71198 226294
rect 70578 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 71198 226226
rect 70578 226102 71198 226170
rect 70578 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 71198 226102
rect 70578 225978 71198 226046
rect 70578 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 71198 225978
rect 70578 208350 71198 225922
rect 70578 208294 70674 208350
rect 70730 208294 70798 208350
rect 70854 208294 70922 208350
rect 70978 208294 71046 208350
rect 71102 208294 71198 208350
rect 70578 208226 71198 208294
rect 70578 208170 70674 208226
rect 70730 208170 70798 208226
rect 70854 208170 70922 208226
rect 70978 208170 71046 208226
rect 71102 208170 71198 208226
rect 70578 208102 71198 208170
rect 70578 208046 70674 208102
rect 70730 208046 70798 208102
rect 70854 208046 70922 208102
rect 70978 208046 71046 208102
rect 71102 208046 71198 208102
rect 70578 207978 71198 208046
rect 70578 207922 70674 207978
rect 70730 207922 70798 207978
rect 70854 207922 70922 207978
rect 70978 207922 71046 207978
rect 71102 207922 71198 207978
rect 70578 190350 71198 207922
rect 70578 190294 70674 190350
rect 70730 190294 70798 190350
rect 70854 190294 70922 190350
rect 70978 190294 71046 190350
rect 71102 190294 71198 190350
rect 70578 190226 71198 190294
rect 70578 190170 70674 190226
rect 70730 190170 70798 190226
rect 70854 190170 70922 190226
rect 70978 190170 71046 190226
rect 71102 190170 71198 190226
rect 70578 190102 71198 190170
rect 70578 190046 70674 190102
rect 70730 190046 70798 190102
rect 70854 190046 70922 190102
rect 70978 190046 71046 190102
rect 71102 190046 71198 190102
rect 70578 189978 71198 190046
rect 70578 189922 70674 189978
rect 70730 189922 70798 189978
rect 70854 189922 70922 189978
rect 70978 189922 71046 189978
rect 71102 189922 71198 189978
rect 70578 172350 71198 189922
rect 70578 172294 70674 172350
rect 70730 172294 70798 172350
rect 70854 172294 70922 172350
rect 70978 172294 71046 172350
rect 71102 172294 71198 172350
rect 70578 172226 71198 172294
rect 70578 172170 70674 172226
rect 70730 172170 70798 172226
rect 70854 172170 70922 172226
rect 70978 172170 71046 172226
rect 71102 172170 71198 172226
rect 70578 172102 71198 172170
rect 70578 172046 70674 172102
rect 70730 172046 70798 172102
rect 70854 172046 70922 172102
rect 70978 172046 71046 172102
rect 71102 172046 71198 172102
rect 70578 171978 71198 172046
rect 70578 171922 70674 171978
rect 70730 171922 70798 171978
rect 70854 171922 70922 171978
rect 70978 171922 71046 171978
rect 71102 171922 71198 171978
rect 70578 154350 71198 171922
rect 72156 276612 72212 276622
rect 72156 275604 72212 276556
rect 72156 195778 72212 275548
rect 72156 165732 72212 195722
rect 72156 165666 72212 165676
rect 73052 157444 73108 276902
rect 84812 276948 84868 276958
rect 73052 157378 73108 157388
rect 74732 276418 74788 276428
rect 70578 154294 70674 154350
rect 70730 154294 70798 154350
rect 70854 154294 70922 154350
rect 70978 154294 71046 154350
rect 71102 154294 71198 154350
rect 70578 154226 71198 154294
rect 70578 154170 70674 154226
rect 70730 154170 70798 154226
rect 70854 154170 70922 154226
rect 70978 154170 71046 154226
rect 71102 154170 71198 154226
rect 70578 154102 71198 154170
rect 70578 154046 70674 154102
rect 70730 154046 70798 154102
rect 70854 154046 70922 154102
rect 70978 154046 71046 154102
rect 71102 154046 71198 154102
rect 70578 153978 71198 154046
rect 70578 153922 70674 153978
rect 70730 153922 70798 153978
rect 70854 153922 70922 153978
rect 70978 153922 71046 153978
rect 71102 153922 71198 153978
rect 66858 148294 66954 148350
rect 67010 148294 67078 148350
rect 67134 148294 67202 148350
rect 67258 148294 67326 148350
rect 67382 148294 67478 148350
rect 66858 148226 67478 148294
rect 66858 148170 66954 148226
rect 67010 148170 67078 148226
rect 67134 148170 67202 148226
rect 67258 148170 67326 148226
rect 67382 148170 67478 148226
rect 66858 148102 67478 148170
rect 66858 148046 66954 148102
rect 67010 148046 67078 148102
rect 67134 148046 67202 148102
rect 67258 148046 67326 148102
rect 67382 148046 67478 148102
rect 66858 147978 67478 148046
rect 66858 147922 66954 147978
rect 67010 147922 67078 147978
rect 67134 147922 67202 147978
rect 67258 147922 67326 147978
rect 67382 147922 67478 147978
rect 66858 130350 67478 147922
rect 66858 130294 66954 130350
rect 67010 130294 67078 130350
rect 67134 130294 67202 130350
rect 67258 130294 67326 130350
rect 67382 130294 67478 130350
rect 66858 130226 67478 130294
rect 66858 130170 66954 130226
rect 67010 130170 67078 130226
rect 67134 130170 67202 130226
rect 67258 130170 67326 130226
rect 67382 130170 67478 130226
rect 66858 130102 67478 130170
rect 66858 130046 66954 130102
rect 67010 130046 67078 130102
rect 67134 130046 67202 130102
rect 67258 130046 67326 130102
rect 67382 130046 67478 130102
rect 66858 129978 67478 130046
rect 66858 129922 66954 129978
rect 67010 129922 67078 129978
rect 67134 129922 67202 129978
rect 67258 129922 67326 129978
rect 67382 129922 67478 129978
rect 66858 112350 67478 129922
rect 66858 112294 66954 112350
rect 67010 112294 67078 112350
rect 67134 112294 67202 112350
rect 67258 112294 67326 112350
rect 67382 112294 67478 112350
rect 66858 112226 67478 112294
rect 66858 112170 66954 112226
rect 67010 112170 67078 112226
rect 67134 112170 67202 112226
rect 67258 112170 67326 112226
rect 67382 112170 67478 112226
rect 66858 112102 67478 112170
rect 66858 112046 66954 112102
rect 67010 112046 67078 112102
rect 67134 112046 67202 112102
rect 67258 112046 67326 112102
rect 67382 112046 67478 112102
rect 66858 111978 67478 112046
rect 66858 111922 66954 111978
rect 67010 111922 67078 111978
rect 67134 111922 67202 111978
rect 67258 111922 67326 111978
rect 67382 111922 67478 111978
rect 66858 94350 67478 111922
rect 66858 94294 66954 94350
rect 67010 94294 67078 94350
rect 67134 94294 67202 94350
rect 67258 94294 67326 94350
rect 67382 94294 67478 94350
rect 66858 94226 67478 94294
rect 66858 94170 66954 94226
rect 67010 94170 67078 94226
rect 67134 94170 67202 94226
rect 67258 94170 67326 94226
rect 67382 94170 67478 94226
rect 66858 94102 67478 94170
rect 66858 94046 66954 94102
rect 67010 94046 67078 94102
rect 67134 94046 67202 94102
rect 67258 94046 67326 94102
rect 67382 94046 67478 94102
rect 66858 93978 67478 94046
rect 66858 93922 66954 93978
rect 67010 93922 67078 93978
rect 67134 93922 67202 93978
rect 67258 93922 67326 93978
rect 67382 93922 67478 93978
rect 66858 76350 67478 93922
rect 66858 76294 66954 76350
rect 67010 76294 67078 76350
rect 67134 76294 67202 76350
rect 67258 76294 67326 76350
rect 67382 76294 67478 76350
rect 66858 76226 67478 76294
rect 66858 76170 66954 76226
rect 67010 76170 67078 76226
rect 67134 76170 67202 76226
rect 67258 76170 67326 76226
rect 67382 76170 67478 76226
rect 66858 76102 67478 76170
rect 66858 76046 66954 76102
rect 67010 76046 67078 76102
rect 67134 76046 67202 76102
rect 67258 76046 67326 76102
rect 67382 76046 67478 76102
rect 66858 75978 67478 76046
rect 66858 75922 66954 75978
rect 67010 75922 67078 75978
rect 67134 75922 67202 75978
rect 67258 75922 67326 75978
rect 67382 75922 67478 75978
rect 66858 58350 67478 75922
rect 66858 58294 66954 58350
rect 67010 58294 67078 58350
rect 67134 58294 67202 58350
rect 67258 58294 67326 58350
rect 67382 58294 67478 58350
rect 66858 58226 67478 58294
rect 66858 58170 66954 58226
rect 67010 58170 67078 58226
rect 67134 58170 67202 58226
rect 67258 58170 67326 58226
rect 67382 58170 67478 58226
rect 66858 58102 67478 58170
rect 66858 58046 66954 58102
rect 67010 58046 67078 58102
rect 67134 58046 67202 58102
rect 67258 58046 67326 58102
rect 67382 58046 67478 58102
rect 66858 57978 67478 58046
rect 66858 57922 66954 57978
rect 67010 57922 67078 57978
rect 67134 57922 67202 57978
rect 67258 57922 67326 57978
rect 67382 57922 67478 57978
rect 66858 40350 67478 57922
rect 66858 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 67478 40350
rect 66858 40226 67478 40294
rect 66858 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 67478 40226
rect 66858 40102 67478 40170
rect 66858 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 67478 40102
rect 66858 39978 67478 40046
rect 66858 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 67478 39978
rect 66858 22350 67478 39922
rect 66858 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 67478 22350
rect 66858 22226 67478 22294
rect 66858 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 67478 22226
rect 66858 22102 67478 22170
rect 66858 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 67478 22102
rect 66858 21978 67478 22046
rect 66858 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 67478 21978
rect 66858 4350 67478 21922
rect 66858 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 67478 4350
rect 66858 4226 67478 4294
rect 66858 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 67478 4226
rect 66858 4102 67478 4170
rect 66858 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 67478 4102
rect 66858 3978 67478 4046
rect 66858 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 67478 3978
rect 66858 -160 67478 3922
rect 66858 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 67478 -160
rect 66858 -284 67478 -216
rect 66858 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 67478 -284
rect 66858 -408 67478 -340
rect 66858 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 67478 -408
rect 66858 -532 67478 -464
rect 66858 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 67478 -532
rect 66858 -1644 67478 -588
rect 70578 136350 71198 153922
rect 74732 152180 74788 276362
rect 82236 276388 82292 276398
rect 82236 276164 82292 276332
rect 74732 152114 74788 152124
rect 79772 272916 79828 272926
rect 72044 149518 72100 149528
rect 72044 147924 72100 149462
rect 79772 148708 79828 272860
rect 82236 199018 82292 276108
rect 84812 274820 84868 276892
rect 82236 165732 82292 198962
rect 82236 165666 82292 165676
rect 83916 266420 83972 266430
rect 79772 148642 79828 148652
rect 81452 149338 81508 149348
rect 72044 147858 72100 147868
rect 81452 147924 81508 149282
rect 81452 147858 81508 147868
rect 83916 147924 83972 266364
rect 84812 201538 84868 274764
rect 84812 165620 84868 201482
rect 84812 165554 84868 165564
rect 94892 276052 94948 276062
rect 94892 274708 94948 275996
rect 94892 204958 94948 274652
rect 100044 271236 100100 271246
rect 99932 268100 99988 268110
rect 98418 256350 98894 256384
rect 98418 256294 98442 256350
rect 98498 256294 98566 256350
rect 98622 256294 98690 256350
rect 98746 256294 98814 256350
rect 98870 256294 98894 256350
rect 98418 256226 98894 256294
rect 98418 256170 98442 256226
rect 98498 256170 98566 256226
rect 98622 256170 98690 256226
rect 98746 256170 98814 256226
rect 98870 256170 98894 256226
rect 98418 256102 98894 256170
rect 98418 256046 98442 256102
rect 98498 256046 98566 256102
rect 98622 256046 98690 256102
rect 98746 256046 98814 256102
rect 98870 256046 98894 256102
rect 98418 255978 98894 256046
rect 98418 255922 98442 255978
rect 98498 255922 98566 255978
rect 98622 255922 98690 255978
rect 98746 255922 98814 255978
rect 98870 255922 98894 255978
rect 98418 255888 98894 255922
rect 97618 244350 98094 244384
rect 97618 244294 97642 244350
rect 97698 244294 97766 244350
rect 97822 244294 97890 244350
rect 97946 244294 98014 244350
rect 98070 244294 98094 244350
rect 97618 244226 98094 244294
rect 97618 244170 97642 244226
rect 97698 244170 97766 244226
rect 97822 244170 97890 244226
rect 97946 244170 98014 244226
rect 98070 244170 98094 244226
rect 97618 244102 98094 244170
rect 97618 244046 97642 244102
rect 97698 244046 97766 244102
rect 97822 244046 97890 244102
rect 97946 244046 98014 244102
rect 98070 244046 98094 244102
rect 97618 243978 98094 244046
rect 97618 243922 97642 243978
rect 97698 243922 97766 243978
rect 97822 243922 97890 243978
rect 97946 243922 98014 243978
rect 98070 243922 98094 243978
rect 97618 243888 98094 243922
rect 98418 238350 98894 238384
rect 98418 238294 98442 238350
rect 98498 238294 98566 238350
rect 98622 238294 98690 238350
rect 98746 238294 98814 238350
rect 98870 238294 98894 238350
rect 98418 238226 98894 238294
rect 98418 238170 98442 238226
rect 98498 238170 98566 238226
rect 98622 238170 98690 238226
rect 98746 238170 98814 238226
rect 98870 238170 98894 238226
rect 98418 238102 98894 238170
rect 98418 238046 98442 238102
rect 98498 238046 98566 238102
rect 98622 238046 98690 238102
rect 98746 238046 98814 238102
rect 98870 238046 98894 238102
rect 98418 237978 98894 238046
rect 98418 237922 98442 237978
rect 98498 237922 98566 237978
rect 98622 237922 98690 237978
rect 98746 237922 98814 237978
rect 98870 237922 98894 237978
rect 98418 237888 98894 237922
rect 97618 226350 98094 226384
rect 97618 226294 97642 226350
rect 97698 226294 97766 226350
rect 97822 226294 97890 226350
rect 97946 226294 98014 226350
rect 98070 226294 98094 226350
rect 97618 226226 98094 226294
rect 97618 226170 97642 226226
rect 97698 226170 97766 226226
rect 97822 226170 97890 226226
rect 97946 226170 98014 226226
rect 98070 226170 98094 226226
rect 97618 226102 98094 226170
rect 97618 226046 97642 226102
rect 97698 226046 97766 226102
rect 97822 226046 97890 226102
rect 97946 226046 98014 226102
rect 98070 226046 98094 226102
rect 97618 225978 98094 226046
rect 97618 225922 97642 225978
rect 97698 225922 97766 225978
rect 97822 225922 97890 225978
rect 97946 225922 98014 225978
rect 98070 225922 98094 225978
rect 97618 225888 98094 225922
rect 98418 220350 98894 220384
rect 98418 220294 98442 220350
rect 98498 220294 98566 220350
rect 98622 220294 98690 220350
rect 98746 220294 98814 220350
rect 98870 220294 98894 220350
rect 98418 220226 98894 220294
rect 98418 220170 98442 220226
rect 98498 220170 98566 220226
rect 98622 220170 98690 220226
rect 98746 220170 98814 220226
rect 98870 220170 98894 220226
rect 98418 220102 98894 220170
rect 98418 220046 98442 220102
rect 98498 220046 98566 220102
rect 98622 220046 98690 220102
rect 98746 220046 98814 220102
rect 98870 220046 98894 220102
rect 98418 219978 98894 220046
rect 98418 219922 98442 219978
rect 98498 219922 98566 219978
rect 98622 219922 98690 219978
rect 98746 219922 98814 219978
rect 98870 219922 98894 219978
rect 98418 219888 98894 219922
rect 97618 208350 98094 208384
rect 97618 208294 97642 208350
rect 97698 208294 97766 208350
rect 97822 208294 97890 208350
rect 97946 208294 98014 208350
rect 98070 208294 98094 208350
rect 97618 208226 98094 208294
rect 97618 208170 97642 208226
rect 97698 208170 97766 208226
rect 97822 208170 97890 208226
rect 97946 208170 98014 208226
rect 98070 208170 98094 208226
rect 97618 208102 98094 208170
rect 97618 208046 97642 208102
rect 97698 208046 97766 208102
rect 97822 208046 97890 208102
rect 97946 208046 98014 208102
rect 98070 208046 98094 208102
rect 97618 207978 98094 208046
rect 97618 207922 97642 207978
rect 97698 207922 97766 207978
rect 97822 207922 97890 207978
rect 97946 207922 98014 207978
rect 98070 207922 98094 207978
rect 97618 207888 98094 207922
rect 94892 164612 94948 204902
rect 98418 202350 98894 202384
rect 98418 202294 98442 202350
rect 98498 202294 98566 202350
rect 98622 202294 98690 202350
rect 98746 202294 98814 202350
rect 98870 202294 98894 202350
rect 98418 202226 98894 202294
rect 98418 202170 98442 202226
rect 98498 202170 98566 202226
rect 98622 202170 98690 202226
rect 98746 202170 98814 202226
rect 98870 202170 98894 202226
rect 98418 202102 98894 202170
rect 98418 202046 98442 202102
rect 98498 202046 98566 202102
rect 98622 202046 98690 202102
rect 98746 202046 98814 202102
rect 98870 202046 98894 202102
rect 98418 201978 98894 202046
rect 98418 201922 98442 201978
rect 98498 201922 98566 201978
rect 98622 201922 98690 201978
rect 98746 201922 98814 201978
rect 98870 201922 98894 201978
rect 98418 201888 98894 201922
rect 97618 190350 98094 190384
rect 97618 190294 97642 190350
rect 97698 190294 97766 190350
rect 97822 190294 97890 190350
rect 97946 190294 98014 190350
rect 98070 190294 98094 190350
rect 97618 190226 98094 190294
rect 97618 190170 97642 190226
rect 97698 190170 97766 190226
rect 97822 190170 97890 190226
rect 97946 190170 98014 190226
rect 98070 190170 98094 190226
rect 97618 190102 98094 190170
rect 97618 190046 97642 190102
rect 97698 190046 97766 190102
rect 97822 190046 97890 190102
rect 97946 190046 98014 190102
rect 98070 190046 98094 190102
rect 97618 189978 98094 190046
rect 97618 189922 97642 189978
rect 97698 189922 97766 189978
rect 97822 189922 97890 189978
rect 97946 189922 98014 189978
rect 98070 189922 98094 189978
rect 97618 189888 98094 189922
rect 98418 184350 98894 184384
rect 98418 184294 98442 184350
rect 98498 184294 98566 184350
rect 98622 184294 98690 184350
rect 98746 184294 98814 184350
rect 98870 184294 98894 184350
rect 98418 184226 98894 184294
rect 98418 184170 98442 184226
rect 98498 184170 98566 184226
rect 98622 184170 98690 184226
rect 98746 184170 98814 184226
rect 98870 184170 98894 184226
rect 98418 184102 98894 184170
rect 98418 184046 98442 184102
rect 98498 184046 98566 184102
rect 98622 184046 98690 184102
rect 98746 184046 98814 184102
rect 98870 184046 98894 184102
rect 98418 183978 98894 184046
rect 98418 183922 98442 183978
rect 98498 183922 98566 183978
rect 98622 183922 98690 183978
rect 98746 183922 98814 183978
rect 98870 183922 98894 183978
rect 98418 183888 98894 183922
rect 99932 173818 99988 268044
rect 100044 178858 100100 271180
rect 100044 178792 100100 178802
rect 101298 262350 101918 279922
rect 106652 279658 106708 279668
rect 105308 279076 105364 279086
rect 105308 277956 105364 279020
rect 105308 277890 105364 277900
rect 103628 275604 103684 275614
rect 103404 274708 103460 274718
rect 101298 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 101918 262350
rect 101298 262226 101918 262294
rect 101298 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 101918 262226
rect 101298 262102 101918 262170
rect 101298 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 101918 262102
rect 101298 261978 101918 262046
rect 101298 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 101918 261978
rect 101298 244350 101918 261922
rect 101298 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 101918 244350
rect 101298 244226 101918 244294
rect 101298 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 101918 244226
rect 101298 244102 101918 244170
rect 101298 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 101918 244102
rect 101298 243978 101918 244046
rect 101298 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 101918 243978
rect 101298 226350 101918 243922
rect 101298 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 101918 226350
rect 101298 226226 101918 226294
rect 101298 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 101918 226226
rect 101298 226102 101918 226170
rect 101298 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 101918 226102
rect 101298 225978 101918 226046
rect 101298 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 101918 225978
rect 101298 208350 101918 225922
rect 101298 208294 101394 208350
rect 101450 208294 101518 208350
rect 101574 208294 101642 208350
rect 101698 208294 101766 208350
rect 101822 208294 101918 208350
rect 101298 208226 101918 208294
rect 101298 208170 101394 208226
rect 101450 208170 101518 208226
rect 101574 208170 101642 208226
rect 101698 208170 101766 208226
rect 101822 208170 101918 208226
rect 101298 208102 101918 208170
rect 101298 208046 101394 208102
rect 101450 208046 101518 208102
rect 101574 208046 101642 208102
rect 101698 208046 101766 208102
rect 101822 208046 101918 208102
rect 101298 207978 101918 208046
rect 101298 207922 101394 207978
rect 101450 207922 101518 207978
rect 101574 207922 101642 207978
rect 101698 207922 101766 207978
rect 101822 207922 101918 207978
rect 101298 190350 101918 207922
rect 101298 190294 101394 190350
rect 101450 190294 101518 190350
rect 101574 190294 101642 190350
rect 101698 190294 101766 190350
rect 101822 190294 101918 190350
rect 101298 190226 101918 190294
rect 101298 190170 101394 190226
rect 101450 190170 101518 190226
rect 101574 190170 101642 190226
rect 101698 190170 101766 190226
rect 101822 190170 101918 190226
rect 101298 190102 101918 190170
rect 101298 190046 101394 190102
rect 101450 190046 101518 190102
rect 101574 190046 101642 190102
rect 101698 190046 101766 190102
rect 101822 190046 101918 190102
rect 101298 189978 101918 190046
rect 101298 189922 101394 189978
rect 101450 189922 101518 189978
rect 101574 189922 101642 189978
rect 101698 189922 101766 189978
rect 101822 189922 101918 189978
rect 99932 173752 99988 173762
rect 97618 172350 98094 172384
rect 97618 172294 97642 172350
rect 97698 172294 97766 172350
rect 97822 172294 97890 172350
rect 97946 172294 98014 172350
rect 98070 172294 98094 172350
rect 97618 172226 98094 172294
rect 97618 172170 97642 172226
rect 97698 172170 97766 172226
rect 97822 172170 97890 172226
rect 97946 172170 98014 172226
rect 98070 172170 98094 172226
rect 97618 172102 98094 172170
rect 97618 172046 97642 172102
rect 97698 172046 97766 172102
rect 97822 172046 97890 172102
rect 97946 172046 98014 172102
rect 98070 172046 98094 172102
rect 97618 171978 98094 172046
rect 97618 171922 97642 171978
rect 97698 171922 97766 171978
rect 97822 171922 97890 171978
rect 97946 171922 98014 171978
rect 98070 171922 98094 171978
rect 97618 171888 98094 171922
rect 101298 172350 101918 189922
rect 101298 172294 101394 172350
rect 101450 172294 101518 172350
rect 101574 172294 101642 172350
rect 101698 172294 101766 172350
rect 101822 172294 101918 172350
rect 101298 172226 101918 172294
rect 101298 172170 101394 172226
rect 101450 172170 101518 172226
rect 101574 172170 101642 172226
rect 101698 172170 101766 172226
rect 101822 172170 101918 172226
rect 101298 172102 101918 172170
rect 101298 172046 101394 172102
rect 101450 172046 101518 172102
rect 101574 172046 101642 172102
rect 101698 172046 101766 172102
rect 101822 172046 101918 172102
rect 101298 171978 101918 172046
rect 101298 171922 101394 171978
rect 101450 171922 101518 171978
rect 101574 171922 101642 171978
rect 101698 171922 101766 171978
rect 101822 171922 101918 171978
rect 94892 164546 94948 164556
rect 97578 166350 98198 166456
rect 97578 166294 97674 166350
rect 97730 166294 97798 166350
rect 97854 166294 97922 166350
rect 97978 166294 98046 166350
rect 98102 166294 98198 166350
rect 97578 166226 98198 166294
rect 97578 166170 97674 166226
rect 97730 166170 97798 166226
rect 97854 166170 97922 166226
rect 97978 166170 98046 166226
rect 98102 166170 98198 166226
rect 97578 166102 98198 166170
rect 97578 166046 97674 166102
rect 97730 166046 97798 166102
rect 97854 166046 97922 166102
rect 97978 166046 98046 166102
rect 98102 166046 98198 166102
rect 97578 165978 98198 166046
rect 97578 165922 97674 165978
rect 97730 165922 97798 165978
rect 97854 165922 97922 165978
rect 97978 165922 98046 165978
rect 98102 165922 98198 165978
rect 83916 147858 83972 147868
rect 97578 148350 98198 165922
rect 97578 148294 97674 148350
rect 97730 148294 97798 148350
rect 97854 148294 97922 148350
rect 97978 148294 98046 148350
rect 98102 148294 98198 148350
rect 97578 148226 98198 148294
rect 97578 148170 97674 148226
rect 97730 148170 97798 148226
rect 97854 148170 97922 148226
rect 97978 148170 98046 148226
rect 98102 148170 98198 148226
rect 97578 148102 98198 148170
rect 97578 148046 97674 148102
rect 97730 148046 97798 148102
rect 97854 148046 97922 148102
rect 97978 148046 98046 148102
rect 98102 148046 98198 148102
rect 97578 147978 98198 148046
rect 97578 147922 97674 147978
rect 97730 147922 97798 147978
rect 97854 147922 97922 147978
rect 97978 147922 98046 147978
rect 98102 147922 98198 147978
rect 70578 136294 70674 136350
rect 70730 136294 70798 136350
rect 70854 136294 70922 136350
rect 70978 136294 71046 136350
rect 71102 136294 71198 136350
rect 70578 136226 71198 136294
rect 70578 136170 70674 136226
rect 70730 136170 70798 136226
rect 70854 136170 70922 136226
rect 70978 136170 71046 136226
rect 71102 136170 71198 136226
rect 70578 136102 71198 136170
rect 70578 136046 70674 136102
rect 70730 136046 70798 136102
rect 70854 136046 70922 136102
rect 70978 136046 71046 136102
rect 71102 136046 71198 136102
rect 70578 135978 71198 136046
rect 70578 135922 70674 135978
rect 70730 135922 70798 135978
rect 70854 135922 70922 135978
rect 70978 135922 71046 135978
rect 71102 135922 71198 135978
rect 70578 118350 71198 135922
rect 96588 136350 97064 136384
rect 96588 136294 96612 136350
rect 96668 136294 96736 136350
rect 96792 136294 96860 136350
rect 96916 136294 96984 136350
rect 97040 136294 97064 136350
rect 96588 136226 97064 136294
rect 96588 136170 96612 136226
rect 96668 136170 96736 136226
rect 96792 136170 96860 136226
rect 96916 136170 96984 136226
rect 97040 136170 97064 136226
rect 96588 136102 97064 136170
rect 96588 136046 96612 136102
rect 96668 136046 96736 136102
rect 96792 136046 96860 136102
rect 96916 136046 96984 136102
rect 97040 136046 97064 136102
rect 96588 135978 97064 136046
rect 96588 135922 96612 135978
rect 96668 135922 96736 135978
rect 96792 135922 96860 135978
rect 96916 135922 96984 135978
rect 97040 135922 97064 135978
rect 96588 135888 97064 135922
rect 95788 130350 96264 130384
rect 95788 130294 95812 130350
rect 95868 130294 95936 130350
rect 95992 130294 96060 130350
rect 96116 130294 96184 130350
rect 96240 130294 96264 130350
rect 95788 130226 96264 130294
rect 95788 130170 95812 130226
rect 95868 130170 95936 130226
rect 95992 130170 96060 130226
rect 96116 130170 96184 130226
rect 96240 130170 96264 130226
rect 95788 130102 96264 130170
rect 95788 130046 95812 130102
rect 95868 130046 95936 130102
rect 95992 130046 96060 130102
rect 96116 130046 96184 130102
rect 96240 130046 96264 130102
rect 95788 129978 96264 130046
rect 95788 129922 95812 129978
rect 95868 129922 95936 129978
rect 95992 129922 96060 129978
rect 96116 129922 96184 129978
rect 96240 129922 96264 129978
rect 95788 129888 96264 129922
rect 97578 130350 98198 147922
rect 97578 130294 97674 130350
rect 97730 130294 97798 130350
rect 97854 130294 97922 130350
rect 97978 130294 98046 130350
rect 98102 130294 98198 130350
rect 97578 130226 98198 130294
rect 97578 130170 97674 130226
rect 97730 130170 97798 130226
rect 97854 130170 97922 130226
rect 97978 130170 98046 130226
rect 98102 130170 98198 130226
rect 97578 130102 98198 130170
rect 97578 130046 97674 130102
rect 97730 130046 97798 130102
rect 97854 130046 97922 130102
rect 97978 130046 98046 130102
rect 98102 130046 98198 130102
rect 97578 129978 98198 130046
rect 97578 129922 97674 129978
rect 97730 129922 97798 129978
rect 97854 129922 97922 129978
rect 97978 129922 98046 129978
rect 98102 129922 98198 129978
rect 70578 118294 70674 118350
rect 70730 118294 70798 118350
rect 70854 118294 70922 118350
rect 70978 118294 71046 118350
rect 71102 118294 71198 118350
rect 70578 118226 71198 118294
rect 70578 118170 70674 118226
rect 70730 118170 70798 118226
rect 70854 118170 70922 118226
rect 70978 118170 71046 118226
rect 71102 118170 71198 118226
rect 70578 118102 71198 118170
rect 70578 118046 70674 118102
rect 70730 118046 70798 118102
rect 70854 118046 70922 118102
rect 70978 118046 71046 118102
rect 71102 118046 71198 118102
rect 70578 117978 71198 118046
rect 70578 117922 70674 117978
rect 70730 117922 70798 117978
rect 70854 117922 70922 117978
rect 70978 117922 71046 117978
rect 71102 117922 71198 117978
rect 70578 100350 71198 117922
rect 96588 118350 97064 118384
rect 96588 118294 96612 118350
rect 96668 118294 96736 118350
rect 96792 118294 96860 118350
rect 96916 118294 96984 118350
rect 97040 118294 97064 118350
rect 96588 118226 97064 118294
rect 96588 118170 96612 118226
rect 96668 118170 96736 118226
rect 96792 118170 96860 118226
rect 96916 118170 96984 118226
rect 97040 118170 97064 118226
rect 96588 118102 97064 118170
rect 96588 118046 96612 118102
rect 96668 118046 96736 118102
rect 96792 118046 96860 118102
rect 96916 118046 96984 118102
rect 97040 118046 97064 118102
rect 96588 117978 97064 118046
rect 96588 117922 96612 117978
rect 96668 117922 96736 117978
rect 96792 117922 96860 117978
rect 96916 117922 96984 117978
rect 97040 117922 97064 117978
rect 96588 117888 97064 117922
rect 95788 112350 96264 112384
rect 95788 112294 95812 112350
rect 95868 112294 95936 112350
rect 95992 112294 96060 112350
rect 96116 112294 96184 112350
rect 96240 112294 96264 112350
rect 95788 112226 96264 112294
rect 95788 112170 95812 112226
rect 95868 112170 95936 112226
rect 95992 112170 96060 112226
rect 96116 112170 96184 112226
rect 96240 112170 96264 112226
rect 95788 112102 96264 112170
rect 95788 112046 95812 112102
rect 95868 112046 95936 112102
rect 95992 112046 96060 112102
rect 96116 112046 96184 112102
rect 96240 112046 96264 112102
rect 95788 111978 96264 112046
rect 95788 111922 95812 111978
rect 95868 111922 95936 111978
rect 95992 111922 96060 111978
rect 96116 111922 96184 111978
rect 96240 111922 96264 111978
rect 95788 111888 96264 111922
rect 97578 112350 98198 129922
rect 97578 112294 97674 112350
rect 97730 112294 97798 112350
rect 97854 112294 97922 112350
rect 97978 112294 98046 112350
rect 98102 112294 98198 112350
rect 97578 112226 98198 112294
rect 97578 112170 97674 112226
rect 97730 112170 97798 112226
rect 97854 112170 97922 112226
rect 97978 112170 98046 112226
rect 98102 112170 98198 112226
rect 97578 112102 98198 112170
rect 97578 112046 97674 112102
rect 97730 112046 97798 112102
rect 97854 112046 97922 112102
rect 97978 112046 98046 112102
rect 98102 112046 98198 112102
rect 97578 111978 98198 112046
rect 97578 111922 97674 111978
rect 97730 111922 97798 111978
rect 97854 111922 97922 111978
rect 97978 111922 98046 111978
rect 98102 111922 98198 111978
rect 70578 100294 70674 100350
rect 70730 100294 70798 100350
rect 70854 100294 70922 100350
rect 70978 100294 71046 100350
rect 71102 100294 71198 100350
rect 70578 100226 71198 100294
rect 70578 100170 70674 100226
rect 70730 100170 70798 100226
rect 70854 100170 70922 100226
rect 70978 100170 71046 100226
rect 71102 100170 71198 100226
rect 70578 100102 71198 100170
rect 70578 100046 70674 100102
rect 70730 100046 70798 100102
rect 70854 100046 70922 100102
rect 70978 100046 71046 100102
rect 71102 100046 71198 100102
rect 70578 99978 71198 100046
rect 70578 99922 70674 99978
rect 70730 99922 70798 99978
rect 70854 99922 70922 99978
rect 70978 99922 71046 99978
rect 71102 99922 71198 99978
rect 70578 82350 71198 99922
rect 96588 100350 97064 100384
rect 96588 100294 96612 100350
rect 96668 100294 96736 100350
rect 96792 100294 96860 100350
rect 96916 100294 96984 100350
rect 97040 100294 97064 100350
rect 96588 100226 97064 100294
rect 96588 100170 96612 100226
rect 96668 100170 96736 100226
rect 96792 100170 96860 100226
rect 96916 100170 96984 100226
rect 97040 100170 97064 100226
rect 96588 100102 97064 100170
rect 96588 100046 96612 100102
rect 96668 100046 96736 100102
rect 96792 100046 96860 100102
rect 96916 100046 96984 100102
rect 97040 100046 97064 100102
rect 96588 99978 97064 100046
rect 96588 99922 96612 99978
rect 96668 99922 96736 99978
rect 96792 99922 96860 99978
rect 96916 99922 96984 99978
rect 97040 99922 97064 99978
rect 96588 99888 97064 99922
rect 95788 94350 96264 94384
rect 95788 94294 95812 94350
rect 95868 94294 95936 94350
rect 95992 94294 96060 94350
rect 96116 94294 96184 94350
rect 96240 94294 96264 94350
rect 95788 94226 96264 94294
rect 95788 94170 95812 94226
rect 95868 94170 95936 94226
rect 95992 94170 96060 94226
rect 96116 94170 96184 94226
rect 96240 94170 96264 94226
rect 95788 94102 96264 94170
rect 95788 94046 95812 94102
rect 95868 94046 95936 94102
rect 95992 94046 96060 94102
rect 96116 94046 96184 94102
rect 96240 94046 96264 94102
rect 95788 93978 96264 94046
rect 95788 93922 95812 93978
rect 95868 93922 95936 93978
rect 95992 93922 96060 93978
rect 96116 93922 96184 93978
rect 96240 93922 96264 93978
rect 95788 93888 96264 93922
rect 97578 94350 98198 111922
rect 97578 94294 97674 94350
rect 97730 94294 97798 94350
rect 97854 94294 97922 94350
rect 97978 94294 98046 94350
rect 98102 94294 98198 94350
rect 97578 94226 98198 94294
rect 97578 94170 97674 94226
rect 97730 94170 97798 94226
rect 97854 94170 97922 94226
rect 97978 94170 98046 94226
rect 98102 94170 98198 94226
rect 97578 94102 98198 94170
rect 97578 94046 97674 94102
rect 97730 94046 97798 94102
rect 97854 94046 97922 94102
rect 97978 94046 98046 94102
rect 98102 94046 98198 94102
rect 97578 93978 98198 94046
rect 97578 93922 97674 93978
rect 97730 93922 97798 93978
rect 97854 93922 97922 93978
rect 97978 93922 98046 93978
rect 98102 93922 98198 93978
rect 70578 82294 70674 82350
rect 70730 82294 70798 82350
rect 70854 82294 70922 82350
rect 70978 82294 71046 82350
rect 71102 82294 71198 82350
rect 70578 82226 71198 82294
rect 70578 82170 70674 82226
rect 70730 82170 70798 82226
rect 70854 82170 70922 82226
rect 70978 82170 71046 82226
rect 71102 82170 71198 82226
rect 70578 82102 71198 82170
rect 70578 82046 70674 82102
rect 70730 82046 70798 82102
rect 70854 82046 70922 82102
rect 70978 82046 71046 82102
rect 71102 82046 71198 82102
rect 70578 81978 71198 82046
rect 70578 81922 70674 81978
rect 70730 81922 70798 81978
rect 70854 81922 70922 81978
rect 70978 81922 71046 81978
rect 71102 81922 71198 81978
rect 70578 64350 71198 81922
rect 96588 82350 97064 82384
rect 96588 82294 96612 82350
rect 96668 82294 96736 82350
rect 96792 82294 96860 82350
rect 96916 82294 96984 82350
rect 97040 82294 97064 82350
rect 96588 82226 97064 82294
rect 96588 82170 96612 82226
rect 96668 82170 96736 82226
rect 96792 82170 96860 82226
rect 96916 82170 96984 82226
rect 97040 82170 97064 82226
rect 96588 82102 97064 82170
rect 96588 82046 96612 82102
rect 96668 82046 96736 82102
rect 96792 82046 96860 82102
rect 96916 82046 96984 82102
rect 97040 82046 97064 82102
rect 96588 81978 97064 82046
rect 96588 81922 96612 81978
rect 96668 81922 96736 81978
rect 96792 81922 96860 81978
rect 96916 81922 96984 81978
rect 97040 81922 97064 81978
rect 96588 81888 97064 81922
rect 95788 76350 96264 76384
rect 95788 76294 95812 76350
rect 95868 76294 95936 76350
rect 95992 76294 96060 76350
rect 96116 76294 96184 76350
rect 96240 76294 96264 76350
rect 95788 76226 96264 76294
rect 95788 76170 95812 76226
rect 95868 76170 95936 76226
rect 95992 76170 96060 76226
rect 96116 76170 96184 76226
rect 96240 76170 96264 76226
rect 95788 76102 96264 76170
rect 95788 76046 95812 76102
rect 95868 76046 95936 76102
rect 95992 76046 96060 76102
rect 96116 76046 96184 76102
rect 96240 76046 96264 76102
rect 95788 75978 96264 76046
rect 95788 75922 95812 75978
rect 95868 75922 95936 75978
rect 95992 75922 96060 75978
rect 96116 75922 96184 75978
rect 96240 75922 96264 75978
rect 95788 75888 96264 75922
rect 97578 76350 98198 93922
rect 97578 76294 97674 76350
rect 97730 76294 97798 76350
rect 97854 76294 97922 76350
rect 97978 76294 98046 76350
rect 98102 76294 98198 76350
rect 97578 76226 98198 76294
rect 97578 76170 97674 76226
rect 97730 76170 97798 76226
rect 97854 76170 97922 76226
rect 97978 76170 98046 76226
rect 98102 76170 98198 76226
rect 97578 76102 98198 76170
rect 97578 76046 97674 76102
rect 97730 76046 97798 76102
rect 97854 76046 97922 76102
rect 97978 76046 98046 76102
rect 98102 76046 98198 76102
rect 97578 75978 98198 76046
rect 97578 75922 97674 75978
rect 97730 75922 97798 75978
rect 97854 75922 97922 75978
rect 97978 75922 98046 75978
rect 98102 75922 98198 75978
rect 70578 64294 70674 64350
rect 70730 64294 70798 64350
rect 70854 64294 70922 64350
rect 70978 64294 71046 64350
rect 71102 64294 71198 64350
rect 70578 64226 71198 64294
rect 70578 64170 70674 64226
rect 70730 64170 70798 64226
rect 70854 64170 70922 64226
rect 70978 64170 71046 64226
rect 71102 64170 71198 64226
rect 70578 64102 71198 64170
rect 70578 64046 70674 64102
rect 70730 64046 70798 64102
rect 70854 64046 70922 64102
rect 70978 64046 71046 64102
rect 71102 64046 71198 64102
rect 70578 63978 71198 64046
rect 70578 63922 70674 63978
rect 70730 63922 70798 63978
rect 70854 63922 70922 63978
rect 70978 63922 71046 63978
rect 71102 63922 71198 63978
rect 70578 46350 71198 63922
rect 96588 64350 97064 64384
rect 96588 64294 96612 64350
rect 96668 64294 96736 64350
rect 96792 64294 96860 64350
rect 96916 64294 96984 64350
rect 97040 64294 97064 64350
rect 96588 64226 97064 64294
rect 96588 64170 96612 64226
rect 96668 64170 96736 64226
rect 96792 64170 96860 64226
rect 96916 64170 96984 64226
rect 97040 64170 97064 64226
rect 96588 64102 97064 64170
rect 96588 64046 96612 64102
rect 96668 64046 96736 64102
rect 96792 64046 96860 64102
rect 96916 64046 96984 64102
rect 97040 64046 97064 64102
rect 96588 63978 97064 64046
rect 96588 63922 96612 63978
rect 96668 63922 96736 63978
rect 96792 63922 96860 63978
rect 96916 63922 96984 63978
rect 97040 63922 97064 63978
rect 96588 63888 97064 63922
rect 95788 58350 96264 58384
rect 95788 58294 95812 58350
rect 95868 58294 95936 58350
rect 95992 58294 96060 58350
rect 96116 58294 96184 58350
rect 96240 58294 96264 58350
rect 95788 58226 96264 58294
rect 95788 58170 95812 58226
rect 95868 58170 95936 58226
rect 95992 58170 96060 58226
rect 96116 58170 96184 58226
rect 96240 58170 96264 58226
rect 95788 58102 96264 58170
rect 95788 58046 95812 58102
rect 95868 58046 95936 58102
rect 95992 58046 96060 58102
rect 96116 58046 96184 58102
rect 96240 58046 96264 58102
rect 95788 57978 96264 58046
rect 95788 57922 95812 57978
rect 95868 57922 95936 57978
rect 95992 57922 96060 57978
rect 96116 57922 96184 57978
rect 96240 57922 96264 57978
rect 95788 57888 96264 57922
rect 97578 58350 98198 75922
rect 97578 58294 97674 58350
rect 97730 58294 97798 58350
rect 97854 58294 97922 58350
rect 97978 58294 98046 58350
rect 98102 58294 98198 58350
rect 97578 58226 98198 58294
rect 97578 58170 97674 58226
rect 97730 58170 97798 58226
rect 97854 58170 97922 58226
rect 97978 58170 98046 58226
rect 98102 58170 98198 58226
rect 97578 58102 98198 58170
rect 97578 58046 97674 58102
rect 97730 58046 97798 58102
rect 97854 58046 97922 58102
rect 97978 58046 98046 58102
rect 98102 58046 98198 58102
rect 97578 57978 98198 58046
rect 97578 57922 97674 57978
rect 97730 57922 97798 57978
rect 97854 57922 97922 57978
rect 97978 57922 98046 57978
rect 98102 57922 98198 57978
rect 70578 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 71198 46350
rect 70578 46226 71198 46294
rect 70578 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 71198 46226
rect 70578 46102 71198 46170
rect 70578 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 71198 46102
rect 70578 45978 71198 46046
rect 70578 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 71198 45978
rect 70578 28350 71198 45922
rect 70578 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 71198 28350
rect 70578 28226 71198 28294
rect 70578 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 71198 28226
rect 70578 28102 71198 28170
rect 70578 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 71198 28102
rect 70578 27978 71198 28046
rect 70578 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 71198 27978
rect 70578 10350 71198 27922
rect 97578 40350 98198 57922
rect 97578 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 98198 40350
rect 97578 40226 98198 40294
rect 97578 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 98198 40226
rect 97578 40102 98198 40170
rect 97578 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 98198 40102
rect 97578 39978 98198 40046
rect 97578 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 98198 39978
rect 85836 22350 86156 22384
rect 85836 22294 85906 22350
rect 85962 22294 86030 22350
rect 86086 22294 86156 22350
rect 85836 22226 86156 22294
rect 85836 22170 85906 22226
rect 85962 22170 86030 22226
rect 86086 22170 86156 22226
rect 85836 22102 86156 22170
rect 85836 22046 85906 22102
rect 85962 22046 86030 22102
rect 86086 22046 86156 22102
rect 85836 21978 86156 22046
rect 85836 21922 85906 21978
rect 85962 21922 86030 21978
rect 86086 21922 86156 21978
rect 85836 21888 86156 21922
rect 97578 22350 98198 39922
rect 97578 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 98198 22350
rect 97578 22226 98198 22294
rect 97578 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 98198 22226
rect 97578 22102 98198 22170
rect 97578 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 98198 22102
rect 97578 21978 98198 22046
rect 97578 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 98198 21978
rect 70578 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 71198 10350
rect 70578 10226 71198 10294
rect 70578 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 71198 10226
rect 70578 10102 71198 10170
rect 70578 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 71198 10102
rect 70578 9978 71198 10046
rect 70578 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 71198 9978
rect 70578 -1120 71198 9922
rect 70578 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 71198 -1120
rect 70578 -1244 71198 -1176
rect 70578 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 71198 -1244
rect 70578 -1368 71198 -1300
rect 70578 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 71198 -1368
rect 70578 -1492 71198 -1424
rect 70578 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 71198 -1492
rect 70578 -1644 71198 -1548
rect 97578 4350 98198 21922
rect 97578 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 98198 4350
rect 97578 4226 98198 4294
rect 97578 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 98198 4226
rect 97578 4102 98198 4170
rect 97578 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 98198 4102
rect 97578 3978 98198 4046
rect 97578 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 98198 3978
rect 97578 -160 98198 3922
rect 97578 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 98198 -160
rect 97578 -284 98198 -216
rect 97578 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 98198 -284
rect 97578 -408 98198 -340
rect 97578 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 98198 -408
rect 97578 -532 98198 -464
rect 97578 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 98198 -532
rect 97578 -1644 98198 -588
rect 101298 154350 101918 171922
rect 101298 154294 101394 154350
rect 101450 154294 101518 154350
rect 101574 154294 101642 154350
rect 101698 154294 101766 154350
rect 101822 154294 101918 154350
rect 101298 154226 101918 154294
rect 101298 154170 101394 154226
rect 101450 154170 101518 154226
rect 101574 154170 101642 154226
rect 101698 154170 101766 154226
rect 101822 154170 101918 154226
rect 101298 154102 101918 154170
rect 101298 154046 101394 154102
rect 101450 154046 101518 154102
rect 101574 154046 101642 154102
rect 101698 154046 101766 154102
rect 101822 154046 101918 154102
rect 101298 153978 101918 154046
rect 101298 153922 101394 153978
rect 101450 153922 101518 153978
rect 101574 153922 101642 153978
rect 101698 153922 101766 153978
rect 101822 153922 101918 153978
rect 101298 136350 101918 153922
rect 103292 264898 103348 264908
rect 103292 149716 103348 264842
rect 103404 162658 103460 274652
rect 103516 271378 103572 271388
rect 103516 177238 103572 271322
rect 103628 205858 103684 275548
rect 103628 205792 103684 205802
rect 104972 264740 105028 264750
rect 104972 181558 105028 264684
rect 104972 181492 105028 181502
rect 103516 177172 103572 177182
rect 106652 162708 106708 279602
rect 106764 276836 106820 326042
rect 106764 276770 106820 276780
rect 108332 273358 108388 544796
rect 110012 431956 110068 431966
rect 109116 365158 109172 365168
rect 108332 273292 108388 273302
rect 108444 357598 108500 357608
rect 108332 266878 108388 266888
rect 108332 163828 108388 266822
rect 108332 163762 108388 163772
rect 106652 162642 106708 162652
rect 103404 162592 103460 162602
rect 108444 152180 108500 357542
rect 108668 339444 108724 339454
rect 108556 279478 108612 279488
rect 108556 162372 108612 279422
rect 108668 276052 108724 339388
rect 109116 337204 109172 365102
rect 109116 336084 109172 337148
rect 109116 336018 109172 336028
rect 110012 278398 110068 431900
rect 110012 278332 110068 278342
rect 110124 366598 110180 366608
rect 108668 275986 108724 275996
rect 108556 162306 108612 162316
rect 110012 268498 110068 268508
rect 108444 152114 108500 152124
rect 103292 149650 103348 149660
rect 101298 136294 101394 136350
rect 101450 136294 101518 136350
rect 101574 136294 101642 136350
rect 101698 136294 101766 136350
rect 101822 136294 101918 136350
rect 101298 136226 101918 136294
rect 101298 136170 101394 136226
rect 101450 136170 101518 136226
rect 101574 136170 101642 136226
rect 101698 136170 101766 136226
rect 101822 136170 101918 136226
rect 101298 136102 101918 136170
rect 101298 136046 101394 136102
rect 101450 136046 101518 136102
rect 101574 136046 101642 136102
rect 101698 136046 101766 136102
rect 101822 136046 101918 136102
rect 101298 135978 101918 136046
rect 101298 135922 101394 135978
rect 101450 135922 101518 135978
rect 101574 135922 101642 135978
rect 101698 135922 101766 135978
rect 101822 135922 101918 135978
rect 101298 118350 101918 135922
rect 101298 118294 101394 118350
rect 101450 118294 101518 118350
rect 101574 118294 101642 118350
rect 101698 118294 101766 118350
rect 101822 118294 101918 118350
rect 101298 118226 101918 118294
rect 101298 118170 101394 118226
rect 101450 118170 101518 118226
rect 101574 118170 101642 118226
rect 101698 118170 101766 118226
rect 101822 118170 101918 118226
rect 101298 118102 101918 118170
rect 101298 118046 101394 118102
rect 101450 118046 101518 118102
rect 101574 118046 101642 118102
rect 101698 118046 101766 118102
rect 101822 118046 101918 118102
rect 101298 117978 101918 118046
rect 101298 117922 101394 117978
rect 101450 117922 101518 117978
rect 101574 117922 101642 117978
rect 101698 117922 101766 117978
rect 101822 117922 101918 117978
rect 101298 100350 101918 117922
rect 101298 100294 101394 100350
rect 101450 100294 101518 100350
rect 101574 100294 101642 100350
rect 101698 100294 101766 100350
rect 101822 100294 101918 100350
rect 101298 100226 101918 100294
rect 101298 100170 101394 100226
rect 101450 100170 101518 100226
rect 101574 100170 101642 100226
rect 101698 100170 101766 100226
rect 101822 100170 101918 100226
rect 101298 100102 101918 100170
rect 101298 100046 101394 100102
rect 101450 100046 101518 100102
rect 101574 100046 101642 100102
rect 101698 100046 101766 100102
rect 101822 100046 101918 100102
rect 101298 99978 101918 100046
rect 101298 99922 101394 99978
rect 101450 99922 101518 99978
rect 101574 99922 101642 99978
rect 101698 99922 101766 99978
rect 101822 99922 101918 99978
rect 101298 82350 101918 99922
rect 101298 82294 101394 82350
rect 101450 82294 101518 82350
rect 101574 82294 101642 82350
rect 101698 82294 101766 82350
rect 101822 82294 101918 82350
rect 101298 82226 101918 82294
rect 101298 82170 101394 82226
rect 101450 82170 101518 82226
rect 101574 82170 101642 82226
rect 101698 82170 101766 82226
rect 101822 82170 101918 82226
rect 101298 82102 101918 82170
rect 101298 82046 101394 82102
rect 101450 82046 101518 82102
rect 101574 82046 101642 82102
rect 101698 82046 101766 82102
rect 101822 82046 101918 82102
rect 101298 81978 101918 82046
rect 101298 81922 101394 81978
rect 101450 81922 101518 81978
rect 101574 81922 101642 81978
rect 101698 81922 101766 81978
rect 101822 81922 101918 81978
rect 101298 64350 101918 81922
rect 101298 64294 101394 64350
rect 101450 64294 101518 64350
rect 101574 64294 101642 64350
rect 101698 64294 101766 64350
rect 101822 64294 101918 64350
rect 101298 64226 101918 64294
rect 101298 64170 101394 64226
rect 101450 64170 101518 64226
rect 101574 64170 101642 64226
rect 101698 64170 101766 64226
rect 101822 64170 101918 64226
rect 101298 64102 101918 64170
rect 101298 64046 101394 64102
rect 101450 64046 101518 64102
rect 101574 64046 101642 64102
rect 101698 64046 101766 64102
rect 101822 64046 101918 64102
rect 101298 63978 101918 64046
rect 101298 63922 101394 63978
rect 101450 63922 101518 63978
rect 101574 63922 101642 63978
rect 101698 63922 101766 63978
rect 101822 63922 101918 63978
rect 101298 46350 101918 63922
rect 101298 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 101918 46350
rect 101298 46226 101918 46294
rect 101298 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 101918 46226
rect 101298 46102 101918 46170
rect 101298 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 101918 46102
rect 101298 45978 101918 46046
rect 101298 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 101918 45978
rect 101298 28350 101918 45922
rect 110012 36820 110068 268442
rect 110124 149518 110180 366542
rect 110124 149452 110180 149462
rect 110236 360118 110292 360128
rect 110236 148596 110292 360062
rect 110348 357958 110404 357968
rect 110348 149338 110404 357902
rect 110908 300916 110964 300926
rect 110908 278908 110964 300860
rect 111132 278964 111188 278974
rect 110908 278852 111188 278908
rect 110908 278218 110964 278852
rect 110908 278152 110964 278162
rect 111692 271738 111748 590940
rect 120092 590772 120148 590782
rect 111692 271672 111748 271682
rect 111804 558964 111860 558974
rect 111804 269938 111860 558908
rect 114268 474292 114324 474302
rect 112476 365540 112532 365550
rect 112364 359938 112420 359948
rect 111916 328468 111972 328478
rect 111916 300020 111972 328412
rect 112252 327908 112308 327918
rect 111916 299954 111972 299964
rect 112028 324436 112084 324446
rect 112028 297668 112084 324380
rect 112252 299124 112308 327852
rect 112252 299058 112308 299068
rect 112028 297602 112084 297612
rect 111804 269872 111860 269882
rect 111916 274618 111972 274628
rect 111692 268100 111748 268110
rect 111692 206578 111748 268044
rect 111692 206512 111748 206522
rect 111916 162838 111972 274562
rect 111916 162772 111972 162782
rect 110348 149272 110404 149282
rect 110236 148530 110292 148540
rect 112364 148596 112420 359882
rect 112476 149518 112532 365484
rect 114156 363412 114212 363422
rect 112588 346948 112644 346958
rect 112588 338772 112644 346892
rect 112588 338706 112644 338716
rect 114156 332038 114212 363356
rect 114156 331044 114212 331982
rect 114156 330978 114212 330988
rect 112588 327796 112644 327806
rect 112588 317492 112644 327740
rect 113484 325780 113540 325790
rect 113260 323428 113316 323438
rect 112588 317426 112644 317436
rect 113036 323092 113092 323102
rect 113036 312598 113092 323036
rect 113036 312532 113092 312542
rect 113148 319732 113204 319742
rect 113148 312228 113204 319676
rect 113148 312162 113204 312172
rect 113260 300244 113316 323372
rect 113372 321748 113428 321758
rect 113372 311108 113428 321692
rect 113372 311042 113428 311052
rect 113260 300178 113316 300188
rect 112700 299124 112756 299134
rect 112588 295652 112644 295662
rect 112588 291508 112644 295596
rect 112588 291442 112644 291452
rect 112700 286132 112756 299068
rect 113484 291956 113540 325724
rect 113820 325108 113876 325118
rect 113708 323764 113764 323774
rect 113596 322420 113652 322430
rect 113596 293188 113652 322364
rect 113596 293122 113652 293132
rect 113484 291890 113540 291900
rect 113708 291396 113764 323708
rect 113820 300580 113876 325052
rect 114268 324212 114324 474236
rect 119196 364978 119252 364988
rect 117516 362278 117572 362288
rect 117404 355908 117460 355918
rect 117180 352548 117236 352558
rect 116620 350308 116676 350318
rect 116620 338884 116676 350252
rect 116620 338818 116676 338828
rect 116732 340228 116788 340238
rect 114268 324146 114324 324156
rect 115052 329812 115108 329822
rect 114828 321188 114884 321198
rect 113820 300514 113876 300524
rect 113932 316372 113988 316382
rect 113708 291330 113764 291340
rect 113932 290948 113988 316316
rect 113932 290882 113988 290892
rect 114044 312564 114100 312574
rect 112700 286066 112756 286076
rect 112812 290836 112868 290846
rect 112812 278908 112868 290780
rect 114044 289492 114100 312508
rect 114268 310996 114324 311016
rect 114268 310912 114324 310922
rect 114828 306292 114884 321132
rect 114828 306226 114884 306236
rect 115052 305508 115108 329756
rect 115948 329028 116004 329038
rect 115948 326098 116004 328972
rect 115948 326032 116004 326042
rect 115276 325668 115332 325678
rect 115052 305442 115108 305452
rect 115164 317716 115220 317726
rect 114716 291956 114772 291966
rect 114044 289426 114100 289436
rect 114268 291396 114324 291406
rect 114268 288708 114324 291340
rect 114716 289828 114772 291900
rect 114716 289762 114772 289772
rect 114268 288642 114324 288652
rect 112700 278852 112868 278908
rect 113372 284564 113428 284574
rect 112700 278180 112756 278852
rect 112700 261658 112756 278124
rect 113372 278292 113428 284508
rect 115164 282324 115220 317660
rect 115276 295652 115332 325612
rect 115500 324548 115556 324558
rect 115276 295586 115332 295596
rect 115388 320068 115444 320078
rect 115388 292852 115444 320012
rect 115500 296212 115556 324492
rect 115612 322308 115668 322318
rect 115612 302932 115668 322252
rect 116620 319060 116676 319070
rect 115948 317044 116004 317054
rect 115836 316708 115892 316718
rect 115724 315700 115780 315710
rect 115724 304388 115780 315644
rect 115836 314356 115892 316652
rect 115836 314290 115892 314300
rect 115948 309988 116004 316988
rect 116620 313348 116676 319004
rect 116620 313282 116676 313292
rect 115948 309922 116004 309932
rect 115724 304322 115780 304332
rect 115612 302866 115668 302876
rect 115500 296146 115556 296156
rect 115836 300580 115892 300590
rect 115836 295428 115892 300524
rect 115836 295362 115892 295372
rect 115388 292786 115444 292796
rect 115164 282258 115220 282268
rect 113372 262918 113428 278236
rect 115164 282100 115220 282110
rect 115052 278180 115108 278190
rect 115052 277318 115108 278124
rect 115052 277252 115108 277262
rect 115164 267148 115220 282044
rect 113372 262852 113428 262862
rect 115052 267092 115220 267148
rect 112700 261592 112756 261602
rect 113736 256350 114212 256384
rect 113736 256294 113760 256350
rect 113816 256294 113884 256350
rect 113940 256294 114008 256350
rect 114064 256294 114132 256350
rect 114188 256294 114212 256350
rect 113736 256226 114212 256294
rect 113736 256170 113760 256226
rect 113816 256170 113884 256226
rect 113940 256170 114008 256226
rect 114064 256170 114132 256226
rect 114188 256170 114212 256226
rect 113736 256102 114212 256170
rect 113736 256046 113760 256102
rect 113816 256046 113884 256102
rect 113940 256046 114008 256102
rect 114064 256046 114132 256102
rect 114188 256046 114212 256102
rect 113736 255978 114212 256046
rect 113736 255922 113760 255978
rect 113816 255922 113884 255978
rect 113940 255922 114008 255978
rect 114064 255922 114132 255978
rect 114188 255922 114212 255978
rect 113736 255888 114212 255922
rect 115052 255358 115108 267092
rect 115052 255292 115108 255302
rect 112936 244350 113412 244384
rect 112936 244294 112960 244350
rect 113016 244294 113084 244350
rect 113140 244294 113208 244350
rect 113264 244294 113332 244350
rect 113388 244294 113412 244350
rect 112936 244226 113412 244294
rect 112936 244170 112960 244226
rect 113016 244170 113084 244226
rect 113140 244170 113208 244226
rect 113264 244170 113332 244226
rect 113388 244170 113412 244226
rect 112936 244102 113412 244170
rect 112936 244046 112960 244102
rect 113016 244046 113084 244102
rect 113140 244046 113208 244102
rect 113264 244046 113332 244102
rect 113388 244046 113412 244102
rect 112936 243978 113412 244046
rect 112936 243922 112960 243978
rect 113016 243922 113084 243978
rect 113140 243922 113208 243978
rect 113264 243922 113332 243978
rect 113388 243922 113412 243978
rect 112936 243888 113412 243922
rect 113736 238350 114212 238384
rect 113736 238294 113760 238350
rect 113816 238294 113884 238350
rect 113940 238294 114008 238350
rect 114064 238294 114132 238350
rect 114188 238294 114212 238350
rect 113736 238226 114212 238294
rect 113736 238170 113760 238226
rect 113816 238170 113884 238226
rect 113940 238170 114008 238226
rect 114064 238170 114132 238226
rect 114188 238170 114212 238226
rect 113736 238102 114212 238170
rect 113736 238046 113760 238102
rect 113816 238046 113884 238102
rect 113940 238046 114008 238102
rect 114064 238046 114132 238102
rect 114188 238046 114212 238102
rect 113736 237978 114212 238046
rect 113736 237922 113760 237978
rect 113816 237922 113884 237978
rect 113940 237922 114008 237978
rect 114064 237922 114132 237978
rect 114188 237922 114212 237978
rect 113736 237888 114212 237922
rect 112936 226350 113412 226384
rect 112936 226294 112960 226350
rect 113016 226294 113084 226350
rect 113140 226294 113208 226350
rect 113264 226294 113332 226350
rect 113388 226294 113412 226350
rect 112936 226226 113412 226294
rect 112936 226170 112960 226226
rect 113016 226170 113084 226226
rect 113140 226170 113208 226226
rect 113264 226170 113332 226226
rect 113388 226170 113412 226226
rect 112936 226102 113412 226170
rect 112936 226046 112960 226102
rect 113016 226046 113084 226102
rect 113140 226046 113208 226102
rect 113264 226046 113332 226102
rect 113388 226046 113412 226102
rect 112936 225978 113412 226046
rect 112936 225922 112960 225978
rect 113016 225922 113084 225978
rect 113140 225922 113208 225978
rect 113264 225922 113332 225978
rect 113388 225922 113412 225978
rect 112936 225888 113412 225922
rect 113736 220350 114212 220384
rect 113736 220294 113760 220350
rect 113816 220294 113884 220350
rect 113940 220294 114008 220350
rect 114064 220294 114132 220350
rect 114188 220294 114212 220350
rect 113736 220226 114212 220294
rect 113736 220170 113760 220226
rect 113816 220170 113884 220226
rect 113940 220170 114008 220226
rect 114064 220170 114132 220226
rect 114188 220170 114212 220226
rect 113736 220102 114212 220170
rect 113736 220046 113760 220102
rect 113816 220046 113884 220102
rect 113940 220046 114008 220102
rect 114064 220046 114132 220102
rect 114188 220046 114212 220102
rect 113736 219978 114212 220046
rect 113736 219922 113760 219978
rect 113816 219922 113884 219978
rect 113940 219922 114008 219978
rect 114064 219922 114132 219978
rect 114188 219922 114212 219978
rect 113736 219888 114212 219922
rect 112936 208350 113412 208384
rect 112936 208294 112960 208350
rect 113016 208294 113084 208350
rect 113140 208294 113208 208350
rect 113264 208294 113332 208350
rect 113388 208294 113412 208350
rect 112936 208226 113412 208294
rect 112936 208170 112960 208226
rect 113016 208170 113084 208226
rect 113140 208170 113208 208226
rect 113264 208170 113332 208226
rect 113388 208170 113412 208226
rect 112936 208102 113412 208170
rect 112936 208046 112960 208102
rect 113016 208046 113084 208102
rect 113140 208046 113208 208102
rect 113264 208046 113332 208102
rect 113388 208046 113412 208102
rect 112936 207978 113412 208046
rect 112936 207922 112960 207978
rect 113016 207922 113084 207978
rect 113140 207922 113208 207978
rect 113264 207922 113332 207978
rect 113388 207922 113412 207978
rect 112936 207888 113412 207922
rect 113736 202350 114212 202384
rect 113736 202294 113760 202350
rect 113816 202294 113884 202350
rect 113940 202294 114008 202350
rect 114064 202294 114132 202350
rect 114188 202294 114212 202350
rect 113736 202226 114212 202294
rect 113736 202170 113760 202226
rect 113816 202170 113884 202226
rect 113940 202170 114008 202226
rect 114064 202170 114132 202226
rect 114188 202170 114212 202226
rect 113736 202102 114212 202170
rect 113736 202046 113760 202102
rect 113816 202046 113884 202102
rect 113940 202046 114008 202102
rect 114064 202046 114132 202102
rect 114188 202046 114212 202102
rect 113736 201978 114212 202046
rect 113736 201922 113760 201978
rect 113816 201922 113884 201978
rect 113940 201922 114008 201978
rect 114064 201922 114132 201978
rect 114188 201922 114212 201978
rect 113736 201888 114212 201922
rect 112936 190350 113412 190384
rect 112936 190294 112960 190350
rect 113016 190294 113084 190350
rect 113140 190294 113208 190350
rect 113264 190294 113332 190350
rect 113388 190294 113412 190350
rect 112936 190226 113412 190294
rect 112936 190170 112960 190226
rect 113016 190170 113084 190226
rect 113140 190170 113208 190226
rect 113264 190170 113332 190226
rect 113388 190170 113412 190226
rect 112936 190102 113412 190170
rect 112936 190046 112960 190102
rect 113016 190046 113084 190102
rect 113140 190046 113208 190102
rect 113264 190046 113332 190102
rect 113388 190046 113412 190102
rect 112936 189978 113412 190046
rect 112936 189922 112960 189978
rect 113016 189922 113084 189978
rect 113140 189922 113208 189978
rect 113264 189922 113332 189978
rect 113388 189922 113412 189978
rect 112936 189888 113412 189922
rect 113736 184350 114212 184384
rect 113736 184294 113760 184350
rect 113816 184294 113884 184350
rect 113940 184294 114008 184350
rect 114064 184294 114132 184350
rect 114188 184294 114212 184350
rect 113736 184226 114212 184294
rect 113736 184170 113760 184226
rect 113816 184170 113884 184226
rect 113940 184170 114008 184226
rect 114064 184170 114132 184226
rect 114188 184170 114212 184226
rect 113736 184102 114212 184170
rect 113736 184046 113760 184102
rect 113816 184046 113884 184102
rect 113940 184046 114008 184102
rect 114064 184046 114132 184102
rect 114188 184046 114212 184102
rect 113736 183978 114212 184046
rect 113736 183922 113760 183978
rect 113816 183922 113884 183978
rect 113940 183922 114008 183978
rect 114064 183922 114132 183978
rect 114188 183922 114212 183978
rect 113736 183888 114212 183922
rect 112936 172350 113412 172384
rect 112936 172294 112960 172350
rect 113016 172294 113084 172350
rect 113140 172294 113208 172350
rect 113264 172294 113332 172350
rect 113388 172294 113412 172350
rect 112936 172226 113412 172294
rect 112936 172170 112960 172226
rect 113016 172170 113084 172226
rect 113140 172170 113208 172226
rect 113264 172170 113332 172226
rect 113388 172170 113412 172226
rect 112936 172102 113412 172170
rect 112936 172046 112960 172102
rect 113016 172046 113084 172102
rect 113140 172046 113208 172102
rect 113264 172046 113332 172102
rect 113388 172046 113412 172102
rect 112936 171978 113412 172046
rect 112936 171922 112960 171978
rect 113016 171922 113084 171978
rect 113140 171922 113208 171978
rect 113264 171922 113332 171978
rect 113388 171922 113412 171978
rect 112936 171888 113412 171922
rect 116732 157444 116788 340172
rect 117068 340228 117124 340238
rect 116732 157378 116788 157388
rect 116844 338660 116900 338670
rect 116844 155652 116900 338604
rect 116956 336084 117012 336094
rect 116956 314020 117012 336028
rect 116956 313954 117012 313964
rect 116844 155586 116900 155596
rect 116956 310772 117012 310782
rect 116956 152180 117012 310716
rect 117068 274596 117124 340172
rect 117180 337316 117236 352492
rect 117180 337250 117236 337260
rect 117404 331138 117460 355852
rect 117516 332668 117572 362222
rect 118636 339332 118692 339342
rect 117516 332612 118468 332668
rect 117516 331858 117572 332612
rect 117516 331792 117572 331802
rect 117404 331082 117684 331138
rect 117404 321076 117460 321086
rect 117292 320404 117348 320414
rect 117180 318388 117236 318398
rect 117180 315588 117236 318332
rect 117180 315522 117236 315532
rect 117180 315028 117236 315038
rect 117180 292068 117236 314972
rect 117292 314468 117348 320348
rect 117292 314402 117348 314412
rect 117404 314188 117460 321020
rect 117292 314132 117460 314188
rect 117292 306628 117348 314132
rect 117292 306562 117348 306572
rect 117404 312598 117460 312608
rect 117404 298788 117460 312542
rect 117404 298722 117460 298732
rect 117628 298228 117684 331082
rect 118412 319078 118468 332612
rect 118412 319012 118468 319022
rect 118524 308420 118580 308430
rect 117628 298162 117684 298172
rect 118412 305060 118468 305070
rect 117180 292002 117236 292012
rect 117068 274530 117124 274540
rect 118412 153748 118468 305004
rect 118524 157556 118580 308364
rect 118636 278578 118692 339276
rect 119196 337540 119252 364922
rect 119196 336980 119252 337484
rect 119196 336914 119252 336924
rect 118636 278512 118692 278522
rect 118748 334852 118804 334862
rect 118748 277138 118804 334796
rect 119196 331716 119252 331726
rect 118860 329140 118916 329150
rect 118860 303268 118916 329084
rect 118860 303202 118916 303212
rect 118748 277072 118804 277082
rect 118860 281428 118916 281438
rect 118860 270118 118916 281372
rect 119196 276598 119252 331660
rect 119868 331604 119924 331614
rect 119644 330036 119700 330046
rect 119308 283978 119364 283988
rect 119308 280084 119364 283922
rect 119308 280018 119364 280028
rect 119644 276778 119700 329980
rect 119868 276958 119924 331548
rect 119980 286498 120036 286508
rect 119980 277172 120036 286442
rect 119980 277106 120036 277116
rect 119868 276892 119924 276902
rect 119644 276712 119700 276722
rect 119196 276532 119252 276542
rect 118860 270052 118916 270062
rect 119196 274820 119252 274830
rect 118524 157490 118580 157500
rect 118636 181558 118692 181568
rect 118412 153682 118468 153692
rect 116956 152114 117012 152124
rect 112476 149452 112532 149462
rect 112364 148530 112420 148540
rect 118636 147924 118692 181502
rect 118748 149518 118804 149528
rect 118748 148148 118804 149462
rect 118748 148082 118804 148092
rect 119196 148036 119252 274764
rect 120092 271558 120148 590716
rect 128298 580350 128918 596784
rect 128298 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 128918 580350
rect 128298 580226 128918 580294
rect 128298 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 128918 580226
rect 128298 580102 128918 580170
rect 128298 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 128918 580102
rect 128298 579978 128918 580046
rect 128298 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 128918 579978
rect 120204 573076 120260 573086
rect 120204 278218 120260 573020
rect 128298 562350 128918 579922
rect 128298 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 128918 562350
rect 128298 562226 128918 562294
rect 128298 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 128918 562226
rect 128298 562102 128918 562170
rect 128298 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 128918 562102
rect 128298 561978 128918 562046
rect 128298 561922 128394 561978
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 128918 561978
rect 128298 544350 128918 561922
rect 128298 544294 128394 544350
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 128918 544350
rect 128298 544226 128918 544294
rect 128298 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 128918 544226
rect 128298 544102 128918 544170
rect 128298 544046 128394 544102
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 128918 544102
rect 128298 543978 128918 544046
rect 128298 543922 128394 543978
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 128918 543978
rect 128298 526350 128918 543922
rect 128298 526294 128394 526350
rect 128450 526294 128518 526350
rect 128574 526294 128642 526350
rect 128698 526294 128766 526350
rect 128822 526294 128918 526350
rect 128298 526226 128918 526294
rect 128298 526170 128394 526226
rect 128450 526170 128518 526226
rect 128574 526170 128642 526226
rect 128698 526170 128766 526226
rect 128822 526170 128918 526226
rect 128298 526102 128918 526170
rect 128298 526046 128394 526102
rect 128450 526046 128518 526102
rect 128574 526046 128642 526102
rect 128698 526046 128766 526102
rect 128822 526046 128918 526102
rect 128298 525978 128918 526046
rect 128298 525922 128394 525978
rect 128450 525922 128518 525978
rect 128574 525922 128642 525978
rect 128698 525922 128766 525978
rect 128822 525922 128918 525978
rect 128298 508350 128918 525922
rect 128298 508294 128394 508350
rect 128450 508294 128518 508350
rect 128574 508294 128642 508350
rect 128698 508294 128766 508350
rect 128822 508294 128918 508350
rect 128298 508226 128918 508294
rect 128298 508170 128394 508226
rect 128450 508170 128518 508226
rect 128574 508170 128642 508226
rect 128698 508170 128766 508226
rect 128822 508170 128918 508226
rect 128298 508102 128918 508170
rect 128298 508046 128394 508102
rect 128450 508046 128518 508102
rect 128574 508046 128642 508102
rect 128698 508046 128766 508102
rect 128822 508046 128918 508102
rect 128298 507978 128918 508046
rect 128298 507922 128394 507978
rect 128450 507922 128518 507978
rect 128574 507922 128642 507978
rect 128698 507922 128766 507978
rect 128822 507922 128918 507978
rect 128298 490350 128918 507922
rect 128298 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 128918 490350
rect 128298 490226 128918 490294
rect 128298 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 128918 490226
rect 128298 490102 128918 490170
rect 128298 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 128918 490102
rect 128298 489978 128918 490046
rect 128298 489922 128394 489978
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 128918 489978
rect 128298 472350 128918 489922
rect 128298 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 128918 472350
rect 128298 472226 128918 472294
rect 128298 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 128918 472226
rect 128298 472102 128918 472170
rect 128298 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 128918 472102
rect 128298 471978 128918 472046
rect 128298 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 128918 471978
rect 128298 454350 128918 471922
rect 128298 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 128918 454350
rect 128298 454226 128918 454294
rect 128298 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 128918 454226
rect 128298 454102 128918 454170
rect 128298 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 128918 454102
rect 128298 453978 128918 454046
rect 128298 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 128918 453978
rect 128298 436350 128918 453922
rect 128298 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 128918 436350
rect 128298 436226 128918 436294
rect 128298 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 128918 436226
rect 128298 436102 128918 436170
rect 128298 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 128918 436102
rect 128298 435978 128918 436046
rect 128298 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 128918 435978
rect 128298 418350 128918 435922
rect 128298 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 128918 418350
rect 128298 418226 128918 418294
rect 128298 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 128918 418226
rect 128298 418102 128918 418170
rect 128298 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 128918 418102
rect 128298 417978 128918 418046
rect 128298 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 128918 417978
rect 128298 400350 128918 417922
rect 128298 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 128918 400350
rect 128298 400226 128918 400294
rect 128298 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 128918 400226
rect 128298 400102 128918 400170
rect 128298 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 128918 400102
rect 128298 399978 128918 400046
rect 128298 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 128918 399978
rect 128298 382350 128918 399922
rect 128298 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 128918 382350
rect 128298 382226 128918 382294
rect 128298 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 128918 382226
rect 128298 382102 128918 382170
rect 128298 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 128918 382102
rect 128298 381978 128918 382046
rect 128298 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 128918 381978
rect 128298 364350 128918 381922
rect 128298 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 128918 364350
rect 128298 364226 128918 364294
rect 128298 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 128918 364226
rect 128298 364102 128918 364170
rect 128298 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 128918 364102
rect 128298 363978 128918 364046
rect 128298 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 128918 363978
rect 128298 358958 128918 363922
rect 132018 598172 132638 598268
rect 132018 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 132638 598172
rect 132018 598048 132638 598116
rect 132018 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 132638 598048
rect 132018 597924 132638 597992
rect 132018 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 132638 597924
rect 132018 597800 132638 597868
rect 132018 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 132638 597800
rect 132018 586350 132638 597744
rect 132018 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 132638 586350
rect 132018 586226 132638 586294
rect 132018 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 132638 586226
rect 132018 586102 132638 586170
rect 132018 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 132638 586102
rect 132018 585978 132638 586046
rect 132018 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 132638 585978
rect 132018 568350 132638 585922
rect 132018 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 132638 568350
rect 132018 568226 132638 568294
rect 132018 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 132638 568226
rect 132018 568102 132638 568170
rect 132018 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 132638 568102
rect 132018 567978 132638 568046
rect 132018 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 132638 567978
rect 132018 550350 132638 567922
rect 132018 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 132638 550350
rect 132018 550226 132638 550294
rect 132018 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 132638 550226
rect 132018 550102 132638 550170
rect 132018 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 132638 550102
rect 132018 549978 132638 550046
rect 132018 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 132638 549978
rect 132018 532350 132638 549922
rect 132018 532294 132114 532350
rect 132170 532294 132238 532350
rect 132294 532294 132362 532350
rect 132418 532294 132486 532350
rect 132542 532294 132638 532350
rect 132018 532226 132638 532294
rect 132018 532170 132114 532226
rect 132170 532170 132238 532226
rect 132294 532170 132362 532226
rect 132418 532170 132486 532226
rect 132542 532170 132638 532226
rect 132018 532102 132638 532170
rect 132018 532046 132114 532102
rect 132170 532046 132238 532102
rect 132294 532046 132362 532102
rect 132418 532046 132486 532102
rect 132542 532046 132638 532102
rect 132018 531978 132638 532046
rect 132018 531922 132114 531978
rect 132170 531922 132238 531978
rect 132294 531922 132362 531978
rect 132418 531922 132486 531978
rect 132542 531922 132638 531978
rect 132018 514350 132638 531922
rect 132018 514294 132114 514350
rect 132170 514294 132238 514350
rect 132294 514294 132362 514350
rect 132418 514294 132486 514350
rect 132542 514294 132638 514350
rect 132018 514226 132638 514294
rect 132018 514170 132114 514226
rect 132170 514170 132238 514226
rect 132294 514170 132362 514226
rect 132418 514170 132486 514226
rect 132542 514170 132638 514226
rect 132018 514102 132638 514170
rect 132018 514046 132114 514102
rect 132170 514046 132238 514102
rect 132294 514046 132362 514102
rect 132418 514046 132486 514102
rect 132542 514046 132638 514102
rect 132018 513978 132638 514046
rect 132018 513922 132114 513978
rect 132170 513922 132238 513978
rect 132294 513922 132362 513978
rect 132418 513922 132486 513978
rect 132542 513922 132638 513978
rect 132018 496350 132638 513922
rect 132018 496294 132114 496350
rect 132170 496294 132238 496350
rect 132294 496294 132362 496350
rect 132418 496294 132486 496350
rect 132542 496294 132638 496350
rect 132018 496226 132638 496294
rect 132018 496170 132114 496226
rect 132170 496170 132238 496226
rect 132294 496170 132362 496226
rect 132418 496170 132486 496226
rect 132542 496170 132638 496226
rect 132018 496102 132638 496170
rect 132018 496046 132114 496102
rect 132170 496046 132238 496102
rect 132294 496046 132362 496102
rect 132418 496046 132486 496102
rect 132542 496046 132638 496102
rect 132018 495978 132638 496046
rect 132018 495922 132114 495978
rect 132170 495922 132238 495978
rect 132294 495922 132362 495978
rect 132418 495922 132486 495978
rect 132542 495922 132638 495978
rect 132018 478350 132638 495922
rect 132018 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 132638 478350
rect 132018 478226 132638 478294
rect 132018 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 132638 478226
rect 132018 478102 132638 478170
rect 132018 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 132638 478102
rect 132018 477978 132638 478046
rect 132018 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 132638 477978
rect 132018 460350 132638 477922
rect 132018 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 132638 460350
rect 132018 460226 132638 460294
rect 132018 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 132638 460226
rect 132018 460102 132638 460170
rect 132018 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 132638 460102
rect 132018 459978 132638 460046
rect 132018 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 132638 459978
rect 132018 442350 132638 459922
rect 132018 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 132638 442350
rect 132018 442226 132638 442294
rect 132018 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 132638 442226
rect 132018 442102 132638 442170
rect 132018 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 132638 442102
rect 132018 441978 132638 442046
rect 132018 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 132638 441978
rect 132018 424350 132638 441922
rect 132018 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 132638 424350
rect 132018 424226 132638 424294
rect 132018 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 132638 424226
rect 132018 424102 132638 424170
rect 132018 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 132638 424102
rect 132018 423978 132638 424046
rect 132018 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 132638 423978
rect 132018 406350 132638 423922
rect 132018 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 132638 406350
rect 132018 406226 132638 406294
rect 132018 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 132638 406226
rect 132018 406102 132638 406170
rect 132018 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 132638 406102
rect 132018 405978 132638 406046
rect 132018 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 132638 405978
rect 132018 388350 132638 405922
rect 132018 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 132638 388350
rect 132018 388226 132638 388294
rect 132018 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 132638 388226
rect 132018 388102 132638 388170
rect 132018 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 132638 388102
rect 132018 387978 132638 388046
rect 132018 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 132638 387978
rect 132018 370350 132638 387922
rect 132018 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 132638 370350
rect 132018 370226 132638 370294
rect 132018 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 132638 370226
rect 132018 370102 132638 370170
rect 132018 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 132638 370102
rect 132018 369978 132638 370046
rect 132018 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 132638 369978
rect 132018 358958 132638 369922
rect 159018 597212 159638 598268
rect 159018 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 159638 597212
rect 159018 597088 159638 597156
rect 159018 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 159638 597088
rect 159018 596964 159638 597032
rect 159018 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 159638 596964
rect 159018 596840 159638 596908
rect 159018 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 159638 596840
rect 159018 580350 159638 596784
rect 159018 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 159638 580350
rect 159018 580226 159638 580294
rect 159018 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 159638 580226
rect 159018 580102 159638 580170
rect 159018 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 159638 580102
rect 159018 579978 159638 580046
rect 159018 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 159638 579978
rect 159018 562350 159638 579922
rect 159018 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 159638 562350
rect 159018 562226 159638 562294
rect 159018 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 159638 562226
rect 159018 562102 159638 562170
rect 159018 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 159638 562102
rect 159018 561978 159638 562046
rect 159018 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 159638 561978
rect 159018 544350 159638 561922
rect 159018 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 159638 544350
rect 159018 544226 159638 544294
rect 159018 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 159638 544226
rect 159018 544102 159638 544170
rect 159018 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 159638 544102
rect 159018 543978 159638 544046
rect 159018 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 159638 543978
rect 159018 526350 159638 543922
rect 159018 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 159638 526350
rect 159018 526226 159638 526294
rect 159018 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 159638 526226
rect 159018 526102 159638 526170
rect 159018 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 159638 526102
rect 159018 525978 159638 526046
rect 159018 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 159638 525978
rect 159018 508350 159638 525922
rect 159018 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 159638 508350
rect 159018 508226 159638 508294
rect 159018 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 159638 508226
rect 159018 508102 159638 508170
rect 159018 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 159638 508102
rect 159018 507978 159638 508046
rect 159018 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 159638 507978
rect 159018 490350 159638 507922
rect 159018 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 159638 490350
rect 159018 490226 159638 490294
rect 159018 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 159638 490226
rect 159018 490102 159638 490170
rect 159018 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 159638 490102
rect 159018 489978 159638 490046
rect 159018 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 159638 489978
rect 159018 472350 159638 489922
rect 159018 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 159638 472350
rect 159018 472226 159638 472294
rect 159018 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 159638 472226
rect 159018 472102 159638 472170
rect 159018 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 159638 472102
rect 159018 471978 159638 472046
rect 159018 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 159638 471978
rect 159018 454350 159638 471922
rect 159018 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 159638 454350
rect 159018 454226 159638 454294
rect 159018 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 159638 454226
rect 159018 454102 159638 454170
rect 159018 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 159638 454102
rect 159018 453978 159638 454046
rect 159018 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 159638 453978
rect 159018 436350 159638 453922
rect 159018 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 159638 436350
rect 159018 436226 159638 436294
rect 159018 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 159638 436226
rect 159018 436102 159638 436170
rect 159018 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 159638 436102
rect 159018 435978 159638 436046
rect 159018 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 159638 435978
rect 159018 418350 159638 435922
rect 159018 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 159638 418350
rect 159018 418226 159638 418294
rect 159018 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 159638 418226
rect 159018 418102 159638 418170
rect 159018 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 159638 418102
rect 159018 417978 159638 418046
rect 159018 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 159638 417978
rect 159018 400350 159638 417922
rect 159018 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 159638 400350
rect 159018 400226 159638 400294
rect 159018 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 159638 400226
rect 159018 400102 159638 400170
rect 159018 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 159638 400102
rect 159018 399978 159638 400046
rect 159018 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 159638 399978
rect 159018 382350 159638 399922
rect 159018 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 159638 382350
rect 159018 382226 159638 382294
rect 159018 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 159638 382226
rect 159018 382102 159638 382170
rect 159018 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 159638 382102
rect 159018 381978 159638 382046
rect 159018 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 159638 381978
rect 156156 364798 156212 364808
rect 151340 363178 151396 363188
rect 151340 362964 151396 363122
rect 151340 362898 151396 362908
rect 152012 362998 152068 363008
rect 152012 362898 152068 362908
rect 156156 362964 156212 364742
rect 156156 362898 156212 362908
rect 157836 364618 157892 364628
rect 157836 362964 157892 364562
rect 157836 362898 157892 362908
rect 159018 364350 159638 381922
rect 162738 598172 163358 598268
rect 162738 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 163358 598172
rect 162738 598048 163358 598116
rect 162738 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 163358 598048
rect 162738 597924 163358 597992
rect 162738 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 163358 597924
rect 162738 597800 163358 597868
rect 162738 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 163358 597800
rect 162738 586350 163358 597744
rect 162738 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 163358 586350
rect 162738 586226 163358 586294
rect 162738 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 163358 586226
rect 162738 586102 163358 586170
rect 162738 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 163358 586102
rect 162738 585978 163358 586046
rect 162738 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 163358 585978
rect 162738 568350 163358 585922
rect 162738 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 163358 568350
rect 162738 568226 163358 568294
rect 162738 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 163358 568226
rect 162738 568102 163358 568170
rect 162738 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 163358 568102
rect 162738 567978 163358 568046
rect 162738 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 163358 567978
rect 162738 550350 163358 567922
rect 162738 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 163358 550350
rect 162738 550226 163358 550294
rect 162738 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 163358 550226
rect 162738 550102 163358 550170
rect 162738 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 163358 550102
rect 162738 549978 163358 550046
rect 162738 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 163358 549978
rect 162738 532350 163358 549922
rect 162738 532294 162834 532350
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 163358 532350
rect 162738 532226 163358 532294
rect 162738 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 163358 532226
rect 162738 532102 163358 532170
rect 162738 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 163358 532102
rect 162738 531978 163358 532046
rect 162738 531922 162834 531978
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 163358 531978
rect 162738 514350 163358 531922
rect 162738 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 163358 514350
rect 162738 514226 163358 514294
rect 162738 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 163358 514226
rect 162738 514102 163358 514170
rect 162738 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 163358 514102
rect 162738 513978 163358 514046
rect 162738 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 163358 513978
rect 162738 496350 163358 513922
rect 162738 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 163358 496350
rect 162738 496226 163358 496294
rect 162738 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 163358 496226
rect 162738 496102 163358 496170
rect 162738 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 163358 496102
rect 162738 495978 163358 496046
rect 162738 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 163358 495978
rect 162738 478350 163358 495922
rect 162738 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 163358 478350
rect 162738 478226 163358 478294
rect 162738 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 163358 478226
rect 162738 478102 163358 478170
rect 162738 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 163358 478102
rect 162738 477978 163358 478046
rect 162738 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 163358 477978
rect 162738 460350 163358 477922
rect 162738 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 163358 460350
rect 162738 460226 163358 460294
rect 162738 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 163358 460226
rect 162738 460102 163358 460170
rect 162738 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 163358 460102
rect 162738 459978 163358 460046
rect 162738 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 163358 459978
rect 162738 442350 163358 459922
rect 162738 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 163358 442350
rect 162738 442226 163358 442294
rect 162738 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 163358 442226
rect 162738 442102 163358 442170
rect 162738 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 163358 442102
rect 162738 441978 163358 442046
rect 162738 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 163358 441978
rect 162738 424350 163358 441922
rect 162738 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 163358 424350
rect 162738 424226 163358 424294
rect 162738 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 163358 424226
rect 162738 424102 163358 424170
rect 162738 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 163358 424102
rect 162738 423978 163358 424046
rect 162738 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 163358 423978
rect 162738 406350 163358 423922
rect 162738 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 163358 406350
rect 162738 406226 163358 406294
rect 162738 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 163358 406226
rect 162738 406102 163358 406170
rect 162738 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 163358 406102
rect 162738 405978 163358 406046
rect 162738 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 163358 405978
rect 162738 388350 163358 405922
rect 162738 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 163358 388350
rect 162738 388226 163358 388294
rect 162738 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 163358 388226
rect 162738 388102 163358 388170
rect 162738 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 163358 388102
rect 162738 387978 163358 388046
rect 162738 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 163358 387978
rect 162738 370350 163358 387922
rect 162738 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 163358 370350
rect 162738 370226 163358 370294
rect 162738 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 163358 370226
rect 162738 370102 163358 370170
rect 162738 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 163358 370102
rect 162738 369978 163358 370046
rect 162738 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 163358 369978
rect 159018 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 159638 364350
rect 159018 364226 159638 364294
rect 159018 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 159638 364226
rect 159018 364102 159638 364170
rect 159018 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 159638 364102
rect 159018 363978 159638 364046
rect 159018 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 159638 363978
rect 150668 362098 150724 362108
rect 150668 361620 150724 362042
rect 150668 361554 150724 361564
rect 155372 361956 155428 361966
rect 155372 361620 155428 361900
rect 155372 361554 155428 361564
rect 159018 358958 159638 363922
rect 160748 365158 160804 365168
rect 160748 363076 160804 365102
rect 160748 363010 160804 363020
rect 161420 361558 161476 361568
rect 161420 361172 161476 361502
rect 161420 361106 161476 361116
rect 162738 358958 163358 369922
rect 189738 597212 190358 598268
rect 189738 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 190358 597212
rect 189738 597088 190358 597156
rect 189738 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 190358 597088
rect 189738 596964 190358 597032
rect 189738 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 190358 596964
rect 189738 596840 190358 596908
rect 189738 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 190358 596840
rect 189738 580350 190358 596784
rect 189738 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 190358 580350
rect 189738 580226 190358 580294
rect 189738 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 190358 580226
rect 189738 580102 190358 580170
rect 189738 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 190358 580102
rect 189738 579978 190358 580046
rect 189738 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 190358 579978
rect 189738 562350 190358 579922
rect 189738 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 190358 562350
rect 189738 562226 190358 562294
rect 189738 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 190358 562226
rect 189738 562102 190358 562170
rect 189738 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 190358 562102
rect 189738 561978 190358 562046
rect 189738 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 190358 561978
rect 189738 544350 190358 561922
rect 189738 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 190358 544350
rect 189738 544226 190358 544294
rect 189738 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 190358 544226
rect 189738 544102 190358 544170
rect 189738 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 190358 544102
rect 189738 543978 190358 544046
rect 189738 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 190358 543978
rect 189738 526350 190358 543922
rect 189738 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 190358 526350
rect 189738 526226 190358 526294
rect 189738 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 190358 526226
rect 189738 526102 190358 526170
rect 189738 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 190358 526102
rect 189738 525978 190358 526046
rect 189738 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 190358 525978
rect 189738 508350 190358 525922
rect 189738 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 190358 508350
rect 189738 508226 190358 508294
rect 189738 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 190358 508226
rect 189738 508102 190358 508170
rect 189738 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 190358 508102
rect 189738 507978 190358 508046
rect 189738 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 190358 507978
rect 189738 490350 190358 507922
rect 189738 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 190358 490350
rect 189738 490226 190358 490294
rect 189738 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 190358 490226
rect 189738 490102 190358 490170
rect 189738 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 190358 490102
rect 189738 489978 190358 490046
rect 189738 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 190358 489978
rect 189738 472350 190358 489922
rect 189738 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 190358 472350
rect 189738 472226 190358 472294
rect 189738 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 190358 472226
rect 189738 472102 190358 472170
rect 189738 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 190358 472102
rect 189738 471978 190358 472046
rect 189738 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 190358 471978
rect 189738 454350 190358 471922
rect 189738 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 190358 454350
rect 189738 454226 190358 454294
rect 189738 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 190358 454226
rect 189738 454102 190358 454170
rect 189738 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 190358 454102
rect 189738 453978 190358 454046
rect 189738 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 190358 453978
rect 189738 436350 190358 453922
rect 189738 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 190358 436350
rect 189738 436226 190358 436294
rect 189738 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 190358 436226
rect 189738 436102 190358 436170
rect 189738 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 190358 436102
rect 189738 435978 190358 436046
rect 189738 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 190358 435978
rect 189738 418350 190358 435922
rect 189738 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 190358 418350
rect 189738 418226 190358 418294
rect 189738 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 190358 418226
rect 189738 418102 190358 418170
rect 189738 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 190358 418102
rect 189738 417978 190358 418046
rect 189738 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 190358 417978
rect 189738 400350 190358 417922
rect 189738 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 190358 400350
rect 189738 400226 190358 400294
rect 189738 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 190358 400226
rect 189738 400102 190358 400170
rect 189738 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 190358 400102
rect 189738 399978 190358 400046
rect 189738 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 190358 399978
rect 189738 382350 190358 399922
rect 189738 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 190358 382350
rect 189738 382226 190358 382294
rect 189738 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 190358 382226
rect 189738 382102 190358 382170
rect 189738 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 190358 382102
rect 189738 381978 190358 382046
rect 189738 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 190358 381978
rect 171276 366778 171332 366788
rect 164668 364978 164724 364988
rect 164668 363076 164724 364922
rect 171276 363748 171332 366722
rect 171276 363682 171332 363692
rect 189738 364350 190358 381922
rect 189738 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 190358 364350
rect 189738 364226 190358 364294
rect 189738 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 190358 364226
rect 189738 364102 190358 364170
rect 189738 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 190358 364102
rect 189738 363978 190358 364046
rect 189738 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 190358 363978
rect 164668 363010 164724 363020
rect 163436 362278 163492 362288
rect 163436 362180 163492 362222
rect 163436 362114 163492 362124
rect 173516 360298 173572 360308
rect 166124 359604 166180 359614
rect 166124 358678 166180 359548
rect 173516 359604 173572 360242
rect 173516 359538 173572 359548
rect 182252 359492 182308 359502
rect 182252 359038 182308 359436
rect 182252 358972 182308 358982
rect 186956 359492 187012 359502
rect 166124 358612 166180 358622
rect 186956 357058 187012 359436
rect 189532 359492 189588 359502
rect 189532 358858 189588 359436
rect 189738 358958 190358 363922
rect 193458 598172 194078 598268
rect 193458 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 194078 598172
rect 193458 598048 194078 598116
rect 193458 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 194078 598048
rect 193458 597924 194078 597992
rect 193458 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 194078 597924
rect 193458 597800 194078 597868
rect 193458 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 194078 597800
rect 193458 586350 194078 597744
rect 220458 597212 221078 598268
rect 220458 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 221078 597212
rect 220458 597088 221078 597156
rect 220458 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 221078 597088
rect 220458 596964 221078 597032
rect 220458 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 221078 596964
rect 220458 596840 221078 596908
rect 220458 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 221078 596840
rect 199948 590772 200004 590782
rect 193458 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 194078 586350
rect 193458 586226 194078 586294
rect 193458 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 194078 586226
rect 193458 586102 194078 586170
rect 193458 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 194078 586102
rect 193458 585978 194078 586046
rect 193458 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 194078 585978
rect 193458 568350 194078 585922
rect 193458 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 194078 568350
rect 193458 568226 194078 568294
rect 193458 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 194078 568226
rect 193458 568102 194078 568170
rect 193458 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 194078 568102
rect 193458 567978 194078 568046
rect 193458 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 194078 567978
rect 193458 550350 194078 567922
rect 193458 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 194078 550350
rect 193458 550226 194078 550294
rect 193458 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 194078 550226
rect 193458 550102 194078 550170
rect 193458 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 194078 550102
rect 193458 549978 194078 550046
rect 193458 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 194078 549978
rect 193458 532350 194078 549922
rect 193458 532294 193554 532350
rect 193610 532294 193678 532350
rect 193734 532294 193802 532350
rect 193858 532294 193926 532350
rect 193982 532294 194078 532350
rect 193458 532226 194078 532294
rect 193458 532170 193554 532226
rect 193610 532170 193678 532226
rect 193734 532170 193802 532226
rect 193858 532170 193926 532226
rect 193982 532170 194078 532226
rect 193458 532102 194078 532170
rect 193458 532046 193554 532102
rect 193610 532046 193678 532102
rect 193734 532046 193802 532102
rect 193858 532046 193926 532102
rect 193982 532046 194078 532102
rect 193458 531978 194078 532046
rect 193458 531922 193554 531978
rect 193610 531922 193678 531978
rect 193734 531922 193802 531978
rect 193858 531922 193926 531978
rect 193982 531922 194078 531978
rect 193458 514350 194078 531922
rect 193458 514294 193554 514350
rect 193610 514294 193678 514350
rect 193734 514294 193802 514350
rect 193858 514294 193926 514350
rect 193982 514294 194078 514350
rect 193458 514226 194078 514294
rect 193458 514170 193554 514226
rect 193610 514170 193678 514226
rect 193734 514170 193802 514226
rect 193858 514170 193926 514226
rect 193982 514170 194078 514226
rect 193458 514102 194078 514170
rect 193458 514046 193554 514102
rect 193610 514046 193678 514102
rect 193734 514046 193802 514102
rect 193858 514046 193926 514102
rect 193982 514046 194078 514102
rect 193458 513978 194078 514046
rect 193458 513922 193554 513978
rect 193610 513922 193678 513978
rect 193734 513922 193802 513978
rect 193858 513922 193926 513978
rect 193982 513922 194078 513978
rect 193458 496350 194078 513922
rect 193458 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 194078 496350
rect 193458 496226 194078 496294
rect 193458 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 194078 496226
rect 193458 496102 194078 496170
rect 193458 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 194078 496102
rect 193458 495978 194078 496046
rect 193458 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 194078 495978
rect 193458 478350 194078 495922
rect 193458 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 194078 478350
rect 193458 478226 194078 478294
rect 193458 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 194078 478226
rect 193458 478102 194078 478170
rect 193458 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 194078 478102
rect 193458 477978 194078 478046
rect 193458 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 194078 477978
rect 193458 460350 194078 477922
rect 193458 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 194078 460350
rect 193458 460226 194078 460294
rect 193458 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 194078 460226
rect 193458 460102 194078 460170
rect 193458 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 194078 460102
rect 193458 459978 194078 460046
rect 193458 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 194078 459978
rect 193458 442350 194078 459922
rect 193458 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 194078 442350
rect 193458 442226 194078 442294
rect 193458 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 194078 442226
rect 193458 442102 194078 442170
rect 193458 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 194078 442102
rect 193458 441978 194078 442046
rect 193458 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 194078 441978
rect 193458 424350 194078 441922
rect 193458 424294 193554 424350
rect 193610 424294 193678 424350
rect 193734 424294 193802 424350
rect 193858 424294 193926 424350
rect 193982 424294 194078 424350
rect 193458 424226 194078 424294
rect 193458 424170 193554 424226
rect 193610 424170 193678 424226
rect 193734 424170 193802 424226
rect 193858 424170 193926 424226
rect 193982 424170 194078 424226
rect 193458 424102 194078 424170
rect 193458 424046 193554 424102
rect 193610 424046 193678 424102
rect 193734 424046 193802 424102
rect 193858 424046 193926 424102
rect 193982 424046 194078 424102
rect 193458 423978 194078 424046
rect 193458 423922 193554 423978
rect 193610 423922 193678 423978
rect 193734 423922 193802 423978
rect 193858 423922 193926 423978
rect 193982 423922 194078 423978
rect 193458 406350 194078 423922
rect 193458 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 194078 406350
rect 193458 406226 194078 406294
rect 193458 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 194078 406226
rect 193458 406102 194078 406170
rect 193458 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 194078 406102
rect 193458 405978 194078 406046
rect 193458 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 194078 405978
rect 193458 388350 194078 405922
rect 193458 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 194078 388350
rect 193458 388226 194078 388294
rect 193458 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 194078 388226
rect 193458 388102 194078 388170
rect 193458 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 194078 388102
rect 193458 387978 194078 388046
rect 193458 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 194078 387978
rect 193458 370350 194078 387922
rect 199836 587188 199892 587198
rect 193458 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 194078 370350
rect 193458 370226 194078 370294
rect 197708 371812 197764 371822
rect 193458 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 194078 370226
rect 193458 370102 194078 370170
rect 196588 370244 196644 370254
rect 193458 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 194078 370102
rect 193458 369978 194078 370046
rect 193458 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 194078 369978
rect 193340 362180 193396 362190
rect 190988 359758 191044 359768
rect 190764 359604 190820 359614
rect 190988 359604 191044 359702
rect 190988 359538 191044 359548
rect 192556 359604 192612 359614
rect 192612 359548 192948 359578
rect 192556 359522 192948 359548
rect 190764 359510 190820 359522
rect 189532 358792 189588 358802
rect 186956 356992 187012 357002
rect 149152 352350 149472 352384
rect 149152 352294 149222 352350
rect 149278 352294 149346 352350
rect 149402 352294 149472 352350
rect 149152 352226 149472 352294
rect 149152 352170 149222 352226
rect 149278 352170 149346 352226
rect 149402 352170 149472 352226
rect 149152 352102 149472 352170
rect 149152 352046 149222 352102
rect 149278 352046 149346 352102
rect 149402 352046 149472 352102
rect 149152 351978 149472 352046
rect 149152 351922 149222 351978
rect 149278 351922 149346 351978
rect 149402 351922 149472 351978
rect 149152 351888 149472 351922
rect 179872 352350 180192 352384
rect 179872 352294 179942 352350
rect 179998 352294 180066 352350
rect 180122 352294 180192 352350
rect 179872 352226 180192 352294
rect 179872 352170 179942 352226
rect 179998 352170 180066 352226
rect 180122 352170 180192 352226
rect 179872 352102 180192 352170
rect 179872 352046 179942 352102
rect 179998 352046 180066 352102
rect 180122 352046 180192 352102
rect 179872 351978 180192 352046
rect 179872 351922 179942 351978
rect 179998 351922 180066 351978
rect 180122 351922 180192 351978
rect 179872 351888 180192 351922
rect 133792 346350 134112 346384
rect 133792 346294 133862 346350
rect 133918 346294 133986 346350
rect 134042 346294 134112 346350
rect 133792 346226 134112 346294
rect 133792 346170 133862 346226
rect 133918 346170 133986 346226
rect 134042 346170 134112 346226
rect 133792 346102 134112 346170
rect 133792 346046 133862 346102
rect 133918 346046 133986 346102
rect 134042 346046 134112 346102
rect 133792 345978 134112 346046
rect 133792 345922 133862 345978
rect 133918 345922 133986 345978
rect 134042 345922 134112 345978
rect 133792 345888 134112 345922
rect 164512 346350 164832 346384
rect 164512 346294 164582 346350
rect 164638 346294 164706 346350
rect 164762 346294 164832 346350
rect 164512 346226 164832 346294
rect 164512 346170 164582 346226
rect 164638 346170 164706 346226
rect 164762 346170 164832 346226
rect 164512 346102 164832 346170
rect 164512 346046 164582 346102
rect 164638 346046 164706 346102
rect 164762 346046 164832 346102
rect 164512 345978 164832 346046
rect 164512 345922 164582 345978
rect 164638 345922 164706 345978
rect 164762 345922 164832 345978
rect 164512 345888 164832 345922
rect 120540 334516 120596 334526
rect 120204 278152 120260 278162
rect 120316 329364 120372 329374
rect 120092 271492 120148 271502
rect 120092 205858 120148 205868
rect 120092 165620 120148 205802
rect 120092 165554 120148 165564
rect 119196 147970 119252 147980
rect 118636 147858 118692 147868
rect 120316 147028 120372 329308
rect 120428 314020 120484 314030
rect 120428 153860 120484 313964
rect 120540 276418 120596 334460
rect 149152 334350 149472 334384
rect 149152 334294 149222 334350
rect 149278 334294 149346 334350
rect 149402 334294 149472 334350
rect 149152 334226 149472 334294
rect 149152 334170 149222 334226
rect 149278 334170 149346 334226
rect 149402 334170 149472 334226
rect 149152 334102 149472 334170
rect 149152 334046 149222 334102
rect 149278 334046 149346 334102
rect 149402 334046 149472 334102
rect 149152 333978 149472 334046
rect 149152 333922 149222 333978
rect 149278 333922 149346 333978
rect 149402 333922 149472 333978
rect 149152 333888 149472 333922
rect 179872 334350 180192 334384
rect 179872 334294 179942 334350
rect 179998 334294 180066 334350
rect 180122 334294 180192 334350
rect 179872 334226 180192 334294
rect 179872 334170 179942 334226
rect 179998 334170 180066 334226
rect 180122 334170 180192 334226
rect 179872 334102 180192 334170
rect 179872 334046 179942 334102
rect 179998 334046 180066 334102
rect 180122 334046 180192 334102
rect 179872 333978 180192 334046
rect 179872 333922 179942 333978
rect 179998 333922 180066 333978
rect 180122 333922 180192 333978
rect 179872 333888 180192 333922
rect 133792 328350 134112 328384
rect 133792 328294 133862 328350
rect 133918 328294 133986 328350
rect 134042 328294 134112 328350
rect 133792 328226 134112 328294
rect 133792 328170 133862 328226
rect 133918 328170 133986 328226
rect 134042 328170 134112 328226
rect 133792 328102 134112 328170
rect 133792 328046 133862 328102
rect 133918 328046 133986 328102
rect 134042 328046 134112 328102
rect 133792 327978 134112 328046
rect 133792 327922 133862 327978
rect 133918 327922 133986 327978
rect 134042 327922 134112 327978
rect 133792 327888 134112 327922
rect 164512 328350 164832 328384
rect 164512 328294 164582 328350
rect 164638 328294 164706 328350
rect 164762 328294 164832 328350
rect 164512 328226 164832 328294
rect 164512 328170 164582 328226
rect 164638 328170 164706 328226
rect 164762 328170 164832 328226
rect 164512 328102 164832 328170
rect 164512 328046 164582 328102
rect 164638 328046 164706 328102
rect 164762 328046 164832 328102
rect 164512 327978 164832 328046
rect 164512 327922 164582 327978
rect 164638 327922 164706 327978
rect 164762 327922 164832 327978
rect 164512 327888 164832 327922
rect 121772 319078 121828 319088
rect 121660 310978 121716 310988
rect 121436 283438 121492 283448
rect 121436 279748 121492 283382
rect 121548 281818 121604 281828
rect 121548 280756 121604 281762
rect 121548 280690 121604 280700
rect 121436 279682 121492 279692
rect 120540 276352 120596 276362
rect 120428 153794 120484 153804
rect 120316 146962 120372 146972
rect 121660 145460 121716 310922
rect 121660 145394 121716 145404
rect 121772 145348 121828 319022
rect 149152 316350 149472 316384
rect 149152 316294 149222 316350
rect 149278 316294 149346 316350
rect 149402 316294 149472 316350
rect 149152 316226 149472 316294
rect 149152 316170 149222 316226
rect 149278 316170 149346 316226
rect 149402 316170 149472 316226
rect 149152 316102 149472 316170
rect 149152 316046 149222 316102
rect 149278 316046 149346 316102
rect 149402 316046 149472 316102
rect 149152 315978 149472 316046
rect 149152 315922 149222 315978
rect 149278 315922 149346 315978
rect 149402 315922 149472 315978
rect 149152 315888 149472 315922
rect 179872 316350 180192 316384
rect 179872 316294 179942 316350
rect 179998 316294 180066 316350
rect 180122 316294 180192 316350
rect 179872 316226 180192 316294
rect 179872 316170 179942 316226
rect 179998 316170 180066 316226
rect 180122 316170 180192 316226
rect 179872 316102 180192 316170
rect 179872 316046 179942 316102
rect 179998 316046 180066 316102
rect 180122 316046 180192 316102
rect 179872 315978 180192 316046
rect 179872 315922 179942 315978
rect 179998 315922 180066 315978
rect 180122 315922 180192 315978
rect 179872 315888 180192 315922
rect 133792 310350 134112 310384
rect 133792 310294 133862 310350
rect 133918 310294 133986 310350
rect 134042 310294 134112 310350
rect 133792 310226 134112 310294
rect 133792 310170 133862 310226
rect 133918 310170 133986 310226
rect 134042 310170 134112 310226
rect 133792 310102 134112 310170
rect 133792 310046 133862 310102
rect 133918 310046 133986 310102
rect 134042 310046 134112 310102
rect 133792 309978 134112 310046
rect 133792 309922 133862 309978
rect 133918 309922 133986 309978
rect 134042 309922 134112 309978
rect 133792 309888 134112 309922
rect 164512 310350 164832 310384
rect 164512 310294 164582 310350
rect 164638 310294 164706 310350
rect 164762 310294 164832 310350
rect 164512 310226 164832 310294
rect 164512 310170 164582 310226
rect 164638 310170 164706 310226
rect 164762 310170 164832 310226
rect 164512 310102 164832 310170
rect 164512 310046 164582 310102
rect 164638 310046 164706 310102
rect 164762 310046 164832 310102
rect 164512 309978 164832 310046
rect 164512 309922 164582 309978
rect 164638 309922 164706 309978
rect 164762 309922 164832 309978
rect 164512 309888 164832 309922
rect 149152 298350 149472 298384
rect 149152 298294 149222 298350
rect 149278 298294 149346 298350
rect 149402 298294 149472 298350
rect 149152 298226 149472 298294
rect 149152 298170 149222 298226
rect 149278 298170 149346 298226
rect 149402 298170 149472 298226
rect 149152 298102 149472 298170
rect 149152 298046 149222 298102
rect 149278 298046 149346 298102
rect 149402 298046 149472 298102
rect 149152 297978 149472 298046
rect 149152 297922 149222 297978
rect 149278 297922 149346 297978
rect 149402 297922 149472 297978
rect 149152 297888 149472 297922
rect 179872 298350 180192 298384
rect 179872 298294 179942 298350
rect 179998 298294 180066 298350
rect 180122 298294 180192 298350
rect 179872 298226 180192 298294
rect 179872 298170 179942 298226
rect 179998 298170 180066 298226
rect 180122 298170 180192 298226
rect 179872 298102 180192 298170
rect 179872 298046 179942 298102
rect 179998 298046 180066 298102
rect 180122 298046 180192 298102
rect 179872 297978 180192 298046
rect 179872 297922 179942 297978
rect 179998 297922 180066 297978
rect 180122 297922 180192 297978
rect 179872 297888 180192 297922
rect 133792 292350 134112 292384
rect 133792 292294 133862 292350
rect 133918 292294 133986 292350
rect 134042 292294 134112 292350
rect 133792 292226 134112 292294
rect 133792 292170 133862 292226
rect 133918 292170 133986 292226
rect 134042 292170 134112 292226
rect 133792 292102 134112 292170
rect 133792 292046 133862 292102
rect 133918 292046 133986 292102
rect 134042 292046 134112 292102
rect 133792 291978 134112 292046
rect 133792 291922 133862 291978
rect 133918 291922 133986 291978
rect 134042 291922 134112 291978
rect 133792 291888 134112 291922
rect 164512 292350 164832 292384
rect 164512 292294 164582 292350
rect 164638 292294 164706 292350
rect 164762 292294 164832 292350
rect 164512 292226 164832 292294
rect 164512 292170 164582 292226
rect 164638 292170 164706 292226
rect 164762 292170 164832 292226
rect 164512 292102 164832 292170
rect 164512 292046 164582 292102
rect 164638 292046 164706 292102
rect 164762 292046 164832 292102
rect 164512 291978 164832 292046
rect 164512 291922 164582 291978
rect 164638 291922 164706 291978
rect 164762 291922 164832 291978
rect 164512 291888 164832 291922
rect 121884 284698 121940 284708
rect 121884 280084 121940 284642
rect 141036 283258 141092 283268
rect 139692 283078 139748 283088
rect 121884 280018 121940 280028
rect 122332 282358 122388 282368
rect 122332 280084 122388 282302
rect 127708 281638 127764 281648
rect 122332 280018 122388 280028
rect 127484 280532 127540 280542
rect 127484 280084 127540 280476
rect 127708 280532 127764 281582
rect 133644 281458 133700 281468
rect 127708 280466 127764 280476
rect 127484 280018 127540 280028
rect 128298 274350 128918 281298
rect 128298 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 128918 274350
rect 128298 274226 128918 274294
rect 128298 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 128918 274226
rect 128298 274102 128918 274170
rect 128298 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 128918 274102
rect 128298 273978 128918 274046
rect 128298 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 128918 273978
rect 122556 266532 122612 266542
rect 122556 165620 122612 266476
rect 127596 265078 127652 265088
rect 122556 165554 122612 165564
rect 126812 178138 126868 178148
rect 126252 162932 126308 162942
rect 126252 162838 126308 162876
rect 126252 162772 126308 162782
rect 126812 147924 126868 178082
rect 127596 165620 127652 265022
rect 127596 165554 127652 165564
rect 128298 256350 128918 273922
rect 128298 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 128918 256350
rect 128298 256226 128918 256294
rect 128298 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 128918 256226
rect 128298 256102 128918 256170
rect 128298 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 128918 256102
rect 128298 255978 128918 256046
rect 128298 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 128918 255978
rect 128298 238350 128918 255922
rect 128298 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 128918 238350
rect 128298 238226 128918 238294
rect 128298 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 128918 238226
rect 128298 238102 128918 238170
rect 128298 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 128918 238102
rect 128298 237978 128918 238046
rect 128298 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 128918 237978
rect 128298 220350 128918 237922
rect 128298 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 128918 220350
rect 128298 220226 128918 220294
rect 128298 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 128918 220226
rect 128298 220102 128918 220170
rect 128298 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 128918 220102
rect 128298 219978 128918 220046
rect 128298 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 128918 219978
rect 128298 202350 128918 219922
rect 128298 202294 128394 202350
rect 128450 202294 128518 202350
rect 128574 202294 128642 202350
rect 128698 202294 128766 202350
rect 128822 202294 128918 202350
rect 128298 202226 128918 202294
rect 128298 202170 128394 202226
rect 128450 202170 128518 202226
rect 128574 202170 128642 202226
rect 128698 202170 128766 202226
rect 128822 202170 128918 202226
rect 128298 202102 128918 202170
rect 128298 202046 128394 202102
rect 128450 202046 128518 202102
rect 128574 202046 128642 202102
rect 128698 202046 128766 202102
rect 128822 202046 128918 202102
rect 128298 201978 128918 202046
rect 128298 201922 128394 201978
rect 128450 201922 128518 201978
rect 128574 201922 128642 201978
rect 128698 201922 128766 201978
rect 128822 201922 128918 201978
rect 128298 184350 128918 201922
rect 128298 184294 128394 184350
rect 128450 184294 128518 184350
rect 128574 184294 128642 184350
rect 128698 184294 128766 184350
rect 128822 184294 128918 184350
rect 128298 184226 128918 184294
rect 128298 184170 128394 184226
rect 128450 184170 128518 184226
rect 128574 184170 128642 184226
rect 128698 184170 128766 184226
rect 128822 184170 128918 184226
rect 128298 184102 128918 184170
rect 128298 184046 128394 184102
rect 128450 184046 128518 184102
rect 128574 184046 128642 184102
rect 128698 184046 128766 184102
rect 128822 184046 128918 184102
rect 128298 183978 128918 184046
rect 128298 183922 128394 183978
rect 128450 183922 128518 183978
rect 128574 183922 128642 183978
rect 128698 183922 128766 183978
rect 128822 183922 128918 183978
rect 128298 166350 128918 183922
rect 132018 280350 132638 281298
rect 133644 280532 133700 281402
rect 133644 280466 133700 280476
rect 139692 280532 139748 283022
rect 139692 280466 139748 280476
rect 141036 280532 141092 283202
rect 141036 280466 141092 280476
rect 146412 282178 146468 282188
rect 146412 280532 146468 282122
rect 163660 281998 163716 282008
rect 146412 280466 146468 280476
rect 157052 280644 157108 280654
rect 132018 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 132638 280350
rect 132018 280226 132638 280294
rect 132018 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 132638 280226
rect 132018 280102 132638 280170
rect 132018 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 132638 280102
rect 132018 279978 132638 280046
rect 132018 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 132638 279978
rect 132018 262350 132638 279922
rect 137676 279748 137732 279758
rect 137004 278292 137060 278302
rect 137004 278038 137060 278236
rect 137004 277972 137060 277982
rect 132018 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 132638 262350
rect 132018 262226 132638 262294
rect 132018 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 132638 262226
rect 132018 262102 132638 262170
rect 132018 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 132638 262102
rect 132018 261978 132638 262046
rect 132018 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 132638 261978
rect 132018 244350 132638 261922
rect 132018 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 132638 244350
rect 132018 244226 132638 244294
rect 132018 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 132638 244226
rect 132018 244102 132638 244170
rect 132018 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 132638 244102
rect 132018 243978 132638 244046
rect 132018 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 132638 243978
rect 132018 226350 132638 243922
rect 132018 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 132638 226350
rect 132018 226226 132638 226294
rect 132018 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 132638 226226
rect 132018 226102 132638 226170
rect 132018 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 132638 226102
rect 132018 225978 132638 226046
rect 132018 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 132638 225978
rect 132018 208350 132638 225922
rect 132018 208294 132114 208350
rect 132170 208294 132238 208350
rect 132294 208294 132362 208350
rect 132418 208294 132486 208350
rect 132542 208294 132638 208350
rect 132018 208226 132638 208294
rect 132018 208170 132114 208226
rect 132170 208170 132238 208226
rect 132294 208170 132362 208226
rect 132418 208170 132486 208226
rect 132542 208170 132638 208226
rect 132018 208102 132638 208170
rect 132018 208046 132114 208102
rect 132170 208046 132238 208102
rect 132294 208046 132362 208102
rect 132418 208046 132486 208102
rect 132542 208046 132638 208102
rect 132018 207978 132638 208046
rect 132018 207922 132114 207978
rect 132170 207922 132238 207978
rect 132294 207922 132362 207978
rect 132418 207922 132486 207978
rect 132542 207922 132638 207978
rect 132018 190350 132638 207922
rect 132018 190294 132114 190350
rect 132170 190294 132238 190350
rect 132294 190294 132362 190350
rect 132418 190294 132486 190350
rect 132542 190294 132638 190350
rect 132018 190226 132638 190294
rect 132018 190170 132114 190226
rect 132170 190170 132238 190226
rect 132294 190170 132362 190226
rect 132418 190170 132486 190226
rect 132542 190170 132638 190226
rect 132018 190102 132638 190170
rect 132018 190046 132114 190102
rect 132170 190046 132238 190102
rect 132294 190046 132362 190102
rect 132418 190046 132486 190102
rect 132542 190046 132638 190102
rect 132018 189978 132638 190046
rect 132018 189922 132114 189978
rect 132170 189922 132238 189978
rect 132294 189922 132362 189978
rect 132418 189922 132486 189978
rect 132542 189922 132638 189978
rect 128298 166294 128394 166350
rect 128450 166294 128518 166350
rect 128574 166294 128642 166350
rect 128698 166294 128766 166350
rect 128822 166294 128918 166350
rect 128298 166226 128918 166294
rect 128298 166170 128394 166226
rect 128450 166170 128518 166226
rect 128574 166170 128642 166226
rect 128698 166170 128766 166226
rect 128822 166170 128918 166226
rect 128298 166102 128918 166170
rect 128298 166046 128394 166102
rect 128450 166046 128518 166102
rect 128574 166046 128642 166102
rect 128698 166046 128766 166102
rect 128822 166046 128918 166102
rect 128298 165978 128918 166046
rect 128298 165922 128394 165978
rect 128450 165922 128518 165978
rect 128574 165922 128642 165978
rect 128698 165922 128766 165978
rect 128822 165922 128918 165978
rect 126812 147858 126868 147868
rect 128298 148350 128918 165922
rect 129052 176518 129108 176528
rect 129052 155316 129108 176462
rect 129052 155250 129108 155260
rect 132018 172350 132638 189922
rect 132018 172294 132114 172350
rect 132170 172294 132238 172350
rect 132294 172294 132362 172350
rect 132418 172294 132486 172350
rect 132542 172294 132638 172350
rect 132018 172226 132638 172294
rect 132018 172170 132114 172226
rect 132170 172170 132238 172226
rect 132294 172170 132362 172226
rect 132418 172170 132486 172226
rect 132542 172170 132638 172226
rect 132018 172102 132638 172170
rect 132018 172046 132114 172102
rect 132170 172046 132238 172102
rect 132294 172046 132362 172102
rect 132418 172046 132486 172102
rect 132542 172046 132638 172102
rect 132018 171978 132638 172046
rect 132018 171922 132114 171978
rect 132170 171922 132238 171978
rect 132294 171922 132362 171978
rect 132418 171922 132486 171978
rect 132542 171922 132638 171978
rect 128298 148294 128394 148350
rect 128450 148294 128518 148350
rect 128574 148294 128642 148350
rect 128698 148294 128766 148350
rect 128822 148294 128918 148350
rect 128298 148226 128918 148294
rect 128298 148170 128394 148226
rect 128450 148170 128518 148226
rect 128574 148170 128642 148226
rect 128698 148170 128766 148226
rect 128822 148170 128918 148226
rect 128298 148102 128918 148170
rect 128298 148046 128394 148102
rect 128450 148046 128518 148102
rect 128574 148046 128642 148102
rect 128698 148046 128766 148102
rect 128822 148046 128918 148102
rect 128298 147978 128918 148046
rect 128298 147922 128394 147978
rect 128450 147922 128518 147978
rect 128574 147922 128642 147978
rect 128698 147922 128766 147978
rect 128822 147922 128918 147978
rect 121772 145282 121828 145292
rect 111906 136350 112382 136384
rect 111906 136294 111930 136350
rect 111986 136294 112054 136350
rect 112110 136294 112178 136350
rect 112234 136294 112302 136350
rect 112358 136294 112382 136350
rect 111906 136226 112382 136294
rect 111906 136170 111930 136226
rect 111986 136170 112054 136226
rect 112110 136170 112178 136226
rect 112234 136170 112302 136226
rect 112358 136170 112382 136226
rect 111906 136102 112382 136170
rect 111906 136046 111930 136102
rect 111986 136046 112054 136102
rect 112110 136046 112178 136102
rect 112234 136046 112302 136102
rect 112358 136046 112382 136102
rect 111906 135978 112382 136046
rect 111906 135922 111930 135978
rect 111986 135922 112054 135978
rect 112110 135922 112178 135978
rect 112234 135922 112302 135978
rect 112358 135922 112382 135978
rect 111906 135888 112382 135922
rect 111106 130350 111582 130384
rect 111106 130294 111130 130350
rect 111186 130294 111254 130350
rect 111310 130294 111378 130350
rect 111434 130294 111502 130350
rect 111558 130294 111582 130350
rect 111106 130226 111582 130294
rect 111106 130170 111130 130226
rect 111186 130170 111254 130226
rect 111310 130170 111378 130226
rect 111434 130170 111502 130226
rect 111558 130170 111582 130226
rect 111106 130102 111582 130170
rect 111106 130046 111130 130102
rect 111186 130046 111254 130102
rect 111310 130046 111378 130102
rect 111434 130046 111502 130102
rect 111558 130046 111582 130102
rect 111106 129978 111582 130046
rect 111106 129922 111130 129978
rect 111186 129922 111254 129978
rect 111310 129922 111378 129978
rect 111434 129922 111502 129978
rect 111558 129922 111582 129978
rect 111106 129888 111582 129922
rect 128298 130350 128918 147922
rect 128298 130294 128394 130350
rect 128450 130294 128518 130350
rect 128574 130294 128642 130350
rect 128698 130294 128766 130350
rect 128822 130294 128918 130350
rect 128298 130226 128918 130294
rect 128298 130170 128394 130226
rect 128450 130170 128518 130226
rect 128574 130170 128642 130226
rect 128698 130170 128766 130226
rect 128822 130170 128918 130226
rect 128298 130102 128918 130170
rect 128298 130046 128394 130102
rect 128450 130046 128518 130102
rect 128574 130046 128642 130102
rect 128698 130046 128766 130102
rect 128822 130046 128918 130102
rect 128298 129978 128918 130046
rect 128298 129922 128394 129978
rect 128450 129922 128518 129978
rect 128574 129922 128642 129978
rect 128698 129922 128766 129978
rect 128822 129922 128918 129978
rect 111906 118350 112382 118384
rect 111906 118294 111930 118350
rect 111986 118294 112054 118350
rect 112110 118294 112178 118350
rect 112234 118294 112302 118350
rect 112358 118294 112382 118350
rect 111906 118226 112382 118294
rect 111906 118170 111930 118226
rect 111986 118170 112054 118226
rect 112110 118170 112178 118226
rect 112234 118170 112302 118226
rect 112358 118170 112382 118226
rect 111906 118102 112382 118170
rect 111906 118046 111930 118102
rect 111986 118046 112054 118102
rect 112110 118046 112178 118102
rect 112234 118046 112302 118102
rect 112358 118046 112382 118102
rect 111906 117978 112382 118046
rect 111906 117922 111930 117978
rect 111986 117922 112054 117978
rect 112110 117922 112178 117978
rect 112234 117922 112302 117978
rect 112358 117922 112382 117978
rect 111906 117888 112382 117922
rect 111106 112350 111582 112384
rect 111106 112294 111130 112350
rect 111186 112294 111254 112350
rect 111310 112294 111378 112350
rect 111434 112294 111502 112350
rect 111558 112294 111582 112350
rect 111106 112226 111582 112294
rect 111106 112170 111130 112226
rect 111186 112170 111254 112226
rect 111310 112170 111378 112226
rect 111434 112170 111502 112226
rect 111558 112170 111582 112226
rect 111106 112102 111582 112170
rect 111106 112046 111130 112102
rect 111186 112046 111254 112102
rect 111310 112046 111378 112102
rect 111434 112046 111502 112102
rect 111558 112046 111582 112102
rect 111106 111978 111582 112046
rect 111106 111922 111130 111978
rect 111186 111922 111254 111978
rect 111310 111922 111378 111978
rect 111434 111922 111502 111978
rect 111558 111922 111582 111978
rect 111106 111888 111582 111922
rect 128298 112350 128918 129922
rect 128298 112294 128394 112350
rect 128450 112294 128518 112350
rect 128574 112294 128642 112350
rect 128698 112294 128766 112350
rect 128822 112294 128918 112350
rect 128298 112226 128918 112294
rect 128298 112170 128394 112226
rect 128450 112170 128518 112226
rect 128574 112170 128642 112226
rect 128698 112170 128766 112226
rect 128822 112170 128918 112226
rect 128298 112102 128918 112170
rect 128298 112046 128394 112102
rect 128450 112046 128518 112102
rect 128574 112046 128642 112102
rect 128698 112046 128766 112102
rect 128822 112046 128918 112102
rect 128298 111978 128918 112046
rect 128298 111922 128394 111978
rect 128450 111922 128518 111978
rect 128574 111922 128642 111978
rect 128698 111922 128766 111978
rect 128822 111922 128918 111978
rect 111906 100350 112382 100384
rect 111906 100294 111930 100350
rect 111986 100294 112054 100350
rect 112110 100294 112178 100350
rect 112234 100294 112302 100350
rect 112358 100294 112382 100350
rect 111906 100226 112382 100294
rect 111906 100170 111930 100226
rect 111986 100170 112054 100226
rect 112110 100170 112178 100226
rect 112234 100170 112302 100226
rect 112358 100170 112382 100226
rect 111906 100102 112382 100170
rect 111906 100046 111930 100102
rect 111986 100046 112054 100102
rect 112110 100046 112178 100102
rect 112234 100046 112302 100102
rect 112358 100046 112382 100102
rect 111906 99978 112382 100046
rect 111906 99922 111930 99978
rect 111986 99922 112054 99978
rect 112110 99922 112178 99978
rect 112234 99922 112302 99978
rect 112358 99922 112382 99978
rect 111906 99888 112382 99922
rect 111106 94350 111582 94384
rect 111106 94294 111130 94350
rect 111186 94294 111254 94350
rect 111310 94294 111378 94350
rect 111434 94294 111502 94350
rect 111558 94294 111582 94350
rect 111106 94226 111582 94294
rect 111106 94170 111130 94226
rect 111186 94170 111254 94226
rect 111310 94170 111378 94226
rect 111434 94170 111502 94226
rect 111558 94170 111582 94226
rect 111106 94102 111582 94170
rect 111106 94046 111130 94102
rect 111186 94046 111254 94102
rect 111310 94046 111378 94102
rect 111434 94046 111502 94102
rect 111558 94046 111582 94102
rect 111106 93978 111582 94046
rect 111106 93922 111130 93978
rect 111186 93922 111254 93978
rect 111310 93922 111378 93978
rect 111434 93922 111502 93978
rect 111558 93922 111582 93978
rect 111106 93888 111582 93922
rect 128298 94350 128918 111922
rect 128298 94294 128394 94350
rect 128450 94294 128518 94350
rect 128574 94294 128642 94350
rect 128698 94294 128766 94350
rect 128822 94294 128918 94350
rect 128298 94226 128918 94294
rect 128298 94170 128394 94226
rect 128450 94170 128518 94226
rect 128574 94170 128642 94226
rect 128698 94170 128766 94226
rect 128822 94170 128918 94226
rect 128298 94102 128918 94170
rect 128298 94046 128394 94102
rect 128450 94046 128518 94102
rect 128574 94046 128642 94102
rect 128698 94046 128766 94102
rect 128822 94046 128918 94102
rect 128298 93978 128918 94046
rect 128298 93922 128394 93978
rect 128450 93922 128518 93978
rect 128574 93922 128642 93978
rect 128698 93922 128766 93978
rect 128822 93922 128918 93978
rect 111906 82350 112382 82384
rect 111906 82294 111930 82350
rect 111986 82294 112054 82350
rect 112110 82294 112178 82350
rect 112234 82294 112302 82350
rect 112358 82294 112382 82350
rect 111906 82226 112382 82294
rect 111906 82170 111930 82226
rect 111986 82170 112054 82226
rect 112110 82170 112178 82226
rect 112234 82170 112302 82226
rect 112358 82170 112382 82226
rect 111906 82102 112382 82170
rect 111906 82046 111930 82102
rect 111986 82046 112054 82102
rect 112110 82046 112178 82102
rect 112234 82046 112302 82102
rect 112358 82046 112382 82102
rect 111906 81978 112382 82046
rect 111906 81922 111930 81978
rect 111986 81922 112054 81978
rect 112110 81922 112178 81978
rect 112234 81922 112302 81978
rect 112358 81922 112382 81978
rect 111906 81888 112382 81922
rect 111106 76350 111582 76384
rect 111106 76294 111130 76350
rect 111186 76294 111254 76350
rect 111310 76294 111378 76350
rect 111434 76294 111502 76350
rect 111558 76294 111582 76350
rect 111106 76226 111582 76294
rect 111106 76170 111130 76226
rect 111186 76170 111254 76226
rect 111310 76170 111378 76226
rect 111434 76170 111502 76226
rect 111558 76170 111582 76226
rect 111106 76102 111582 76170
rect 111106 76046 111130 76102
rect 111186 76046 111254 76102
rect 111310 76046 111378 76102
rect 111434 76046 111502 76102
rect 111558 76046 111582 76102
rect 111106 75978 111582 76046
rect 111106 75922 111130 75978
rect 111186 75922 111254 75978
rect 111310 75922 111378 75978
rect 111434 75922 111502 75978
rect 111558 75922 111582 75978
rect 111106 75888 111582 75922
rect 128298 76350 128918 93922
rect 128298 76294 128394 76350
rect 128450 76294 128518 76350
rect 128574 76294 128642 76350
rect 128698 76294 128766 76350
rect 128822 76294 128918 76350
rect 128298 76226 128918 76294
rect 128298 76170 128394 76226
rect 128450 76170 128518 76226
rect 128574 76170 128642 76226
rect 128698 76170 128766 76226
rect 128822 76170 128918 76226
rect 128298 76102 128918 76170
rect 128298 76046 128394 76102
rect 128450 76046 128518 76102
rect 128574 76046 128642 76102
rect 128698 76046 128766 76102
rect 128822 76046 128918 76102
rect 128298 75978 128918 76046
rect 128298 75922 128394 75978
rect 128450 75922 128518 75978
rect 128574 75922 128642 75978
rect 128698 75922 128766 75978
rect 128822 75922 128918 75978
rect 111906 64350 112382 64384
rect 111906 64294 111930 64350
rect 111986 64294 112054 64350
rect 112110 64294 112178 64350
rect 112234 64294 112302 64350
rect 112358 64294 112382 64350
rect 111906 64226 112382 64294
rect 111906 64170 111930 64226
rect 111986 64170 112054 64226
rect 112110 64170 112178 64226
rect 112234 64170 112302 64226
rect 112358 64170 112382 64226
rect 111906 64102 112382 64170
rect 111906 64046 111930 64102
rect 111986 64046 112054 64102
rect 112110 64046 112178 64102
rect 112234 64046 112302 64102
rect 112358 64046 112382 64102
rect 111906 63978 112382 64046
rect 111906 63922 111930 63978
rect 111986 63922 112054 63978
rect 112110 63922 112178 63978
rect 112234 63922 112302 63978
rect 112358 63922 112382 63978
rect 111906 63888 112382 63922
rect 111106 58350 111582 58384
rect 111106 58294 111130 58350
rect 111186 58294 111254 58350
rect 111310 58294 111378 58350
rect 111434 58294 111502 58350
rect 111558 58294 111582 58350
rect 111106 58226 111582 58294
rect 111106 58170 111130 58226
rect 111186 58170 111254 58226
rect 111310 58170 111378 58226
rect 111434 58170 111502 58226
rect 111558 58170 111582 58226
rect 111106 58102 111582 58170
rect 111106 58046 111130 58102
rect 111186 58046 111254 58102
rect 111310 58046 111378 58102
rect 111434 58046 111502 58102
rect 111558 58046 111582 58102
rect 111106 57978 111582 58046
rect 111106 57922 111130 57978
rect 111186 57922 111254 57978
rect 111310 57922 111378 57978
rect 111434 57922 111502 57978
rect 111558 57922 111582 57978
rect 111106 57888 111582 57922
rect 128298 58350 128918 75922
rect 128298 58294 128394 58350
rect 128450 58294 128518 58350
rect 128574 58294 128642 58350
rect 128698 58294 128766 58350
rect 128822 58294 128918 58350
rect 128298 58226 128918 58294
rect 128298 58170 128394 58226
rect 128450 58170 128518 58226
rect 128574 58170 128642 58226
rect 128698 58170 128766 58226
rect 128822 58170 128918 58226
rect 128298 58102 128918 58170
rect 128298 58046 128394 58102
rect 128450 58046 128518 58102
rect 128574 58046 128642 58102
rect 128698 58046 128766 58102
rect 128822 58046 128918 58102
rect 128298 57978 128918 58046
rect 128298 57922 128394 57978
rect 128450 57922 128518 57978
rect 128574 57922 128642 57978
rect 128698 57922 128766 57978
rect 128822 57922 128918 57978
rect 110012 36754 110068 36764
rect 128298 40350 128918 57922
rect 128298 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 128918 40350
rect 128298 40226 128918 40294
rect 128298 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 128918 40226
rect 128298 40102 128918 40170
rect 128298 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 128918 40102
rect 128298 39978 128918 40046
rect 128298 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 128918 39978
rect 101298 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 101918 28350
rect 101298 28226 101918 28294
rect 101298 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 101918 28226
rect 101298 28102 101918 28170
rect 101298 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 101918 28102
rect 101298 27978 101918 28046
rect 101298 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 101918 27978
rect 101298 10350 101918 27922
rect 101298 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 101918 10350
rect 101298 10226 101918 10294
rect 101298 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 101918 10226
rect 101298 10102 101918 10170
rect 101298 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 101918 10102
rect 101298 9978 101918 10046
rect 101298 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 101918 9978
rect 101298 -1120 101918 9922
rect 101298 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 101918 -1120
rect 101298 -1244 101918 -1176
rect 101298 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 101918 -1244
rect 101298 -1368 101918 -1300
rect 101298 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 101918 -1368
rect 101298 -1492 101918 -1424
rect 101298 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 101918 -1492
rect 101298 -1644 101918 -1548
rect 128298 22350 128918 39922
rect 128298 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 128918 22350
rect 128298 22226 128918 22294
rect 128298 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 128918 22226
rect 128298 22102 128918 22170
rect 128298 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 128918 22102
rect 128298 21978 128918 22046
rect 128298 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 128918 21978
rect 128298 4350 128918 21922
rect 128298 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 128918 4350
rect 128298 4226 128918 4294
rect 128298 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 128918 4226
rect 128298 4102 128918 4170
rect 128298 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 128918 4102
rect 128298 3978 128918 4046
rect 128298 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 128918 3978
rect 128298 -160 128918 3922
rect 128298 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 128918 -160
rect 128298 -284 128918 -216
rect 128298 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 128918 -284
rect 128298 -408 128918 -340
rect 128298 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 128918 -408
rect 128298 -532 128918 -464
rect 128298 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 128918 -532
rect 128298 -1644 128918 -588
rect 132018 154350 132638 171922
rect 132018 154294 132114 154350
rect 132170 154294 132238 154350
rect 132294 154294 132362 154350
rect 132418 154294 132486 154350
rect 132542 154294 132638 154350
rect 132018 154226 132638 154294
rect 132018 154170 132114 154226
rect 132170 154170 132238 154226
rect 132294 154170 132362 154226
rect 132418 154170 132486 154226
rect 132542 154170 132638 154226
rect 132018 154102 132638 154170
rect 132018 154046 132114 154102
rect 132170 154046 132238 154102
rect 132294 154046 132362 154102
rect 132418 154046 132486 154102
rect 132542 154046 132638 154102
rect 132018 153978 132638 154046
rect 132018 153922 132114 153978
rect 132170 153922 132238 153978
rect 132294 153922 132362 153978
rect 132418 153922 132486 153978
rect 132542 153922 132638 153978
rect 132018 136350 132638 153922
rect 137452 149044 137508 149054
rect 137452 148596 137508 148988
rect 137452 148530 137508 148540
rect 137676 148484 137732 279692
rect 155372 278578 155428 278588
rect 154476 278180 154532 278190
rect 151116 277172 151172 277182
rect 151116 276418 151172 277116
rect 151116 276352 151172 276362
rect 150332 274596 150388 274606
rect 139356 268436 139412 268446
rect 138572 173098 138628 173108
rect 138572 161308 138628 173042
rect 138572 161252 138740 161308
rect 138684 150388 138740 161252
rect 138684 150322 138740 150332
rect 139356 149044 139412 268380
rect 139356 148978 139412 148988
rect 137676 148418 137732 148428
rect 150332 147140 150388 274540
rect 154476 165620 154532 278124
rect 154476 165554 154532 165564
rect 155372 147364 155428 278522
rect 157052 162820 157108 280588
rect 157948 277172 158004 277182
rect 157948 276598 158004 277116
rect 157948 276532 158004 276542
rect 157052 162754 157108 162764
rect 159018 274350 159638 281298
rect 162738 280350 163358 281298
rect 163660 280532 163716 281942
rect 163660 280466 163716 280476
rect 186396 280532 186452 280542
rect 162738 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 163358 280350
rect 162738 280226 163358 280294
rect 162738 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 163358 280226
rect 162738 280102 163358 280170
rect 162738 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 163358 280102
rect 162738 279978 163358 280046
rect 162738 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 163358 279978
rect 159964 277172 160020 277182
rect 159964 276778 160020 277116
rect 159964 276712 160020 276722
rect 160412 276948 160468 276958
rect 159018 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 159638 274350
rect 159018 274226 159638 274294
rect 159018 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 159638 274226
rect 159018 274102 159638 274170
rect 159018 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 159638 274102
rect 159018 273978 159638 274046
rect 159018 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 159638 273978
rect 159018 256350 159638 273922
rect 159018 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 159638 256350
rect 159018 256226 159638 256294
rect 159018 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 159638 256226
rect 159018 256102 159638 256170
rect 159018 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 159638 256102
rect 159018 255978 159638 256046
rect 159018 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 159638 255978
rect 159018 238350 159638 255922
rect 159018 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 159638 238350
rect 159018 238226 159638 238294
rect 159018 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 159638 238226
rect 159018 238102 159638 238170
rect 159018 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 159638 238102
rect 159018 237978 159638 238046
rect 159018 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 159638 237978
rect 159018 220350 159638 237922
rect 159018 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 159638 220350
rect 159018 220226 159638 220294
rect 159018 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 159638 220226
rect 159018 220102 159638 220170
rect 159018 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 159638 220102
rect 159018 219978 159638 220046
rect 159018 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 159638 219978
rect 159018 202350 159638 219922
rect 159018 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 159638 202350
rect 159018 202226 159638 202294
rect 159018 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 159638 202226
rect 159018 202102 159638 202170
rect 159018 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 159638 202102
rect 159018 201978 159638 202046
rect 159018 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 159638 201978
rect 159018 184350 159638 201922
rect 159018 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 159638 184350
rect 159018 184226 159638 184294
rect 159018 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 159638 184226
rect 159018 184102 159638 184170
rect 159018 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 159638 184102
rect 159018 183978 159638 184046
rect 159018 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 159638 183978
rect 159018 166350 159638 183922
rect 159018 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 159638 166350
rect 159018 166226 159638 166294
rect 159018 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 159638 166226
rect 159018 166102 159638 166170
rect 159018 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 159638 166102
rect 159018 165978 159638 166046
rect 159018 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 159638 165978
rect 155372 147298 155428 147308
rect 159018 148350 159638 165922
rect 160412 158900 160468 276892
rect 160524 276724 160580 276734
rect 160524 257878 160580 276668
rect 160524 257812 160580 257822
rect 162738 262350 163358 279922
rect 186284 280420 186340 280430
rect 165676 279860 165732 279870
rect 165228 277172 165284 277182
rect 165228 276958 165284 277116
rect 165228 276892 165284 276902
rect 163772 276836 163828 276846
rect 163772 266698 163828 276780
rect 163772 266632 163828 266642
rect 162738 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 163358 262350
rect 162738 262226 163358 262294
rect 162738 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 163358 262226
rect 162738 262102 163358 262170
rect 162738 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 163358 262102
rect 162738 261978 163358 262046
rect 162738 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 163358 261978
rect 162738 244350 163358 261922
rect 162738 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 163358 244350
rect 162738 244226 163358 244294
rect 162738 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 163358 244226
rect 162738 244102 163358 244170
rect 162738 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 163358 244102
rect 162738 243978 163358 244046
rect 162738 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 163358 243978
rect 162738 226350 163358 243922
rect 162738 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 163358 226350
rect 162738 226226 163358 226294
rect 162738 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 163358 226226
rect 162738 226102 163358 226170
rect 162738 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 163358 226102
rect 162738 225978 163358 226046
rect 162738 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 163358 225978
rect 160524 214138 160580 214148
rect 160524 164612 160580 214082
rect 160524 164546 160580 164556
rect 162738 208350 163358 225922
rect 162738 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 163358 208350
rect 162738 208226 163358 208294
rect 162738 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 163358 208226
rect 162738 208102 163358 208170
rect 162738 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 163358 208102
rect 162738 207978 163358 208046
rect 162738 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 163358 207978
rect 162738 190350 163358 207922
rect 162738 190294 162834 190350
rect 162890 190294 162958 190350
rect 163014 190294 163082 190350
rect 163138 190294 163206 190350
rect 163262 190294 163358 190350
rect 162738 190226 163358 190294
rect 162738 190170 162834 190226
rect 162890 190170 162958 190226
rect 163014 190170 163082 190226
rect 163138 190170 163206 190226
rect 163262 190170 163358 190226
rect 162738 190102 163358 190170
rect 162738 190046 162834 190102
rect 162890 190046 162958 190102
rect 163014 190046 163082 190102
rect 163138 190046 163206 190102
rect 163262 190046 163358 190102
rect 162738 189978 163358 190046
rect 162738 189922 162834 189978
rect 162890 189922 162958 189978
rect 163014 189922 163082 189978
rect 163138 189922 163206 189978
rect 163262 189922 163358 189978
rect 162738 172350 163358 189922
rect 162738 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 163358 172350
rect 162738 172226 163358 172294
rect 162738 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 163358 172226
rect 162738 172102 163358 172170
rect 162738 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 163358 172102
rect 162738 171978 163358 172046
rect 162738 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 163358 171978
rect 160412 158834 160468 158844
rect 159018 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 159638 148350
rect 159018 148226 159638 148294
rect 159018 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 159638 148226
rect 159018 148102 159638 148170
rect 159018 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 159638 148102
rect 159018 147978 159638 148046
rect 159018 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 159638 147978
rect 150332 147074 150388 147084
rect 132018 136294 132114 136350
rect 132170 136294 132238 136350
rect 132294 136294 132362 136350
rect 132418 136294 132486 136350
rect 132542 136294 132638 136350
rect 132018 136226 132638 136294
rect 132018 136170 132114 136226
rect 132170 136170 132238 136226
rect 132294 136170 132362 136226
rect 132418 136170 132486 136226
rect 132542 136170 132638 136226
rect 132018 136102 132638 136170
rect 132018 136046 132114 136102
rect 132170 136046 132238 136102
rect 132294 136046 132362 136102
rect 132418 136046 132486 136102
rect 132542 136046 132638 136102
rect 132018 135978 132638 136046
rect 132018 135922 132114 135978
rect 132170 135922 132238 135978
rect 132294 135922 132362 135978
rect 132418 135922 132486 135978
rect 132542 135922 132638 135978
rect 132018 118350 132638 135922
rect 132018 118294 132114 118350
rect 132170 118294 132238 118350
rect 132294 118294 132362 118350
rect 132418 118294 132486 118350
rect 132542 118294 132638 118350
rect 132018 118226 132638 118294
rect 132018 118170 132114 118226
rect 132170 118170 132238 118226
rect 132294 118170 132362 118226
rect 132418 118170 132486 118226
rect 132542 118170 132638 118226
rect 132018 118102 132638 118170
rect 132018 118046 132114 118102
rect 132170 118046 132238 118102
rect 132294 118046 132362 118102
rect 132418 118046 132486 118102
rect 132542 118046 132638 118102
rect 132018 117978 132638 118046
rect 132018 117922 132114 117978
rect 132170 117922 132238 117978
rect 132294 117922 132362 117978
rect 132418 117922 132486 117978
rect 132542 117922 132638 117978
rect 132018 100350 132638 117922
rect 132018 100294 132114 100350
rect 132170 100294 132238 100350
rect 132294 100294 132362 100350
rect 132418 100294 132486 100350
rect 132542 100294 132638 100350
rect 132018 100226 132638 100294
rect 132018 100170 132114 100226
rect 132170 100170 132238 100226
rect 132294 100170 132362 100226
rect 132418 100170 132486 100226
rect 132542 100170 132638 100226
rect 132018 100102 132638 100170
rect 132018 100046 132114 100102
rect 132170 100046 132238 100102
rect 132294 100046 132362 100102
rect 132418 100046 132486 100102
rect 132542 100046 132638 100102
rect 132018 99978 132638 100046
rect 132018 99922 132114 99978
rect 132170 99922 132238 99978
rect 132294 99922 132362 99978
rect 132418 99922 132486 99978
rect 132542 99922 132638 99978
rect 132018 82350 132638 99922
rect 132018 82294 132114 82350
rect 132170 82294 132238 82350
rect 132294 82294 132362 82350
rect 132418 82294 132486 82350
rect 132542 82294 132638 82350
rect 132018 82226 132638 82294
rect 132018 82170 132114 82226
rect 132170 82170 132238 82226
rect 132294 82170 132362 82226
rect 132418 82170 132486 82226
rect 132542 82170 132638 82226
rect 132018 82102 132638 82170
rect 132018 82046 132114 82102
rect 132170 82046 132238 82102
rect 132294 82046 132362 82102
rect 132418 82046 132486 82102
rect 132542 82046 132638 82102
rect 132018 81978 132638 82046
rect 132018 81922 132114 81978
rect 132170 81922 132238 81978
rect 132294 81922 132362 81978
rect 132418 81922 132486 81978
rect 132542 81922 132638 81978
rect 132018 64350 132638 81922
rect 132018 64294 132114 64350
rect 132170 64294 132238 64350
rect 132294 64294 132362 64350
rect 132418 64294 132486 64350
rect 132542 64294 132638 64350
rect 132018 64226 132638 64294
rect 132018 64170 132114 64226
rect 132170 64170 132238 64226
rect 132294 64170 132362 64226
rect 132418 64170 132486 64226
rect 132542 64170 132638 64226
rect 132018 64102 132638 64170
rect 132018 64046 132114 64102
rect 132170 64046 132238 64102
rect 132294 64046 132362 64102
rect 132418 64046 132486 64102
rect 132542 64046 132638 64102
rect 132018 63978 132638 64046
rect 132018 63922 132114 63978
rect 132170 63922 132238 63978
rect 132294 63922 132362 63978
rect 132418 63922 132486 63978
rect 132542 63922 132638 63978
rect 132018 46350 132638 63922
rect 132018 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 132638 46350
rect 132018 46226 132638 46294
rect 132018 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 132638 46226
rect 132018 46102 132638 46170
rect 132018 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 132638 46102
rect 132018 45978 132638 46046
rect 132018 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 132638 45978
rect 132018 28350 132638 45922
rect 159018 130350 159638 147922
rect 159018 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 159638 130350
rect 159018 130226 159638 130294
rect 159018 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 159638 130226
rect 159018 130102 159638 130170
rect 159018 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 159638 130102
rect 159018 129978 159638 130046
rect 159018 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 159638 129978
rect 159018 112350 159638 129922
rect 159018 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 159638 112350
rect 159018 112226 159638 112294
rect 159018 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 159638 112226
rect 159018 112102 159638 112170
rect 159018 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 159638 112102
rect 159018 111978 159638 112046
rect 159018 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 159638 111978
rect 159018 94350 159638 111922
rect 159018 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 159638 94350
rect 159018 94226 159638 94294
rect 159018 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 159638 94226
rect 159018 94102 159638 94170
rect 159018 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 159638 94102
rect 159018 93978 159638 94046
rect 159018 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 159638 93978
rect 159018 76350 159638 93922
rect 159018 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 159638 76350
rect 159018 76226 159638 76294
rect 159018 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 159638 76226
rect 159018 76102 159638 76170
rect 159018 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 159638 76102
rect 159018 75978 159638 76046
rect 159018 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 159638 75978
rect 159018 58350 159638 75922
rect 159018 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 159638 58350
rect 159018 58226 159638 58294
rect 159018 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 159638 58226
rect 159018 58102 159638 58170
rect 159018 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 159638 58102
rect 159018 57978 159638 58046
rect 159018 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 159638 57978
rect 159018 40350 159638 57922
rect 159018 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 159638 40350
rect 159018 40226 159638 40294
rect 159018 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 159638 40226
rect 159018 40102 159638 40170
rect 159018 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 159638 40102
rect 159018 39978 159638 40046
rect 159018 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 159638 39978
rect 132018 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 132638 28350
rect 132018 28226 132638 28294
rect 132018 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 132638 28226
rect 132018 28102 132638 28170
rect 132018 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 132638 28102
rect 132018 27978 132638 28046
rect 132018 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 132638 27978
rect 132018 10350 132638 27922
rect 150488 28350 150808 28384
rect 150488 28294 150558 28350
rect 150614 28294 150682 28350
rect 150738 28294 150808 28350
rect 150488 28226 150808 28294
rect 150488 28170 150558 28226
rect 150614 28170 150682 28226
rect 150738 28170 150808 28226
rect 150488 28102 150808 28170
rect 150488 28046 150558 28102
rect 150614 28046 150682 28102
rect 150738 28046 150808 28102
rect 150488 27978 150808 28046
rect 150488 27922 150558 27978
rect 150614 27922 150682 27978
rect 150738 27922 150808 27978
rect 150488 27888 150808 27922
rect 159018 22350 159638 39922
rect 159018 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 159638 22350
rect 159018 22226 159638 22294
rect 159018 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 159638 22226
rect 159018 22102 159638 22170
rect 159018 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 159638 22102
rect 159018 21978 159638 22046
rect 159018 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 159638 21978
rect 132018 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 132638 10350
rect 132018 10226 132638 10294
rect 132018 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 132638 10226
rect 132018 10102 132638 10170
rect 132018 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 132638 10102
rect 132018 9978 132638 10046
rect 132018 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 132638 9978
rect 132018 -1120 132638 9922
rect 150488 10350 150808 10384
rect 150488 10294 150558 10350
rect 150614 10294 150682 10350
rect 150738 10294 150808 10350
rect 150488 10226 150808 10294
rect 150488 10170 150558 10226
rect 150614 10170 150682 10226
rect 150738 10170 150808 10226
rect 150488 10102 150808 10170
rect 150488 10046 150558 10102
rect 150614 10046 150682 10102
rect 150738 10046 150808 10102
rect 150488 9978 150808 10046
rect 150488 9922 150558 9978
rect 150614 9922 150682 9978
rect 150738 9922 150808 9978
rect 150488 9888 150808 9922
rect 132018 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 132638 -1120
rect 132018 -1244 132638 -1176
rect 132018 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 132638 -1244
rect 132018 -1368 132638 -1300
rect 132018 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 132638 -1368
rect 132018 -1492 132638 -1424
rect 132018 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 132638 -1492
rect 132018 -1644 132638 -1548
rect 159018 4350 159638 21922
rect 159018 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 159638 4350
rect 159018 4226 159638 4294
rect 159018 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 159638 4226
rect 159018 4102 159638 4170
rect 159018 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 159638 4102
rect 159018 3978 159638 4046
rect 159018 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 159638 3978
rect 159018 -160 159638 3922
rect 159018 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 159638 -160
rect 159018 -284 159638 -216
rect 159018 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 159638 -284
rect 159018 -408 159638 -340
rect 159018 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 159638 -408
rect 159018 -532 159638 -464
rect 159018 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 159638 -532
rect 159018 -1644 159638 -588
rect 162738 154350 163358 171922
rect 165676 163940 165732 279804
rect 174636 278740 174692 278750
rect 170492 278628 170548 278638
rect 168812 278292 168868 278302
rect 165900 277172 165956 277182
rect 165900 277072 165956 277082
rect 168140 275604 168196 275614
rect 165676 163874 165732 163884
rect 167132 271348 167188 271358
rect 167132 159460 167188 271292
rect 168140 266518 168196 275548
rect 168140 266452 168196 266462
rect 168812 255388 168868 278236
rect 169260 275604 169316 275614
rect 169260 268318 169316 275548
rect 169260 268252 169316 268262
rect 169708 275604 169764 275614
rect 169708 264718 169764 275548
rect 169708 264652 169764 264662
rect 168028 255358 168868 255388
rect 168084 255332 168868 255358
rect 168028 214138 168084 255302
rect 168028 214072 168084 214082
rect 170492 162932 170548 278572
rect 174636 278398 174692 278684
rect 174636 278332 174692 278342
rect 186172 278404 186228 278414
rect 175308 277318 175364 277328
rect 175308 277172 175364 277262
rect 175308 277106 175364 277116
rect 178892 277172 178948 277182
rect 178892 276612 178948 277116
rect 173852 276418 173908 276428
rect 172172 270004 172228 270014
rect 172172 164500 172228 269948
rect 172172 164434 172228 164444
rect 173852 261658 173908 276362
rect 175980 276276 176036 276286
rect 175980 273538 176036 276220
rect 175980 273472 176036 273482
rect 176540 275604 176596 275614
rect 173852 212518 173908 261602
rect 176428 270564 176484 270574
rect 176428 218278 176484 270508
rect 176540 269938 176596 275548
rect 177324 275604 177380 275614
rect 177324 271558 177380 275548
rect 177324 271492 177380 271502
rect 178108 275604 178164 275614
rect 176540 269872 176596 269882
rect 178108 267958 178164 275548
rect 178108 267892 178164 267902
rect 176428 216838 176484 218222
rect 170492 162866 170548 162876
rect 173852 160804 173908 212462
rect 176316 216782 176484 216838
rect 176316 196588 176372 216782
rect 175532 196532 176372 196588
rect 177212 209998 177268 210008
rect 175532 164612 175588 196532
rect 175532 164546 175588 164556
rect 177212 160916 177268 209942
rect 178892 209998 178948 276556
rect 181356 277060 181412 277070
rect 180012 275828 180068 275838
rect 179788 275716 179844 275726
rect 179788 264898 179844 275660
rect 179900 275604 179956 275614
rect 179900 266338 179956 275548
rect 180012 268138 180068 275772
rect 180012 268072 180068 268082
rect 179900 266272 179956 266282
rect 179788 264832 179844 264842
rect 178892 209932 178948 209942
rect 179228 164388 179284 164398
rect 179228 163156 179284 164332
rect 179228 163090 179284 163100
rect 177212 160850 177268 160860
rect 173852 160738 173908 160748
rect 167132 159394 167188 159404
rect 181356 159572 181412 277004
rect 184716 275828 184772 275838
rect 183148 275716 183204 275726
rect 181468 275604 181524 275614
rect 181468 264538 181524 275548
rect 183148 270298 183204 275660
rect 184716 271918 184772 275772
rect 184716 271852 184772 271862
rect 184828 275604 184884 275614
rect 184828 270478 184884 275548
rect 184828 270412 184884 270422
rect 183148 270232 183204 270242
rect 181468 264472 181524 264482
rect 183036 265412 183092 265422
rect 183036 219178 183092 265356
rect 183932 262918 183988 262928
rect 183932 222598 183988 262862
rect 186172 260398 186228 278348
rect 186172 260332 186228 260342
rect 183932 222532 183988 222542
rect 184716 222598 184772 222608
rect 183036 165620 183092 219122
rect 184716 173068 184772 222542
rect 186284 201538 186340 280364
rect 186284 201472 186340 201482
rect 186396 191458 186452 280476
rect 187404 278516 187460 278526
rect 187404 278218 187460 278460
rect 187404 278152 187460 278162
rect 189532 276778 189588 276788
rect 189420 276722 189532 276778
rect 189420 276500 189476 276722
rect 189532 276712 189588 276722
rect 188972 276388 189028 276398
rect 186732 276276 186788 276286
rect 186732 273718 186788 276220
rect 186732 273652 186788 273662
rect 188076 275716 188132 275726
rect 188076 272098 188132 275660
rect 188076 272032 188132 272042
rect 188748 275604 188804 275614
rect 188748 271738 188804 275548
rect 188748 271672 188804 271682
rect 187404 265524 187460 265534
rect 186396 191392 186452 191402
rect 187292 260398 187348 260408
rect 183036 165554 183092 165564
rect 184492 173012 184772 173068
rect 184492 165620 184548 173012
rect 184492 165554 184548 165564
rect 187292 172738 187348 260342
rect 187404 225118 187460 265468
rect 187404 225052 187460 225062
rect 181356 158004 181412 159516
rect 187292 159236 187348 172682
rect 188972 165620 189028 276332
rect 189420 275878 189476 276444
rect 189532 276598 189588 276608
rect 189532 276388 189588 276542
rect 189532 276322 189588 276332
rect 189420 275822 189588 275878
rect 189420 275604 189476 275614
rect 189420 268498 189476 275548
rect 189420 268432 189476 268442
rect 188972 165554 189028 165564
rect 189084 264180 189140 264190
rect 189084 168778 189140 264124
rect 189532 173068 189588 275822
rect 189084 160692 189140 168722
rect 189420 173012 189588 173068
rect 189738 274350 190358 281298
rect 189738 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 190358 274350
rect 189738 274226 190358 274294
rect 189738 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 190358 274226
rect 189738 274102 190358 274170
rect 189738 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 190358 274102
rect 189738 273978 190358 274046
rect 189738 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 190358 273978
rect 189738 256350 190358 273922
rect 190428 275604 190484 275614
rect 190428 266878 190484 275548
rect 190428 266812 190484 266822
rect 189738 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 190358 256350
rect 189738 256226 190358 256294
rect 189738 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 190358 256226
rect 189738 256102 190358 256170
rect 189738 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 190358 256102
rect 189738 255978 190358 256046
rect 189738 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 190358 255978
rect 189738 238350 190358 255922
rect 189738 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 190358 238350
rect 189738 238226 190358 238294
rect 189738 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 190358 238226
rect 189738 238102 190358 238170
rect 189738 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 190358 238102
rect 189738 237978 190358 238046
rect 189738 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 190358 237978
rect 189738 220350 190358 237922
rect 189738 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 190358 220350
rect 189738 220226 190358 220294
rect 189738 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 190358 220226
rect 189738 220102 190358 220170
rect 189738 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 190358 220102
rect 189738 219978 190358 220046
rect 189738 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 190358 219978
rect 189738 202350 190358 219922
rect 189738 202294 189834 202350
rect 189890 202294 189958 202350
rect 190014 202294 190082 202350
rect 190138 202294 190206 202350
rect 190262 202294 190358 202350
rect 189738 202226 190358 202294
rect 189738 202170 189834 202226
rect 189890 202170 189958 202226
rect 190014 202170 190082 202226
rect 190138 202170 190206 202226
rect 190262 202170 190358 202226
rect 189738 202102 190358 202170
rect 189738 202046 189834 202102
rect 189890 202046 189958 202102
rect 190014 202046 190082 202102
rect 190138 202046 190206 202102
rect 190262 202046 190358 202102
rect 189738 201978 190358 202046
rect 189738 201922 189834 201978
rect 189890 201922 189958 201978
rect 190014 201922 190082 201978
rect 190138 201922 190206 201978
rect 190262 201922 190358 201978
rect 189738 184350 190358 201922
rect 189738 184294 189834 184350
rect 189890 184294 189958 184350
rect 190014 184294 190082 184350
rect 190138 184294 190206 184350
rect 190262 184294 190358 184350
rect 189738 184226 190358 184294
rect 189738 184170 189834 184226
rect 189890 184170 189958 184226
rect 190014 184170 190082 184226
rect 190138 184170 190206 184226
rect 190262 184170 190358 184226
rect 189738 184102 190358 184170
rect 189738 184046 189834 184102
rect 189890 184046 189958 184102
rect 190014 184046 190082 184102
rect 190138 184046 190206 184102
rect 190262 184046 190358 184102
rect 189738 183978 190358 184046
rect 189738 183922 189834 183978
rect 189890 183922 189958 183978
rect 190014 183922 190082 183978
rect 190138 183922 190206 183978
rect 190262 183922 190358 183978
rect 189420 164500 189476 173012
rect 189738 166350 190358 183922
rect 189738 166294 189834 166350
rect 189890 166294 189958 166350
rect 190014 166294 190082 166350
rect 190138 166294 190206 166350
rect 190262 166294 190358 166350
rect 189738 166226 190358 166294
rect 189738 166170 189834 166226
rect 189890 166170 189958 166226
rect 190014 166170 190082 166226
rect 190138 166170 190206 166226
rect 190262 166170 190358 166226
rect 189738 166102 190358 166170
rect 189738 166046 189834 166102
rect 189890 166046 189958 166102
rect 190014 166046 190082 166102
rect 190138 166046 190206 166102
rect 190262 166046 190358 166102
rect 189738 165978 190358 166046
rect 189738 165922 189834 165978
rect 189890 165922 189958 165978
rect 190014 165922 190082 165978
rect 190138 165922 190206 165978
rect 190262 165922 190358 165978
rect 189532 165620 189588 165630
rect 189532 164948 189588 165564
rect 189532 164882 189588 164892
rect 189420 164434 189476 164444
rect 189084 160626 189140 160636
rect 187292 159170 187348 159180
rect 181356 157938 181412 157948
rect 162738 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 163358 154350
rect 162738 154226 163358 154294
rect 162738 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 163358 154226
rect 162738 154102 163358 154170
rect 162738 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 163358 154102
rect 162738 153978 163358 154046
rect 162738 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 163358 153978
rect 162738 136350 163358 153922
rect 162738 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 163358 136350
rect 162738 136226 163358 136294
rect 162738 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 163358 136226
rect 162738 136102 163358 136170
rect 162738 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 163358 136102
rect 162738 135978 163358 136046
rect 162738 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 163358 135978
rect 162738 118350 163358 135922
rect 162738 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 163358 118350
rect 162738 118226 163358 118294
rect 162738 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 163358 118226
rect 162738 118102 163358 118170
rect 162738 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 163358 118102
rect 162738 117978 163358 118046
rect 162738 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 163358 117978
rect 162738 100350 163358 117922
rect 162738 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 163358 100350
rect 162738 100226 163358 100294
rect 162738 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 163358 100226
rect 162738 100102 163358 100170
rect 162738 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 163358 100102
rect 162738 99978 163358 100046
rect 162738 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99922 163358 99978
rect 162738 82350 163358 99922
rect 162738 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 163358 82350
rect 162738 82226 163358 82294
rect 162738 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 163358 82226
rect 162738 82102 163358 82170
rect 162738 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 163358 82102
rect 162738 81978 163358 82046
rect 162738 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 163358 81978
rect 162738 64350 163358 81922
rect 162738 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 163358 64350
rect 162738 64226 163358 64294
rect 162738 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 163358 64226
rect 162738 64102 163358 64170
rect 162738 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 163358 64102
rect 162738 63978 163358 64046
rect 162738 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 163358 63978
rect 162738 46350 163358 63922
rect 162738 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 163358 46350
rect 162738 46226 163358 46294
rect 162738 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 163358 46226
rect 162738 46102 163358 46170
rect 162738 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 163358 46102
rect 162738 45978 163358 46046
rect 162738 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 163358 45978
rect 162738 28350 163358 45922
rect 162738 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 163358 28350
rect 162738 28226 163358 28294
rect 162738 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 163358 28226
rect 162738 28102 163358 28170
rect 162738 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 163358 28102
rect 162738 27978 163358 28046
rect 162738 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 163358 27978
rect 162738 10350 163358 27922
rect 162738 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 163358 10350
rect 162738 10226 163358 10294
rect 162738 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 163358 10226
rect 162738 10102 163358 10170
rect 162738 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 163358 10102
rect 162738 9978 163358 10046
rect 162738 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 163358 9978
rect 162738 -1120 163358 9922
rect 162738 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 163358 -1120
rect 162738 -1244 163358 -1176
rect 162738 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 163358 -1244
rect 162738 -1368 163358 -1300
rect 162738 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 163358 -1368
rect 162738 -1492 163358 -1424
rect 162738 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 163358 -1492
rect 162738 -1644 163358 -1548
rect 189738 148350 190358 165922
rect 192332 225118 192388 225128
rect 192332 223498 192388 225062
rect 192332 165620 192388 223442
rect 192892 184828 192948 359522
rect 193004 359492 193060 359502
rect 193004 357418 193060 359436
rect 193004 357352 193060 357362
rect 193116 282178 193172 282188
rect 192892 184772 193060 184828
rect 192332 165554 192388 165564
rect 191548 156212 191604 156222
rect 191548 155316 191604 156156
rect 191548 155250 191604 155260
rect 193004 155316 193060 184772
rect 193004 155250 193060 155260
rect 193116 152852 193172 282122
rect 193340 278628 193396 362124
rect 193458 358958 194078 369922
rect 194908 370132 194964 370142
rect 194572 363076 194628 363086
rect 194236 359604 194292 359614
rect 193340 278562 193396 278572
rect 193458 280350 194078 281298
rect 193458 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 194078 280350
rect 193458 280226 194078 280294
rect 193458 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 194078 280226
rect 193458 280102 194078 280170
rect 193458 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 194078 280102
rect 193458 279978 194078 280046
rect 193458 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 194078 279978
rect 193116 152786 193172 152796
rect 193458 262350 194078 279922
rect 193458 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 194078 262350
rect 193458 262226 194078 262294
rect 193458 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 194078 262226
rect 193458 262102 194078 262170
rect 193458 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 194078 262102
rect 193458 261978 194078 262046
rect 193458 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 194078 261978
rect 193458 244350 194078 261922
rect 193458 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 194078 244350
rect 193458 244226 194078 244294
rect 193458 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 194078 244226
rect 193458 244102 194078 244170
rect 193458 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 194078 244102
rect 193458 243978 194078 244046
rect 193458 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 194078 243978
rect 193458 226350 194078 243922
rect 193458 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 194078 226350
rect 193458 226226 194078 226294
rect 193458 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 194078 226226
rect 193458 226102 194078 226170
rect 193458 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 194078 226102
rect 193458 225978 194078 226046
rect 193458 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 194078 225978
rect 193458 208350 194078 225922
rect 193458 208294 193554 208350
rect 193610 208294 193678 208350
rect 193734 208294 193802 208350
rect 193858 208294 193926 208350
rect 193982 208294 194078 208350
rect 193458 208226 194078 208294
rect 193458 208170 193554 208226
rect 193610 208170 193678 208226
rect 193734 208170 193802 208226
rect 193858 208170 193926 208226
rect 193982 208170 194078 208226
rect 193458 208102 194078 208170
rect 193458 208046 193554 208102
rect 193610 208046 193678 208102
rect 193734 208046 193802 208102
rect 193858 208046 193926 208102
rect 193982 208046 194078 208102
rect 193458 207978 194078 208046
rect 193458 207922 193554 207978
rect 193610 207922 193678 207978
rect 193734 207922 193802 207978
rect 193858 207922 193926 207978
rect 193982 207922 194078 207978
rect 193458 190350 194078 207922
rect 193458 190294 193554 190350
rect 193610 190294 193678 190350
rect 193734 190294 193802 190350
rect 193858 190294 193926 190350
rect 193982 190294 194078 190350
rect 193458 190226 194078 190294
rect 193458 190170 193554 190226
rect 193610 190170 193678 190226
rect 193734 190170 193802 190226
rect 193858 190170 193926 190226
rect 193982 190170 194078 190226
rect 193458 190102 194078 190170
rect 193458 190046 193554 190102
rect 193610 190046 193678 190102
rect 193734 190046 193802 190102
rect 193858 190046 193926 190102
rect 193982 190046 194078 190102
rect 193458 189978 194078 190046
rect 193458 189922 193554 189978
rect 193610 189922 193678 189978
rect 193734 189922 193802 189978
rect 193858 189922 193926 189978
rect 193982 189922 194078 189978
rect 193458 172350 194078 189922
rect 193458 172294 193554 172350
rect 193610 172294 193678 172350
rect 193734 172294 193802 172350
rect 193858 172294 193926 172350
rect 193982 172294 194078 172350
rect 193458 172226 194078 172294
rect 193458 172170 193554 172226
rect 193610 172170 193678 172226
rect 193734 172170 193802 172226
rect 193858 172170 193926 172226
rect 193982 172170 194078 172226
rect 193458 172102 194078 172170
rect 193458 172046 193554 172102
rect 193610 172046 193678 172102
rect 193734 172046 193802 172102
rect 193858 172046 193926 172102
rect 193982 172046 194078 172102
rect 193458 171978 194078 172046
rect 193458 171922 193554 171978
rect 193610 171922 193678 171978
rect 193734 171922 193802 171978
rect 193858 171922 193926 171978
rect 193982 171922 194078 171978
rect 193458 154350 194078 171922
rect 193458 154294 193554 154350
rect 193610 154294 193678 154350
rect 193734 154294 193802 154350
rect 193858 154294 193926 154350
rect 193982 154294 194078 154350
rect 193458 154226 194078 154294
rect 193458 154170 193554 154226
rect 193610 154170 193678 154226
rect 193734 154170 193802 154226
rect 193858 154170 193926 154226
rect 193982 154170 194078 154226
rect 193458 154102 194078 154170
rect 193458 154046 193554 154102
rect 193610 154046 193678 154102
rect 193734 154046 193802 154102
rect 193858 154046 193926 154102
rect 193982 154046 194078 154102
rect 193458 153978 194078 154046
rect 193458 153922 193554 153978
rect 193610 153922 193678 153978
rect 193734 153922 193802 153978
rect 193858 153922 193926 153978
rect 193982 153922 194078 153978
rect 189738 148294 189834 148350
rect 189890 148294 189958 148350
rect 190014 148294 190082 148350
rect 190138 148294 190206 148350
rect 190262 148294 190358 148350
rect 189738 148226 190358 148294
rect 189738 148170 189834 148226
rect 189890 148170 189958 148226
rect 190014 148170 190082 148226
rect 190138 148170 190206 148226
rect 190262 148170 190358 148226
rect 189738 148102 190358 148170
rect 189738 148046 189834 148102
rect 189890 148046 189958 148102
rect 190014 148046 190082 148102
rect 190138 148046 190206 148102
rect 190262 148046 190358 148102
rect 189738 147978 190358 148046
rect 189738 147922 189834 147978
rect 189890 147922 189958 147978
rect 190014 147922 190082 147978
rect 190138 147922 190206 147978
rect 190262 147922 190358 147978
rect 189738 130350 190358 147922
rect 189738 130294 189834 130350
rect 189890 130294 189958 130350
rect 190014 130294 190082 130350
rect 190138 130294 190206 130350
rect 190262 130294 190358 130350
rect 189738 130226 190358 130294
rect 189738 130170 189834 130226
rect 189890 130170 189958 130226
rect 190014 130170 190082 130226
rect 190138 130170 190206 130226
rect 190262 130170 190358 130226
rect 189738 130102 190358 130170
rect 189738 130046 189834 130102
rect 189890 130046 189958 130102
rect 190014 130046 190082 130102
rect 190138 130046 190206 130102
rect 190262 130046 190358 130102
rect 189738 129978 190358 130046
rect 189738 129922 189834 129978
rect 189890 129922 189958 129978
rect 190014 129922 190082 129978
rect 190138 129922 190206 129978
rect 190262 129922 190358 129978
rect 189738 112350 190358 129922
rect 189738 112294 189834 112350
rect 189890 112294 189958 112350
rect 190014 112294 190082 112350
rect 190138 112294 190206 112350
rect 190262 112294 190358 112350
rect 189738 112226 190358 112294
rect 189738 112170 189834 112226
rect 189890 112170 189958 112226
rect 190014 112170 190082 112226
rect 190138 112170 190206 112226
rect 190262 112170 190358 112226
rect 189738 112102 190358 112170
rect 189738 112046 189834 112102
rect 189890 112046 189958 112102
rect 190014 112046 190082 112102
rect 190138 112046 190206 112102
rect 190262 112046 190358 112102
rect 189738 111978 190358 112046
rect 189738 111922 189834 111978
rect 189890 111922 189958 111978
rect 190014 111922 190082 111978
rect 190138 111922 190206 111978
rect 190262 111922 190358 111978
rect 189738 94350 190358 111922
rect 189738 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 190358 94350
rect 189738 94226 190358 94294
rect 189738 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 190358 94226
rect 189738 94102 190358 94170
rect 189738 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 190358 94102
rect 189738 93978 190358 94046
rect 189738 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 190358 93978
rect 189738 76350 190358 93922
rect 189738 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 190358 76350
rect 189738 76226 190358 76294
rect 189738 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 190358 76226
rect 189738 76102 190358 76170
rect 189738 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 190358 76102
rect 189738 75978 190358 76046
rect 189738 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 190358 75978
rect 189738 58350 190358 75922
rect 189738 58294 189834 58350
rect 189890 58294 189958 58350
rect 190014 58294 190082 58350
rect 190138 58294 190206 58350
rect 190262 58294 190358 58350
rect 189738 58226 190358 58294
rect 189738 58170 189834 58226
rect 189890 58170 189958 58226
rect 190014 58170 190082 58226
rect 190138 58170 190206 58226
rect 190262 58170 190358 58226
rect 189738 58102 190358 58170
rect 189738 58046 189834 58102
rect 189890 58046 189958 58102
rect 190014 58046 190082 58102
rect 190138 58046 190206 58102
rect 190262 58046 190358 58102
rect 189738 57978 190358 58046
rect 189738 57922 189834 57978
rect 189890 57922 189958 57978
rect 190014 57922 190082 57978
rect 190138 57922 190206 57978
rect 190262 57922 190358 57978
rect 189738 40350 190358 57922
rect 189738 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 190358 40350
rect 189738 40226 190358 40294
rect 189738 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 190358 40226
rect 189738 40102 190358 40170
rect 189738 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 190358 40102
rect 189738 39978 190358 40046
rect 189738 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 190358 39978
rect 189738 22350 190358 39922
rect 189738 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 190358 22350
rect 189738 22226 190358 22294
rect 189738 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 190358 22226
rect 189738 22102 190358 22170
rect 189738 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 190358 22102
rect 189738 21978 190358 22046
rect 189738 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 190358 21978
rect 189738 4350 190358 21922
rect 189738 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 190358 4350
rect 189738 4226 190358 4294
rect 189738 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 190358 4226
rect 189738 4102 190358 4170
rect 189738 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 190358 4102
rect 189738 3978 190358 4046
rect 189738 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 190358 3978
rect 189738 -160 190358 3922
rect 189738 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 190358 -160
rect 189738 -284 190358 -216
rect 189738 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 190358 -284
rect 189738 -408 190358 -340
rect 189738 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 190358 -408
rect 189738 -532 190358 -464
rect 189738 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 190358 -532
rect 189738 -1644 190358 -588
rect 193458 136350 194078 153922
rect 194236 148708 194292 359548
rect 194348 359492 194404 359502
rect 194348 349468 194404 359436
rect 194348 349412 194516 349468
rect 194348 296758 194404 296768
rect 194348 271348 194404 296702
rect 194348 271282 194404 271292
rect 194460 149492 194516 349412
rect 194572 280532 194628 363020
rect 194796 360298 194852 360308
rect 194684 360164 194740 360174
rect 194684 282178 194740 360108
rect 194684 282112 194740 282122
rect 194572 280466 194628 280476
rect 194796 280084 194852 360242
rect 194796 280018 194852 280028
rect 194572 270118 194628 270154
rect 194572 270050 194628 270060
rect 194460 148820 194516 149436
rect 194460 148754 194516 148764
rect 194236 148642 194292 148652
rect 194908 148260 194964 370076
rect 195020 366436 195076 366446
rect 195020 280420 195076 366380
rect 195916 359758 195972 359768
rect 195692 359604 195748 359614
rect 195232 346350 195552 346384
rect 195232 346294 195302 346350
rect 195358 346294 195426 346350
rect 195482 346294 195552 346350
rect 195232 346226 195552 346294
rect 195232 346170 195302 346226
rect 195358 346170 195426 346226
rect 195482 346170 195552 346226
rect 195232 346102 195552 346170
rect 195232 346046 195302 346102
rect 195358 346046 195426 346102
rect 195482 346046 195552 346102
rect 195232 345978 195552 346046
rect 195232 345922 195302 345978
rect 195358 345922 195426 345978
rect 195482 345922 195552 345978
rect 195232 345888 195552 345922
rect 195232 328350 195552 328384
rect 195232 328294 195302 328350
rect 195358 328294 195426 328350
rect 195482 328294 195552 328350
rect 195232 328226 195552 328294
rect 195232 328170 195302 328226
rect 195358 328170 195426 328226
rect 195482 328170 195552 328226
rect 195232 328102 195552 328170
rect 195232 328046 195302 328102
rect 195358 328046 195426 328102
rect 195482 328046 195552 328102
rect 195232 327978 195552 328046
rect 195232 327922 195302 327978
rect 195358 327922 195426 327978
rect 195482 327922 195552 327978
rect 195232 327888 195552 327922
rect 195232 310350 195552 310384
rect 195232 310294 195302 310350
rect 195358 310294 195426 310350
rect 195482 310294 195552 310350
rect 195232 310226 195552 310294
rect 195232 310170 195302 310226
rect 195358 310170 195426 310226
rect 195482 310170 195552 310226
rect 195232 310102 195552 310170
rect 195232 310046 195302 310102
rect 195358 310046 195426 310102
rect 195482 310046 195552 310102
rect 195232 309978 195552 310046
rect 195232 309922 195302 309978
rect 195358 309922 195426 309978
rect 195482 309922 195552 309978
rect 195232 309888 195552 309922
rect 195232 292350 195552 292384
rect 195232 292294 195302 292350
rect 195358 292294 195426 292350
rect 195482 292294 195552 292350
rect 195232 292226 195552 292294
rect 195232 292170 195302 292226
rect 195358 292170 195426 292226
rect 195482 292170 195552 292226
rect 195232 292102 195552 292170
rect 195232 292046 195302 292102
rect 195358 292046 195426 292102
rect 195482 292046 195552 292102
rect 195232 291978 195552 292046
rect 195232 291922 195302 291978
rect 195358 291922 195426 291978
rect 195482 291922 195552 291978
rect 195232 291888 195552 291922
rect 195020 280354 195076 280364
rect 195692 149380 195748 359548
rect 195804 296398 195860 296408
rect 195804 162932 195860 296342
rect 195916 277060 195972 359702
rect 196476 359578 196532 359588
rect 196476 357598 196532 359522
rect 196476 357532 196532 357542
rect 196588 277172 196644 370188
rect 196700 363412 196756 363422
rect 196700 278404 196756 363356
rect 197372 360612 197428 360622
rect 197372 359604 197428 360556
rect 197372 359538 197428 359548
rect 196700 278338 196756 278348
rect 197372 336358 197428 336368
rect 196588 277106 196644 277116
rect 195916 276994 195972 277004
rect 197036 276164 197092 276174
rect 197036 273358 197092 276108
rect 197036 273292 197092 273302
rect 197372 270004 197428 336302
rect 197372 269938 197428 269948
rect 197484 330238 197540 330248
rect 197484 266532 197540 330182
rect 197596 317818 197652 317828
rect 197596 278180 197652 317762
rect 197596 278114 197652 278124
rect 197708 275604 197764 371756
rect 199500 368676 199556 368686
rect 199276 359578 199332 359588
rect 199276 357700 199332 359522
rect 199276 357634 199332 357644
rect 199388 357958 199444 357968
rect 199276 357238 199332 357248
rect 199276 357140 199332 357182
rect 199276 357074 199332 357084
rect 199388 356020 199444 357902
rect 199388 355954 199444 355964
rect 199276 336420 199332 336430
rect 199276 336358 199332 336364
rect 199276 336292 199332 336302
rect 199276 330260 199332 330270
rect 199276 330166 199332 330182
rect 199276 325220 199332 325230
rect 199276 317998 199332 325164
rect 199164 317942 199332 317998
rect 199388 324100 199444 324110
rect 199164 314188 199220 317942
rect 199276 317828 199332 317838
rect 199276 317734 199332 317762
rect 199164 314132 199332 314188
rect 198156 305758 198212 305768
rect 197708 275538 197764 275548
rect 197820 287578 197876 287588
rect 197484 266466 197540 266476
rect 197820 265078 197876 287522
rect 198156 280532 198212 305702
rect 199276 301252 199332 314132
rect 199276 301186 199332 301196
rect 199276 300580 199332 300590
rect 199276 297478 199332 300524
rect 198716 297422 199332 297478
rect 198716 294028 198772 297422
rect 199276 296772 199332 296782
rect 199276 296678 199332 296702
rect 199276 296436 199332 296446
rect 199276 294028 199332 296380
rect 198716 293972 198884 294028
rect 198828 287218 198884 293972
rect 199164 293972 199332 294028
rect 199164 287218 199220 293972
rect 199276 287588 199332 287598
rect 199276 287494 199332 287522
rect 198828 287162 199108 287218
rect 199164 287162 199332 287218
rect 198156 280466 198212 280476
rect 199052 274820 199108 287162
rect 199052 274754 199108 274764
rect 197820 265012 197876 265022
rect 198418 256350 198894 256384
rect 198418 256294 198442 256350
rect 198498 256294 198566 256350
rect 198622 256294 198690 256350
rect 198746 256294 198814 256350
rect 198870 256294 198894 256350
rect 198418 256226 198894 256294
rect 198418 256170 198442 256226
rect 198498 256170 198566 256226
rect 198622 256170 198690 256226
rect 198746 256170 198814 256226
rect 198870 256170 198894 256226
rect 198418 256102 198894 256170
rect 198418 256046 198442 256102
rect 198498 256046 198566 256102
rect 198622 256046 198690 256102
rect 198746 256046 198814 256102
rect 198870 256046 198894 256102
rect 198418 255978 198894 256046
rect 198418 255922 198442 255978
rect 198498 255922 198566 255978
rect 198622 255922 198690 255978
rect 198746 255922 198814 255978
rect 198870 255922 198894 255978
rect 198418 255888 198894 255922
rect 197618 244350 198094 244384
rect 197618 244294 197642 244350
rect 197698 244294 197766 244350
rect 197822 244294 197890 244350
rect 197946 244294 198014 244350
rect 198070 244294 198094 244350
rect 197618 244226 198094 244294
rect 197618 244170 197642 244226
rect 197698 244170 197766 244226
rect 197822 244170 197890 244226
rect 197946 244170 198014 244226
rect 198070 244170 198094 244226
rect 197618 244102 198094 244170
rect 197618 244046 197642 244102
rect 197698 244046 197766 244102
rect 197822 244046 197890 244102
rect 197946 244046 198014 244102
rect 198070 244046 198094 244102
rect 197618 243978 198094 244046
rect 197618 243922 197642 243978
rect 197698 243922 197766 243978
rect 197822 243922 197890 243978
rect 197946 243922 198014 243978
rect 198070 243922 198094 243978
rect 197618 243888 198094 243922
rect 198418 238350 198894 238384
rect 198418 238294 198442 238350
rect 198498 238294 198566 238350
rect 198622 238294 198690 238350
rect 198746 238294 198814 238350
rect 198870 238294 198894 238350
rect 198418 238226 198894 238294
rect 198418 238170 198442 238226
rect 198498 238170 198566 238226
rect 198622 238170 198690 238226
rect 198746 238170 198814 238226
rect 198870 238170 198894 238226
rect 198418 238102 198894 238170
rect 198418 238046 198442 238102
rect 198498 238046 198566 238102
rect 198622 238046 198690 238102
rect 198746 238046 198814 238102
rect 198870 238046 198894 238102
rect 198418 237978 198894 238046
rect 198418 237922 198442 237978
rect 198498 237922 198566 237978
rect 198622 237922 198690 237978
rect 198746 237922 198814 237978
rect 198870 237922 198894 237978
rect 198418 237888 198894 237922
rect 197618 226350 198094 226384
rect 197618 226294 197642 226350
rect 197698 226294 197766 226350
rect 197822 226294 197890 226350
rect 197946 226294 198014 226350
rect 198070 226294 198094 226350
rect 197618 226226 198094 226294
rect 197618 226170 197642 226226
rect 197698 226170 197766 226226
rect 197822 226170 197890 226226
rect 197946 226170 198014 226226
rect 198070 226170 198094 226226
rect 197618 226102 198094 226170
rect 197618 226046 197642 226102
rect 197698 226046 197766 226102
rect 197822 226046 197890 226102
rect 197946 226046 198014 226102
rect 198070 226046 198094 226102
rect 197618 225978 198094 226046
rect 197618 225922 197642 225978
rect 197698 225922 197766 225978
rect 197822 225922 197890 225978
rect 197946 225922 198014 225978
rect 198070 225922 198094 225978
rect 197618 225888 198094 225922
rect 198418 220350 198894 220384
rect 198418 220294 198442 220350
rect 198498 220294 198566 220350
rect 198622 220294 198690 220350
rect 198746 220294 198814 220350
rect 198870 220294 198894 220350
rect 198418 220226 198894 220294
rect 198418 220170 198442 220226
rect 198498 220170 198566 220226
rect 198622 220170 198690 220226
rect 198746 220170 198814 220226
rect 198870 220170 198894 220226
rect 198418 220102 198894 220170
rect 198418 220046 198442 220102
rect 198498 220046 198566 220102
rect 198622 220046 198690 220102
rect 198746 220046 198814 220102
rect 198870 220046 198894 220102
rect 198418 219978 198894 220046
rect 198418 219922 198442 219978
rect 198498 219922 198566 219978
rect 198622 219922 198690 219978
rect 198746 219922 198814 219978
rect 198870 219922 198894 219978
rect 198418 219888 198894 219922
rect 197618 208350 198094 208384
rect 197618 208294 197642 208350
rect 197698 208294 197766 208350
rect 197822 208294 197890 208350
rect 197946 208294 198014 208350
rect 198070 208294 198094 208350
rect 197618 208226 198094 208294
rect 197618 208170 197642 208226
rect 197698 208170 197766 208226
rect 197822 208170 197890 208226
rect 197946 208170 198014 208226
rect 198070 208170 198094 208226
rect 197618 208102 198094 208170
rect 197618 208046 197642 208102
rect 197698 208046 197766 208102
rect 197822 208046 197890 208102
rect 197946 208046 198014 208102
rect 198070 208046 198094 208102
rect 197618 207978 198094 208046
rect 197618 207922 197642 207978
rect 197698 207922 197766 207978
rect 197822 207922 197890 207978
rect 197946 207922 198014 207978
rect 198070 207922 198094 207978
rect 197618 207888 198094 207922
rect 198418 202350 198894 202384
rect 198418 202294 198442 202350
rect 198498 202294 198566 202350
rect 198622 202294 198690 202350
rect 198746 202294 198814 202350
rect 198870 202294 198894 202350
rect 198418 202226 198894 202294
rect 198418 202170 198442 202226
rect 198498 202170 198566 202226
rect 198622 202170 198690 202226
rect 198746 202170 198814 202226
rect 198870 202170 198894 202226
rect 198418 202102 198894 202170
rect 198418 202046 198442 202102
rect 198498 202046 198566 202102
rect 198622 202046 198690 202102
rect 198746 202046 198814 202102
rect 198870 202046 198894 202102
rect 198418 201978 198894 202046
rect 198418 201922 198442 201978
rect 198498 201922 198566 201978
rect 198622 201922 198690 201978
rect 198746 201922 198814 201978
rect 198870 201922 198894 201978
rect 198418 201888 198894 201922
rect 197618 190350 198094 190384
rect 197618 190294 197642 190350
rect 197698 190294 197766 190350
rect 197822 190294 197890 190350
rect 197946 190294 198014 190350
rect 198070 190294 198094 190350
rect 197618 190226 198094 190294
rect 197618 190170 197642 190226
rect 197698 190170 197766 190226
rect 197822 190170 197890 190226
rect 197946 190170 198014 190226
rect 198070 190170 198094 190226
rect 197618 190102 198094 190170
rect 197618 190046 197642 190102
rect 197698 190046 197766 190102
rect 197822 190046 197890 190102
rect 197946 190046 198014 190102
rect 198070 190046 198094 190102
rect 197618 189978 198094 190046
rect 197618 189922 197642 189978
rect 197698 189922 197766 189978
rect 197822 189922 197890 189978
rect 197946 189922 198014 189978
rect 198070 189922 198094 189978
rect 197618 189888 198094 189922
rect 198418 184350 198894 184384
rect 198418 184294 198442 184350
rect 198498 184294 198566 184350
rect 198622 184294 198690 184350
rect 198746 184294 198814 184350
rect 198870 184294 198894 184350
rect 198418 184226 198894 184294
rect 198418 184170 198442 184226
rect 198498 184170 198566 184226
rect 198622 184170 198690 184226
rect 198746 184170 198814 184226
rect 198870 184170 198894 184226
rect 198418 184102 198894 184170
rect 198418 184046 198442 184102
rect 198498 184046 198566 184102
rect 198622 184046 198690 184102
rect 198746 184046 198814 184102
rect 198870 184046 198894 184102
rect 198418 183978 198894 184046
rect 198418 183922 198442 183978
rect 198498 183922 198566 183978
rect 198622 183922 198690 183978
rect 198746 183922 198814 183978
rect 198870 183922 198894 183978
rect 198418 183888 198894 183922
rect 197618 172350 198094 172384
rect 197618 172294 197642 172350
rect 197698 172294 197766 172350
rect 197822 172294 197890 172350
rect 197946 172294 198014 172350
rect 198070 172294 198094 172350
rect 197618 172226 198094 172294
rect 197618 172170 197642 172226
rect 197698 172170 197766 172226
rect 197822 172170 197890 172226
rect 197946 172170 198014 172226
rect 198070 172170 198094 172226
rect 197618 172102 198094 172170
rect 197618 172046 197642 172102
rect 197698 172046 197766 172102
rect 197822 172046 197890 172102
rect 197946 172046 198014 172102
rect 198070 172046 198094 172102
rect 197618 171978 198094 172046
rect 197618 171922 197642 171978
rect 197698 171922 197766 171978
rect 197822 171922 197890 171978
rect 197946 171922 198014 171978
rect 198070 171922 198094 171978
rect 197618 171888 198094 171922
rect 199164 164388 199220 164398
rect 199164 163558 199220 164332
rect 199276 163940 199332 287162
rect 199388 164612 199444 324044
rect 199388 164546 199444 164556
rect 199276 163874 199332 163884
rect 199164 163502 199332 163558
rect 195804 162866 195860 162876
rect 199276 163044 199332 163502
rect 199276 161364 199332 162988
rect 199276 161298 199332 161308
rect 199500 149548 199556 368620
rect 199724 364644 199780 364654
rect 199612 315140 199668 315150
rect 199612 266420 199668 315084
rect 199724 275828 199780 364588
rect 199836 305758 199892 587132
rect 199948 362180 200004 590716
rect 220458 580350 221078 596784
rect 220458 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 221078 580350
rect 220458 580226 221078 580294
rect 220458 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 221078 580226
rect 220458 580102 221078 580170
rect 220458 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 221078 580102
rect 220458 579978 221078 580046
rect 220458 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 221078 579978
rect 220458 562350 221078 579922
rect 220458 562294 220554 562350
rect 220610 562294 220678 562350
rect 220734 562294 220802 562350
rect 220858 562294 220926 562350
rect 220982 562294 221078 562350
rect 220458 562226 221078 562294
rect 220458 562170 220554 562226
rect 220610 562170 220678 562226
rect 220734 562170 220802 562226
rect 220858 562170 220926 562226
rect 220982 562170 221078 562226
rect 220458 562102 221078 562170
rect 220458 562046 220554 562102
rect 220610 562046 220678 562102
rect 220734 562046 220802 562102
rect 220858 562046 220926 562102
rect 220982 562046 221078 562102
rect 220458 561978 221078 562046
rect 220458 561922 220554 561978
rect 220610 561922 220678 561978
rect 220734 561922 220802 561978
rect 220858 561922 220926 561978
rect 220982 561922 221078 561978
rect 220458 544350 221078 561922
rect 220458 544294 220554 544350
rect 220610 544294 220678 544350
rect 220734 544294 220802 544350
rect 220858 544294 220926 544350
rect 220982 544294 221078 544350
rect 220458 544226 221078 544294
rect 220458 544170 220554 544226
rect 220610 544170 220678 544226
rect 220734 544170 220802 544226
rect 220858 544170 220926 544226
rect 220982 544170 221078 544226
rect 220458 544102 221078 544170
rect 220458 544046 220554 544102
rect 220610 544046 220678 544102
rect 220734 544046 220802 544102
rect 220858 544046 220926 544102
rect 220982 544046 221078 544102
rect 220458 543978 221078 544046
rect 220458 543922 220554 543978
rect 220610 543922 220678 543978
rect 220734 543922 220802 543978
rect 220858 543922 220926 543978
rect 220982 543922 221078 543978
rect 220458 526350 221078 543922
rect 220458 526294 220554 526350
rect 220610 526294 220678 526350
rect 220734 526294 220802 526350
rect 220858 526294 220926 526350
rect 220982 526294 221078 526350
rect 220458 526226 221078 526294
rect 220458 526170 220554 526226
rect 220610 526170 220678 526226
rect 220734 526170 220802 526226
rect 220858 526170 220926 526226
rect 220982 526170 221078 526226
rect 220458 526102 221078 526170
rect 220458 526046 220554 526102
rect 220610 526046 220678 526102
rect 220734 526046 220802 526102
rect 220858 526046 220926 526102
rect 220982 526046 221078 526102
rect 220458 525978 221078 526046
rect 220458 525922 220554 525978
rect 220610 525922 220678 525978
rect 220734 525922 220802 525978
rect 220858 525922 220926 525978
rect 220982 525922 221078 525978
rect 200060 511588 200116 511598
rect 200060 364588 200116 511532
rect 220458 508350 221078 525922
rect 220458 508294 220554 508350
rect 220610 508294 220678 508350
rect 220734 508294 220802 508350
rect 220858 508294 220926 508350
rect 220982 508294 221078 508350
rect 220458 508226 221078 508294
rect 220458 508170 220554 508226
rect 220610 508170 220678 508226
rect 220734 508170 220802 508226
rect 220858 508170 220926 508226
rect 220982 508170 221078 508226
rect 220458 508102 221078 508170
rect 220458 508046 220554 508102
rect 220610 508046 220678 508102
rect 220734 508046 220802 508102
rect 220858 508046 220926 508102
rect 220982 508046 221078 508102
rect 220458 507978 221078 508046
rect 220458 507922 220554 507978
rect 220610 507922 220678 507978
rect 220734 507922 220802 507978
rect 220858 507922 220926 507978
rect 220982 507922 221078 507978
rect 220458 490350 221078 507922
rect 220458 490294 220554 490350
rect 220610 490294 220678 490350
rect 220734 490294 220802 490350
rect 220858 490294 220926 490350
rect 220982 490294 221078 490350
rect 220458 490226 221078 490294
rect 220458 490170 220554 490226
rect 220610 490170 220678 490226
rect 220734 490170 220802 490226
rect 220858 490170 220926 490226
rect 220982 490170 221078 490226
rect 220458 490102 221078 490170
rect 220458 490046 220554 490102
rect 220610 490046 220678 490102
rect 220734 490046 220802 490102
rect 220858 490046 220926 490102
rect 220982 490046 221078 490102
rect 220458 489978 221078 490046
rect 220458 489922 220554 489978
rect 220610 489922 220678 489978
rect 220734 489922 220802 489978
rect 220858 489922 220926 489978
rect 220982 489922 221078 489978
rect 220458 472350 221078 489922
rect 220458 472294 220554 472350
rect 220610 472294 220678 472350
rect 220734 472294 220802 472350
rect 220858 472294 220926 472350
rect 220982 472294 221078 472350
rect 220458 472226 221078 472294
rect 220458 472170 220554 472226
rect 220610 472170 220678 472226
rect 220734 472170 220802 472226
rect 220858 472170 220926 472226
rect 220982 472170 221078 472226
rect 220458 472102 221078 472170
rect 220458 472046 220554 472102
rect 220610 472046 220678 472102
rect 220734 472046 220802 472102
rect 220858 472046 220926 472102
rect 220982 472046 221078 472102
rect 220458 471978 221078 472046
rect 220458 471922 220554 471978
rect 220610 471922 220678 471978
rect 220734 471922 220802 471978
rect 220858 471922 220926 471978
rect 220982 471922 221078 471978
rect 220458 454350 221078 471922
rect 220458 454294 220554 454350
rect 220610 454294 220678 454350
rect 220734 454294 220802 454350
rect 220858 454294 220926 454350
rect 220982 454294 221078 454350
rect 220458 454226 221078 454294
rect 220458 454170 220554 454226
rect 220610 454170 220678 454226
rect 220734 454170 220802 454226
rect 220858 454170 220926 454226
rect 220982 454170 221078 454226
rect 220458 454102 221078 454170
rect 220458 454046 220554 454102
rect 220610 454046 220678 454102
rect 220734 454046 220802 454102
rect 220858 454046 220926 454102
rect 220982 454046 221078 454102
rect 220458 453978 221078 454046
rect 220458 453922 220554 453978
rect 220610 453922 220678 453978
rect 220734 453922 220802 453978
rect 220858 453922 220926 453978
rect 220982 453922 221078 453978
rect 220458 436350 221078 453922
rect 220458 436294 220554 436350
rect 220610 436294 220678 436350
rect 220734 436294 220802 436350
rect 220858 436294 220926 436350
rect 220982 436294 221078 436350
rect 220458 436226 221078 436294
rect 220458 436170 220554 436226
rect 220610 436170 220678 436226
rect 220734 436170 220802 436226
rect 220858 436170 220926 436226
rect 220982 436170 221078 436226
rect 220458 436102 221078 436170
rect 220458 436046 220554 436102
rect 220610 436046 220678 436102
rect 220734 436046 220802 436102
rect 220858 436046 220926 436102
rect 220982 436046 221078 436102
rect 220458 435978 221078 436046
rect 220458 435922 220554 435978
rect 220610 435922 220678 435978
rect 220734 435922 220802 435978
rect 220858 435922 220926 435978
rect 220982 435922 221078 435978
rect 220458 418350 221078 435922
rect 220458 418294 220554 418350
rect 220610 418294 220678 418350
rect 220734 418294 220802 418350
rect 220858 418294 220926 418350
rect 220982 418294 221078 418350
rect 220458 418226 221078 418294
rect 220458 418170 220554 418226
rect 220610 418170 220678 418226
rect 220734 418170 220802 418226
rect 220858 418170 220926 418226
rect 220982 418170 221078 418226
rect 220458 418102 221078 418170
rect 220458 418046 220554 418102
rect 220610 418046 220678 418102
rect 220734 418046 220802 418102
rect 220858 418046 220926 418102
rect 220982 418046 221078 418102
rect 220458 417978 221078 418046
rect 220458 417922 220554 417978
rect 220610 417922 220678 417978
rect 220734 417922 220802 417978
rect 220858 417922 220926 417978
rect 220982 417922 221078 417978
rect 220458 400350 221078 417922
rect 220458 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 221078 400350
rect 220458 400226 221078 400294
rect 220458 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 221078 400226
rect 220458 400102 221078 400170
rect 220458 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 221078 400102
rect 220458 399978 221078 400046
rect 220458 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 221078 399978
rect 203420 390628 203476 390638
rect 202412 366778 202468 366788
rect 202076 366598 202132 366608
rect 201852 366418 201908 366428
rect 200060 364532 200452 364588
rect 199948 362114 200004 362124
rect 200284 362180 200340 362190
rect 200060 358708 200116 358718
rect 200060 329308 200116 358652
rect 200284 337708 200340 362124
rect 200396 358708 200452 364532
rect 200396 358642 200452 358652
rect 201852 349860 201908 366362
rect 201852 349794 201908 349804
rect 201964 361378 202020 361388
rect 200060 329242 200116 329252
rect 200172 337652 200340 337708
rect 200620 344260 200676 344270
rect 200172 327178 200228 337652
rect 199836 305692 199892 305702
rect 199948 327122 200228 327178
rect 200284 329252 200340 329262
rect 199724 275762 199780 275772
rect 199836 303940 199892 303950
rect 199836 268436 199892 303884
rect 199948 280756 200004 327122
rect 200284 326998 200340 329196
rect 200284 326942 200452 326998
rect 200396 317548 200452 326942
rect 199948 280690 200004 280700
rect 200060 317492 200452 317548
rect 200060 278852 200116 317492
rect 200060 278786 200116 278796
rect 200172 316260 200228 316270
rect 199836 268370 199892 268380
rect 199612 266354 199668 266364
rect 200172 157332 200228 316204
rect 200508 312900 200564 312910
rect 200172 157266 200228 157276
rect 200284 310660 200340 310670
rect 200284 150500 200340 310604
rect 200396 309540 200452 309550
rect 200396 155428 200452 309484
rect 200508 158788 200564 312844
rect 200620 302428 200676 344204
rect 201964 339780 202020 361322
rect 202076 354340 202132 366542
rect 202076 354274 202132 354284
rect 202188 359578 202244 359588
rect 202188 342020 202244 359522
rect 202188 341954 202244 341964
rect 201964 339714 202020 339724
rect 202076 334180 202132 334190
rect 201964 331940 202020 331950
rect 201852 322980 201908 322990
rect 200620 302372 200788 302428
rect 200732 279748 200788 302372
rect 201852 296398 201908 322924
rect 201852 296332 201908 296342
rect 201852 296100 201908 296110
rect 200732 279682 200788 279692
rect 201740 293860 201796 293870
rect 201740 279658 201796 293804
rect 201740 279592 201796 279602
rect 201516 168778 201572 168794
rect 201516 168690 201572 168700
rect 201852 164052 201908 296044
rect 201964 269780 202020 331884
rect 202076 279478 202132 334124
rect 202300 317380 202356 317390
rect 202076 279412 202132 279422
rect 202188 299460 202244 299470
rect 202188 274618 202244 299404
rect 202188 274552 202244 274562
rect 201964 269714 202020 269724
rect 201852 163986 201908 163996
rect 200508 158722 200564 158732
rect 202300 155540 202356 317324
rect 202412 284788 202468 366722
rect 203308 333060 203364 333070
rect 202412 284722 202468 284732
rect 202524 314020 202580 314030
rect 202412 206612 202468 206622
rect 202412 205138 202468 206556
rect 202412 205072 202468 205082
rect 202300 155474 202356 155484
rect 200396 155362 200452 155372
rect 202524 152068 202580 313964
rect 202636 298340 202692 298350
rect 202636 274708 202692 298284
rect 202636 274642 202692 274652
rect 203308 165732 203364 333004
rect 203420 275940 203476 390572
rect 220458 382350 221078 399922
rect 220458 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 221078 382350
rect 220458 382226 221078 382294
rect 220458 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 221078 382226
rect 220458 382102 221078 382170
rect 220458 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 221078 382102
rect 220458 381978 221078 382046
rect 220458 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 221078 381978
rect 212156 373380 212212 373390
rect 211932 373268 211988 373278
rect 211708 371700 211764 371710
rect 210252 371476 210308 371486
rect 210140 370356 210196 370366
rect 204204 366884 204260 366894
rect 203420 275874 203476 275884
rect 204092 364798 204148 364808
rect 203420 187572 203476 187582
rect 203420 187318 203476 187516
rect 203420 187252 203476 187262
rect 203420 182868 203476 182878
rect 203420 181558 203476 182812
rect 203420 181492 203476 181502
rect 203308 165666 203364 165676
rect 202524 152002 202580 152012
rect 200284 150434 200340 150444
rect 195692 149314 195748 149324
rect 199052 149492 199556 149548
rect 194908 147476 194964 148204
rect 194908 147410 194964 147420
rect 199052 147252 199108 149492
rect 193458 136294 193554 136350
rect 193610 136294 193678 136350
rect 193734 136294 193802 136350
rect 193858 136294 193926 136350
rect 193982 136294 194078 136350
rect 193458 136226 194078 136294
rect 193458 136170 193554 136226
rect 193610 136170 193678 136226
rect 193734 136170 193802 136226
rect 193858 136170 193926 136226
rect 193982 136170 194078 136226
rect 193458 136102 194078 136170
rect 193458 136046 193554 136102
rect 193610 136046 193678 136102
rect 193734 136046 193802 136102
rect 193858 136046 193926 136102
rect 193982 136046 194078 136102
rect 193458 135978 194078 136046
rect 193458 135922 193554 135978
rect 193610 135922 193678 135978
rect 193734 135922 193802 135978
rect 193858 135922 193926 135978
rect 193982 135922 194078 135978
rect 193458 118350 194078 135922
rect 196588 136350 197064 136384
rect 196588 136294 196612 136350
rect 196668 136294 196736 136350
rect 196792 136294 196860 136350
rect 196916 136294 196984 136350
rect 197040 136294 197064 136350
rect 196588 136226 197064 136294
rect 196588 136170 196612 136226
rect 196668 136170 196736 136226
rect 196792 136170 196860 136226
rect 196916 136170 196984 136226
rect 197040 136170 197064 136226
rect 196588 136102 197064 136170
rect 196588 136046 196612 136102
rect 196668 136046 196736 136102
rect 196792 136046 196860 136102
rect 196916 136046 196984 136102
rect 197040 136046 197064 136102
rect 196588 135978 197064 136046
rect 196588 135922 196612 135978
rect 196668 135922 196736 135978
rect 196792 135922 196860 135978
rect 196916 135922 196984 135978
rect 197040 135922 197064 135978
rect 196588 135888 197064 135922
rect 195788 130350 196264 130384
rect 195788 130294 195812 130350
rect 195868 130294 195936 130350
rect 195992 130294 196060 130350
rect 196116 130294 196184 130350
rect 196240 130294 196264 130350
rect 195788 130226 196264 130294
rect 195788 130170 195812 130226
rect 195868 130170 195936 130226
rect 195992 130170 196060 130226
rect 196116 130170 196184 130226
rect 196240 130170 196264 130226
rect 195788 130102 196264 130170
rect 195788 130046 195812 130102
rect 195868 130046 195936 130102
rect 195992 130046 196060 130102
rect 196116 130046 196184 130102
rect 196240 130046 196264 130102
rect 195788 129978 196264 130046
rect 195788 129922 195812 129978
rect 195868 129922 195936 129978
rect 195992 129922 196060 129978
rect 196116 129922 196184 129978
rect 196240 129922 196264 129978
rect 195788 129888 196264 129922
rect 193458 118294 193554 118350
rect 193610 118294 193678 118350
rect 193734 118294 193802 118350
rect 193858 118294 193926 118350
rect 193982 118294 194078 118350
rect 193458 118226 194078 118294
rect 193458 118170 193554 118226
rect 193610 118170 193678 118226
rect 193734 118170 193802 118226
rect 193858 118170 193926 118226
rect 193982 118170 194078 118226
rect 193458 118102 194078 118170
rect 193458 118046 193554 118102
rect 193610 118046 193678 118102
rect 193734 118046 193802 118102
rect 193858 118046 193926 118102
rect 193982 118046 194078 118102
rect 193458 117978 194078 118046
rect 193458 117922 193554 117978
rect 193610 117922 193678 117978
rect 193734 117922 193802 117978
rect 193858 117922 193926 117978
rect 193982 117922 194078 117978
rect 193458 100350 194078 117922
rect 196588 118350 197064 118384
rect 196588 118294 196612 118350
rect 196668 118294 196736 118350
rect 196792 118294 196860 118350
rect 196916 118294 196984 118350
rect 197040 118294 197064 118350
rect 196588 118226 197064 118294
rect 196588 118170 196612 118226
rect 196668 118170 196736 118226
rect 196792 118170 196860 118226
rect 196916 118170 196984 118226
rect 197040 118170 197064 118226
rect 196588 118102 197064 118170
rect 196588 118046 196612 118102
rect 196668 118046 196736 118102
rect 196792 118046 196860 118102
rect 196916 118046 196984 118102
rect 197040 118046 197064 118102
rect 196588 117978 197064 118046
rect 196588 117922 196612 117978
rect 196668 117922 196736 117978
rect 196792 117922 196860 117978
rect 196916 117922 196984 117978
rect 197040 117922 197064 117978
rect 196588 117888 197064 117922
rect 195788 112350 196264 112384
rect 195788 112294 195812 112350
rect 195868 112294 195936 112350
rect 195992 112294 196060 112350
rect 196116 112294 196184 112350
rect 196240 112294 196264 112350
rect 195788 112226 196264 112294
rect 195788 112170 195812 112226
rect 195868 112170 195936 112226
rect 195992 112170 196060 112226
rect 196116 112170 196184 112226
rect 196240 112170 196264 112226
rect 195788 112102 196264 112170
rect 195788 112046 195812 112102
rect 195868 112046 195936 112102
rect 195992 112046 196060 112102
rect 196116 112046 196184 112102
rect 196240 112046 196264 112102
rect 195788 111978 196264 112046
rect 195788 111922 195812 111978
rect 195868 111922 195936 111978
rect 195992 111922 196060 111978
rect 196116 111922 196184 111978
rect 196240 111922 196264 111978
rect 195788 111888 196264 111922
rect 193458 100294 193554 100350
rect 193610 100294 193678 100350
rect 193734 100294 193802 100350
rect 193858 100294 193926 100350
rect 193982 100294 194078 100350
rect 193458 100226 194078 100294
rect 193458 100170 193554 100226
rect 193610 100170 193678 100226
rect 193734 100170 193802 100226
rect 193858 100170 193926 100226
rect 193982 100170 194078 100226
rect 193458 100102 194078 100170
rect 193458 100046 193554 100102
rect 193610 100046 193678 100102
rect 193734 100046 193802 100102
rect 193858 100046 193926 100102
rect 193982 100046 194078 100102
rect 193458 99978 194078 100046
rect 193458 99922 193554 99978
rect 193610 99922 193678 99978
rect 193734 99922 193802 99978
rect 193858 99922 193926 99978
rect 193982 99922 194078 99978
rect 193458 82350 194078 99922
rect 196588 100350 197064 100384
rect 196588 100294 196612 100350
rect 196668 100294 196736 100350
rect 196792 100294 196860 100350
rect 196916 100294 196984 100350
rect 197040 100294 197064 100350
rect 196588 100226 197064 100294
rect 196588 100170 196612 100226
rect 196668 100170 196736 100226
rect 196792 100170 196860 100226
rect 196916 100170 196984 100226
rect 197040 100170 197064 100226
rect 196588 100102 197064 100170
rect 196588 100046 196612 100102
rect 196668 100046 196736 100102
rect 196792 100046 196860 100102
rect 196916 100046 196984 100102
rect 197040 100046 197064 100102
rect 196588 99978 197064 100046
rect 196588 99922 196612 99978
rect 196668 99922 196736 99978
rect 196792 99922 196860 99978
rect 196916 99922 196984 99978
rect 197040 99922 197064 99978
rect 196588 99888 197064 99922
rect 195788 94350 196264 94384
rect 195788 94294 195812 94350
rect 195868 94294 195936 94350
rect 195992 94294 196060 94350
rect 196116 94294 196184 94350
rect 196240 94294 196264 94350
rect 195788 94226 196264 94294
rect 195788 94170 195812 94226
rect 195868 94170 195936 94226
rect 195992 94170 196060 94226
rect 196116 94170 196184 94226
rect 196240 94170 196264 94226
rect 195788 94102 196264 94170
rect 195788 94046 195812 94102
rect 195868 94046 195936 94102
rect 195992 94046 196060 94102
rect 196116 94046 196184 94102
rect 196240 94046 196264 94102
rect 195788 93978 196264 94046
rect 195788 93922 195812 93978
rect 195868 93922 195936 93978
rect 195992 93922 196060 93978
rect 196116 93922 196184 93978
rect 196240 93922 196264 93978
rect 195788 93888 196264 93922
rect 199052 82740 199108 147196
rect 204092 125748 204148 364742
rect 204204 139188 204260 366828
rect 210028 366660 210084 366670
rect 209692 365428 209748 365438
rect 209244 365316 209300 365326
rect 205884 364618 205940 364628
rect 204316 363524 204372 363534
rect 204316 249508 204372 363468
rect 205100 359038 205156 359048
rect 204988 357418 205044 357428
rect 204316 249442 204372 249452
rect 204876 306658 204932 306668
rect 204876 204958 204932 306602
rect 204988 225298 205044 357362
rect 205100 225478 205156 358982
rect 205772 358678 205828 358688
rect 205100 225422 205380 225478
rect 204988 225242 205156 225298
rect 204988 225092 205044 225102
rect 204988 223498 205044 225036
rect 204988 223432 205044 223442
rect 204988 222598 205044 222608
rect 204988 222516 205044 222542
rect 204988 222450 205044 222460
rect 205100 222418 205156 225242
rect 205100 222362 205268 222418
rect 205212 222058 205268 222362
rect 204876 203700 204932 204902
rect 204876 203634 204932 203644
rect 204988 222002 205268 222058
rect 204988 202438 205044 222002
rect 205324 220258 205380 225422
rect 205100 220202 205380 220258
rect 205100 208348 205156 220202
rect 205100 208292 205268 208348
rect 204988 202382 205156 202438
rect 204988 201538 205044 201548
rect 204988 201012 205044 201482
rect 204988 200946 205044 200956
rect 204988 191458 205044 191468
rect 204988 190260 205044 191402
rect 204988 190194 205044 190204
rect 204988 185698 205044 185708
rect 204988 184996 205044 185642
rect 204988 184930 205044 184940
rect 204988 179508 205044 179518
rect 204988 178138 205044 179452
rect 204988 178072 205044 178082
rect 204988 172738 205044 172748
rect 204988 171444 205044 172682
rect 204988 171378 205044 171388
rect 205100 161252 205156 202382
rect 205212 193078 205268 208292
rect 205212 192948 205268 193022
rect 205212 192882 205268 192892
rect 205100 160692 205156 161196
rect 205100 160626 205156 160636
rect 204204 139122 204260 139132
rect 204092 125682 204148 125692
rect 205772 85428 205828 358622
rect 205884 120372 205940 364562
rect 206108 363178 206164 363188
rect 205996 361956 206052 361966
rect 205996 136500 206052 361900
rect 206108 252084 206164 363122
rect 207452 362098 207508 362108
rect 206892 335300 206948 335310
rect 206108 252018 206164 252028
rect 206668 321860 206724 321870
rect 206668 220108 206724 321804
rect 206780 300804 206836 300814
rect 206780 231868 206836 300748
rect 206892 279860 206948 335244
rect 206892 279794 206948 279804
rect 206780 231812 206948 231868
rect 206668 220052 206836 220108
rect 206668 219828 206724 219838
rect 206668 219178 206724 219772
rect 206668 219112 206724 219122
rect 206668 218278 206724 218288
rect 206668 217140 206724 218222
rect 206668 217074 206724 217084
rect 206668 215038 206724 215048
rect 206668 214452 206724 214982
rect 206668 214386 206724 214396
rect 206668 212518 206724 212528
rect 206668 211764 206724 212462
rect 206668 211698 206724 211708
rect 206668 209998 206724 210008
rect 206668 209076 206724 209942
rect 206668 209010 206724 209020
rect 206668 199108 206724 199118
rect 206668 199018 206724 199052
rect 206668 198952 206724 198962
rect 206780 198838 206836 220052
rect 206668 198782 206836 198838
rect 206668 177058 206724 198782
rect 206892 196588 206948 231812
rect 206780 196532 206948 196588
rect 206780 184828 206836 196532
rect 206892 195778 206948 195788
rect 206892 195636 206948 195722
rect 206892 195570 206948 195580
rect 206780 184772 206948 184828
rect 206668 177002 206836 177058
rect 206668 176820 206724 176830
rect 206668 176518 206724 176764
rect 206668 176452 206724 176462
rect 206780 176338 206836 177002
rect 206668 176282 206836 176338
rect 206668 157220 206724 176282
rect 206892 176158 206948 184772
rect 206780 176102 206948 176158
rect 206780 162838 206836 176102
rect 206892 174132 206948 174142
rect 206892 173098 206948 174076
rect 206892 173032 206948 173042
rect 206780 162772 206836 162782
rect 206668 157154 206724 157164
rect 205996 136434 206052 136444
rect 205884 120306 205940 120316
rect 205772 85362 205828 85372
rect 199052 82674 199108 82684
rect 193458 82294 193554 82350
rect 193610 82294 193678 82350
rect 193734 82294 193802 82350
rect 193858 82294 193926 82350
rect 193982 82294 194078 82350
rect 193458 82226 194078 82294
rect 193458 82170 193554 82226
rect 193610 82170 193678 82226
rect 193734 82170 193802 82226
rect 193858 82170 193926 82226
rect 193982 82170 194078 82226
rect 193458 82102 194078 82170
rect 193458 82046 193554 82102
rect 193610 82046 193678 82102
rect 193734 82046 193802 82102
rect 193858 82046 193926 82102
rect 193982 82046 194078 82102
rect 193458 81978 194078 82046
rect 193458 81922 193554 81978
rect 193610 81922 193678 81978
rect 193734 81922 193802 81978
rect 193858 81922 193926 81978
rect 193982 81922 194078 81978
rect 193458 64350 194078 81922
rect 196588 82350 197064 82384
rect 196588 82294 196612 82350
rect 196668 82294 196736 82350
rect 196792 82294 196860 82350
rect 196916 82294 196984 82350
rect 197040 82294 197064 82350
rect 196588 82226 197064 82294
rect 196588 82170 196612 82226
rect 196668 82170 196736 82226
rect 196792 82170 196860 82226
rect 196916 82170 196984 82226
rect 197040 82170 197064 82226
rect 196588 82102 197064 82170
rect 196588 82046 196612 82102
rect 196668 82046 196736 82102
rect 196792 82046 196860 82102
rect 196916 82046 196984 82102
rect 197040 82046 197064 82102
rect 196588 81978 197064 82046
rect 196588 81922 196612 81978
rect 196668 81922 196736 81978
rect 196792 81922 196860 81978
rect 196916 81922 196984 81978
rect 197040 81922 197064 81978
rect 196588 81888 197064 81922
rect 195788 76350 196264 76384
rect 195788 76294 195812 76350
rect 195868 76294 195936 76350
rect 195992 76294 196060 76350
rect 196116 76294 196184 76350
rect 196240 76294 196264 76350
rect 195788 76226 196264 76294
rect 195788 76170 195812 76226
rect 195868 76170 195936 76226
rect 195992 76170 196060 76226
rect 196116 76170 196184 76226
rect 196240 76170 196264 76226
rect 195788 76102 196264 76170
rect 195788 76046 195812 76102
rect 195868 76046 195936 76102
rect 195992 76046 196060 76102
rect 196116 76046 196184 76102
rect 196240 76046 196264 76102
rect 195788 75978 196264 76046
rect 195788 75922 195812 75978
rect 195868 75922 195936 75978
rect 195992 75922 196060 75978
rect 196116 75922 196184 75978
rect 196240 75922 196264 75978
rect 195788 75888 196264 75922
rect 193458 64294 193554 64350
rect 193610 64294 193678 64350
rect 193734 64294 193802 64350
rect 193858 64294 193926 64350
rect 193982 64294 194078 64350
rect 193458 64226 194078 64294
rect 193458 64170 193554 64226
rect 193610 64170 193678 64226
rect 193734 64170 193802 64226
rect 193858 64170 193926 64226
rect 193982 64170 194078 64226
rect 193458 64102 194078 64170
rect 193458 64046 193554 64102
rect 193610 64046 193678 64102
rect 193734 64046 193802 64102
rect 193858 64046 193926 64102
rect 193982 64046 194078 64102
rect 193458 63978 194078 64046
rect 193458 63922 193554 63978
rect 193610 63922 193678 63978
rect 193734 63922 193802 63978
rect 193858 63922 193926 63978
rect 193982 63922 194078 63978
rect 193458 46350 194078 63922
rect 196588 64350 197064 64384
rect 196588 64294 196612 64350
rect 196668 64294 196736 64350
rect 196792 64294 196860 64350
rect 196916 64294 196984 64350
rect 197040 64294 197064 64350
rect 196588 64226 197064 64294
rect 196588 64170 196612 64226
rect 196668 64170 196736 64226
rect 196792 64170 196860 64226
rect 196916 64170 196984 64226
rect 197040 64170 197064 64226
rect 196588 64102 197064 64170
rect 196588 64046 196612 64102
rect 196668 64046 196736 64102
rect 196792 64046 196860 64102
rect 196916 64046 196984 64102
rect 197040 64046 197064 64102
rect 196588 63978 197064 64046
rect 196588 63922 196612 63978
rect 196668 63922 196736 63978
rect 196792 63922 196860 63978
rect 196916 63922 196984 63978
rect 197040 63922 197064 63978
rect 196588 63888 197064 63922
rect 195788 58350 196264 58384
rect 195788 58294 195812 58350
rect 195868 58294 195936 58350
rect 195992 58294 196060 58350
rect 196116 58294 196184 58350
rect 196240 58294 196264 58350
rect 195788 58226 196264 58294
rect 195788 58170 195812 58226
rect 195868 58170 195936 58226
rect 195992 58170 196060 58226
rect 196116 58170 196184 58226
rect 196240 58170 196264 58226
rect 195788 58102 196264 58170
rect 195788 58046 195812 58102
rect 195868 58046 195936 58102
rect 195992 58046 196060 58102
rect 196116 58046 196184 58102
rect 196240 58046 196264 58102
rect 195788 57978 196264 58046
rect 195788 57922 195812 57978
rect 195868 57922 195936 57978
rect 195992 57922 196060 57978
rect 196116 57922 196184 57978
rect 196240 57922 196264 57978
rect 195788 57888 196264 57922
rect 207452 53172 207508 362042
rect 207564 361844 207620 361854
rect 207564 233268 207620 361788
rect 209132 361558 209188 361568
rect 208348 357238 208404 357248
rect 208124 325108 208180 325118
rect 207564 233202 207620 233212
rect 207676 284788 207732 284798
rect 207676 58548 207732 284732
rect 207676 58482 207732 58492
rect 207452 53106 207508 53116
rect 208124 47796 208180 325052
rect 208348 150612 208404 357182
rect 208460 357058 208516 357068
rect 208460 174132 208516 357002
rect 208460 174066 208516 174076
rect 208348 150546 208404 150556
rect 209132 104244 209188 361502
rect 209244 123060 209300 365260
rect 209468 365204 209524 365214
rect 209468 128436 209524 365148
rect 209580 277138 209636 277148
rect 209580 276598 209636 277082
rect 209580 276532 209636 276542
rect 209692 133812 209748 365372
rect 210028 238644 210084 366604
rect 210140 260148 210196 370300
rect 210252 270900 210308 371420
rect 210252 270834 210308 270844
rect 210364 337540 210420 337550
rect 210140 260082 210196 260092
rect 210028 238578 210084 238588
rect 210364 161140 210420 337484
rect 210476 328580 210532 328590
rect 210476 164276 210532 328524
rect 210476 164210 210532 164220
rect 210588 320068 210644 320078
rect 210588 161364 210644 320012
rect 210700 276418 210756 276428
rect 210700 276276 210756 276362
rect 210700 276210 210756 276220
rect 210700 257878 210756 257888
rect 210700 257460 210756 257822
rect 210700 257394 210756 257404
rect 210700 236098 210756 236108
rect 210700 235956 210756 236042
rect 211708 236098 211764 371644
rect 211820 361620 211876 361630
rect 211820 257878 211876 361564
rect 211932 276598 211988 373212
rect 212044 358858 212100 358868
rect 212044 276778 212100 358802
rect 212156 306658 212212 373324
rect 213388 368004 213444 368014
rect 212268 362998 212324 363008
rect 212268 325108 212324 362942
rect 212268 325042 212324 325052
rect 212156 306592 212212 306602
rect 213388 277138 213444 367948
rect 213388 277072 213444 277082
rect 213500 364868 213556 364878
rect 212044 276712 212100 276722
rect 211932 276532 211988 276542
rect 213500 276418 213556 364812
rect 220458 364350 221078 381922
rect 220458 364294 220554 364350
rect 220610 364294 220678 364350
rect 220734 364294 220802 364350
rect 220858 364294 220926 364350
rect 220982 364294 221078 364350
rect 220458 364226 221078 364294
rect 220458 364170 220554 364226
rect 220610 364170 220678 364226
rect 220734 364170 220802 364226
rect 220858 364170 220926 364226
rect 220982 364170 221078 364226
rect 220458 364102 221078 364170
rect 220458 364046 220554 364102
rect 220610 364046 220678 364102
rect 220734 364046 220802 364102
rect 220858 364046 220926 364102
rect 220982 364046 221078 364102
rect 220458 363978 221078 364046
rect 220458 363922 220554 363978
rect 220610 363922 220678 363978
rect 220734 363922 220802 363978
rect 220858 363922 220926 363978
rect 220982 363922 221078 363978
rect 220458 346350 221078 363922
rect 220458 346294 220554 346350
rect 220610 346294 220678 346350
rect 220734 346294 220802 346350
rect 220858 346294 220926 346350
rect 220982 346294 221078 346350
rect 220458 346226 221078 346294
rect 220458 346170 220554 346226
rect 220610 346170 220678 346226
rect 220734 346170 220802 346226
rect 220858 346170 220926 346226
rect 220982 346170 221078 346226
rect 220458 346102 221078 346170
rect 220458 346046 220554 346102
rect 220610 346046 220678 346102
rect 220734 346046 220802 346102
rect 220858 346046 220926 346102
rect 220982 346046 221078 346102
rect 220458 345978 221078 346046
rect 220458 345922 220554 345978
rect 220610 345922 220678 345978
rect 220734 345922 220802 345978
rect 220858 345922 220926 345978
rect 220982 345922 221078 345978
rect 220458 328350 221078 345922
rect 220458 328294 220554 328350
rect 220610 328294 220678 328350
rect 220734 328294 220802 328350
rect 220858 328294 220926 328350
rect 220982 328294 221078 328350
rect 220458 328226 221078 328294
rect 220458 328170 220554 328226
rect 220610 328170 220678 328226
rect 220734 328170 220802 328226
rect 220858 328170 220926 328226
rect 220982 328170 221078 328226
rect 220458 328102 221078 328170
rect 220458 328046 220554 328102
rect 220610 328046 220678 328102
rect 220734 328046 220802 328102
rect 220858 328046 220926 328102
rect 220982 328046 221078 328102
rect 220458 327978 221078 328046
rect 220458 327922 220554 327978
rect 220610 327922 220678 327978
rect 220734 327922 220802 327978
rect 220858 327922 220926 327978
rect 220982 327922 221078 327978
rect 220458 321718 221078 327922
rect 224178 598172 224798 598268
rect 224178 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 224798 598172
rect 224178 598048 224798 598116
rect 224178 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 224798 598048
rect 224178 597924 224798 597992
rect 224178 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 224798 597924
rect 224178 597800 224798 597868
rect 224178 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 224798 597800
rect 224178 586350 224798 597744
rect 224178 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 224798 586350
rect 224178 586226 224798 586294
rect 224178 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 224798 586226
rect 224178 586102 224798 586170
rect 224178 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 224798 586102
rect 224178 585978 224798 586046
rect 224178 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 224798 585978
rect 224178 568350 224798 585922
rect 224178 568294 224274 568350
rect 224330 568294 224398 568350
rect 224454 568294 224522 568350
rect 224578 568294 224646 568350
rect 224702 568294 224798 568350
rect 224178 568226 224798 568294
rect 224178 568170 224274 568226
rect 224330 568170 224398 568226
rect 224454 568170 224522 568226
rect 224578 568170 224646 568226
rect 224702 568170 224798 568226
rect 224178 568102 224798 568170
rect 224178 568046 224274 568102
rect 224330 568046 224398 568102
rect 224454 568046 224522 568102
rect 224578 568046 224646 568102
rect 224702 568046 224798 568102
rect 224178 567978 224798 568046
rect 224178 567922 224274 567978
rect 224330 567922 224398 567978
rect 224454 567922 224522 567978
rect 224578 567922 224646 567978
rect 224702 567922 224798 567978
rect 224178 550350 224798 567922
rect 224178 550294 224274 550350
rect 224330 550294 224398 550350
rect 224454 550294 224522 550350
rect 224578 550294 224646 550350
rect 224702 550294 224798 550350
rect 224178 550226 224798 550294
rect 224178 550170 224274 550226
rect 224330 550170 224398 550226
rect 224454 550170 224522 550226
rect 224578 550170 224646 550226
rect 224702 550170 224798 550226
rect 224178 550102 224798 550170
rect 224178 550046 224274 550102
rect 224330 550046 224398 550102
rect 224454 550046 224522 550102
rect 224578 550046 224646 550102
rect 224702 550046 224798 550102
rect 224178 549978 224798 550046
rect 224178 549922 224274 549978
rect 224330 549922 224398 549978
rect 224454 549922 224522 549978
rect 224578 549922 224646 549978
rect 224702 549922 224798 549978
rect 224178 532350 224798 549922
rect 224178 532294 224274 532350
rect 224330 532294 224398 532350
rect 224454 532294 224522 532350
rect 224578 532294 224646 532350
rect 224702 532294 224798 532350
rect 224178 532226 224798 532294
rect 224178 532170 224274 532226
rect 224330 532170 224398 532226
rect 224454 532170 224522 532226
rect 224578 532170 224646 532226
rect 224702 532170 224798 532226
rect 224178 532102 224798 532170
rect 224178 532046 224274 532102
rect 224330 532046 224398 532102
rect 224454 532046 224522 532102
rect 224578 532046 224646 532102
rect 224702 532046 224798 532102
rect 224178 531978 224798 532046
rect 224178 531922 224274 531978
rect 224330 531922 224398 531978
rect 224454 531922 224522 531978
rect 224578 531922 224646 531978
rect 224702 531922 224798 531978
rect 224178 514350 224798 531922
rect 224178 514294 224274 514350
rect 224330 514294 224398 514350
rect 224454 514294 224522 514350
rect 224578 514294 224646 514350
rect 224702 514294 224798 514350
rect 224178 514226 224798 514294
rect 224178 514170 224274 514226
rect 224330 514170 224398 514226
rect 224454 514170 224522 514226
rect 224578 514170 224646 514226
rect 224702 514170 224798 514226
rect 224178 514102 224798 514170
rect 224178 514046 224274 514102
rect 224330 514046 224398 514102
rect 224454 514046 224522 514102
rect 224578 514046 224646 514102
rect 224702 514046 224798 514102
rect 224178 513978 224798 514046
rect 224178 513922 224274 513978
rect 224330 513922 224398 513978
rect 224454 513922 224522 513978
rect 224578 513922 224646 513978
rect 224702 513922 224798 513978
rect 224178 496350 224798 513922
rect 224178 496294 224274 496350
rect 224330 496294 224398 496350
rect 224454 496294 224522 496350
rect 224578 496294 224646 496350
rect 224702 496294 224798 496350
rect 224178 496226 224798 496294
rect 224178 496170 224274 496226
rect 224330 496170 224398 496226
rect 224454 496170 224522 496226
rect 224578 496170 224646 496226
rect 224702 496170 224798 496226
rect 224178 496102 224798 496170
rect 224178 496046 224274 496102
rect 224330 496046 224398 496102
rect 224454 496046 224522 496102
rect 224578 496046 224646 496102
rect 224702 496046 224798 496102
rect 224178 495978 224798 496046
rect 224178 495922 224274 495978
rect 224330 495922 224398 495978
rect 224454 495922 224522 495978
rect 224578 495922 224646 495978
rect 224702 495922 224798 495978
rect 224178 478350 224798 495922
rect 224178 478294 224274 478350
rect 224330 478294 224398 478350
rect 224454 478294 224522 478350
rect 224578 478294 224646 478350
rect 224702 478294 224798 478350
rect 224178 478226 224798 478294
rect 224178 478170 224274 478226
rect 224330 478170 224398 478226
rect 224454 478170 224522 478226
rect 224578 478170 224646 478226
rect 224702 478170 224798 478226
rect 224178 478102 224798 478170
rect 224178 478046 224274 478102
rect 224330 478046 224398 478102
rect 224454 478046 224522 478102
rect 224578 478046 224646 478102
rect 224702 478046 224798 478102
rect 224178 477978 224798 478046
rect 224178 477922 224274 477978
rect 224330 477922 224398 477978
rect 224454 477922 224522 477978
rect 224578 477922 224646 477978
rect 224702 477922 224798 477978
rect 224178 460350 224798 477922
rect 224178 460294 224274 460350
rect 224330 460294 224398 460350
rect 224454 460294 224522 460350
rect 224578 460294 224646 460350
rect 224702 460294 224798 460350
rect 224178 460226 224798 460294
rect 224178 460170 224274 460226
rect 224330 460170 224398 460226
rect 224454 460170 224522 460226
rect 224578 460170 224646 460226
rect 224702 460170 224798 460226
rect 224178 460102 224798 460170
rect 224178 460046 224274 460102
rect 224330 460046 224398 460102
rect 224454 460046 224522 460102
rect 224578 460046 224646 460102
rect 224702 460046 224798 460102
rect 224178 459978 224798 460046
rect 224178 459922 224274 459978
rect 224330 459922 224398 459978
rect 224454 459922 224522 459978
rect 224578 459922 224646 459978
rect 224702 459922 224798 459978
rect 224178 442350 224798 459922
rect 224178 442294 224274 442350
rect 224330 442294 224398 442350
rect 224454 442294 224522 442350
rect 224578 442294 224646 442350
rect 224702 442294 224798 442350
rect 224178 442226 224798 442294
rect 224178 442170 224274 442226
rect 224330 442170 224398 442226
rect 224454 442170 224522 442226
rect 224578 442170 224646 442226
rect 224702 442170 224798 442226
rect 224178 442102 224798 442170
rect 224178 442046 224274 442102
rect 224330 442046 224398 442102
rect 224454 442046 224522 442102
rect 224578 442046 224646 442102
rect 224702 442046 224798 442102
rect 224178 441978 224798 442046
rect 224178 441922 224274 441978
rect 224330 441922 224398 441978
rect 224454 441922 224522 441978
rect 224578 441922 224646 441978
rect 224702 441922 224798 441978
rect 224178 424350 224798 441922
rect 224178 424294 224274 424350
rect 224330 424294 224398 424350
rect 224454 424294 224522 424350
rect 224578 424294 224646 424350
rect 224702 424294 224798 424350
rect 224178 424226 224798 424294
rect 224178 424170 224274 424226
rect 224330 424170 224398 424226
rect 224454 424170 224522 424226
rect 224578 424170 224646 424226
rect 224702 424170 224798 424226
rect 224178 424102 224798 424170
rect 224178 424046 224274 424102
rect 224330 424046 224398 424102
rect 224454 424046 224522 424102
rect 224578 424046 224646 424102
rect 224702 424046 224798 424102
rect 224178 423978 224798 424046
rect 224178 423922 224274 423978
rect 224330 423922 224398 423978
rect 224454 423922 224522 423978
rect 224578 423922 224646 423978
rect 224702 423922 224798 423978
rect 224178 406350 224798 423922
rect 224178 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 224798 406350
rect 224178 406226 224798 406294
rect 224178 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 224798 406226
rect 224178 406102 224798 406170
rect 224178 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 224798 406102
rect 224178 405978 224798 406046
rect 224178 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 224798 405978
rect 224178 388350 224798 405922
rect 224178 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 224798 388350
rect 224178 388226 224798 388294
rect 224178 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 224798 388226
rect 224178 388102 224798 388170
rect 224178 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 224798 388102
rect 224178 387978 224798 388046
rect 224178 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 224798 387978
rect 224178 370350 224798 387922
rect 224178 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 224798 370350
rect 224178 370226 224798 370294
rect 224178 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 224798 370226
rect 224178 370102 224798 370170
rect 224178 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 224798 370102
rect 224178 369978 224798 370046
rect 224178 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 224798 369978
rect 224178 352350 224798 369922
rect 224178 352294 224274 352350
rect 224330 352294 224398 352350
rect 224454 352294 224522 352350
rect 224578 352294 224646 352350
rect 224702 352294 224798 352350
rect 224178 352226 224798 352294
rect 224178 352170 224274 352226
rect 224330 352170 224398 352226
rect 224454 352170 224522 352226
rect 224578 352170 224646 352226
rect 224702 352170 224798 352226
rect 224178 352102 224798 352170
rect 224178 352046 224274 352102
rect 224330 352046 224398 352102
rect 224454 352046 224522 352102
rect 224578 352046 224646 352102
rect 224702 352046 224798 352102
rect 224178 351978 224798 352046
rect 224178 351922 224274 351978
rect 224330 351922 224398 351978
rect 224454 351922 224522 351978
rect 224578 351922 224646 351978
rect 224702 351922 224798 351978
rect 224178 334350 224798 351922
rect 224178 334294 224274 334350
rect 224330 334294 224398 334350
rect 224454 334294 224522 334350
rect 224578 334294 224646 334350
rect 224702 334294 224798 334350
rect 224178 334226 224798 334294
rect 224178 334170 224274 334226
rect 224330 334170 224398 334226
rect 224454 334170 224522 334226
rect 224578 334170 224646 334226
rect 224702 334170 224798 334226
rect 224178 334102 224798 334170
rect 224178 334046 224274 334102
rect 224330 334046 224398 334102
rect 224454 334046 224522 334102
rect 224578 334046 224646 334102
rect 224702 334046 224798 334102
rect 224178 333978 224798 334046
rect 224178 333922 224274 333978
rect 224330 333922 224398 333978
rect 224454 333922 224522 333978
rect 224578 333922 224646 333978
rect 224702 333922 224798 333978
rect 224178 321718 224798 333922
rect 251178 597212 251798 598268
rect 251178 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 251798 597212
rect 251178 597088 251798 597156
rect 251178 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 251798 597088
rect 251178 596964 251798 597032
rect 251178 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 251798 596964
rect 251178 596840 251798 596908
rect 251178 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 251798 596840
rect 251178 580350 251798 596784
rect 251178 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 251798 580350
rect 251178 580226 251798 580294
rect 251178 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 251798 580226
rect 251178 580102 251798 580170
rect 251178 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 251798 580102
rect 251178 579978 251798 580046
rect 251178 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 251798 579978
rect 251178 562350 251798 579922
rect 251178 562294 251274 562350
rect 251330 562294 251398 562350
rect 251454 562294 251522 562350
rect 251578 562294 251646 562350
rect 251702 562294 251798 562350
rect 251178 562226 251798 562294
rect 251178 562170 251274 562226
rect 251330 562170 251398 562226
rect 251454 562170 251522 562226
rect 251578 562170 251646 562226
rect 251702 562170 251798 562226
rect 251178 562102 251798 562170
rect 251178 562046 251274 562102
rect 251330 562046 251398 562102
rect 251454 562046 251522 562102
rect 251578 562046 251646 562102
rect 251702 562046 251798 562102
rect 251178 561978 251798 562046
rect 251178 561922 251274 561978
rect 251330 561922 251398 561978
rect 251454 561922 251522 561978
rect 251578 561922 251646 561978
rect 251702 561922 251798 561978
rect 251178 544350 251798 561922
rect 251178 544294 251274 544350
rect 251330 544294 251398 544350
rect 251454 544294 251522 544350
rect 251578 544294 251646 544350
rect 251702 544294 251798 544350
rect 251178 544226 251798 544294
rect 251178 544170 251274 544226
rect 251330 544170 251398 544226
rect 251454 544170 251522 544226
rect 251578 544170 251646 544226
rect 251702 544170 251798 544226
rect 251178 544102 251798 544170
rect 251178 544046 251274 544102
rect 251330 544046 251398 544102
rect 251454 544046 251522 544102
rect 251578 544046 251646 544102
rect 251702 544046 251798 544102
rect 251178 543978 251798 544046
rect 251178 543922 251274 543978
rect 251330 543922 251398 543978
rect 251454 543922 251522 543978
rect 251578 543922 251646 543978
rect 251702 543922 251798 543978
rect 251178 526350 251798 543922
rect 251178 526294 251274 526350
rect 251330 526294 251398 526350
rect 251454 526294 251522 526350
rect 251578 526294 251646 526350
rect 251702 526294 251798 526350
rect 251178 526226 251798 526294
rect 251178 526170 251274 526226
rect 251330 526170 251398 526226
rect 251454 526170 251522 526226
rect 251578 526170 251646 526226
rect 251702 526170 251798 526226
rect 251178 526102 251798 526170
rect 251178 526046 251274 526102
rect 251330 526046 251398 526102
rect 251454 526046 251522 526102
rect 251578 526046 251646 526102
rect 251702 526046 251798 526102
rect 251178 525978 251798 526046
rect 251178 525922 251274 525978
rect 251330 525922 251398 525978
rect 251454 525922 251522 525978
rect 251578 525922 251646 525978
rect 251702 525922 251798 525978
rect 251178 508350 251798 525922
rect 251178 508294 251274 508350
rect 251330 508294 251398 508350
rect 251454 508294 251522 508350
rect 251578 508294 251646 508350
rect 251702 508294 251798 508350
rect 251178 508226 251798 508294
rect 251178 508170 251274 508226
rect 251330 508170 251398 508226
rect 251454 508170 251522 508226
rect 251578 508170 251646 508226
rect 251702 508170 251798 508226
rect 251178 508102 251798 508170
rect 251178 508046 251274 508102
rect 251330 508046 251398 508102
rect 251454 508046 251522 508102
rect 251578 508046 251646 508102
rect 251702 508046 251798 508102
rect 251178 507978 251798 508046
rect 251178 507922 251274 507978
rect 251330 507922 251398 507978
rect 251454 507922 251522 507978
rect 251578 507922 251646 507978
rect 251702 507922 251798 507978
rect 251178 490350 251798 507922
rect 251178 490294 251274 490350
rect 251330 490294 251398 490350
rect 251454 490294 251522 490350
rect 251578 490294 251646 490350
rect 251702 490294 251798 490350
rect 251178 490226 251798 490294
rect 251178 490170 251274 490226
rect 251330 490170 251398 490226
rect 251454 490170 251522 490226
rect 251578 490170 251646 490226
rect 251702 490170 251798 490226
rect 251178 490102 251798 490170
rect 251178 490046 251274 490102
rect 251330 490046 251398 490102
rect 251454 490046 251522 490102
rect 251578 490046 251646 490102
rect 251702 490046 251798 490102
rect 251178 489978 251798 490046
rect 251178 489922 251274 489978
rect 251330 489922 251398 489978
rect 251454 489922 251522 489978
rect 251578 489922 251646 489978
rect 251702 489922 251798 489978
rect 251178 472350 251798 489922
rect 251178 472294 251274 472350
rect 251330 472294 251398 472350
rect 251454 472294 251522 472350
rect 251578 472294 251646 472350
rect 251702 472294 251798 472350
rect 251178 472226 251798 472294
rect 251178 472170 251274 472226
rect 251330 472170 251398 472226
rect 251454 472170 251522 472226
rect 251578 472170 251646 472226
rect 251702 472170 251798 472226
rect 251178 472102 251798 472170
rect 251178 472046 251274 472102
rect 251330 472046 251398 472102
rect 251454 472046 251522 472102
rect 251578 472046 251646 472102
rect 251702 472046 251798 472102
rect 251178 471978 251798 472046
rect 251178 471922 251274 471978
rect 251330 471922 251398 471978
rect 251454 471922 251522 471978
rect 251578 471922 251646 471978
rect 251702 471922 251798 471978
rect 251178 454350 251798 471922
rect 251178 454294 251274 454350
rect 251330 454294 251398 454350
rect 251454 454294 251522 454350
rect 251578 454294 251646 454350
rect 251702 454294 251798 454350
rect 251178 454226 251798 454294
rect 251178 454170 251274 454226
rect 251330 454170 251398 454226
rect 251454 454170 251522 454226
rect 251578 454170 251646 454226
rect 251702 454170 251798 454226
rect 251178 454102 251798 454170
rect 251178 454046 251274 454102
rect 251330 454046 251398 454102
rect 251454 454046 251522 454102
rect 251578 454046 251646 454102
rect 251702 454046 251798 454102
rect 251178 453978 251798 454046
rect 251178 453922 251274 453978
rect 251330 453922 251398 453978
rect 251454 453922 251522 453978
rect 251578 453922 251646 453978
rect 251702 453922 251798 453978
rect 251178 436350 251798 453922
rect 251178 436294 251274 436350
rect 251330 436294 251398 436350
rect 251454 436294 251522 436350
rect 251578 436294 251646 436350
rect 251702 436294 251798 436350
rect 251178 436226 251798 436294
rect 251178 436170 251274 436226
rect 251330 436170 251398 436226
rect 251454 436170 251522 436226
rect 251578 436170 251646 436226
rect 251702 436170 251798 436226
rect 251178 436102 251798 436170
rect 251178 436046 251274 436102
rect 251330 436046 251398 436102
rect 251454 436046 251522 436102
rect 251578 436046 251646 436102
rect 251702 436046 251798 436102
rect 251178 435978 251798 436046
rect 251178 435922 251274 435978
rect 251330 435922 251398 435978
rect 251454 435922 251522 435978
rect 251578 435922 251646 435978
rect 251702 435922 251798 435978
rect 251178 418350 251798 435922
rect 251178 418294 251274 418350
rect 251330 418294 251398 418350
rect 251454 418294 251522 418350
rect 251578 418294 251646 418350
rect 251702 418294 251798 418350
rect 251178 418226 251798 418294
rect 251178 418170 251274 418226
rect 251330 418170 251398 418226
rect 251454 418170 251522 418226
rect 251578 418170 251646 418226
rect 251702 418170 251798 418226
rect 251178 418102 251798 418170
rect 251178 418046 251274 418102
rect 251330 418046 251398 418102
rect 251454 418046 251522 418102
rect 251578 418046 251646 418102
rect 251702 418046 251798 418102
rect 251178 417978 251798 418046
rect 251178 417922 251274 417978
rect 251330 417922 251398 417978
rect 251454 417922 251522 417978
rect 251578 417922 251646 417978
rect 251702 417922 251798 417978
rect 251178 400350 251798 417922
rect 251178 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 251798 400350
rect 251178 400226 251798 400294
rect 251178 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 251798 400226
rect 251178 400102 251798 400170
rect 251178 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 251798 400102
rect 251178 399978 251798 400046
rect 251178 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 251798 399978
rect 251178 382350 251798 399922
rect 251178 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 251798 382350
rect 251178 382226 251798 382294
rect 251178 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 251798 382226
rect 251178 382102 251798 382170
rect 251178 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 251798 382102
rect 251178 381978 251798 382046
rect 251178 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 251798 381978
rect 251178 364350 251798 381922
rect 251178 364294 251274 364350
rect 251330 364294 251398 364350
rect 251454 364294 251522 364350
rect 251578 364294 251646 364350
rect 251702 364294 251798 364350
rect 251178 364226 251798 364294
rect 251178 364170 251274 364226
rect 251330 364170 251398 364226
rect 251454 364170 251522 364226
rect 251578 364170 251646 364226
rect 251702 364170 251798 364226
rect 251178 364102 251798 364170
rect 251178 364046 251274 364102
rect 251330 364046 251398 364102
rect 251454 364046 251522 364102
rect 251578 364046 251646 364102
rect 251702 364046 251798 364102
rect 251178 363978 251798 364046
rect 251178 363922 251274 363978
rect 251330 363922 251398 363978
rect 251454 363922 251522 363978
rect 251578 363922 251646 363978
rect 251702 363922 251798 363978
rect 251178 346350 251798 363922
rect 251178 346294 251274 346350
rect 251330 346294 251398 346350
rect 251454 346294 251522 346350
rect 251578 346294 251646 346350
rect 251702 346294 251798 346350
rect 251178 346226 251798 346294
rect 251178 346170 251274 346226
rect 251330 346170 251398 346226
rect 251454 346170 251522 346226
rect 251578 346170 251646 346226
rect 251702 346170 251798 346226
rect 251178 346102 251798 346170
rect 251178 346046 251274 346102
rect 251330 346046 251398 346102
rect 251454 346046 251522 346102
rect 251578 346046 251646 346102
rect 251702 346046 251798 346102
rect 251178 345978 251798 346046
rect 251178 345922 251274 345978
rect 251330 345922 251398 345978
rect 251454 345922 251522 345978
rect 251578 345922 251646 345978
rect 251702 345922 251798 345978
rect 251178 328350 251798 345922
rect 251178 328294 251274 328350
rect 251330 328294 251398 328350
rect 251454 328294 251522 328350
rect 251578 328294 251646 328350
rect 251702 328294 251798 328350
rect 251178 328226 251798 328294
rect 251178 328170 251274 328226
rect 251330 328170 251398 328226
rect 251454 328170 251522 328226
rect 251578 328170 251646 328226
rect 251702 328170 251798 328226
rect 251178 328102 251798 328170
rect 251178 328046 251274 328102
rect 251330 328046 251398 328102
rect 251454 328046 251522 328102
rect 251578 328046 251646 328102
rect 251702 328046 251798 328102
rect 251178 327978 251798 328046
rect 251178 327922 251274 327978
rect 251330 327922 251398 327978
rect 251454 327922 251522 327978
rect 251578 327922 251646 327978
rect 251702 327922 251798 327978
rect 251178 321718 251798 327922
rect 254898 598172 255518 598268
rect 254898 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 255518 598172
rect 254898 598048 255518 598116
rect 254898 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 255518 598048
rect 254898 597924 255518 597992
rect 254898 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 255518 597924
rect 254898 597800 255518 597868
rect 254898 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 255518 597800
rect 254898 586350 255518 597744
rect 254898 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 255518 586350
rect 254898 586226 255518 586294
rect 254898 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 255518 586226
rect 254898 586102 255518 586170
rect 254898 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 255518 586102
rect 254898 585978 255518 586046
rect 254898 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 255518 585978
rect 254898 568350 255518 585922
rect 254898 568294 254994 568350
rect 255050 568294 255118 568350
rect 255174 568294 255242 568350
rect 255298 568294 255366 568350
rect 255422 568294 255518 568350
rect 254898 568226 255518 568294
rect 254898 568170 254994 568226
rect 255050 568170 255118 568226
rect 255174 568170 255242 568226
rect 255298 568170 255366 568226
rect 255422 568170 255518 568226
rect 254898 568102 255518 568170
rect 254898 568046 254994 568102
rect 255050 568046 255118 568102
rect 255174 568046 255242 568102
rect 255298 568046 255366 568102
rect 255422 568046 255518 568102
rect 254898 567978 255518 568046
rect 254898 567922 254994 567978
rect 255050 567922 255118 567978
rect 255174 567922 255242 567978
rect 255298 567922 255366 567978
rect 255422 567922 255518 567978
rect 254898 550350 255518 567922
rect 254898 550294 254994 550350
rect 255050 550294 255118 550350
rect 255174 550294 255242 550350
rect 255298 550294 255366 550350
rect 255422 550294 255518 550350
rect 254898 550226 255518 550294
rect 254898 550170 254994 550226
rect 255050 550170 255118 550226
rect 255174 550170 255242 550226
rect 255298 550170 255366 550226
rect 255422 550170 255518 550226
rect 254898 550102 255518 550170
rect 254898 550046 254994 550102
rect 255050 550046 255118 550102
rect 255174 550046 255242 550102
rect 255298 550046 255366 550102
rect 255422 550046 255518 550102
rect 254898 549978 255518 550046
rect 254898 549922 254994 549978
rect 255050 549922 255118 549978
rect 255174 549922 255242 549978
rect 255298 549922 255366 549978
rect 255422 549922 255518 549978
rect 254898 532350 255518 549922
rect 254898 532294 254994 532350
rect 255050 532294 255118 532350
rect 255174 532294 255242 532350
rect 255298 532294 255366 532350
rect 255422 532294 255518 532350
rect 254898 532226 255518 532294
rect 254898 532170 254994 532226
rect 255050 532170 255118 532226
rect 255174 532170 255242 532226
rect 255298 532170 255366 532226
rect 255422 532170 255518 532226
rect 254898 532102 255518 532170
rect 254898 532046 254994 532102
rect 255050 532046 255118 532102
rect 255174 532046 255242 532102
rect 255298 532046 255366 532102
rect 255422 532046 255518 532102
rect 254898 531978 255518 532046
rect 254898 531922 254994 531978
rect 255050 531922 255118 531978
rect 255174 531922 255242 531978
rect 255298 531922 255366 531978
rect 255422 531922 255518 531978
rect 254898 514350 255518 531922
rect 254898 514294 254994 514350
rect 255050 514294 255118 514350
rect 255174 514294 255242 514350
rect 255298 514294 255366 514350
rect 255422 514294 255518 514350
rect 254898 514226 255518 514294
rect 254898 514170 254994 514226
rect 255050 514170 255118 514226
rect 255174 514170 255242 514226
rect 255298 514170 255366 514226
rect 255422 514170 255518 514226
rect 254898 514102 255518 514170
rect 254898 514046 254994 514102
rect 255050 514046 255118 514102
rect 255174 514046 255242 514102
rect 255298 514046 255366 514102
rect 255422 514046 255518 514102
rect 254898 513978 255518 514046
rect 254898 513922 254994 513978
rect 255050 513922 255118 513978
rect 255174 513922 255242 513978
rect 255298 513922 255366 513978
rect 255422 513922 255518 513978
rect 254898 496350 255518 513922
rect 254898 496294 254994 496350
rect 255050 496294 255118 496350
rect 255174 496294 255242 496350
rect 255298 496294 255366 496350
rect 255422 496294 255518 496350
rect 254898 496226 255518 496294
rect 254898 496170 254994 496226
rect 255050 496170 255118 496226
rect 255174 496170 255242 496226
rect 255298 496170 255366 496226
rect 255422 496170 255518 496226
rect 254898 496102 255518 496170
rect 254898 496046 254994 496102
rect 255050 496046 255118 496102
rect 255174 496046 255242 496102
rect 255298 496046 255366 496102
rect 255422 496046 255518 496102
rect 254898 495978 255518 496046
rect 254898 495922 254994 495978
rect 255050 495922 255118 495978
rect 255174 495922 255242 495978
rect 255298 495922 255366 495978
rect 255422 495922 255518 495978
rect 254898 478350 255518 495922
rect 254898 478294 254994 478350
rect 255050 478294 255118 478350
rect 255174 478294 255242 478350
rect 255298 478294 255366 478350
rect 255422 478294 255518 478350
rect 254898 478226 255518 478294
rect 254898 478170 254994 478226
rect 255050 478170 255118 478226
rect 255174 478170 255242 478226
rect 255298 478170 255366 478226
rect 255422 478170 255518 478226
rect 254898 478102 255518 478170
rect 254898 478046 254994 478102
rect 255050 478046 255118 478102
rect 255174 478046 255242 478102
rect 255298 478046 255366 478102
rect 255422 478046 255518 478102
rect 254898 477978 255518 478046
rect 254898 477922 254994 477978
rect 255050 477922 255118 477978
rect 255174 477922 255242 477978
rect 255298 477922 255366 477978
rect 255422 477922 255518 477978
rect 254898 460350 255518 477922
rect 254898 460294 254994 460350
rect 255050 460294 255118 460350
rect 255174 460294 255242 460350
rect 255298 460294 255366 460350
rect 255422 460294 255518 460350
rect 254898 460226 255518 460294
rect 254898 460170 254994 460226
rect 255050 460170 255118 460226
rect 255174 460170 255242 460226
rect 255298 460170 255366 460226
rect 255422 460170 255518 460226
rect 254898 460102 255518 460170
rect 254898 460046 254994 460102
rect 255050 460046 255118 460102
rect 255174 460046 255242 460102
rect 255298 460046 255366 460102
rect 255422 460046 255518 460102
rect 254898 459978 255518 460046
rect 254898 459922 254994 459978
rect 255050 459922 255118 459978
rect 255174 459922 255242 459978
rect 255298 459922 255366 459978
rect 255422 459922 255518 459978
rect 254898 442350 255518 459922
rect 254898 442294 254994 442350
rect 255050 442294 255118 442350
rect 255174 442294 255242 442350
rect 255298 442294 255366 442350
rect 255422 442294 255518 442350
rect 254898 442226 255518 442294
rect 254898 442170 254994 442226
rect 255050 442170 255118 442226
rect 255174 442170 255242 442226
rect 255298 442170 255366 442226
rect 255422 442170 255518 442226
rect 254898 442102 255518 442170
rect 254898 442046 254994 442102
rect 255050 442046 255118 442102
rect 255174 442046 255242 442102
rect 255298 442046 255366 442102
rect 255422 442046 255518 442102
rect 254898 441978 255518 442046
rect 254898 441922 254994 441978
rect 255050 441922 255118 441978
rect 255174 441922 255242 441978
rect 255298 441922 255366 441978
rect 255422 441922 255518 441978
rect 254898 424350 255518 441922
rect 254898 424294 254994 424350
rect 255050 424294 255118 424350
rect 255174 424294 255242 424350
rect 255298 424294 255366 424350
rect 255422 424294 255518 424350
rect 254898 424226 255518 424294
rect 254898 424170 254994 424226
rect 255050 424170 255118 424226
rect 255174 424170 255242 424226
rect 255298 424170 255366 424226
rect 255422 424170 255518 424226
rect 254898 424102 255518 424170
rect 254898 424046 254994 424102
rect 255050 424046 255118 424102
rect 255174 424046 255242 424102
rect 255298 424046 255366 424102
rect 255422 424046 255518 424102
rect 254898 423978 255518 424046
rect 254898 423922 254994 423978
rect 255050 423922 255118 423978
rect 255174 423922 255242 423978
rect 255298 423922 255366 423978
rect 255422 423922 255518 423978
rect 254898 406350 255518 423922
rect 254898 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 255518 406350
rect 254898 406226 255518 406294
rect 254898 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 255518 406226
rect 254898 406102 255518 406170
rect 254898 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 255518 406102
rect 254898 405978 255518 406046
rect 254898 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 255518 405978
rect 254898 388350 255518 405922
rect 254898 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 255518 388350
rect 254898 388226 255518 388294
rect 254898 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 255518 388226
rect 254898 388102 255518 388170
rect 254898 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 255518 388102
rect 254898 387978 255518 388046
rect 254898 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 255518 387978
rect 254898 370350 255518 387922
rect 254898 370294 254994 370350
rect 255050 370294 255118 370350
rect 255174 370294 255242 370350
rect 255298 370294 255366 370350
rect 255422 370294 255518 370350
rect 254898 370226 255518 370294
rect 254898 370170 254994 370226
rect 255050 370170 255118 370226
rect 255174 370170 255242 370226
rect 255298 370170 255366 370226
rect 255422 370170 255518 370226
rect 254898 370102 255518 370170
rect 254898 370046 254994 370102
rect 255050 370046 255118 370102
rect 255174 370046 255242 370102
rect 255298 370046 255366 370102
rect 255422 370046 255518 370102
rect 254898 369978 255518 370046
rect 254898 369922 254994 369978
rect 255050 369922 255118 369978
rect 255174 369922 255242 369978
rect 255298 369922 255366 369978
rect 255422 369922 255518 369978
rect 254898 352350 255518 369922
rect 254898 352294 254994 352350
rect 255050 352294 255118 352350
rect 255174 352294 255242 352350
rect 255298 352294 255366 352350
rect 255422 352294 255518 352350
rect 254898 352226 255518 352294
rect 254898 352170 254994 352226
rect 255050 352170 255118 352226
rect 255174 352170 255242 352226
rect 255298 352170 255366 352226
rect 255422 352170 255518 352226
rect 254898 352102 255518 352170
rect 254898 352046 254994 352102
rect 255050 352046 255118 352102
rect 255174 352046 255242 352102
rect 255298 352046 255366 352102
rect 255422 352046 255518 352102
rect 254898 351978 255518 352046
rect 254898 351922 254994 351978
rect 255050 351922 255118 351978
rect 255174 351922 255242 351978
rect 255298 351922 255366 351978
rect 255422 351922 255518 351978
rect 254898 334350 255518 351922
rect 254898 334294 254994 334350
rect 255050 334294 255118 334350
rect 255174 334294 255242 334350
rect 255298 334294 255366 334350
rect 255422 334294 255518 334350
rect 254898 334226 255518 334294
rect 254898 334170 254994 334226
rect 255050 334170 255118 334226
rect 255174 334170 255242 334226
rect 255298 334170 255366 334226
rect 255422 334170 255518 334226
rect 254898 334102 255518 334170
rect 254898 334046 254994 334102
rect 255050 334046 255118 334102
rect 255174 334046 255242 334102
rect 255298 334046 255366 334102
rect 255422 334046 255518 334102
rect 254898 333978 255518 334046
rect 254898 333922 254994 333978
rect 255050 333922 255118 333978
rect 255174 333922 255242 333978
rect 255298 333922 255366 333978
rect 255422 333922 255518 333978
rect 254898 321718 255518 333922
rect 281898 597212 282518 598268
rect 281898 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 282518 597212
rect 281898 597088 282518 597156
rect 281898 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 282518 597088
rect 281898 596964 282518 597032
rect 281898 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 282518 596964
rect 281898 596840 282518 596908
rect 281898 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 282518 596840
rect 281898 580350 282518 596784
rect 281898 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 282518 580350
rect 281898 580226 282518 580294
rect 281898 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 282518 580226
rect 281898 580102 282518 580170
rect 281898 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 282518 580102
rect 281898 579978 282518 580046
rect 281898 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 282518 579978
rect 281898 562350 282518 579922
rect 281898 562294 281994 562350
rect 282050 562294 282118 562350
rect 282174 562294 282242 562350
rect 282298 562294 282366 562350
rect 282422 562294 282518 562350
rect 281898 562226 282518 562294
rect 281898 562170 281994 562226
rect 282050 562170 282118 562226
rect 282174 562170 282242 562226
rect 282298 562170 282366 562226
rect 282422 562170 282518 562226
rect 281898 562102 282518 562170
rect 281898 562046 281994 562102
rect 282050 562046 282118 562102
rect 282174 562046 282242 562102
rect 282298 562046 282366 562102
rect 282422 562046 282518 562102
rect 281898 561978 282518 562046
rect 281898 561922 281994 561978
rect 282050 561922 282118 561978
rect 282174 561922 282242 561978
rect 282298 561922 282366 561978
rect 282422 561922 282518 561978
rect 281898 544350 282518 561922
rect 281898 544294 281994 544350
rect 282050 544294 282118 544350
rect 282174 544294 282242 544350
rect 282298 544294 282366 544350
rect 282422 544294 282518 544350
rect 281898 544226 282518 544294
rect 281898 544170 281994 544226
rect 282050 544170 282118 544226
rect 282174 544170 282242 544226
rect 282298 544170 282366 544226
rect 282422 544170 282518 544226
rect 281898 544102 282518 544170
rect 281898 544046 281994 544102
rect 282050 544046 282118 544102
rect 282174 544046 282242 544102
rect 282298 544046 282366 544102
rect 282422 544046 282518 544102
rect 281898 543978 282518 544046
rect 281898 543922 281994 543978
rect 282050 543922 282118 543978
rect 282174 543922 282242 543978
rect 282298 543922 282366 543978
rect 282422 543922 282518 543978
rect 281898 526350 282518 543922
rect 281898 526294 281994 526350
rect 282050 526294 282118 526350
rect 282174 526294 282242 526350
rect 282298 526294 282366 526350
rect 282422 526294 282518 526350
rect 281898 526226 282518 526294
rect 281898 526170 281994 526226
rect 282050 526170 282118 526226
rect 282174 526170 282242 526226
rect 282298 526170 282366 526226
rect 282422 526170 282518 526226
rect 281898 526102 282518 526170
rect 281898 526046 281994 526102
rect 282050 526046 282118 526102
rect 282174 526046 282242 526102
rect 282298 526046 282366 526102
rect 282422 526046 282518 526102
rect 281898 525978 282518 526046
rect 281898 525922 281994 525978
rect 282050 525922 282118 525978
rect 282174 525922 282242 525978
rect 282298 525922 282366 525978
rect 282422 525922 282518 525978
rect 281898 508350 282518 525922
rect 281898 508294 281994 508350
rect 282050 508294 282118 508350
rect 282174 508294 282242 508350
rect 282298 508294 282366 508350
rect 282422 508294 282518 508350
rect 281898 508226 282518 508294
rect 281898 508170 281994 508226
rect 282050 508170 282118 508226
rect 282174 508170 282242 508226
rect 282298 508170 282366 508226
rect 282422 508170 282518 508226
rect 281898 508102 282518 508170
rect 281898 508046 281994 508102
rect 282050 508046 282118 508102
rect 282174 508046 282242 508102
rect 282298 508046 282366 508102
rect 282422 508046 282518 508102
rect 281898 507978 282518 508046
rect 281898 507922 281994 507978
rect 282050 507922 282118 507978
rect 282174 507922 282242 507978
rect 282298 507922 282366 507978
rect 282422 507922 282518 507978
rect 281898 490350 282518 507922
rect 281898 490294 281994 490350
rect 282050 490294 282118 490350
rect 282174 490294 282242 490350
rect 282298 490294 282366 490350
rect 282422 490294 282518 490350
rect 281898 490226 282518 490294
rect 281898 490170 281994 490226
rect 282050 490170 282118 490226
rect 282174 490170 282242 490226
rect 282298 490170 282366 490226
rect 282422 490170 282518 490226
rect 281898 490102 282518 490170
rect 281898 490046 281994 490102
rect 282050 490046 282118 490102
rect 282174 490046 282242 490102
rect 282298 490046 282366 490102
rect 282422 490046 282518 490102
rect 281898 489978 282518 490046
rect 281898 489922 281994 489978
rect 282050 489922 282118 489978
rect 282174 489922 282242 489978
rect 282298 489922 282366 489978
rect 282422 489922 282518 489978
rect 281898 472350 282518 489922
rect 281898 472294 281994 472350
rect 282050 472294 282118 472350
rect 282174 472294 282242 472350
rect 282298 472294 282366 472350
rect 282422 472294 282518 472350
rect 281898 472226 282518 472294
rect 281898 472170 281994 472226
rect 282050 472170 282118 472226
rect 282174 472170 282242 472226
rect 282298 472170 282366 472226
rect 282422 472170 282518 472226
rect 281898 472102 282518 472170
rect 281898 472046 281994 472102
rect 282050 472046 282118 472102
rect 282174 472046 282242 472102
rect 282298 472046 282366 472102
rect 282422 472046 282518 472102
rect 281898 471978 282518 472046
rect 281898 471922 281994 471978
rect 282050 471922 282118 471978
rect 282174 471922 282242 471978
rect 282298 471922 282366 471978
rect 282422 471922 282518 471978
rect 281898 454350 282518 471922
rect 281898 454294 281994 454350
rect 282050 454294 282118 454350
rect 282174 454294 282242 454350
rect 282298 454294 282366 454350
rect 282422 454294 282518 454350
rect 281898 454226 282518 454294
rect 281898 454170 281994 454226
rect 282050 454170 282118 454226
rect 282174 454170 282242 454226
rect 282298 454170 282366 454226
rect 282422 454170 282518 454226
rect 281898 454102 282518 454170
rect 281898 454046 281994 454102
rect 282050 454046 282118 454102
rect 282174 454046 282242 454102
rect 282298 454046 282366 454102
rect 282422 454046 282518 454102
rect 281898 453978 282518 454046
rect 281898 453922 281994 453978
rect 282050 453922 282118 453978
rect 282174 453922 282242 453978
rect 282298 453922 282366 453978
rect 282422 453922 282518 453978
rect 281898 436350 282518 453922
rect 281898 436294 281994 436350
rect 282050 436294 282118 436350
rect 282174 436294 282242 436350
rect 282298 436294 282366 436350
rect 282422 436294 282518 436350
rect 281898 436226 282518 436294
rect 281898 436170 281994 436226
rect 282050 436170 282118 436226
rect 282174 436170 282242 436226
rect 282298 436170 282366 436226
rect 282422 436170 282518 436226
rect 281898 436102 282518 436170
rect 281898 436046 281994 436102
rect 282050 436046 282118 436102
rect 282174 436046 282242 436102
rect 282298 436046 282366 436102
rect 282422 436046 282518 436102
rect 281898 435978 282518 436046
rect 281898 435922 281994 435978
rect 282050 435922 282118 435978
rect 282174 435922 282242 435978
rect 282298 435922 282366 435978
rect 282422 435922 282518 435978
rect 281898 418350 282518 435922
rect 281898 418294 281994 418350
rect 282050 418294 282118 418350
rect 282174 418294 282242 418350
rect 282298 418294 282366 418350
rect 282422 418294 282518 418350
rect 281898 418226 282518 418294
rect 281898 418170 281994 418226
rect 282050 418170 282118 418226
rect 282174 418170 282242 418226
rect 282298 418170 282366 418226
rect 282422 418170 282518 418226
rect 281898 418102 282518 418170
rect 281898 418046 281994 418102
rect 282050 418046 282118 418102
rect 282174 418046 282242 418102
rect 282298 418046 282366 418102
rect 282422 418046 282518 418102
rect 281898 417978 282518 418046
rect 281898 417922 281994 417978
rect 282050 417922 282118 417978
rect 282174 417922 282242 417978
rect 282298 417922 282366 417978
rect 282422 417922 282518 417978
rect 281898 400350 282518 417922
rect 281898 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 282518 400350
rect 281898 400226 282518 400294
rect 281898 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 282518 400226
rect 281898 400102 282518 400170
rect 281898 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 282518 400102
rect 281898 399978 282518 400046
rect 281898 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 282518 399978
rect 281898 382350 282518 399922
rect 281898 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 282518 382350
rect 281898 382226 282518 382294
rect 281898 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 282518 382226
rect 281898 382102 282518 382170
rect 281898 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 282518 382102
rect 281898 381978 282518 382046
rect 281898 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 282518 381978
rect 281898 364350 282518 381922
rect 281898 364294 281994 364350
rect 282050 364294 282118 364350
rect 282174 364294 282242 364350
rect 282298 364294 282366 364350
rect 282422 364294 282518 364350
rect 281898 364226 282518 364294
rect 281898 364170 281994 364226
rect 282050 364170 282118 364226
rect 282174 364170 282242 364226
rect 282298 364170 282366 364226
rect 282422 364170 282518 364226
rect 281898 364102 282518 364170
rect 281898 364046 281994 364102
rect 282050 364046 282118 364102
rect 282174 364046 282242 364102
rect 282298 364046 282366 364102
rect 282422 364046 282518 364102
rect 281898 363978 282518 364046
rect 281898 363922 281994 363978
rect 282050 363922 282118 363978
rect 282174 363922 282242 363978
rect 282298 363922 282366 363978
rect 282422 363922 282518 363978
rect 281898 346350 282518 363922
rect 281898 346294 281994 346350
rect 282050 346294 282118 346350
rect 282174 346294 282242 346350
rect 282298 346294 282366 346350
rect 282422 346294 282518 346350
rect 281898 346226 282518 346294
rect 281898 346170 281994 346226
rect 282050 346170 282118 346226
rect 282174 346170 282242 346226
rect 282298 346170 282366 346226
rect 282422 346170 282518 346226
rect 281898 346102 282518 346170
rect 281898 346046 281994 346102
rect 282050 346046 282118 346102
rect 282174 346046 282242 346102
rect 282298 346046 282366 346102
rect 282422 346046 282518 346102
rect 281898 345978 282518 346046
rect 281898 345922 281994 345978
rect 282050 345922 282118 345978
rect 282174 345922 282242 345978
rect 282298 345922 282366 345978
rect 282422 345922 282518 345978
rect 281898 328350 282518 345922
rect 281898 328294 281994 328350
rect 282050 328294 282118 328350
rect 282174 328294 282242 328350
rect 282298 328294 282366 328350
rect 282422 328294 282518 328350
rect 281898 328226 282518 328294
rect 281898 328170 281994 328226
rect 282050 328170 282118 328226
rect 282174 328170 282242 328226
rect 282298 328170 282366 328226
rect 282422 328170 282518 328226
rect 281898 328102 282518 328170
rect 281898 328046 281994 328102
rect 282050 328046 282118 328102
rect 282174 328046 282242 328102
rect 282298 328046 282366 328102
rect 282422 328046 282518 328102
rect 281898 327978 282518 328046
rect 281898 327922 281994 327978
rect 282050 327922 282118 327978
rect 282174 327922 282242 327978
rect 282298 327922 282366 327978
rect 282422 327922 282518 327978
rect 281898 321718 282518 327922
rect 285618 598172 286238 598268
rect 285618 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 286238 598172
rect 285618 598048 286238 598116
rect 285618 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 286238 598048
rect 285618 597924 286238 597992
rect 285618 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 286238 597924
rect 285618 597800 286238 597868
rect 285618 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 286238 597800
rect 285618 586350 286238 597744
rect 285618 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 286238 586350
rect 285618 586226 286238 586294
rect 285618 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 286238 586226
rect 285618 586102 286238 586170
rect 285618 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 286238 586102
rect 285618 585978 286238 586046
rect 285618 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 286238 585978
rect 285618 568350 286238 585922
rect 285618 568294 285714 568350
rect 285770 568294 285838 568350
rect 285894 568294 285962 568350
rect 286018 568294 286086 568350
rect 286142 568294 286238 568350
rect 285618 568226 286238 568294
rect 285618 568170 285714 568226
rect 285770 568170 285838 568226
rect 285894 568170 285962 568226
rect 286018 568170 286086 568226
rect 286142 568170 286238 568226
rect 285618 568102 286238 568170
rect 285618 568046 285714 568102
rect 285770 568046 285838 568102
rect 285894 568046 285962 568102
rect 286018 568046 286086 568102
rect 286142 568046 286238 568102
rect 285618 567978 286238 568046
rect 285618 567922 285714 567978
rect 285770 567922 285838 567978
rect 285894 567922 285962 567978
rect 286018 567922 286086 567978
rect 286142 567922 286238 567978
rect 285618 550350 286238 567922
rect 285618 550294 285714 550350
rect 285770 550294 285838 550350
rect 285894 550294 285962 550350
rect 286018 550294 286086 550350
rect 286142 550294 286238 550350
rect 285618 550226 286238 550294
rect 285618 550170 285714 550226
rect 285770 550170 285838 550226
rect 285894 550170 285962 550226
rect 286018 550170 286086 550226
rect 286142 550170 286238 550226
rect 285618 550102 286238 550170
rect 285618 550046 285714 550102
rect 285770 550046 285838 550102
rect 285894 550046 285962 550102
rect 286018 550046 286086 550102
rect 286142 550046 286238 550102
rect 285618 549978 286238 550046
rect 285618 549922 285714 549978
rect 285770 549922 285838 549978
rect 285894 549922 285962 549978
rect 286018 549922 286086 549978
rect 286142 549922 286238 549978
rect 285618 532350 286238 549922
rect 285618 532294 285714 532350
rect 285770 532294 285838 532350
rect 285894 532294 285962 532350
rect 286018 532294 286086 532350
rect 286142 532294 286238 532350
rect 285618 532226 286238 532294
rect 285618 532170 285714 532226
rect 285770 532170 285838 532226
rect 285894 532170 285962 532226
rect 286018 532170 286086 532226
rect 286142 532170 286238 532226
rect 285618 532102 286238 532170
rect 285618 532046 285714 532102
rect 285770 532046 285838 532102
rect 285894 532046 285962 532102
rect 286018 532046 286086 532102
rect 286142 532046 286238 532102
rect 285618 531978 286238 532046
rect 285618 531922 285714 531978
rect 285770 531922 285838 531978
rect 285894 531922 285962 531978
rect 286018 531922 286086 531978
rect 286142 531922 286238 531978
rect 285618 514350 286238 531922
rect 285618 514294 285714 514350
rect 285770 514294 285838 514350
rect 285894 514294 285962 514350
rect 286018 514294 286086 514350
rect 286142 514294 286238 514350
rect 285618 514226 286238 514294
rect 285618 514170 285714 514226
rect 285770 514170 285838 514226
rect 285894 514170 285962 514226
rect 286018 514170 286086 514226
rect 286142 514170 286238 514226
rect 285618 514102 286238 514170
rect 285618 514046 285714 514102
rect 285770 514046 285838 514102
rect 285894 514046 285962 514102
rect 286018 514046 286086 514102
rect 286142 514046 286238 514102
rect 285618 513978 286238 514046
rect 285618 513922 285714 513978
rect 285770 513922 285838 513978
rect 285894 513922 285962 513978
rect 286018 513922 286086 513978
rect 286142 513922 286238 513978
rect 285618 496350 286238 513922
rect 285618 496294 285714 496350
rect 285770 496294 285838 496350
rect 285894 496294 285962 496350
rect 286018 496294 286086 496350
rect 286142 496294 286238 496350
rect 285618 496226 286238 496294
rect 285618 496170 285714 496226
rect 285770 496170 285838 496226
rect 285894 496170 285962 496226
rect 286018 496170 286086 496226
rect 286142 496170 286238 496226
rect 285618 496102 286238 496170
rect 285618 496046 285714 496102
rect 285770 496046 285838 496102
rect 285894 496046 285962 496102
rect 286018 496046 286086 496102
rect 286142 496046 286238 496102
rect 285618 495978 286238 496046
rect 285618 495922 285714 495978
rect 285770 495922 285838 495978
rect 285894 495922 285962 495978
rect 286018 495922 286086 495978
rect 286142 495922 286238 495978
rect 285618 478350 286238 495922
rect 285618 478294 285714 478350
rect 285770 478294 285838 478350
rect 285894 478294 285962 478350
rect 286018 478294 286086 478350
rect 286142 478294 286238 478350
rect 285618 478226 286238 478294
rect 285618 478170 285714 478226
rect 285770 478170 285838 478226
rect 285894 478170 285962 478226
rect 286018 478170 286086 478226
rect 286142 478170 286238 478226
rect 285618 478102 286238 478170
rect 285618 478046 285714 478102
rect 285770 478046 285838 478102
rect 285894 478046 285962 478102
rect 286018 478046 286086 478102
rect 286142 478046 286238 478102
rect 285618 477978 286238 478046
rect 285618 477922 285714 477978
rect 285770 477922 285838 477978
rect 285894 477922 285962 477978
rect 286018 477922 286086 477978
rect 286142 477922 286238 477978
rect 285618 460350 286238 477922
rect 285618 460294 285714 460350
rect 285770 460294 285838 460350
rect 285894 460294 285962 460350
rect 286018 460294 286086 460350
rect 286142 460294 286238 460350
rect 285618 460226 286238 460294
rect 285618 460170 285714 460226
rect 285770 460170 285838 460226
rect 285894 460170 285962 460226
rect 286018 460170 286086 460226
rect 286142 460170 286238 460226
rect 285618 460102 286238 460170
rect 285618 460046 285714 460102
rect 285770 460046 285838 460102
rect 285894 460046 285962 460102
rect 286018 460046 286086 460102
rect 286142 460046 286238 460102
rect 285618 459978 286238 460046
rect 285618 459922 285714 459978
rect 285770 459922 285838 459978
rect 285894 459922 285962 459978
rect 286018 459922 286086 459978
rect 286142 459922 286238 459978
rect 285618 442350 286238 459922
rect 285618 442294 285714 442350
rect 285770 442294 285838 442350
rect 285894 442294 285962 442350
rect 286018 442294 286086 442350
rect 286142 442294 286238 442350
rect 285618 442226 286238 442294
rect 285618 442170 285714 442226
rect 285770 442170 285838 442226
rect 285894 442170 285962 442226
rect 286018 442170 286086 442226
rect 286142 442170 286238 442226
rect 285618 442102 286238 442170
rect 285618 442046 285714 442102
rect 285770 442046 285838 442102
rect 285894 442046 285962 442102
rect 286018 442046 286086 442102
rect 286142 442046 286238 442102
rect 285618 441978 286238 442046
rect 285618 441922 285714 441978
rect 285770 441922 285838 441978
rect 285894 441922 285962 441978
rect 286018 441922 286086 441978
rect 286142 441922 286238 441978
rect 285618 424350 286238 441922
rect 285618 424294 285714 424350
rect 285770 424294 285838 424350
rect 285894 424294 285962 424350
rect 286018 424294 286086 424350
rect 286142 424294 286238 424350
rect 285618 424226 286238 424294
rect 285618 424170 285714 424226
rect 285770 424170 285838 424226
rect 285894 424170 285962 424226
rect 286018 424170 286086 424226
rect 286142 424170 286238 424226
rect 285618 424102 286238 424170
rect 285618 424046 285714 424102
rect 285770 424046 285838 424102
rect 285894 424046 285962 424102
rect 286018 424046 286086 424102
rect 286142 424046 286238 424102
rect 285618 423978 286238 424046
rect 285618 423922 285714 423978
rect 285770 423922 285838 423978
rect 285894 423922 285962 423978
rect 286018 423922 286086 423978
rect 286142 423922 286238 423978
rect 285618 406350 286238 423922
rect 285618 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 286238 406350
rect 285618 406226 286238 406294
rect 285618 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 286238 406226
rect 285618 406102 286238 406170
rect 285618 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 286238 406102
rect 285618 405978 286238 406046
rect 285618 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 286238 405978
rect 285618 388350 286238 405922
rect 285618 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 286238 388350
rect 285618 388226 286238 388294
rect 285618 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 286238 388226
rect 285618 388102 286238 388170
rect 285618 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 286238 388102
rect 285618 387978 286238 388046
rect 285618 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 286238 387978
rect 285618 370350 286238 387922
rect 285618 370294 285714 370350
rect 285770 370294 285838 370350
rect 285894 370294 285962 370350
rect 286018 370294 286086 370350
rect 286142 370294 286238 370350
rect 285618 370226 286238 370294
rect 285618 370170 285714 370226
rect 285770 370170 285838 370226
rect 285894 370170 285962 370226
rect 286018 370170 286086 370226
rect 286142 370170 286238 370226
rect 285618 370102 286238 370170
rect 285618 370046 285714 370102
rect 285770 370046 285838 370102
rect 285894 370046 285962 370102
rect 286018 370046 286086 370102
rect 286142 370046 286238 370102
rect 285618 369978 286238 370046
rect 285618 369922 285714 369978
rect 285770 369922 285838 369978
rect 285894 369922 285962 369978
rect 286018 369922 286086 369978
rect 286142 369922 286238 369978
rect 285618 352350 286238 369922
rect 285618 352294 285714 352350
rect 285770 352294 285838 352350
rect 285894 352294 285962 352350
rect 286018 352294 286086 352350
rect 286142 352294 286238 352350
rect 285618 352226 286238 352294
rect 285618 352170 285714 352226
rect 285770 352170 285838 352226
rect 285894 352170 285962 352226
rect 286018 352170 286086 352226
rect 286142 352170 286238 352226
rect 285618 352102 286238 352170
rect 285618 352046 285714 352102
rect 285770 352046 285838 352102
rect 285894 352046 285962 352102
rect 286018 352046 286086 352102
rect 286142 352046 286238 352102
rect 285618 351978 286238 352046
rect 285618 351922 285714 351978
rect 285770 351922 285838 351978
rect 285894 351922 285962 351978
rect 286018 351922 286086 351978
rect 286142 351922 286238 351978
rect 285618 334350 286238 351922
rect 285618 334294 285714 334350
rect 285770 334294 285838 334350
rect 285894 334294 285962 334350
rect 286018 334294 286086 334350
rect 286142 334294 286238 334350
rect 285618 334226 286238 334294
rect 285618 334170 285714 334226
rect 285770 334170 285838 334226
rect 285894 334170 285962 334226
rect 286018 334170 286086 334226
rect 286142 334170 286238 334226
rect 285618 334102 286238 334170
rect 285618 334046 285714 334102
rect 285770 334046 285838 334102
rect 285894 334046 285962 334102
rect 286018 334046 286086 334102
rect 286142 334046 286238 334102
rect 285618 333978 286238 334046
rect 285618 333922 285714 333978
rect 285770 333922 285838 333978
rect 285894 333922 285962 333978
rect 286018 333922 286086 333978
rect 286142 333922 286238 333978
rect 285618 321718 286238 333922
rect 312618 597212 313238 598268
rect 312618 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 313238 597212
rect 312618 597088 313238 597156
rect 312618 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 313238 597088
rect 312618 596964 313238 597032
rect 312618 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 313238 596964
rect 312618 596840 313238 596908
rect 312618 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 313238 596840
rect 312618 580350 313238 596784
rect 312618 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 313238 580350
rect 312618 580226 313238 580294
rect 312618 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 313238 580226
rect 312618 580102 313238 580170
rect 312618 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 313238 580102
rect 312618 579978 313238 580046
rect 312618 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 313238 579978
rect 312618 562350 313238 579922
rect 312618 562294 312714 562350
rect 312770 562294 312838 562350
rect 312894 562294 312962 562350
rect 313018 562294 313086 562350
rect 313142 562294 313238 562350
rect 312618 562226 313238 562294
rect 312618 562170 312714 562226
rect 312770 562170 312838 562226
rect 312894 562170 312962 562226
rect 313018 562170 313086 562226
rect 313142 562170 313238 562226
rect 312618 562102 313238 562170
rect 312618 562046 312714 562102
rect 312770 562046 312838 562102
rect 312894 562046 312962 562102
rect 313018 562046 313086 562102
rect 313142 562046 313238 562102
rect 312618 561978 313238 562046
rect 312618 561922 312714 561978
rect 312770 561922 312838 561978
rect 312894 561922 312962 561978
rect 313018 561922 313086 561978
rect 313142 561922 313238 561978
rect 312618 544350 313238 561922
rect 312618 544294 312714 544350
rect 312770 544294 312838 544350
rect 312894 544294 312962 544350
rect 313018 544294 313086 544350
rect 313142 544294 313238 544350
rect 312618 544226 313238 544294
rect 312618 544170 312714 544226
rect 312770 544170 312838 544226
rect 312894 544170 312962 544226
rect 313018 544170 313086 544226
rect 313142 544170 313238 544226
rect 312618 544102 313238 544170
rect 312618 544046 312714 544102
rect 312770 544046 312838 544102
rect 312894 544046 312962 544102
rect 313018 544046 313086 544102
rect 313142 544046 313238 544102
rect 312618 543978 313238 544046
rect 312618 543922 312714 543978
rect 312770 543922 312838 543978
rect 312894 543922 312962 543978
rect 313018 543922 313086 543978
rect 313142 543922 313238 543978
rect 312618 526350 313238 543922
rect 312618 526294 312714 526350
rect 312770 526294 312838 526350
rect 312894 526294 312962 526350
rect 313018 526294 313086 526350
rect 313142 526294 313238 526350
rect 312618 526226 313238 526294
rect 312618 526170 312714 526226
rect 312770 526170 312838 526226
rect 312894 526170 312962 526226
rect 313018 526170 313086 526226
rect 313142 526170 313238 526226
rect 312618 526102 313238 526170
rect 312618 526046 312714 526102
rect 312770 526046 312838 526102
rect 312894 526046 312962 526102
rect 313018 526046 313086 526102
rect 313142 526046 313238 526102
rect 312618 525978 313238 526046
rect 312618 525922 312714 525978
rect 312770 525922 312838 525978
rect 312894 525922 312962 525978
rect 313018 525922 313086 525978
rect 313142 525922 313238 525978
rect 312618 508350 313238 525922
rect 312618 508294 312714 508350
rect 312770 508294 312838 508350
rect 312894 508294 312962 508350
rect 313018 508294 313086 508350
rect 313142 508294 313238 508350
rect 312618 508226 313238 508294
rect 312618 508170 312714 508226
rect 312770 508170 312838 508226
rect 312894 508170 312962 508226
rect 313018 508170 313086 508226
rect 313142 508170 313238 508226
rect 312618 508102 313238 508170
rect 312618 508046 312714 508102
rect 312770 508046 312838 508102
rect 312894 508046 312962 508102
rect 313018 508046 313086 508102
rect 313142 508046 313238 508102
rect 312618 507978 313238 508046
rect 312618 507922 312714 507978
rect 312770 507922 312838 507978
rect 312894 507922 312962 507978
rect 313018 507922 313086 507978
rect 313142 507922 313238 507978
rect 312618 490350 313238 507922
rect 312618 490294 312714 490350
rect 312770 490294 312838 490350
rect 312894 490294 312962 490350
rect 313018 490294 313086 490350
rect 313142 490294 313238 490350
rect 312618 490226 313238 490294
rect 312618 490170 312714 490226
rect 312770 490170 312838 490226
rect 312894 490170 312962 490226
rect 313018 490170 313086 490226
rect 313142 490170 313238 490226
rect 312618 490102 313238 490170
rect 312618 490046 312714 490102
rect 312770 490046 312838 490102
rect 312894 490046 312962 490102
rect 313018 490046 313086 490102
rect 313142 490046 313238 490102
rect 312618 489978 313238 490046
rect 312618 489922 312714 489978
rect 312770 489922 312838 489978
rect 312894 489922 312962 489978
rect 313018 489922 313086 489978
rect 313142 489922 313238 489978
rect 312618 472350 313238 489922
rect 312618 472294 312714 472350
rect 312770 472294 312838 472350
rect 312894 472294 312962 472350
rect 313018 472294 313086 472350
rect 313142 472294 313238 472350
rect 312618 472226 313238 472294
rect 312618 472170 312714 472226
rect 312770 472170 312838 472226
rect 312894 472170 312962 472226
rect 313018 472170 313086 472226
rect 313142 472170 313238 472226
rect 312618 472102 313238 472170
rect 312618 472046 312714 472102
rect 312770 472046 312838 472102
rect 312894 472046 312962 472102
rect 313018 472046 313086 472102
rect 313142 472046 313238 472102
rect 312618 471978 313238 472046
rect 312618 471922 312714 471978
rect 312770 471922 312838 471978
rect 312894 471922 312962 471978
rect 313018 471922 313086 471978
rect 313142 471922 313238 471978
rect 312618 454350 313238 471922
rect 312618 454294 312714 454350
rect 312770 454294 312838 454350
rect 312894 454294 312962 454350
rect 313018 454294 313086 454350
rect 313142 454294 313238 454350
rect 312618 454226 313238 454294
rect 312618 454170 312714 454226
rect 312770 454170 312838 454226
rect 312894 454170 312962 454226
rect 313018 454170 313086 454226
rect 313142 454170 313238 454226
rect 312618 454102 313238 454170
rect 312618 454046 312714 454102
rect 312770 454046 312838 454102
rect 312894 454046 312962 454102
rect 313018 454046 313086 454102
rect 313142 454046 313238 454102
rect 312618 453978 313238 454046
rect 312618 453922 312714 453978
rect 312770 453922 312838 453978
rect 312894 453922 312962 453978
rect 313018 453922 313086 453978
rect 313142 453922 313238 453978
rect 312618 436350 313238 453922
rect 312618 436294 312714 436350
rect 312770 436294 312838 436350
rect 312894 436294 312962 436350
rect 313018 436294 313086 436350
rect 313142 436294 313238 436350
rect 312618 436226 313238 436294
rect 312618 436170 312714 436226
rect 312770 436170 312838 436226
rect 312894 436170 312962 436226
rect 313018 436170 313086 436226
rect 313142 436170 313238 436226
rect 312618 436102 313238 436170
rect 312618 436046 312714 436102
rect 312770 436046 312838 436102
rect 312894 436046 312962 436102
rect 313018 436046 313086 436102
rect 313142 436046 313238 436102
rect 312618 435978 313238 436046
rect 312618 435922 312714 435978
rect 312770 435922 312838 435978
rect 312894 435922 312962 435978
rect 313018 435922 313086 435978
rect 313142 435922 313238 435978
rect 312618 418350 313238 435922
rect 312618 418294 312714 418350
rect 312770 418294 312838 418350
rect 312894 418294 312962 418350
rect 313018 418294 313086 418350
rect 313142 418294 313238 418350
rect 312618 418226 313238 418294
rect 312618 418170 312714 418226
rect 312770 418170 312838 418226
rect 312894 418170 312962 418226
rect 313018 418170 313086 418226
rect 313142 418170 313238 418226
rect 312618 418102 313238 418170
rect 312618 418046 312714 418102
rect 312770 418046 312838 418102
rect 312894 418046 312962 418102
rect 313018 418046 313086 418102
rect 313142 418046 313238 418102
rect 312618 417978 313238 418046
rect 312618 417922 312714 417978
rect 312770 417922 312838 417978
rect 312894 417922 312962 417978
rect 313018 417922 313086 417978
rect 313142 417922 313238 417978
rect 312618 400350 313238 417922
rect 312618 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 313238 400350
rect 312618 400226 313238 400294
rect 312618 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 313238 400226
rect 312618 400102 313238 400170
rect 312618 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 313238 400102
rect 312618 399978 313238 400046
rect 312618 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 313238 399978
rect 312618 382350 313238 399922
rect 312618 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 313238 382350
rect 312618 382226 313238 382294
rect 312618 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 313238 382226
rect 312618 382102 313238 382170
rect 312618 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 313238 382102
rect 312618 381978 313238 382046
rect 312618 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 313238 381978
rect 312618 364350 313238 381922
rect 312618 364294 312714 364350
rect 312770 364294 312838 364350
rect 312894 364294 312962 364350
rect 313018 364294 313086 364350
rect 313142 364294 313238 364350
rect 312618 364226 313238 364294
rect 312618 364170 312714 364226
rect 312770 364170 312838 364226
rect 312894 364170 312962 364226
rect 313018 364170 313086 364226
rect 313142 364170 313238 364226
rect 312618 364102 313238 364170
rect 312618 364046 312714 364102
rect 312770 364046 312838 364102
rect 312894 364046 312962 364102
rect 313018 364046 313086 364102
rect 313142 364046 313238 364102
rect 312618 363978 313238 364046
rect 312618 363922 312714 363978
rect 312770 363922 312838 363978
rect 312894 363922 312962 363978
rect 313018 363922 313086 363978
rect 313142 363922 313238 363978
rect 312618 346350 313238 363922
rect 312618 346294 312714 346350
rect 312770 346294 312838 346350
rect 312894 346294 312962 346350
rect 313018 346294 313086 346350
rect 313142 346294 313238 346350
rect 312618 346226 313238 346294
rect 312618 346170 312714 346226
rect 312770 346170 312838 346226
rect 312894 346170 312962 346226
rect 313018 346170 313086 346226
rect 313142 346170 313238 346226
rect 312618 346102 313238 346170
rect 312618 346046 312714 346102
rect 312770 346046 312838 346102
rect 312894 346046 312962 346102
rect 313018 346046 313086 346102
rect 313142 346046 313238 346102
rect 312618 345978 313238 346046
rect 312618 345922 312714 345978
rect 312770 345922 312838 345978
rect 312894 345922 312962 345978
rect 313018 345922 313086 345978
rect 313142 345922 313238 345978
rect 312618 328350 313238 345922
rect 312618 328294 312714 328350
rect 312770 328294 312838 328350
rect 312894 328294 312962 328350
rect 313018 328294 313086 328350
rect 313142 328294 313238 328350
rect 312618 328226 313238 328294
rect 312618 328170 312714 328226
rect 312770 328170 312838 328226
rect 312894 328170 312962 328226
rect 313018 328170 313086 328226
rect 313142 328170 313238 328226
rect 312618 328102 313238 328170
rect 312618 328046 312714 328102
rect 312770 328046 312838 328102
rect 312894 328046 312962 328102
rect 313018 328046 313086 328102
rect 313142 328046 313238 328102
rect 312618 327978 313238 328046
rect 312618 327922 312714 327978
rect 312770 327922 312838 327978
rect 312894 327922 312962 327978
rect 313018 327922 313086 327978
rect 313142 327922 313238 327978
rect 312618 321718 313238 327922
rect 316338 598172 316958 598268
rect 316338 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 316958 598172
rect 316338 598048 316958 598116
rect 316338 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 316958 598048
rect 316338 597924 316958 597992
rect 316338 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 316958 597924
rect 316338 597800 316958 597868
rect 316338 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 316958 597800
rect 316338 586350 316958 597744
rect 316338 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 316958 586350
rect 316338 586226 316958 586294
rect 316338 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 316958 586226
rect 316338 586102 316958 586170
rect 316338 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 316958 586102
rect 316338 585978 316958 586046
rect 316338 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 316958 585978
rect 316338 568350 316958 585922
rect 316338 568294 316434 568350
rect 316490 568294 316558 568350
rect 316614 568294 316682 568350
rect 316738 568294 316806 568350
rect 316862 568294 316958 568350
rect 316338 568226 316958 568294
rect 316338 568170 316434 568226
rect 316490 568170 316558 568226
rect 316614 568170 316682 568226
rect 316738 568170 316806 568226
rect 316862 568170 316958 568226
rect 316338 568102 316958 568170
rect 316338 568046 316434 568102
rect 316490 568046 316558 568102
rect 316614 568046 316682 568102
rect 316738 568046 316806 568102
rect 316862 568046 316958 568102
rect 316338 567978 316958 568046
rect 316338 567922 316434 567978
rect 316490 567922 316558 567978
rect 316614 567922 316682 567978
rect 316738 567922 316806 567978
rect 316862 567922 316958 567978
rect 316338 550350 316958 567922
rect 316338 550294 316434 550350
rect 316490 550294 316558 550350
rect 316614 550294 316682 550350
rect 316738 550294 316806 550350
rect 316862 550294 316958 550350
rect 316338 550226 316958 550294
rect 316338 550170 316434 550226
rect 316490 550170 316558 550226
rect 316614 550170 316682 550226
rect 316738 550170 316806 550226
rect 316862 550170 316958 550226
rect 316338 550102 316958 550170
rect 316338 550046 316434 550102
rect 316490 550046 316558 550102
rect 316614 550046 316682 550102
rect 316738 550046 316806 550102
rect 316862 550046 316958 550102
rect 316338 549978 316958 550046
rect 316338 549922 316434 549978
rect 316490 549922 316558 549978
rect 316614 549922 316682 549978
rect 316738 549922 316806 549978
rect 316862 549922 316958 549978
rect 316338 532350 316958 549922
rect 316338 532294 316434 532350
rect 316490 532294 316558 532350
rect 316614 532294 316682 532350
rect 316738 532294 316806 532350
rect 316862 532294 316958 532350
rect 316338 532226 316958 532294
rect 316338 532170 316434 532226
rect 316490 532170 316558 532226
rect 316614 532170 316682 532226
rect 316738 532170 316806 532226
rect 316862 532170 316958 532226
rect 316338 532102 316958 532170
rect 316338 532046 316434 532102
rect 316490 532046 316558 532102
rect 316614 532046 316682 532102
rect 316738 532046 316806 532102
rect 316862 532046 316958 532102
rect 316338 531978 316958 532046
rect 316338 531922 316434 531978
rect 316490 531922 316558 531978
rect 316614 531922 316682 531978
rect 316738 531922 316806 531978
rect 316862 531922 316958 531978
rect 316338 514350 316958 531922
rect 316338 514294 316434 514350
rect 316490 514294 316558 514350
rect 316614 514294 316682 514350
rect 316738 514294 316806 514350
rect 316862 514294 316958 514350
rect 316338 514226 316958 514294
rect 316338 514170 316434 514226
rect 316490 514170 316558 514226
rect 316614 514170 316682 514226
rect 316738 514170 316806 514226
rect 316862 514170 316958 514226
rect 316338 514102 316958 514170
rect 316338 514046 316434 514102
rect 316490 514046 316558 514102
rect 316614 514046 316682 514102
rect 316738 514046 316806 514102
rect 316862 514046 316958 514102
rect 316338 513978 316958 514046
rect 316338 513922 316434 513978
rect 316490 513922 316558 513978
rect 316614 513922 316682 513978
rect 316738 513922 316806 513978
rect 316862 513922 316958 513978
rect 316338 496350 316958 513922
rect 316338 496294 316434 496350
rect 316490 496294 316558 496350
rect 316614 496294 316682 496350
rect 316738 496294 316806 496350
rect 316862 496294 316958 496350
rect 316338 496226 316958 496294
rect 316338 496170 316434 496226
rect 316490 496170 316558 496226
rect 316614 496170 316682 496226
rect 316738 496170 316806 496226
rect 316862 496170 316958 496226
rect 316338 496102 316958 496170
rect 316338 496046 316434 496102
rect 316490 496046 316558 496102
rect 316614 496046 316682 496102
rect 316738 496046 316806 496102
rect 316862 496046 316958 496102
rect 316338 495978 316958 496046
rect 316338 495922 316434 495978
rect 316490 495922 316558 495978
rect 316614 495922 316682 495978
rect 316738 495922 316806 495978
rect 316862 495922 316958 495978
rect 316338 478350 316958 495922
rect 316338 478294 316434 478350
rect 316490 478294 316558 478350
rect 316614 478294 316682 478350
rect 316738 478294 316806 478350
rect 316862 478294 316958 478350
rect 316338 478226 316958 478294
rect 316338 478170 316434 478226
rect 316490 478170 316558 478226
rect 316614 478170 316682 478226
rect 316738 478170 316806 478226
rect 316862 478170 316958 478226
rect 316338 478102 316958 478170
rect 316338 478046 316434 478102
rect 316490 478046 316558 478102
rect 316614 478046 316682 478102
rect 316738 478046 316806 478102
rect 316862 478046 316958 478102
rect 316338 477978 316958 478046
rect 316338 477922 316434 477978
rect 316490 477922 316558 477978
rect 316614 477922 316682 477978
rect 316738 477922 316806 477978
rect 316862 477922 316958 477978
rect 316338 460350 316958 477922
rect 316338 460294 316434 460350
rect 316490 460294 316558 460350
rect 316614 460294 316682 460350
rect 316738 460294 316806 460350
rect 316862 460294 316958 460350
rect 316338 460226 316958 460294
rect 316338 460170 316434 460226
rect 316490 460170 316558 460226
rect 316614 460170 316682 460226
rect 316738 460170 316806 460226
rect 316862 460170 316958 460226
rect 316338 460102 316958 460170
rect 316338 460046 316434 460102
rect 316490 460046 316558 460102
rect 316614 460046 316682 460102
rect 316738 460046 316806 460102
rect 316862 460046 316958 460102
rect 316338 459978 316958 460046
rect 316338 459922 316434 459978
rect 316490 459922 316558 459978
rect 316614 459922 316682 459978
rect 316738 459922 316806 459978
rect 316862 459922 316958 459978
rect 316338 442350 316958 459922
rect 316338 442294 316434 442350
rect 316490 442294 316558 442350
rect 316614 442294 316682 442350
rect 316738 442294 316806 442350
rect 316862 442294 316958 442350
rect 316338 442226 316958 442294
rect 316338 442170 316434 442226
rect 316490 442170 316558 442226
rect 316614 442170 316682 442226
rect 316738 442170 316806 442226
rect 316862 442170 316958 442226
rect 316338 442102 316958 442170
rect 316338 442046 316434 442102
rect 316490 442046 316558 442102
rect 316614 442046 316682 442102
rect 316738 442046 316806 442102
rect 316862 442046 316958 442102
rect 316338 441978 316958 442046
rect 316338 441922 316434 441978
rect 316490 441922 316558 441978
rect 316614 441922 316682 441978
rect 316738 441922 316806 441978
rect 316862 441922 316958 441978
rect 316338 424350 316958 441922
rect 316338 424294 316434 424350
rect 316490 424294 316558 424350
rect 316614 424294 316682 424350
rect 316738 424294 316806 424350
rect 316862 424294 316958 424350
rect 316338 424226 316958 424294
rect 316338 424170 316434 424226
rect 316490 424170 316558 424226
rect 316614 424170 316682 424226
rect 316738 424170 316806 424226
rect 316862 424170 316958 424226
rect 316338 424102 316958 424170
rect 316338 424046 316434 424102
rect 316490 424046 316558 424102
rect 316614 424046 316682 424102
rect 316738 424046 316806 424102
rect 316862 424046 316958 424102
rect 316338 423978 316958 424046
rect 316338 423922 316434 423978
rect 316490 423922 316558 423978
rect 316614 423922 316682 423978
rect 316738 423922 316806 423978
rect 316862 423922 316958 423978
rect 316338 406350 316958 423922
rect 316338 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 316958 406350
rect 316338 406226 316958 406294
rect 316338 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 316958 406226
rect 316338 406102 316958 406170
rect 316338 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 316958 406102
rect 316338 405978 316958 406046
rect 316338 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 316958 405978
rect 316338 388350 316958 405922
rect 316338 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 316958 388350
rect 316338 388226 316958 388294
rect 316338 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 316958 388226
rect 316338 388102 316958 388170
rect 316338 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 316958 388102
rect 316338 387978 316958 388046
rect 316338 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 316958 387978
rect 316338 370350 316958 387922
rect 316338 370294 316434 370350
rect 316490 370294 316558 370350
rect 316614 370294 316682 370350
rect 316738 370294 316806 370350
rect 316862 370294 316958 370350
rect 316338 370226 316958 370294
rect 316338 370170 316434 370226
rect 316490 370170 316558 370226
rect 316614 370170 316682 370226
rect 316738 370170 316806 370226
rect 316862 370170 316958 370226
rect 316338 370102 316958 370170
rect 316338 370046 316434 370102
rect 316490 370046 316558 370102
rect 316614 370046 316682 370102
rect 316738 370046 316806 370102
rect 316862 370046 316958 370102
rect 316338 369978 316958 370046
rect 316338 369922 316434 369978
rect 316490 369922 316558 369978
rect 316614 369922 316682 369978
rect 316738 369922 316806 369978
rect 316862 369922 316958 369978
rect 316338 352350 316958 369922
rect 316338 352294 316434 352350
rect 316490 352294 316558 352350
rect 316614 352294 316682 352350
rect 316738 352294 316806 352350
rect 316862 352294 316958 352350
rect 316338 352226 316958 352294
rect 316338 352170 316434 352226
rect 316490 352170 316558 352226
rect 316614 352170 316682 352226
rect 316738 352170 316806 352226
rect 316862 352170 316958 352226
rect 316338 352102 316958 352170
rect 316338 352046 316434 352102
rect 316490 352046 316558 352102
rect 316614 352046 316682 352102
rect 316738 352046 316806 352102
rect 316862 352046 316958 352102
rect 316338 351978 316958 352046
rect 316338 351922 316434 351978
rect 316490 351922 316558 351978
rect 316614 351922 316682 351978
rect 316738 351922 316806 351978
rect 316862 351922 316958 351978
rect 316338 334350 316958 351922
rect 316338 334294 316434 334350
rect 316490 334294 316558 334350
rect 316614 334294 316682 334350
rect 316738 334294 316806 334350
rect 316862 334294 316958 334350
rect 316338 334226 316958 334294
rect 316338 334170 316434 334226
rect 316490 334170 316558 334226
rect 316614 334170 316682 334226
rect 316738 334170 316806 334226
rect 316862 334170 316958 334226
rect 316338 334102 316958 334170
rect 316338 334046 316434 334102
rect 316490 334046 316558 334102
rect 316614 334046 316682 334102
rect 316738 334046 316806 334102
rect 316862 334046 316958 334102
rect 316338 333978 316958 334046
rect 316338 333922 316434 333978
rect 316490 333922 316558 333978
rect 316614 333922 316682 333978
rect 316738 333922 316806 333978
rect 316862 333922 316958 333978
rect 316338 321718 316958 333922
rect 343338 597212 343958 598268
rect 343338 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 343958 597212
rect 343338 597088 343958 597156
rect 343338 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 343958 597088
rect 343338 596964 343958 597032
rect 343338 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 343958 596964
rect 343338 596840 343958 596908
rect 343338 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 343958 596840
rect 343338 580350 343958 596784
rect 343338 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 343958 580350
rect 343338 580226 343958 580294
rect 343338 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 343958 580226
rect 343338 580102 343958 580170
rect 343338 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 343958 580102
rect 343338 579978 343958 580046
rect 343338 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 343958 579978
rect 343338 562350 343958 579922
rect 343338 562294 343434 562350
rect 343490 562294 343558 562350
rect 343614 562294 343682 562350
rect 343738 562294 343806 562350
rect 343862 562294 343958 562350
rect 343338 562226 343958 562294
rect 343338 562170 343434 562226
rect 343490 562170 343558 562226
rect 343614 562170 343682 562226
rect 343738 562170 343806 562226
rect 343862 562170 343958 562226
rect 343338 562102 343958 562170
rect 343338 562046 343434 562102
rect 343490 562046 343558 562102
rect 343614 562046 343682 562102
rect 343738 562046 343806 562102
rect 343862 562046 343958 562102
rect 343338 561978 343958 562046
rect 343338 561922 343434 561978
rect 343490 561922 343558 561978
rect 343614 561922 343682 561978
rect 343738 561922 343806 561978
rect 343862 561922 343958 561978
rect 343338 544350 343958 561922
rect 343338 544294 343434 544350
rect 343490 544294 343558 544350
rect 343614 544294 343682 544350
rect 343738 544294 343806 544350
rect 343862 544294 343958 544350
rect 343338 544226 343958 544294
rect 343338 544170 343434 544226
rect 343490 544170 343558 544226
rect 343614 544170 343682 544226
rect 343738 544170 343806 544226
rect 343862 544170 343958 544226
rect 343338 544102 343958 544170
rect 343338 544046 343434 544102
rect 343490 544046 343558 544102
rect 343614 544046 343682 544102
rect 343738 544046 343806 544102
rect 343862 544046 343958 544102
rect 343338 543978 343958 544046
rect 343338 543922 343434 543978
rect 343490 543922 343558 543978
rect 343614 543922 343682 543978
rect 343738 543922 343806 543978
rect 343862 543922 343958 543978
rect 343338 526350 343958 543922
rect 343338 526294 343434 526350
rect 343490 526294 343558 526350
rect 343614 526294 343682 526350
rect 343738 526294 343806 526350
rect 343862 526294 343958 526350
rect 343338 526226 343958 526294
rect 343338 526170 343434 526226
rect 343490 526170 343558 526226
rect 343614 526170 343682 526226
rect 343738 526170 343806 526226
rect 343862 526170 343958 526226
rect 343338 526102 343958 526170
rect 343338 526046 343434 526102
rect 343490 526046 343558 526102
rect 343614 526046 343682 526102
rect 343738 526046 343806 526102
rect 343862 526046 343958 526102
rect 343338 525978 343958 526046
rect 343338 525922 343434 525978
rect 343490 525922 343558 525978
rect 343614 525922 343682 525978
rect 343738 525922 343806 525978
rect 343862 525922 343958 525978
rect 343338 508350 343958 525922
rect 343338 508294 343434 508350
rect 343490 508294 343558 508350
rect 343614 508294 343682 508350
rect 343738 508294 343806 508350
rect 343862 508294 343958 508350
rect 343338 508226 343958 508294
rect 343338 508170 343434 508226
rect 343490 508170 343558 508226
rect 343614 508170 343682 508226
rect 343738 508170 343806 508226
rect 343862 508170 343958 508226
rect 343338 508102 343958 508170
rect 343338 508046 343434 508102
rect 343490 508046 343558 508102
rect 343614 508046 343682 508102
rect 343738 508046 343806 508102
rect 343862 508046 343958 508102
rect 343338 507978 343958 508046
rect 343338 507922 343434 507978
rect 343490 507922 343558 507978
rect 343614 507922 343682 507978
rect 343738 507922 343806 507978
rect 343862 507922 343958 507978
rect 343338 490350 343958 507922
rect 343338 490294 343434 490350
rect 343490 490294 343558 490350
rect 343614 490294 343682 490350
rect 343738 490294 343806 490350
rect 343862 490294 343958 490350
rect 343338 490226 343958 490294
rect 343338 490170 343434 490226
rect 343490 490170 343558 490226
rect 343614 490170 343682 490226
rect 343738 490170 343806 490226
rect 343862 490170 343958 490226
rect 343338 490102 343958 490170
rect 343338 490046 343434 490102
rect 343490 490046 343558 490102
rect 343614 490046 343682 490102
rect 343738 490046 343806 490102
rect 343862 490046 343958 490102
rect 343338 489978 343958 490046
rect 343338 489922 343434 489978
rect 343490 489922 343558 489978
rect 343614 489922 343682 489978
rect 343738 489922 343806 489978
rect 343862 489922 343958 489978
rect 343338 472350 343958 489922
rect 343338 472294 343434 472350
rect 343490 472294 343558 472350
rect 343614 472294 343682 472350
rect 343738 472294 343806 472350
rect 343862 472294 343958 472350
rect 343338 472226 343958 472294
rect 343338 472170 343434 472226
rect 343490 472170 343558 472226
rect 343614 472170 343682 472226
rect 343738 472170 343806 472226
rect 343862 472170 343958 472226
rect 343338 472102 343958 472170
rect 343338 472046 343434 472102
rect 343490 472046 343558 472102
rect 343614 472046 343682 472102
rect 343738 472046 343806 472102
rect 343862 472046 343958 472102
rect 343338 471978 343958 472046
rect 343338 471922 343434 471978
rect 343490 471922 343558 471978
rect 343614 471922 343682 471978
rect 343738 471922 343806 471978
rect 343862 471922 343958 471978
rect 343338 454350 343958 471922
rect 343338 454294 343434 454350
rect 343490 454294 343558 454350
rect 343614 454294 343682 454350
rect 343738 454294 343806 454350
rect 343862 454294 343958 454350
rect 343338 454226 343958 454294
rect 343338 454170 343434 454226
rect 343490 454170 343558 454226
rect 343614 454170 343682 454226
rect 343738 454170 343806 454226
rect 343862 454170 343958 454226
rect 343338 454102 343958 454170
rect 343338 454046 343434 454102
rect 343490 454046 343558 454102
rect 343614 454046 343682 454102
rect 343738 454046 343806 454102
rect 343862 454046 343958 454102
rect 343338 453978 343958 454046
rect 343338 453922 343434 453978
rect 343490 453922 343558 453978
rect 343614 453922 343682 453978
rect 343738 453922 343806 453978
rect 343862 453922 343958 453978
rect 343338 436350 343958 453922
rect 343338 436294 343434 436350
rect 343490 436294 343558 436350
rect 343614 436294 343682 436350
rect 343738 436294 343806 436350
rect 343862 436294 343958 436350
rect 343338 436226 343958 436294
rect 343338 436170 343434 436226
rect 343490 436170 343558 436226
rect 343614 436170 343682 436226
rect 343738 436170 343806 436226
rect 343862 436170 343958 436226
rect 343338 436102 343958 436170
rect 343338 436046 343434 436102
rect 343490 436046 343558 436102
rect 343614 436046 343682 436102
rect 343738 436046 343806 436102
rect 343862 436046 343958 436102
rect 343338 435978 343958 436046
rect 343338 435922 343434 435978
rect 343490 435922 343558 435978
rect 343614 435922 343682 435978
rect 343738 435922 343806 435978
rect 343862 435922 343958 435978
rect 343338 418350 343958 435922
rect 343338 418294 343434 418350
rect 343490 418294 343558 418350
rect 343614 418294 343682 418350
rect 343738 418294 343806 418350
rect 343862 418294 343958 418350
rect 343338 418226 343958 418294
rect 343338 418170 343434 418226
rect 343490 418170 343558 418226
rect 343614 418170 343682 418226
rect 343738 418170 343806 418226
rect 343862 418170 343958 418226
rect 343338 418102 343958 418170
rect 343338 418046 343434 418102
rect 343490 418046 343558 418102
rect 343614 418046 343682 418102
rect 343738 418046 343806 418102
rect 343862 418046 343958 418102
rect 343338 417978 343958 418046
rect 343338 417922 343434 417978
rect 343490 417922 343558 417978
rect 343614 417922 343682 417978
rect 343738 417922 343806 417978
rect 343862 417922 343958 417978
rect 343338 400350 343958 417922
rect 343338 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 343958 400350
rect 343338 400226 343958 400294
rect 343338 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 343958 400226
rect 343338 400102 343958 400170
rect 343338 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 343958 400102
rect 343338 399978 343958 400046
rect 343338 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 343958 399978
rect 343338 382350 343958 399922
rect 343338 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 343958 382350
rect 343338 382226 343958 382294
rect 343338 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 343958 382226
rect 343338 382102 343958 382170
rect 343338 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 343958 382102
rect 343338 381978 343958 382046
rect 343338 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 343958 381978
rect 343338 364350 343958 381922
rect 343338 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 343958 364350
rect 343338 364226 343958 364294
rect 343338 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 343958 364226
rect 343338 364102 343958 364170
rect 343338 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 343958 364102
rect 343338 363978 343958 364046
rect 343338 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 343958 363978
rect 343338 346350 343958 363922
rect 343338 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 343958 346350
rect 343338 346226 343958 346294
rect 343338 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 343958 346226
rect 343338 346102 343958 346170
rect 343338 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 343958 346102
rect 343338 345978 343958 346046
rect 343338 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 343958 345978
rect 343338 328350 343958 345922
rect 343338 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 343958 328350
rect 343338 328226 343958 328294
rect 343338 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 343958 328226
rect 343338 328102 343958 328170
rect 343338 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 343958 328102
rect 343338 327978 343958 328046
rect 343338 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 343958 327978
rect 343338 321718 343958 327922
rect 347058 598172 347678 598268
rect 347058 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 347678 598172
rect 347058 598048 347678 598116
rect 347058 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 347678 598048
rect 347058 597924 347678 597992
rect 347058 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 347678 597924
rect 347058 597800 347678 597868
rect 347058 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 347678 597800
rect 347058 586350 347678 597744
rect 347058 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 347678 586350
rect 347058 586226 347678 586294
rect 347058 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 347678 586226
rect 347058 586102 347678 586170
rect 347058 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 347678 586102
rect 347058 585978 347678 586046
rect 347058 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 347678 585978
rect 347058 568350 347678 585922
rect 347058 568294 347154 568350
rect 347210 568294 347278 568350
rect 347334 568294 347402 568350
rect 347458 568294 347526 568350
rect 347582 568294 347678 568350
rect 347058 568226 347678 568294
rect 347058 568170 347154 568226
rect 347210 568170 347278 568226
rect 347334 568170 347402 568226
rect 347458 568170 347526 568226
rect 347582 568170 347678 568226
rect 347058 568102 347678 568170
rect 347058 568046 347154 568102
rect 347210 568046 347278 568102
rect 347334 568046 347402 568102
rect 347458 568046 347526 568102
rect 347582 568046 347678 568102
rect 347058 567978 347678 568046
rect 347058 567922 347154 567978
rect 347210 567922 347278 567978
rect 347334 567922 347402 567978
rect 347458 567922 347526 567978
rect 347582 567922 347678 567978
rect 347058 550350 347678 567922
rect 347058 550294 347154 550350
rect 347210 550294 347278 550350
rect 347334 550294 347402 550350
rect 347458 550294 347526 550350
rect 347582 550294 347678 550350
rect 347058 550226 347678 550294
rect 347058 550170 347154 550226
rect 347210 550170 347278 550226
rect 347334 550170 347402 550226
rect 347458 550170 347526 550226
rect 347582 550170 347678 550226
rect 347058 550102 347678 550170
rect 347058 550046 347154 550102
rect 347210 550046 347278 550102
rect 347334 550046 347402 550102
rect 347458 550046 347526 550102
rect 347582 550046 347678 550102
rect 347058 549978 347678 550046
rect 347058 549922 347154 549978
rect 347210 549922 347278 549978
rect 347334 549922 347402 549978
rect 347458 549922 347526 549978
rect 347582 549922 347678 549978
rect 347058 532350 347678 549922
rect 347058 532294 347154 532350
rect 347210 532294 347278 532350
rect 347334 532294 347402 532350
rect 347458 532294 347526 532350
rect 347582 532294 347678 532350
rect 347058 532226 347678 532294
rect 347058 532170 347154 532226
rect 347210 532170 347278 532226
rect 347334 532170 347402 532226
rect 347458 532170 347526 532226
rect 347582 532170 347678 532226
rect 347058 532102 347678 532170
rect 347058 532046 347154 532102
rect 347210 532046 347278 532102
rect 347334 532046 347402 532102
rect 347458 532046 347526 532102
rect 347582 532046 347678 532102
rect 347058 531978 347678 532046
rect 347058 531922 347154 531978
rect 347210 531922 347278 531978
rect 347334 531922 347402 531978
rect 347458 531922 347526 531978
rect 347582 531922 347678 531978
rect 347058 514350 347678 531922
rect 347058 514294 347154 514350
rect 347210 514294 347278 514350
rect 347334 514294 347402 514350
rect 347458 514294 347526 514350
rect 347582 514294 347678 514350
rect 347058 514226 347678 514294
rect 347058 514170 347154 514226
rect 347210 514170 347278 514226
rect 347334 514170 347402 514226
rect 347458 514170 347526 514226
rect 347582 514170 347678 514226
rect 347058 514102 347678 514170
rect 347058 514046 347154 514102
rect 347210 514046 347278 514102
rect 347334 514046 347402 514102
rect 347458 514046 347526 514102
rect 347582 514046 347678 514102
rect 347058 513978 347678 514046
rect 347058 513922 347154 513978
rect 347210 513922 347278 513978
rect 347334 513922 347402 513978
rect 347458 513922 347526 513978
rect 347582 513922 347678 513978
rect 347058 496350 347678 513922
rect 347058 496294 347154 496350
rect 347210 496294 347278 496350
rect 347334 496294 347402 496350
rect 347458 496294 347526 496350
rect 347582 496294 347678 496350
rect 347058 496226 347678 496294
rect 347058 496170 347154 496226
rect 347210 496170 347278 496226
rect 347334 496170 347402 496226
rect 347458 496170 347526 496226
rect 347582 496170 347678 496226
rect 347058 496102 347678 496170
rect 347058 496046 347154 496102
rect 347210 496046 347278 496102
rect 347334 496046 347402 496102
rect 347458 496046 347526 496102
rect 347582 496046 347678 496102
rect 347058 495978 347678 496046
rect 347058 495922 347154 495978
rect 347210 495922 347278 495978
rect 347334 495922 347402 495978
rect 347458 495922 347526 495978
rect 347582 495922 347678 495978
rect 347058 478350 347678 495922
rect 347058 478294 347154 478350
rect 347210 478294 347278 478350
rect 347334 478294 347402 478350
rect 347458 478294 347526 478350
rect 347582 478294 347678 478350
rect 347058 478226 347678 478294
rect 347058 478170 347154 478226
rect 347210 478170 347278 478226
rect 347334 478170 347402 478226
rect 347458 478170 347526 478226
rect 347582 478170 347678 478226
rect 347058 478102 347678 478170
rect 347058 478046 347154 478102
rect 347210 478046 347278 478102
rect 347334 478046 347402 478102
rect 347458 478046 347526 478102
rect 347582 478046 347678 478102
rect 347058 477978 347678 478046
rect 347058 477922 347154 477978
rect 347210 477922 347278 477978
rect 347334 477922 347402 477978
rect 347458 477922 347526 477978
rect 347582 477922 347678 477978
rect 347058 460350 347678 477922
rect 347058 460294 347154 460350
rect 347210 460294 347278 460350
rect 347334 460294 347402 460350
rect 347458 460294 347526 460350
rect 347582 460294 347678 460350
rect 347058 460226 347678 460294
rect 347058 460170 347154 460226
rect 347210 460170 347278 460226
rect 347334 460170 347402 460226
rect 347458 460170 347526 460226
rect 347582 460170 347678 460226
rect 347058 460102 347678 460170
rect 347058 460046 347154 460102
rect 347210 460046 347278 460102
rect 347334 460046 347402 460102
rect 347458 460046 347526 460102
rect 347582 460046 347678 460102
rect 347058 459978 347678 460046
rect 347058 459922 347154 459978
rect 347210 459922 347278 459978
rect 347334 459922 347402 459978
rect 347458 459922 347526 459978
rect 347582 459922 347678 459978
rect 347058 442350 347678 459922
rect 347058 442294 347154 442350
rect 347210 442294 347278 442350
rect 347334 442294 347402 442350
rect 347458 442294 347526 442350
rect 347582 442294 347678 442350
rect 347058 442226 347678 442294
rect 347058 442170 347154 442226
rect 347210 442170 347278 442226
rect 347334 442170 347402 442226
rect 347458 442170 347526 442226
rect 347582 442170 347678 442226
rect 347058 442102 347678 442170
rect 347058 442046 347154 442102
rect 347210 442046 347278 442102
rect 347334 442046 347402 442102
rect 347458 442046 347526 442102
rect 347582 442046 347678 442102
rect 347058 441978 347678 442046
rect 347058 441922 347154 441978
rect 347210 441922 347278 441978
rect 347334 441922 347402 441978
rect 347458 441922 347526 441978
rect 347582 441922 347678 441978
rect 347058 424350 347678 441922
rect 347058 424294 347154 424350
rect 347210 424294 347278 424350
rect 347334 424294 347402 424350
rect 347458 424294 347526 424350
rect 347582 424294 347678 424350
rect 347058 424226 347678 424294
rect 347058 424170 347154 424226
rect 347210 424170 347278 424226
rect 347334 424170 347402 424226
rect 347458 424170 347526 424226
rect 347582 424170 347678 424226
rect 347058 424102 347678 424170
rect 347058 424046 347154 424102
rect 347210 424046 347278 424102
rect 347334 424046 347402 424102
rect 347458 424046 347526 424102
rect 347582 424046 347678 424102
rect 347058 423978 347678 424046
rect 347058 423922 347154 423978
rect 347210 423922 347278 423978
rect 347334 423922 347402 423978
rect 347458 423922 347526 423978
rect 347582 423922 347678 423978
rect 347058 406350 347678 423922
rect 347058 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 347678 406350
rect 347058 406226 347678 406294
rect 347058 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 347678 406226
rect 347058 406102 347678 406170
rect 347058 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 347678 406102
rect 347058 405978 347678 406046
rect 347058 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 347678 405978
rect 347058 388350 347678 405922
rect 347058 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 347678 388350
rect 347058 388226 347678 388294
rect 347058 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 347678 388226
rect 347058 388102 347678 388170
rect 347058 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 347678 388102
rect 347058 387978 347678 388046
rect 347058 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 347678 387978
rect 347058 370350 347678 387922
rect 347058 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 347678 370350
rect 347058 370226 347678 370294
rect 347058 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 347678 370226
rect 347058 370102 347678 370170
rect 347058 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 347678 370102
rect 347058 369978 347678 370046
rect 347058 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 347678 369978
rect 347058 352350 347678 369922
rect 347058 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 347678 352350
rect 347058 352226 347678 352294
rect 347058 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 347678 352226
rect 347058 352102 347678 352170
rect 347058 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 347678 352102
rect 347058 351978 347678 352046
rect 347058 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 347678 351978
rect 347058 334350 347678 351922
rect 347058 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 347678 334350
rect 347058 334226 347678 334294
rect 347058 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 347678 334226
rect 347058 334102 347678 334170
rect 347058 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 347678 334102
rect 347058 333978 347678 334046
rect 347058 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 347678 333978
rect 347058 321718 347678 333922
rect 374058 597212 374678 598268
rect 374058 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 374678 597212
rect 374058 597088 374678 597156
rect 374058 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 374678 597088
rect 374058 596964 374678 597032
rect 374058 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 374678 596964
rect 374058 596840 374678 596908
rect 374058 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 374678 596840
rect 374058 580350 374678 596784
rect 374058 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 374678 580350
rect 374058 580226 374678 580294
rect 374058 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 374678 580226
rect 374058 580102 374678 580170
rect 374058 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 374678 580102
rect 374058 579978 374678 580046
rect 374058 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 374678 579978
rect 374058 562350 374678 579922
rect 374058 562294 374154 562350
rect 374210 562294 374278 562350
rect 374334 562294 374402 562350
rect 374458 562294 374526 562350
rect 374582 562294 374678 562350
rect 374058 562226 374678 562294
rect 374058 562170 374154 562226
rect 374210 562170 374278 562226
rect 374334 562170 374402 562226
rect 374458 562170 374526 562226
rect 374582 562170 374678 562226
rect 374058 562102 374678 562170
rect 374058 562046 374154 562102
rect 374210 562046 374278 562102
rect 374334 562046 374402 562102
rect 374458 562046 374526 562102
rect 374582 562046 374678 562102
rect 374058 561978 374678 562046
rect 374058 561922 374154 561978
rect 374210 561922 374278 561978
rect 374334 561922 374402 561978
rect 374458 561922 374526 561978
rect 374582 561922 374678 561978
rect 374058 544350 374678 561922
rect 374058 544294 374154 544350
rect 374210 544294 374278 544350
rect 374334 544294 374402 544350
rect 374458 544294 374526 544350
rect 374582 544294 374678 544350
rect 374058 544226 374678 544294
rect 374058 544170 374154 544226
rect 374210 544170 374278 544226
rect 374334 544170 374402 544226
rect 374458 544170 374526 544226
rect 374582 544170 374678 544226
rect 374058 544102 374678 544170
rect 374058 544046 374154 544102
rect 374210 544046 374278 544102
rect 374334 544046 374402 544102
rect 374458 544046 374526 544102
rect 374582 544046 374678 544102
rect 374058 543978 374678 544046
rect 374058 543922 374154 543978
rect 374210 543922 374278 543978
rect 374334 543922 374402 543978
rect 374458 543922 374526 543978
rect 374582 543922 374678 543978
rect 374058 526350 374678 543922
rect 374058 526294 374154 526350
rect 374210 526294 374278 526350
rect 374334 526294 374402 526350
rect 374458 526294 374526 526350
rect 374582 526294 374678 526350
rect 374058 526226 374678 526294
rect 374058 526170 374154 526226
rect 374210 526170 374278 526226
rect 374334 526170 374402 526226
rect 374458 526170 374526 526226
rect 374582 526170 374678 526226
rect 374058 526102 374678 526170
rect 374058 526046 374154 526102
rect 374210 526046 374278 526102
rect 374334 526046 374402 526102
rect 374458 526046 374526 526102
rect 374582 526046 374678 526102
rect 374058 525978 374678 526046
rect 374058 525922 374154 525978
rect 374210 525922 374278 525978
rect 374334 525922 374402 525978
rect 374458 525922 374526 525978
rect 374582 525922 374678 525978
rect 374058 508350 374678 525922
rect 374058 508294 374154 508350
rect 374210 508294 374278 508350
rect 374334 508294 374402 508350
rect 374458 508294 374526 508350
rect 374582 508294 374678 508350
rect 374058 508226 374678 508294
rect 374058 508170 374154 508226
rect 374210 508170 374278 508226
rect 374334 508170 374402 508226
rect 374458 508170 374526 508226
rect 374582 508170 374678 508226
rect 374058 508102 374678 508170
rect 374058 508046 374154 508102
rect 374210 508046 374278 508102
rect 374334 508046 374402 508102
rect 374458 508046 374526 508102
rect 374582 508046 374678 508102
rect 374058 507978 374678 508046
rect 374058 507922 374154 507978
rect 374210 507922 374278 507978
rect 374334 507922 374402 507978
rect 374458 507922 374526 507978
rect 374582 507922 374678 507978
rect 374058 490350 374678 507922
rect 374058 490294 374154 490350
rect 374210 490294 374278 490350
rect 374334 490294 374402 490350
rect 374458 490294 374526 490350
rect 374582 490294 374678 490350
rect 374058 490226 374678 490294
rect 374058 490170 374154 490226
rect 374210 490170 374278 490226
rect 374334 490170 374402 490226
rect 374458 490170 374526 490226
rect 374582 490170 374678 490226
rect 374058 490102 374678 490170
rect 374058 490046 374154 490102
rect 374210 490046 374278 490102
rect 374334 490046 374402 490102
rect 374458 490046 374526 490102
rect 374582 490046 374678 490102
rect 374058 489978 374678 490046
rect 374058 489922 374154 489978
rect 374210 489922 374278 489978
rect 374334 489922 374402 489978
rect 374458 489922 374526 489978
rect 374582 489922 374678 489978
rect 374058 472350 374678 489922
rect 374058 472294 374154 472350
rect 374210 472294 374278 472350
rect 374334 472294 374402 472350
rect 374458 472294 374526 472350
rect 374582 472294 374678 472350
rect 374058 472226 374678 472294
rect 374058 472170 374154 472226
rect 374210 472170 374278 472226
rect 374334 472170 374402 472226
rect 374458 472170 374526 472226
rect 374582 472170 374678 472226
rect 374058 472102 374678 472170
rect 374058 472046 374154 472102
rect 374210 472046 374278 472102
rect 374334 472046 374402 472102
rect 374458 472046 374526 472102
rect 374582 472046 374678 472102
rect 374058 471978 374678 472046
rect 374058 471922 374154 471978
rect 374210 471922 374278 471978
rect 374334 471922 374402 471978
rect 374458 471922 374526 471978
rect 374582 471922 374678 471978
rect 374058 454350 374678 471922
rect 374058 454294 374154 454350
rect 374210 454294 374278 454350
rect 374334 454294 374402 454350
rect 374458 454294 374526 454350
rect 374582 454294 374678 454350
rect 374058 454226 374678 454294
rect 374058 454170 374154 454226
rect 374210 454170 374278 454226
rect 374334 454170 374402 454226
rect 374458 454170 374526 454226
rect 374582 454170 374678 454226
rect 374058 454102 374678 454170
rect 374058 454046 374154 454102
rect 374210 454046 374278 454102
rect 374334 454046 374402 454102
rect 374458 454046 374526 454102
rect 374582 454046 374678 454102
rect 374058 453978 374678 454046
rect 374058 453922 374154 453978
rect 374210 453922 374278 453978
rect 374334 453922 374402 453978
rect 374458 453922 374526 453978
rect 374582 453922 374678 453978
rect 374058 436350 374678 453922
rect 374058 436294 374154 436350
rect 374210 436294 374278 436350
rect 374334 436294 374402 436350
rect 374458 436294 374526 436350
rect 374582 436294 374678 436350
rect 374058 436226 374678 436294
rect 374058 436170 374154 436226
rect 374210 436170 374278 436226
rect 374334 436170 374402 436226
rect 374458 436170 374526 436226
rect 374582 436170 374678 436226
rect 374058 436102 374678 436170
rect 374058 436046 374154 436102
rect 374210 436046 374278 436102
rect 374334 436046 374402 436102
rect 374458 436046 374526 436102
rect 374582 436046 374678 436102
rect 374058 435978 374678 436046
rect 374058 435922 374154 435978
rect 374210 435922 374278 435978
rect 374334 435922 374402 435978
rect 374458 435922 374526 435978
rect 374582 435922 374678 435978
rect 374058 418350 374678 435922
rect 374058 418294 374154 418350
rect 374210 418294 374278 418350
rect 374334 418294 374402 418350
rect 374458 418294 374526 418350
rect 374582 418294 374678 418350
rect 374058 418226 374678 418294
rect 374058 418170 374154 418226
rect 374210 418170 374278 418226
rect 374334 418170 374402 418226
rect 374458 418170 374526 418226
rect 374582 418170 374678 418226
rect 374058 418102 374678 418170
rect 374058 418046 374154 418102
rect 374210 418046 374278 418102
rect 374334 418046 374402 418102
rect 374458 418046 374526 418102
rect 374582 418046 374678 418102
rect 374058 417978 374678 418046
rect 374058 417922 374154 417978
rect 374210 417922 374278 417978
rect 374334 417922 374402 417978
rect 374458 417922 374526 417978
rect 374582 417922 374678 417978
rect 374058 400350 374678 417922
rect 374058 400294 374154 400350
rect 374210 400294 374278 400350
rect 374334 400294 374402 400350
rect 374458 400294 374526 400350
rect 374582 400294 374678 400350
rect 374058 400226 374678 400294
rect 374058 400170 374154 400226
rect 374210 400170 374278 400226
rect 374334 400170 374402 400226
rect 374458 400170 374526 400226
rect 374582 400170 374678 400226
rect 374058 400102 374678 400170
rect 374058 400046 374154 400102
rect 374210 400046 374278 400102
rect 374334 400046 374402 400102
rect 374458 400046 374526 400102
rect 374582 400046 374678 400102
rect 374058 399978 374678 400046
rect 374058 399922 374154 399978
rect 374210 399922 374278 399978
rect 374334 399922 374402 399978
rect 374458 399922 374526 399978
rect 374582 399922 374678 399978
rect 374058 382350 374678 399922
rect 374058 382294 374154 382350
rect 374210 382294 374278 382350
rect 374334 382294 374402 382350
rect 374458 382294 374526 382350
rect 374582 382294 374678 382350
rect 374058 382226 374678 382294
rect 374058 382170 374154 382226
rect 374210 382170 374278 382226
rect 374334 382170 374402 382226
rect 374458 382170 374526 382226
rect 374582 382170 374678 382226
rect 374058 382102 374678 382170
rect 374058 382046 374154 382102
rect 374210 382046 374278 382102
rect 374334 382046 374402 382102
rect 374458 382046 374526 382102
rect 374582 382046 374678 382102
rect 374058 381978 374678 382046
rect 374058 381922 374154 381978
rect 374210 381922 374278 381978
rect 374334 381922 374402 381978
rect 374458 381922 374526 381978
rect 374582 381922 374678 381978
rect 374058 364350 374678 381922
rect 374058 364294 374154 364350
rect 374210 364294 374278 364350
rect 374334 364294 374402 364350
rect 374458 364294 374526 364350
rect 374582 364294 374678 364350
rect 374058 364226 374678 364294
rect 374058 364170 374154 364226
rect 374210 364170 374278 364226
rect 374334 364170 374402 364226
rect 374458 364170 374526 364226
rect 374582 364170 374678 364226
rect 374058 364102 374678 364170
rect 374058 364046 374154 364102
rect 374210 364046 374278 364102
rect 374334 364046 374402 364102
rect 374458 364046 374526 364102
rect 374582 364046 374678 364102
rect 374058 363978 374678 364046
rect 374058 363922 374154 363978
rect 374210 363922 374278 363978
rect 374334 363922 374402 363978
rect 374458 363922 374526 363978
rect 374582 363922 374678 363978
rect 374058 346350 374678 363922
rect 374058 346294 374154 346350
rect 374210 346294 374278 346350
rect 374334 346294 374402 346350
rect 374458 346294 374526 346350
rect 374582 346294 374678 346350
rect 374058 346226 374678 346294
rect 374058 346170 374154 346226
rect 374210 346170 374278 346226
rect 374334 346170 374402 346226
rect 374458 346170 374526 346226
rect 374582 346170 374678 346226
rect 374058 346102 374678 346170
rect 374058 346046 374154 346102
rect 374210 346046 374278 346102
rect 374334 346046 374402 346102
rect 374458 346046 374526 346102
rect 374582 346046 374678 346102
rect 374058 345978 374678 346046
rect 374058 345922 374154 345978
rect 374210 345922 374278 345978
rect 374334 345922 374402 345978
rect 374458 345922 374526 345978
rect 374582 345922 374678 345978
rect 374058 328350 374678 345922
rect 374058 328294 374154 328350
rect 374210 328294 374278 328350
rect 374334 328294 374402 328350
rect 374458 328294 374526 328350
rect 374582 328294 374678 328350
rect 374058 328226 374678 328294
rect 374058 328170 374154 328226
rect 374210 328170 374278 328226
rect 374334 328170 374402 328226
rect 374458 328170 374526 328226
rect 374582 328170 374678 328226
rect 374058 328102 374678 328170
rect 374058 328046 374154 328102
rect 374210 328046 374278 328102
rect 374334 328046 374402 328102
rect 374458 328046 374526 328102
rect 374582 328046 374678 328102
rect 374058 327978 374678 328046
rect 374058 327922 374154 327978
rect 374210 327922 374278 327978
rect 374334 327922 374402 327978
rect 374458 327922 374526 327978
rect 374582 327922 374678 327978
rect 370636 327684 370692 327694
rect 229808 316350 230128 316384
rect 229808 316294 229878 316350
rect 229934 316294 230002 316350
rect 230058 316294 230128 316350
rect 229808 316226 230128 316294
rect 229808 316170 229878 316226
rect 229934 316170 230002 316226
rect 230058 316170 230128 316226
rect 229808 316102 230128 316170
rect 229808 316046 229878 316102
rect 229934 316046 230002 316102
rect 230058 316046 230128 316102
rect 229808 315978 230128 316046
rect 229808 315922 229878 315978
rect 229934 315922 230002 315978
rect 230058 315922 230128 315978
rect 229808 315888 230128 315922
rect 260528 316350 260848 316384
rect 260528 316294 260598 316350
rect 260654 316294 260722 316350
rect 260778 316294 260848 316350
rect 260528 316226 260848 316294
rect 260528 316170 260598 316226
rect 260654 316170 260722 316226
rect 260778 316170 260848 316226
rect 260528 316102 260848 316170
rect 260528 316046 260598 316102
rect 260654 316046 260722 316102
rect 260778 316046 260848 316102
rect 260528 315978 260848 316046
rect 260528 315922 260598 315978
rect 260654 315922 260722 315978
rect 260778 315922 260848 315978
rect 260528 315888 260848 315922
rect 291248 316350 291568 316384
rect 291248 316294 291318 316350
rect 291374 316294 291442 316350
rect 291498 316294 291568 316350
rect 291248 316226 291568 316294
rect 291248 316170 291318 316226
rect 291374 316170 291442 316226
rect 291498 316170 291568 316226
rect 291248 316102 291568 316170
rect 291248 316046 291318 316102
rect 291374 316046 291442 316102
rect 291498 316046 291568 316102
rect 291248 315978 291568 316046
rect 291248 315922 291318 315978
rect 291374 315922 291442 315978
rect 291498 315922 291568 315978
rect 291248 315888 291568 315922
rect 321968 316350 322288 316384
rect 321968 316294 322038 316350
rect 322094 316294 322162 316350
rect 322218 316294 322288 316350
rect 321968 316226 322288 316294
rect 321968 316170 322038 316226
rect 322094 316170 322162 316226
rect 322218 316170 322288 316226
rect 321968 316102 322288 316170
rect 321968 316046 322038 316102
rect 322094 316046 322162 316102
rect 322218 316046 322288 316102
rect 321968 315978 322288 316046
rect 321968 315922 322038 315978
rect 322094 315922 322162 315978
rect 322218 315922 322288 315978
rect 321968 315888 322288 315922
rect 352688 316350 353008 316384
rect 352688 316294 352758 316350
rect 352814 316294 352882 316350
rect 352938 316294 353008 316350
rect 352688 316226 353008 316294
rect 352688 316170 352758 316226
rect 352814 316170 352882 316226
rect 352938 316170 353008 316226
rect 352688 316102 353008 316170
rect 352688 316046 352758 316102
rect 352814 316046 352882 316102
rect 352938 316046 353008 316102
rect 352688 315978 353008 316046
rect 352688 315922 352758 315978
rect 352814 315922 352882 315978
rect 352938 315922 353008 315978
rect 352688 315888 353008 315922
rect 214448 310350 214768 310384
rect 214448 310294 214518 310350
rect 214574 310294 214642 310350
rect 214698 310294 214768 310350
rect 214448 310226 214768 310294
rect 214448 310170 214518 310226
rect 214574 310170 214642 310226
rect 214698 310170 214768 310226
rect 214448 310102 214768 310170
rect 214448 310046 214518 310102
rect 214574 310046 214642 310102
rect 214698 310046 214768 310102
rect 214448 309978 214768 310046
rect 214448 309922 214518 309978
rect 214574 309922 214642 309978
rect 214698 309922 214768 309978
rect 214448 309888 214768 309922
rect 245168 310350 245488 310384
rect 245168 310294 245238 310350
rect 245294 310294 245362 310350
rect 245418 310294 245488 310350
rect 245168 310226 245488 310294
rect 245168 310170 245238 310226
rect 245294 310170 245362 310226
rect 245418 310170 245488 310226
rect 245168 310102 245488 310170
rect 245168 310046 245238 310102
rect 245294 310046 245362 310102
rect 245418 310046 245488 310102
rect 245168 309978 245488 310046
rect 245168 309922 245238 309978
rect 245294 309922 245362 309978
rect 245418 309922 245488 309978
rect 245168 309888 245488 309922
rect 275888 310350 276208 310384
rect 275888 310294 275958 310350
rect 276014 310294 276082 310350
rect 276138 310294 276208 310350
rect 275888 310226 276208 310294
rect 275888 310170 275958 310226
rect 276014 310170 276082 310226
rect 276138 310170 276208 310226
rect 275888 310102 276208 310170
rect 275888 310046 275958 310102
rect 276014 310046 276082 310102
rect 276138 310046 276208 310102
rect 275888 309978 276208 310046
rect 275888 309922 275958 309978
rect 276014 309922 276082 309978
rect 276138 309922 276208 309978
rect 275888 309888 276208 309922
rect 306608 310350 306928 310384
rect 306608 310294 306678 310350
rect 306734 310294 306802 310350
rect 306858 310294 306928 310350
rect 306608 310226 306928 310294
rect 306608 310170 306678 310226
rect 306734 310170 306802 310226
rect 306858 310170 306928 310226
rect 306608 310102 306928 310170
rect 306608 310046 306678 310102
rect 306734 310046 306802 310102
rect 306858 310046 306928 310102
rect 306608 309978 306928 310046
rect 306608 309922 306678 309978
rect 306734 309922 306802 309978
rect 306858 309922 306928 309978
rect 306608 309888 306928 309922
rect 337328 310350 337648 310384
rect 337328 310294 337398 310350
rect 337454 310294 337522 310350
rect 337578 310294 337648 310350
rect 337328 310226 337648 310294
rect 337328 310170 337398 310226
rect 337454 310170 337522 310226
rect 337578 310170 337648 310226
rect 337328 310102 337648 310170
rect 337328 310046 337398 310102
rect 337454 310046 337522 310102
rect 337578 310046 337648 310102
rect 337328 309978 337648 310046
rect 337328 309922 337398 309978
rect 337454 309922 337522 309978
rect 337578 309922 337648 309978
rect 337328 309888 337648 309922
rect 368048 310350 368368 310384
rect 368048 310294 368118 310350
rect 368174 310294 368242 310350
rect 368298 310294 368368 310350
rect 368048 310226 368368 310294
rect 368048 310170 368118 310226
rect 368174 310170 368242 310226
rect 368298 310170 368368 310226
rect 368048 310102 368368 310170
rect 368048 310046 368118 310102
rect 368174 310046 368242 310102
rect 368298 310046 368368 310102
rect 368048 309978 368368 310046
rect 368048 309922 368118 309978
rect 368174 309922 368242 309978
rect 368298 309922 368368 309978
rect 368048 309888 368368 309922
rect 229808 298350 230128 298384
rect 229808 298294 229878 298350
rect 229934 298294 230002 298350
rect 230058 298294 230128 298350
rect 229808 298226 230128 298294
rect 229808 298170 229878 298226
rect 229934 298170 230002 298226
rect 230058 298170 230128 298226
rect 229808 298102 230128 298170
rect 229808 298046 229878 298102
rect 229934 298046 230002 298102
rect 230058 298046 230128 298102
rect 229808 297978 230128 298046
rect 229808 297922 229878 297978
rect 229934 297922 230002 297978
rect 230058 297922 230128 297978
rect 229808 297888 230128 297922
rect 260528 298350 260848 298384
rect 260528 298294 260598 298350
rect 260654 298294 260722 298350
rect 260778 298294 260848 298350
rect 260528 298226 260848 298294
rect 260528 298170 260598 298226
rect 260654 298170 260722 298226
rect 260778 298170 260848 298226
rect 260528 298102 260848 298170
rect 260528 298046 260598 298102
rect 260654 298046 260722 298102
rect 260778 298046 260848 298102
rect 260528 297978 260848 298046
rect 260528 297922 260598 297978
rect 260654 297922 260722 297978
rect 260778 297922 260848 297978
rect 260528 297888 260848 297922
rect 291248 298350 291568 298384
rect 291248 298294 291318 298350
rect 291374 298294 291442 298350
rect 291498 298294 291568 298350
rect 291248 298226 291568 298294
rect 291248 298170 291318 298226
rect 291374 298170 291442 298226
rect 291498 298170 291568 298226
rect 291248 298102 291568 298170
rect 291248 298046 291318 298102
rect 291374 298046 291442 298102
rect 291498 298046 291568 298102
rect 291248 297978 291568 298046
rect 291248 297922 291318 297978
rect 291374 297922 291442 297978
rect 291498 297922 291568 297978
rect 291248 297888 291568 297922
rect 321968 298350 322288 298384
rect 321968 298294 322038 298350
rect 322094 298294 322162 298350
rect 322218 298294 322288 298350
rect 321968 298226 322288 298294
rect 321968 298170 322038 298226
rect 322094 298170 322162 298226
rect 322218 298170 322288 298226
rect 321968 298102 322288 298170
rect 321968 298046 322038 298102
rect 322094 298046 322162 298102
rect 322218 298046 322288 298102
rect 321968 297978 322288 298046
rect 321968 297922 322038 297978
rect 322094 297922 322162 297978
rect 322218 297922 322288 297978
rect 321968 297888 322288 297922
rect 352688 298350 353008 298384
rect 352688 298294 352758 298350
rect 352814 298294 352882 298350
rect 352938 298294 353008 298350
rect 352688 298226 353008 298294
rect 352688 298170 352758 298226
rect 352814 298170 352882 298226
rect 352938 298170 353008 298226
rect 352688 298102 353008 298170
rect 352688 298046 352758 298102
rect 352814 298046 352882 298102
rect 352938 298046 353008 298102
rect 352688 297978 353008 298046
rect 352688 297922 352758 297978
rect 352814 297922 352882 297978
rect 352938 297922 353008 297978
rect 352688 297888 353008 297922
rect 214448 292350 214768 292384
rect 214448 292294 214518 292350
rect 214574 292294 214642 292350
rect 214698 292294 214768 292350
rect 214448 292226 214768 292294
rect 214448 292170 214518 292226
rect 214574 292170 214642 292226
rect 214698 292170 214768 292226
rect 214448 292102 214768 292170
rect 214448 292046 214518 292102
rect 214574 292046 214642 292102
rect 214698 292046 214768 292102
rect 214448 291978 214768 292046
rect 214448 291922 214518 291978
rect 214574 291922 214642 291978
rect 214698 291922 214768 291978
rect 214448 291888 214768 291922
rect 245168 292350 245488 292384
rect 245168 292294 245238 292350
rect 245294 292294 245362 292350
rect 245418 292294 245488 292350
rect 245168 292226 245488 292294
rect 245168 292170 245238 292226
rect 245294 292170 245362 292226
rect 245418 292170 245488 292226
rect 245168 292102 245488 292170
rect 245168 292046 245238 292102
rect 245294 292046 245362 292102
rect 245418 292046 245488 292102
rect 245168 291978 245488 292046
rect 245168 291922 245238 291978
rect 245294 291922 245362 291978
rect 245418 291922 245488 291978
rect 245168 291888 245488 291922
rect 275888 292350 276208 292384
rect 275888 292294 275958 292350
rect 276014 292294 276082 292350
rect 276138 292294 276208 292350
rect 275888 292226 276208 292294
rect 275888 292170 275958 292226
rect 276014 292170 276082 292226
rect 276138 292170 276208 292226
rect 275888 292102 276208 292170
rect 275888 292046 275958 292102
rect 276014 292046 276082 292102
rect 276138 292046 276208 292102
rect 275888 291978 276208 292046
rect 275888 291922 275958 291978
rect 276014 291922 276082 291978
rect 276138 291922 276208 291978
rect 275888 291888 276208 291922
rect 306608 292350 306928 292384
rect 306608 292294 306678 292350
rect 306734 292294 306802 292350
rect 306858 292294 306928 292350
rect 306608 292226 306928 292294
rect 306608 292170 306678 292226
rect 306734 292170 306802 292226
rect 306858 292170 306928 292226
rect 306608 292102 306928 292170
rect 306608 292046 306678 292102
rect 306734 292046 306802 292102
rect 306858 292046 306928 292102
rect 306608 291978 306928 292046
rect 306608 291922 306678 291978
rect 306734 291922 306802 291978
rect 306858 291922 306928 291978
rect 306608 291888 306928 291922
rect 337328 292350 337648 292384
rect 337328 292294 337398 292350
rect 337454 292294 337522 292350
rect 337578 292294 337648 292350
rect 337328 292226 337648 292294
rect 337328 292170 337398 292226
rect 337454 292170 337522 292226
rect 337578 292170 337648 292226
rect 337328 292102 337648 292170
rect 337328 292046 337398 292102
rect 337454 292046 337522 292102
rect 337578 292046 337648 292102
rect 337328 291978 337648 292046
rect 337328 291922 337398 291978
rect 337454 291922 337522 291978
rect 337578 291922 337648 291978
rect 337328 291888 337648 291922
rect 368048 292350 368368 292384
rect 368048 292294 368118 292350
rect 368174 292294 368242 292350
rect 368298 292294 368368 292350
rect 368048 292226 368368 292294
rect 368048 292170 368118 292226
rect 368174 292170 368242 292226
rect 368298 292170 368368 292226
rect 368048 292102 368368 292170
rect 368048 292046 368118 292102
rect 368174 292046 368242 292102
rect 368298 292046 368368 292102
rect 368048 291978 368368 292046
rect 368048 291922 368118 291978
rect 368174 291922 368242 291978
rect 368298 291922 368368 291978
rect 368048 291888 368368 291922
rect 229808 280350 230128 280384
rect 229808 280294 229878 280350
rect 229934 280294 230002 280350
rect 230058 280294 230128 280350
rect 229808 280226 230128 280294
rect 229808 280170 229878 280226
rect 229934 280170 230002 280226
rect 230058 280170 230128 280226
rect 229808 280102 230128 280170
rect 229808 280046 229878 280102
rect 229934 280046 230002 280102
rect 230058 280046 230128 280102
rect 229808 279978 230128 280046
rect 229808 279922 229878 279978
rect 229934 279922 230002 279978
rect 230058 279922 230128 279978
rect 229808 279888 230128 279922
rect 260528 280350 260848 280384
rect 260528 280294 260598 280350
rect 260654 280294 260722 280350
rect 260778 280294 260848 280350
rect 260528 280226 260848 280294
rect 260528 280170 260598 280226
rect 260654 280170 260722 280226
rect 260778 280170 260848 280226
rect 260528 280102 260848 280170
rect 260528 280046 260598 280102
rect 260654 280046 260722 280102
rect 260778 280046 260848 280102
rect 260528 279978 260848 280046
rect 260528 279922 260598 279978
rect 260654 279922 260722 279978
rect 260778 279922 260848 279978
rect 260528 279888 260848 279922
rect 291248 280350 291568 280384
rect 291248 280294 291318 280350
rect 291374 280294 291442 280350
rect 291498 280294 291568 280350
rect 291248 280226 291568 280294
rect 291248 280170 291318 280226
rect 291374 280170 291442 280226
rect 291498 280170 291568 280226
rect 291248 280102 291568 280170
rect 291248 280046 291318 280102
rect 291374 280046 291442 280102
rect 291498 280046 291568 280102
rect 291248 279978 291568 280046
rect 291248 279922 291318 279978
rect 291374 279922 291442 279978
rect 291498 279922 291568 279978
rect 291248 279888 291568 279922
rect 321968 280350 322288 280384
rect 321968 280294 322038 280350
rect 322094 280294 322162 280350
rect 322218 280294 322288 280350
rect 321968 280226 322288 280294
rect 321968 280170 322038 280226
rect 322094 280170 322162 280226
rect 322218 280170 322288 280226
rect 321968 280102 322288 280170
rect 321968 280046 322038 280102
rect 322094 280046 322162 280102
rect 322218 280046 322288 280102
rect 321968 279978 322288 280046
rect 321968 279922 322038 279978
rect 322094 279922 322162 279978
rect 322218 279922 322288 279978
rect 321968 279888 322288 279922
rect 352688 280350 353008 280384
rect 352688 280294 352758 280350
rect 352814 280294 352882 280350
rect 352938 280294 353008 280350
rect 352688 280226 353008 280294
rect 352688 280170 352758 280226
rect 352814 280170 352882 280226
rect 352938 280170 353008 280226
rect 352688 280102 353008 280170
rect 352688 280046 352758 280102
rect 352814 280046 352882 280102
rect 352938 280046 353008 280102
rect 352688 279978 353008 280046
rect 352688 279922 352758 279978
rect 352814 279922 352882 279978
rect 352938 279922 353008 279978
rect 352688 279888 353008 279922
rect 213500 276352 213556 276362
rect 214448 274350 214768 274384
rect 214448 274294 214518 274350
rect 214574 274294 214642 274350
rect 214698 274294 214768 274350
rect 214448 274226 214768 274294
rect 214448 274170 214518 274226
rect 214574 274170 214642 274226
rect 214698 274170 214768 274226
rect 214448 274102 214768 274170
rect 214448 274046 214518 274102
rect 214574 274046 214642 274102
rect 214698 274046 214768 274102
rect 214448 273978 214768 274046
rect 214448 273922 214518 273978
rect 214574 273922 214642 273978
rect 214698 273922 214768 273978
rect 214448 273888 214768 273922
rect 245168 274350 245488 274384
rect 245168 274294 245238 274350
rect 245294 274294 245362 274350
rect 245418 274294 245488 274350
rect 245168 274226 245488 274294
rect 245168 274170 245238 274226
rect 245294 274170 245362 274226
rect 245418 274170 245488 274226
rect 245168 274102 245488 274170
rect 245168 274046 245238 274102
rect 245294 274046 245362 274102
rect 245418 274046 245488 274102
rect 245168 273978 245488 274046
rect 245168 273922 245238 273978
rect 245294 273922 245362 273978
rect 245418 273922 245488 273978
rect 245168 273888 245488 273922
rect 275888 274350 276208 274384
rect 275888 274294 275958 274350
rect 276014 274294 276082 274350
rect 276138 274294 276208 274350
rect 275888 274226 276208 274294
rect 275888 274170 275958 274226
rect 276014 274170 276082 274226
rect 276138 274170 276208 274226
rect 275888 274102 276208 274170
rect 275888 274046 275958 274102
rect 276014 274046 276082 274102
rect 276138 274046 276208 274102
rect 275888 273978 276208 274046
rect 275888 273922 275958 273978
rect 276014 273922 276082 273978
rect 276138 273922 276208 273978
rect 275888 273888 276208 273922
rect 306608 274350 306928 274384
rect 306608 274294 306678 274350
rect 306734 274294 306802 274350
rect 306858 274294 306928 274350
rect 306608 274226 306928 274294
rect 306608 274170 306678 274226
rect 306734 274170 306802 274226
rect 306858 274170 306928 274226
rect 306608 274102 306928 274170
rect 306608 274046 306678 274102
rect 306734 274046 306802 274102
rect 306858 274046 306928 274102
rect 306608 273978 306928 274046
rect 306608 273922 306678 273978
rect 306734 273922 306802 273978
rect 306858 273922 306928 273978
rect 306608 273888 306928 273922
rect 337328 274350 337648 274384
rect 337328 274294 337398 274350
rect 337454 274294 337522 274350
rect 337578 274294 337648 274350
rect 337328 274226 337648 274294
rect 337328 274170 337398 274226
rect 337454 274170 337522 274226
rect 337578 274170 337648 274226
rect 337328 274102 337648 274170
rect 337328 274046 337398 274102
rect 337454 274046 337522 274102
rect 337578 274046 337648 274102
rect 337328 273978 337648 274046
rect 337328 273922 337398 273978
rect 337454 273922 337522 273978
rect 337578 273922 337648 273978
rect 337328 273888 337648 273922
rect 368048 274350 368368 274384
rect 368048 274294 368118 274350
rect 368174 274294 368242 274350
rect 368298 274294 368368 274350
rect 368048 274226 368368 274294
rect 368048 274170 368118 274226
rect 368174 274170 368242 274226
rect 368298 274170 368368 274226
rect 368048 274102 368368 274170
rect 368048 274046 368118 274102
rect 368174 274046 368242 274102
rect 368298 274046 368368 274102
rect 368048 273978 368368 274046
rect 368048 273922 368118 273978
rect 368174 273922 368242 273978
rect 368298 273922 368368 273978
rect 368048 273888 368368 273922
rect 229808 262350 230128 262384
rect 229808 262294 229878 262350
rect 229934 262294 230002 262350
rect 230058 262294 230128 262350
rect 229808 262226 230128 262294
rect 229808 262170 229878 262226
rect 229934 262170 230002 262226
rect 230058 262170 230128 262226
rect 229808 262102 230128 262170
rect 229808 262046 229878 262102
rect 229934 262046 230002 262102
rect 230058 262046 230128 262102
rect 229808 261978 230128 262046
rect 229808 261922 229878 261978
rect 229934 261922 230002 261978
rect 230058 261922 230128 261978
rect 229808 261888 230128 261922
rect 260528 262350 260848 262384
rect 260528 262294 260598 262350
rect 260654 262294 260722 262350
rect 260778 262294 260848 262350
rect 260528 262226 260848 262294
rect 260528 262170 260598 262226
rect 260654 262170 260722 262226
rect 260778 262170 260848 262226
rect 260528 262102 260848 262170
rect 260528 262046 260598 262102
rect 260654 262046 260722 262102
rect 260778 262046 260848 262102
rect 260528 261978 260848 262046
rect 260528 261922 260598 261978
rect 260654 261922 260722 261978
rect 260778 261922 260848 261978
rect 260528 261888 260848 261922
rect 291248 262350 291568 262384
rect 291248 262294 291318 262350
rect 291374 262294 291442 262350
rect 291498 262294 291568 262350
rect 291248 262226 291568 262294
rect 291248 262170 291318 262226
rect 291374 262170 291442 262226
rect 291498 262170 291568 262226
rect 291248 262102 291568 262170
rect 291248 262046 291318 262102
rect 291374 262046 291442 262102
rect 291498 262046 291568 262102
rect 291248 261978 291568 262046
rect 291248 261922 291318 261978
rect 291374 261922 291442 261978
rect 291498 261922 291568 261978
rect 291248 261888 291568 261922
rect 321968 262350 322288 262384
rect 321968 262294 322038 262350
rect 322094 262294 322162 262350
rect 322218 262294 322288 262350
rect 321968 262226 322288 262294
rect 321968 262170 322038 262226
rect 322094 262170 322162 262226
rect 322218 262170 322288 262226
rect 321968 262102 322288 262170
rect 321968 262046 322038 262102
rect 322094 262046 322162 262102
rect 322218 262046 322288 262102
rect 321968 261978 322288 262046
rect 321968 261922 322038 261978
rect 322094 261922 322162 261978
rect 322218 261922 322288 261978
rect 321968 261888 322288 261922
rect 352688 262350 353008 262384
rect 352688 262294 352758 262350
rect 352814 262294 352882 262350
rect 352938 262294 353008 262350
rect 352688 262226 353008 262294
rect 352688 262170 352758 262226
rect 352814 262170 352882 262226
rect 352938 262170 353008 262226
rect 352688 262102 353008 262170
rect 352688 262046 352758 262102
rect 352814 262046 352882 262102
rect 352938 262046 353008 262102
rect 352688 261978 353008 262046
rect 352688 261922 352758 261978
rect 352814 261922 352882 261978
rect 352938 261922 353008 261978
rect 352688 261888 353008 261922
rect 211820 257812 211876 257822
rect 214448 256350 214768 256384
rect 214448 256294 214518 256350
rect 214574 256294 214642 256350
rect 214698 256294 214768 256350
rect 214448 256226 214768 256294
rect 214448 256170 214518 256226
rect 214574 256170 214642 256226
rect 214698 256170 214768 256226
rect 214448 256102 214768 256170
rect 214448 256046 214518 256102
rect 214574 256046 214642 256102
rect 214698 256046 214768 256102
rect 214448 255978 214768 256046
rect 214448 255922 214518 255978
rect 214574 255922 214642 255978
rect 214698 255922 214768 255978
rect 214448 255888 214768 255922
rect 245168 256350 245488 256384
rect 245168 256294 245238 256350
rect 245294 256294 245362 256350
rect 245418 256294 245488 256350
rect 245168 256226 245488 256294
rect 245168 256170 245238 256226
rect 245294 256170 245362 256226
rect 245418 256170 245488 256226
rect 245168 256102 245488 256170
rect 245168 256046 245238 256102
rect 245294 256046 245362 256102
rect 245418 256046 245488 256102
rect 245168 255978 245488 256046
rect 245168 255922 245238 255978
rect 245294 255922 245362 255978
rect 245418 255922 245488 255978
rect 245168 255888 245488 255922
rect 275888 256350 276208 256384
rect 275888 256294 275958 256350
rect 276014 256294 276082 256350
rect 276138 256294 276208 256350
rect 275888 256226 276208 256294
rect 275888 256170 275958 256226
rect 276014 256170 276082 256226
rect 276138 256170 276208 256226
rect 275888 256102 276208 256170
rect 275888 256046 275958 256102
rect 276014 256046 276082 256102
rect 276138 256046 276208 256102
rect 275888 255978 276208 256046
rect 275888 255922 275958 255978
rect 276014 255922 276082 255978
rect 276138 255922 276208 255978
rect 275888 255888 276208 255922
rect 306608 256350 306928 256384
rect 306608 256294 306678 256350
rect 306734 256294 306802 256350
rect 306858 256294 306928 256350
rect 306608 256226 306928 256294
rect 306608 256170 306678 256226
rect 306734 256170 306802 256226
rect 306858 256170 306928 256226
rect 306608 256102 306928 256170
rect 306608 256046 306678 256102
rect 306734 256046 306802 256102
rect 306858 256046 306928 256102
rect 306608 255978 306928 256046
rect 306608 255922 306678 255978
rect 306734 255922 306802 255978
rect 306858 255922 306928 255978
rect 306608 255888 306928 255922
rect 337328 256350 337648 256384
rect 337328 256294 337398 256350
rect 337454 256294 337522 256350
rect 337578 256294 337648 256350
rect 337328 256226 337648 256294
rect 337328 256170 337398 256226
rect 337454 256170 337522 256226
rect 337578 256170 337648 256226
rect 337328 256102 337648 256170
rect 337328 256046 337398 256102
rect 337454 256046 337522 256102
rect 337578 256046 337648 256102
rect 337328 255978 337648 256046
rect 337328 255922 337398 255978
rect 337454 255922 337522 255978
rect 337578 255922 337648 255978
rect 337328 255888 337648 255922
rect 368048 256350 368368 256384
rect 368048 256294 368118 256350
rect 368174 256294 368242 256350
rect 368298 256294 368368 256350
rect 368048 256226 368368 256294
rect 368048 256170 368118 256226
rect 368174 256170 368242 256226
rect 368298 256170 368368 256226
rect 368048 256102 368368 256170
rect 368048 256046 368118 256102
rect 368174 256046 368242 256102
rect 368298 256046 368368 256102
rect 368048 255978 368368 256046
rect 368048 255922 368118 255978
rect 368174 255922 368242 255978
rect 368298 255922 368368 255978
rect 368048 255888 368368 255922
rect 229808 244350 230128 244384
rect 229808 244294 229878 244350
rect 229934 244294 230002 244350
rect 230058 244294 230128 244350
rect 229808 244226 230128 244294
rect 229808 244170 229878 244226
rect 229934 244170 230002 244226
rect 230058 244170 230128 244226
rect 229808 244102 230128 244170
rect 229808 244046 229878 244102
rect 229934 244046 230002 244102
rect 230058 244046 230128 244102
rect 229808 243978 230128 244046
rect 229808 243922 229878 243978
rect 229934 243922 230002 243978
rect 230058 243922 230128 243978
rect 229808 243888 230128 243922
rect 260528 244350 260848 244384
rect 260528 244294 260598 244350
rect 260654 244294 260722 244350
rect 260778 244294 260848 244350
rect 260528 244226 260848 244294
rect 260528 244170 260598 244226
rect 260654 244170 260722 244226
rect 260778 244170 260848 244226
rect 260528 244102 260848 244170
rect 260528 244046 260598 244102
rect 260654 244046 260722 244102
rect 260778 244046 260848 244102
rect 260528 243978 260848 244046
rect 260528 243922 260598 243978
rect 260654 243922 260722 243978
rect 260778 243922 260848 243978
rect 260528 243888 260848 243922
rect 291248 244350 291568 244384
rect 291248 244294 291318 244350
rect 291374 244294 291442 244350
rect 291498 244294 291568 244350
rect 291248 244226 291568 244294
rect 291248 244170 291318 244226
rect 291374 244170 291442 244226
rect 291498 244170 291568 244226
rect 291248 244102 291568 244170
rect 291248 244046 291318 244102
rect 291374 244046 291442 244102
rect 291498 244046 291568 244102
rect 291248 243978 291568 244046
rect 291248 243922 291318 243978
rect 291374 243922 291442 243978
rect 291498 243922 291568 243978
rect 291248 243888 291568 243922
rect 321968 244350 322288 244384
rect 321968 244294 322038 244350
rect 322094 244294 322162 244350
rect 322218 244294 322288 244350
rect 321968 244226 322288 244294
rect 321968 244170 322038 244226
rect 322094 244170 322162 244226
rect 322218 244170 322288 244226
rect 321968 244102 322288 244170
rect 321968 244046 322038 244102
rect 322094 244046 322162 244102
rect 322218 244046 322288 244102
rect 321968 243978 322288 244046
rect 321968 243922 322038 243978
rect 322094 243922 322162 243978
rect 322218 243922 322288 243978
rect 321968 243888 322288 243922
rect 352688 244350 353008 244384
rect 352688 244294 352758 244350
rect 352814 244294 352882 244350
rect 352938 244294 353008 244350
rect 352688 244226 353008 244294
rect 352688 244170 352758 244226
rect 352814 244170 352882 244226
rect 352938 244170 353008 244226
rect 352688 244102 353008 244170
rect 352688 244046 352758 244102
rect 352814 244046 352882 244102
rect 352938 244046 353008 244102
rect 352688 243978 353008 244046
rect 352688 243922 352758 243978
rect 352814 243922 352882 243978
rect 352938 243922 353008 243978
rect 352688 243888 353008 243922
rect 370076 239764 370132 239774
rect 214448 238350 214768 238384
rect 214448 238294 214518 238350
rect 214574 238294 214642 238350
rect 214698 238294 214768 238350
rect 214448 238226 214768 238294
rect 214448 238170 214518 238226
rect 214574 238170 214642 238226
rect 214698 238170 214768 238226
rect 214448 238102 214768 238170
rect 214448 238046 214518 238102
rect 214574 238046 214642 238102
rect 214698 238046 214768 238102
rect 214448 237978 214768 238046
rect 214448 237922 214518 237978
rect 214574 237922 214642 237978
rect 214698 237922 214768 237978
rect 214448 237888 214768 237922
rect 245168 238350 245488 238384
rect 245168 238294 245238 238350
rect 245294 238294 245362 238350
rect 245418 238294 245488 238350
rect 245168 238226 245488 238294
rect 245168 238170 245238 238226
rect 245294 238170 245362 238226
rect 245418 238170 245488 238226
rect 245168 238102 245488 238170
rect 245168 238046 245238 238102
rect 245294 238046 245362 238102
rect 245418 238046 245488 238102
rect 245168 237978 245488 238046
rect 245168 237922 245238 237978
rect 245294 237922 245362 237978
rect 245418 237922 245488 237978
rect 245168 237888 245488 237922
rect 275888 238350 276208 238384
rect 275888 238294 275958 238350
rect 276014 238294 276082 238350
rect 276138 238294 276208 238350
rect 275888 238226 276208 238294
rect 275888 238170 275958 238226
rect 276014 238170 276082 238226
rect 276138 238170 276208 238226
rect 275888 238102 276208 238170
rect 275888 238046 275958 238102
rect 276014 238046 276082 238102
rect 276138 238046 276208 238102
rect 275888 237978 276208 238046
rect 275888 237922 275958 237978
rect 276014 237922 276082 237978
rect 276138 237922 276208 237978
rect 275888 237888 276208 237922
rect 306608 238350 306928 238384
rect 306608 238294 306678 238350
rect 306734 238294 306802 238350
rect 306858 238294 306928 238350
rect 306608 238226 306928 238294
rect 306608 238170 306678 238226
rect 306734 238170 306802 238226
rect 306858 238170 306928 238226
rect 306608 238102 306928 238170
rect 306608 238046 306678 238102
rect 306734 238046 306802 238102
rect 306858 238046 306928 238102
rect 306608 237978 306928 238046
rect 306608 237922 306678 237978
rect 306734 237922 306802 237978
rect 306858 237922 306928 237978
rect 306608 237888 306928 237922
rect 337328 238350 337648 238384
rect 337328 238294 337398 238350
rect 337454 238294 337522 238350
rect 337578 238294 337648 238350
rect 337328 238226 337648 238294
rect 337328 238170 337398 238226
rect 337454 238170 337522 238226
rect 337578 238170 337648 238226
rect 337328 238102 337648 238170
rect 337328 238046 337398 238102
rect 337454 238046 337522 238102
rect 337578 238046 337648 238102
rect 337328 237978 337648 238046
rect 337328 237922 337398 237978
rect 337454 237922 337522 237978
rect 337578 237922 337648 237978
rect 337328 237888 337648 237922
rect 368048 238350 368368 238384
rect 368048 238294 368118 238350
rect 368174 238294 368242 238350
rect 368298 238294 368368 238350
rect 368048 238226 368368 238294
rect 368048 238170 368118 238226
rect 368174 238170 368242 238226
rect 368298 238170 368368 238226
rect 368048 238102 368368 238170
rect 368048 238046 368118 238102
rect 368174 238046 368242 238102
rect 368298 238046 368368 238102
rect 368048 237978 368368 238046
rect 368048 237922 368118 237978
rect 368174 237922 368242 237978
rect 368298 237922 368368 237978
rect 368048 237888 368368 237922
rect 211708 236032 211764 236042
rect 210700 235890 210756 235900
rect 229808 226350 230128 226384
rect 229808 226294 229878 226350
rect 229934 226294 230002 226350
rect 230058 226294 230128 226350
rect 229808 226226 230128 226294
rect 229808 226170 229878 226226
rect 229934 226170 230002 226226
rect 230058 226170 230128 226226
rect 229808 226102 230128 226170
rect 229808 226046 229878 226102
rect 229934 226046 230002 226102
rect 230058 226046 230128 226102
rect 229808 225978 230128 226046
rect 229808 225922 229878 225978
rect 229934 225922 230002 225978
rect 230058 225922 230128 225978
rect 229808 225888 230128 225922
rect 260528 226350 260848 226384
rect 260528 226294 260598 226350
rect 260654 226294 260722 226350
rect 260778 226294 260848 226350
rect 260528 226226 260848 226294
rect 260528 226170 260598 226226
rect 260654 226170 260722 226226
rect 260778 226170 260848 226226
rect 260528 226102 260848 226170
rect 260528 226046 260598 226102
rect 260654 226046 260722 226102
rect 260778 226046 260848 226102
rect 260528 225978 260848 226046
rect 260528 225922 260598 225978
rect 260654 225922 260722 225978
rect 260778 225922 260848 225978
rect 260528 225888 260848 225922
rect 291248 226350 291568 226384
rect 291248 226294 291318 226350
rect 291374 226294 291442 226350
rect 291498 226294 291568 226350
rect 291248 226226 291568 226294
rect 291248 226170 291318 226226
rect 291374 226170 291442 226226
rect 291498 226170 291568 226226
rect 291248 226102 291568 226170
rect 291248 226046 291318 226102
rect 291374 226046 291442 226102
rect 291498 226046 291568 226102
rect 291248 225978 291568 226046
rect 291248 225922 291318 225978
rect 291374 225922 291442 225978
rect 291498 225922 291568 225978
rect 291248 225888 291568 225922
rect 321968 226350 322288 226384
rect 321968 226294 322038 226350
rect 322094 226294 322162 226350
rect 322218 226294 322288 226350
rect 321968 226226 322288 226294
rect 321968 226170 322038 226226
rect 322094 226170 322162 226226
rect 322218 226170 322288 226226
rect 321968 226102 322288 226170
rect 321968 226046 322038 226102
rect 322094 226046 322162 226102
rect 322218 226046 322288 226102
rect 321968 225978 322288 226046
rect 321968 225922 322038 225978
rect 322094 225922 322162 225978
rect 322218 225922 322288 225978
rect 321968 225888 322288 225922
rect 352688 226350 353008 226384
rect 352688 226294 352758 226350
rect 352814 226294 352882 226350
rect 352938 226294 353008 226350
rect 352688 226226 353008 226294
rect 352688 226170 352758 226226
rect 352814 226170 352882 226226
rect 352938 226170 353008 226226
rect 352688 226102 353008 226170
rect 352688 226046 352758 226102
rect 352814 226046 352882 226102
rect 352938 226046 353008 226102
rect 352688 225978 353008 226046
rect 352688 225922 352758 225978
rect 352814 225922 352882 225978
rect 352938 225922 353008 225978
rect 352688 225888 353008 225922
rect 369404 221844 369460 221854
rect 214448 220350 214768 220384
rect 214448 220294 214518 220350
rect 214574 220294 214642 220350
rect 214698 220294 214768 220350
rect 214448 220226 214768 220294
rect 214448 220170 214518 220226
rect 214574 220170 214642 220226
rect 214698 220170 214768 220226
rect 214448 220102 214768 220170
rect 214448 220046 214518 220102
rect 214574 220046 214642 220102
rect 214698 220046 214768 220102
rect 214448 219978 214768 220046
rect 214448 219922 214518 219978
rect 214574 219922 214642 219978
rect 214698 219922 214768 219978
rect 214448 219888 214768 219922
rect 245168 220350 245488 220384
rect 245168 220294 245238 220350
rect 245294 220294 245362 220350
rect 245418 220294 245488 220350
rect 245168 220226 245488 220294
rect 245168 220170 245238 220226
rect 245294 220170 245362 220226
rect 245418 220170 245488 220226
rect 245168 220102 245488 220170
rect 245168 220046 245238 220102
rect 245294 220046 245362 220102
rect 245418 220046 245488 220102
rect 245168 219978 245488 220046
rect 245168 219922 245238 219978
rect 245294 219922 245362 219978
rect 245418 219922 245488 219978
rect 245168 219888 245488 219922
rect 275888 220350 276208 220384
rect 275888 220294 275958 220350
rect 276014 220294 276082 220350
rect 276138 220294 276208 220350
rect 275888 220226 276208 220294
rect 275888 220170 275958 220226
rect 276014 220170 276082 220226
rect 276138 220170 276208 220226
rect 275888 220102 276208 220170
rect 275888 220046 275958 220102
rect 276014 220046 276082 220102
rect 276138 220046 276208 220102
rect 275888 219978 276208 220046
rect 275888 219922 275958 219978
rect 276014 219922 276082 219978
rect 276138 219922 276208 219978
rect 275888 219888 276208 219922
rect 306608 220350 306928 220384
rect 306608 220294 306678 220350
rect 306734 220294 306802 220350
rect 306858 220294 306928 220350
rect 306608 220226 306928 220294
rect 306608 220170 306678 220226
rect 306734 220170 306802 220226
rect 306858 220170 306928 220226
rect 306608 220102 306928 220170
rect 306608 220046 306678 220102
rect 306734 220046 306802 220102
rect 306858 220046 306928 220102
rect 306608 219978 306928 220046
rect 306608 219922 306678 219978
rect 306734 219922 306802 219978
rect 306858 219922 306928 219978
rect 306608 219888 306928 219922
rect 337328 220350 337648 220384
rect 337328 220294 337398 220350
rect 337454 220294 337522 220350
rect 337578 220294 337648 220350
rect 337328 220226 337648 220294
rect 337328 220170 337398 220226
rect 337454 220170 337522 220226
rect 337578 220170 337648 220226
rect 337328 220102 337648 220170
rect 337328 220046 337398 220102
rect 337454 220046 337522 220102
rect 337578 220046 337648 220102
rect 337328 219978 337648 220046
rect 337328 219922 337398 219978
rect 337454 219922 337522 219978
rect 337578 219922 337648 219978
rect 337328 219888 337648 219922
rect 368048 220350 368368 220384
rect 368048 220294 368118 220350
rect 368174 220294 368242 220350
rect 368298 220294 368368 220350
rect 368048 220226 368368 220294
rect 368048 220170 368118 220226
rect 368174 220170 368242 220226
rect 368298 220170 368368 220226
rect 368048 220102 368368 220170
rect 368048 220046 368118 220102
rect 368174 220046 368242 220102
rect 368298 220046 368368 220102
rect 368048 219978 368368 220046
rect 368048 219922 368118 219978
rect 368174 219922 368242 219978
rect 368298 219922 368368 219978
rect 368048 219888 368368 219922
rect 369404 216658 369460 221788
rect 369404 216592 369460 216602
rect 369516 220724 369572 220734
rect 229808 208350 230128 208384
rect 229808 208294 229878 208350
rect 229934 208294 230002 208350
rect 230058 208294 230128 208350
rect 229808 208226 230128 208294
rect 229808 208170 229878 208226
rect 229934 208170 230002 208226
rect 230058 208170 230128 208226
rect 229808 208102 230128 208170
rect 229808 208046 229878 208102
rect 229934 208046 230002 208102
rect 230058 208046 230128 208102
rect 229808 207978 230128 208046
rect 229808 207922 229878 207978
rect 229934 207922 230002 207978
rect 230058 207922 230128 207978
rect 229808 207888 230128 207922
rect 260528 208350 260848 208384
rect 260528 208294 260598 208350
rect 260654 208294 260722 208350
rect 260778 208294 260848 208350
rect 260528 208226 260848 208294
rect 260528 208170 260598 208226
rect 260654 208170 260722 208226
rect 260778 208170 260848 208226
rect 260528 208102 260848 208170
rect 260528 208046 260598 208102
rect 260654 208046 260722 208102
rect 260778 208046 260848 208102
rect 260528 207978 260848 208046
rect 260528 207922 260598 207978
rect 260654 207922 260722 207978
rect 260778 207922 260848 207978
rect 260528 207888 260848 207922
rect 291248 208350 291568 208384
rect 291248 208294 291318 208350
rect 291374 208294 291442 208350
rect 291498 208294 291568 208350
rect 291248 208226 291568 208294
rect 291248 208170 291318 208226
rect 291374 208170 291442 208226
rect 291498 208170 291568 208226
rect 291248 208102 291568 208170
rect 291248 208046 291318 208102
rect 291374 208046 291442 208102
rect 291498 208046 291568 208102
rect 291248 207978 291568 208046
rect 291248 207922 291318 207978
rect 291374 207922 291442 207978
rect 291498 207922 291568 207978
rect 291248 207888 291568 207922
rect 321968 208350 322288 208384
rect 321968 208294 322038 208350
rect 322094 208294 322162 208350
rect 322218 208294 322288 208350
rect 321968 208226 322288 208294
rect 321968 208170 322038 208226
rect 322094 208170 322162 208226
rect 322218 208170 322288 208226
rect 321968 208102 322288 208170
rect 321968 208046 322038 208102
rect 322094 208046 322162 208102
rect 322218 208046 322288 208102
rect 321968 207978 322288 208046
rect 321968 207922 322038 207978
rect 322094 207922 322162 207978
rect 322218 207922 322288 207978
rect 321968 207888 322288 207922
rect 352688 208350 353008 208384
rect 352688 208294 352758 208350
rect 352814 208294 352882 208350
rect 352938 208294 353008 208350
rect 352688 208226 353008 208294
rect 352688 208170 352758 208226
rect 352814 208170 352882 208226
rect 352938 208170 353008 208226
rect 352688 208102 353008 208170
rect 352688 208046 352758 208102
rect 352814 208046 352882 208102
rect 352938 208046 353008 208102
rect 352688 207978 353008 208046
rect 352688 207922 352758 207978
rect 352814 207922 352882 207978
rect 352938 207922 353008 207978
rect 352688 207888 353008 207922
rect 214448 202350 214768 202384
rect 214448 202294 214518 202350
rect 214574 202294 214642 202350
rect 214698 202294 214768 202350
rect 214448 202226 214768 202294
rect 214448 202170 214518 202226
rect 214574 202170 214642 202226
rect 214698 202170 214768 202226
rect 214448 202102 214768 202170
rect 214448 202046 214518 202102
rect 214574 202046 214642 202102
rect 214698 202046 214768 202102
rect 214448 201978 214768 202046
rect 214448 201922 214518 201978
rect 214574 201922 214642 201978
rect 214698 201922 214768 201978
rect 214448 201888 214768 201922
rect 245168 202350 245488 202384
rect 245168 202294 245238 202350
rect 245294 202294 245362 202350
rect 245418 202294 245488 202350
rect 245168 202226 245488 202294
rect 245168 202170 245238 202226
rect 245294 202170 245362 202226
rect 245418 202170 245488 202226
rect 245168 202102 245488 202170
rect 245168 202046 245238 202102
rect 245294 202046 245362 202102
rect 245418 202046 245488 202102
rect 245168 201978 245488 202046
rect 245168 201922 245238 201978
rect 245294 201922 245362 201978
rect 245418 201922 245488 201978
rect 245168 201888 245488 201922
rect 275888 202350 276208 202384
rect 275888 202294 275958 202350
rect 276014 202294 276082 202350
rect 276138 202294 276208 202350
rect 275888 202226 276208 202294
rect 275888 202170 275958 202226
rect 276014 202170 276082 202226
rect 276138 202170 276208 202226
rect 275888 202102 276208 202170
rect 275888 202046 275958 202102
rect 276014 202046 276082 202102
rect 276138 202046 276208 202102
rect 275888 201978 276208 202046
rect 275888 201922 275958 201978
rect 276014 201922 276082 201978
rect 276138 201922 276208 201978
rect 275888 201888 276208 201922
rect 306608 202350 306928 202384
rect 306608 202294 306678 202350
rect 306734 202294 306802 202350
rect 306858 202294 306928 202350
rect 306608 202226 306928 202294
rect 306608 202170 306678 202226
rect 306734 202170 306802 202226
rect 306858 202170 306928 202226
rect 306608 202102 306928 202170
rect 306608 202046 306678 202102
rect 306734 202046 306802 202102
rect 306858 202046 306928 202102
rect 306608 201978 306928 202046
rect 306608 201922 306678 201978
rect 306734 201922 306802 201978
rect 306858 201922 306928 201978
rect 306608 201888 306928 201922
rect 337328 202350 337648 202384
rect 337328 202294 337398 202350
rect 337454 202294 337522 202350
rect 337578 202294 337648 202350
rect 337328 202226 337648 202294
rect 337328 202170 337398 202226
rect 337454 202170 337522 202226
rect 337578 202170 337648 202226
rect 337328 202102 337648 202170
rect 337328 202046 337398 202102
rect 337454 202046 337522 202102
rect 337578 202046 337648 202102
rect 337328 201978 337648 202046
rect 337328 201922 337398 201978
rect 337454 201922 337522 201978
rect 337578 201922 337648 201978
rect 337328 201888 337648 201922
rect 368048 202350 368368 202384
rect 368048 202294 368118 202350
rect 368174 202294 368242 202350
rect 368298 202294 368368 202350
rect 368048 202226 368368 202294
rect 368048 202170 368118 202226
rect 368174 202170 368242 202226
rect 368298 202170 368368 202226
rect 368048 202102 368368 202170
rect 368048 202046 368118 202102
rect 368174 202046 368242 202102
rect 368298 202046 368368 202102
rect 368048 201978 368368 202046
rect 368048 201922 368118 201978
rect 368174 201922 368242 201978
rect 368298 201922 368368 201978
rect 368048 201888 368368 201922
rect 369516 193978 369572 220668
rect 369516 193912 369572 193922
rect 229808 190350 230128 190384
rect 229808 190294 229878 190350
rect 229934 190294 230002 190350
rect 230058 190294 230128 190350
rect 229808 190226 230128 190294
rect 229808 190170 229878 190226
rect 229934 190170 230002 190226
rect 230058 190170 230128 190226
rect 229808 190102 230128 190170
rect 229808 190046 229878 190102
rect 229934 190046 230002 190102
rect 230058 190046 230128 190102
rect 229808 189978 230128 190046
rect 229808 189922 229878 189978
rect 229934 189922 230002 189978
rect 230058 189922 230128 189978
rect 229808 189888 230128 189922
rect 260528 190350 260848 190384
rect 260528 190294 260598 190350
rect 260654 190294 260722 190350
rect 260778 190294 260848 190350
rect 260528 190226 260848 190294
rect 260528 190170 260598 190226
rect 260654 190170 260722 190226
rect 260778 190170 260848 190226
rect 260528 190102 260848 190170
rect 260528 190046 260598 190102
rect 260654 190046 260722 190102
rect 260778 190046 260848 190102
rect 260528 189978 260848 190046
rect 260528 189922 260598 189978
rect 260654 189922 260722 189978
rect 260778 189922 260848 189978
rect 260528 189888 260848 189922
rect 291248 190350 291568 190384
rect 291248 190294 291318 190350
rect 291374 190294 291442 190350
rect 291498 190294 291568 190350
rect 291248 190226 291568 190294
rect 291248 190170 291318 190226
rect 291374 190170 291442 190226
rect 291498 190170 291568 190226
rect 291248 190102 291568 190170
rect 291248 190046 291318 190102
rect 291374 190046 291442 190102
rect 291498 190046 291568 190102
rect 291248 189978 291568 190046
rect 291248 189922 291318 189978
rect 291374 189922 291442 189978
rect 291498 189922 291568 189978
rect 291248 189888 291568 189922
rect 321968 190350 322288 190384
rect 321968 190294 322038 190350
rect 322094 190294 322162 190350
rect 322218 190294 322288 190350
rect 321968 190226 322288 190294
rect 321968 190170 322038 190226
rect 322094 190170 322162 190226
rect 322218 190170 322288 190226
rect 321968 190102 322288 190170
rect 321968 190046 322038 190102
rect 322094 190046 322162 190102
rect 322218 190046 322288 190102
rect 321968 189978 322288 190046
rect 321968 189922 322038 189978
rect 322094 189922 322162 189978
rect 322218 189922 322288 189978
rect 321968 189888 322288 189922
rect 352688 190350 353008 190384
rect 352688 190294 352758 190350
rect 352814 190294 352882 190350
rect 352938 190294 353008 190350
rect 352688 190226 353008 190294
rect 352688 190170 352758 190226
rect 352814 190170 352882 190226
rect 352938 190170 353008 190226
rect 352688 190102 353008 190170
rect 352688 190046 352758 190102
rect 352814 190046 352882 190102
rect 352938 190046 353008 190102
rect 352688 189978 353008 190046
rect 352688 189922 352758 189978
rect 352814 189922 352882 189978
rect 352938 189922 353008 189978
rect 352688 189888 353008 189922
rect 370076 184772 370132 239708
rect 370300 230804 370356 230814
rect 370188 226324 370244 226334
rect 370188 192388 370244 226268
rect 370300 200788 370356 230748
rect 370300 200722 370356 200732
rect 370412 227444 370468 227454
rect 370412 199108 370468 227388
rect 370636 224420 370692 327628
rect 373884 324660 373940 324670
rect 373660 322756 373716 322766
rect 373660 314188 373716 322700
rect 373772 322644 373828 322654
rect 373772 314804 373828 322588
rect 373884 318164 373940 324604
rect 373884 318098 373940 318108
rect 373772 314738 373828 314748
rect 373660 314132 373828 314188
rect 373772 312564 373828 314132
rect 373772 312498 373828 312508
rect 373772 310978 373828 310988
rect 373660 306964 373716 306974
rect 373660 299236 373716 306908
rect 373660 299170 373716 299180
rect 373772 295764 373828 310922
rect 374058 310350 374678 327922
rect 377778 598172 378398 598268
rect 377778 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 378398 598172
rect 377778 598048 378398 598116
rect 377778 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 378398 598048
rect 377778 597924 378398 597992
rect 377778 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 378398 597924
rect 377778 597800 378398 597868
rect 377778 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 378398 597800
rect 377778 586350 378398 597744
rect 377778 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 378398 586350
rect 377778 586226 378398 586294
rect 377778 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 378398 586226
rect 377778 586102 378398 586170
rect 377778 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 378398 586102
rect 377778 585978 378398 586046
rect 377778 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 378398 585978
rect 377778 568350 378398 585922
rect 377778 568294 377874 568350
rect 377930 568294 377998 568350
rect 378054 568294 378122 568350
rect 378178 568294 378246 568350
rect 378302 568294 378398 568350
rect 377778 568226 378398 568294
rect 377778 568170 377874 568226
rect 377930 568170 377998 568226
rect 378054 568170 378122 568226
rect 378178 568170 378246 568226
rect 378302 568170 378398 568226
rect 377778 568102 378398 568170
rect 377778 568046 377874 568102
rect 377930 568046 377998 568102
rect 378054 568046 378122 568102
rect 378178 568046 378246 568102
rect 378302 568046 378398 568102
rect 377778 567978 378398 568046
rect 377778 567922 377874 567978
rect 377930 567922 377998 567978
rect 378054 567922 378122 567978
rect 378178 567922 378246 567978
rect 378302 567922 378398 567978
rect 377778 550350 378398 567922
rect 377778 550294 377874 550350
rect 377930 550294 377998 550350
rect 378054 550294 378122 550350
rect 378178 550294 378246 550350
rect 378302 550294 378398 550350
rect 377778 550226 378398 550294
rect 377778 550170 377874 550226
rect 377930 550170 377998 550226
rect 378054 550170 378122 550226
rect 378178 550170 378246 550226
rect 378302 550170 378398 550226
rect 377778 550102 378398 550170
rect 377778 550046 377874 550102
rect 377930 550046 377998 550102
rect 378054 550046 378122 550102
rect 378178 550046 378246 550102
rect 378302 550046 378398 550102
rect 377778 549978 378398 550046
rect 377778 549922 377874 549978
rect 377930 549922 377998 549978
rect 378054 549922 378122 549978
rect 378178 549922 378246 549978
rect 378302 549922 378398 549978
rect 377778 532350 378398 549922
rect 377778 532294 377874 532350
rect 377930 532294 377998 532350
rect 378054 532294 378122 532350
rect 378178 532294 378246 532350
rect 378302 532294 378398 532350
rect 377778 532226 378398 532294
rect 377778 532170 377874 532226
rect 377930 532170 377998 532226
rect 378054 532170 378122 532226
rect 378178 532170 378246 532226
rect 378302 532170 378398 532226
rect 377778 532102 378398 532170
rect 377778 532046 377874 532102
rect 377930 532046 377998 532102
rect 378054 532046 378122 532102
rect 378178 532046 378246 532102
rect 378302 532046 378398 532102
rect 377778 531978 378398 532046
rect 377778 531922 377874 531978
rect 377930 531922 377998 531978
rect 378054 531922 378122 531978
rect 378178 531922 378246 531978
rect 378302 531922 378398 531978
rect 377778 514350 378398 531922
rect 377778 514294 377874 514350
rect 377930 514294 377998 514350
rect 378054 514294 378122 514350
rect 378178 514294 378246 514350
rect 378302 514294 378398 514350
rect 377778 514226 378398 514294
rect 377778 514170 377874 514226
rect 377930 514170 377998 514226
rect 378054 514170 378122 514226
rect 378178 514170 378246 514226
rect 378302 514170 378398 514226
rect 377778 514102 378398 514170
rect 377778 514046 377874 514102
rect 377930 514046 377998 514102
rect 378054 514046 378122 514102
rect 378178 514046 378246 514102
rect 378302 514046 378398 514102
rect 377778 513978 378398 514046
rect 377778 513922 377874 513978
rect 377930 513922 377998 513978
rect 378054 513922 378122 513978
rect 378178 513922 378246 513978
rect 378302 513922 378398 513978
rect 377778 496350 378398 513922
rect 377778 496294 377874 496350
rect 377930 496294 377998 496350
rect 378054 496294 378122 496350
rect 378178 496294 378246 496350
rect 378302 496294 378398 496350
rect 377778 496226 378398 496294
rect 377778 496170 377874 496226
rect 377930 496170 377998 496226
rect 378054 496170 378122 496226
rect 378178 496170 378246 496226
rect 378302 496170 378398 496226
rect 377778 496102 378398 496170
rect 377778 496046 377874 496102
rect 377930 496046 377998 496102
rect 378054 496046 378122 496102
rect 378178 496046 378246 496102
rect 378302 496046 378398 496102
rect 377778 495978 378398 496046
rect 377778 495922 377874 495978
rect 377930 495922 377998 495978
rect 378054 495922 378122 495978
rect 378178 495922 378246 495978
rect 378302 495922 378398 495978
rect 377778 478350 378398 495922
rect 377778 478294 377874 478350
rect 377930 478294 377998 478350
rect 378054 478294 378122 478350
rect 378178 478294 378246 478350
rect 378302 478294 378398 478350
rect 377778 478226 378398 478294
rect 377778 478170 377874 478226
rect 377930 478170 377998 478226
rect 378054 478170 378122 478226
rect 378178 478170 378246 478226
rect 378302 478170 378398 478226
rect 377778 478102 378398 478170
rect 377778 478046 377874 478102
rect 377930 478046 377998 478102
rect 378054 478046 378122 478102
rect 378178 478046 378246 478102
rect 378302 478046 378398 478102
rect 377778 477978 378398 478046
rect 377778 477922 377874 477978
rect 377930 477922 377998 477978
rect 378054 477922 378122 477978
rect 378178 477922 378246 477978
rect 378302 477922 378398 477978
rect 377778 460350 378398 477922
rect 377778 460294 377874 460350
rect 377930 460294 377998 460350
rect 378054 460294 378122 460350
rect 378178 460294 378246 460350
rect 378302 460294 378398 460350
rect 377778 460226 378398 460294
rect 377778 460170 377874 460226
rect 377930 460170 377998 460226
rect 378054 460170 378122 460226
rect 378178 460170 378246 460226
rect 378302 460170 378398 460226
rect 377778 460102 378398 460170
rect 377778 460046 377874 460102
rect 377930 460046 377998 460102
rect 378054 460046 378122 460102
rect 378178 460046 378246 460102
rect 378302 460046 378398 460102
rect 377778 459978 378398 460046
rect 377778 459922 377874 459978
rect 377930 459922 377998 459978
rect 378054 459922 378122 459978
rect 378178 459922 378246 459978
rect 378302 459922 378398 459978
rect 377778 442350 378398 459922
rect 377778 442294 377874 442350
rect 377930 442294 377998 442350
rect 378054 442294 378122 442350
rect 378178 442294 378246 442350
rect 378302 442294 378398 442350
rect 377778 442226 378398 442294
rect 377778 442170 377874 442226
rect 377930 442170 377998 442226
rect 378054 442170 378122 442226
rect 378178 442170 378246 442226
rect 378302 442170 378398 442226
rect 377778 442102 378398 442170
rect 377778 442046 377874 442102
rect 377930 442046 377998 442102
rect 378054 442046 378122 442102
rect 378178 442046 378246 442102
rect 378302 442046 378398 442102
rect 377778 441978 378398 442046
rect 377778 441922 377874 441978
rect 377930 441922 377998 441978
rect 378054 441922 378122 441978
rect 378178 441922 378246 441978
rect 378302 441922 378398 441978
rect 377778 424350 378398 441922
rect 377778 424294 377874 424350
rect 377930 424294 377998 424350
rect 378054 424294 378122 424350
rect 378178 424294 378246 424350
rect 378302 424294 378398 424350
rect 377778 424226 378398 424294
rect 377778 424170 377874 424226
rect 377930 424170 377998 424226
rect 378054 424170 378122 424226
rect 378178 424170 378246 424226
rect 378302 424170 378398 424226
rect 377778 424102 378398 424170
rect 377778 424046 377874 424102
rect 377930 424046 377998 424102
rect 378054 424046 378122 424102
rect 378178 424046 378246 424102
rect 378302 424046 378398 424102
rect 377778 423978 378398 424046
rect 377778 423922 377874 423978
rect 377930 423922 377998 423978
rect 378054 423922 378122 423978
rect 378178 423922 378246 423978
rect 378302 423922 378398 423978
rect 377778 406350 378398 423922
rect 377778 406294 377874 406350
rect 377930 406294 377998 406350
rect 378054 406294 378122 406350
rect 378178 406294 378246 406350
rect 378302 406294 378398 406350
rect 377778 406226 378398 406294
rect 377778 406170 377874 406226
rect 377930 406170 377998 406226
rect 378054 406170 378122 406226
rect 378178 406170 378246 406226
rect 378302 406170 378398 406226
rect 377778 406102 378398 406170
rect 377778 406046 377874 406102
rect 377930 406046 377998 406102
rect 378054 406046 378122 406102
rect 378178 406046 378246 406102
rect 378302 406046 378398 406102
rect 377778 405978 378398 406046
rect 377778 405922 377874 405978
rect 377930 405922 377998 405978
rect 378054 405922 378122 405978
rect 378178 405922 378246 405978
rect 378302 405922 378398 405978
rect 377778 388350 378398 405922
rect 377778 388294 377874 388350
rect 377930 388294 377998 388350
rect 378054 388294 378122 388350
rect 378178 388294 378246 388350
rect 378302 388294 378398 388350
rect 377778 388226 378398 388294
rect 377778 388170 377874 388226
rect 377930 388170 377998 388226
rect 378054 388170 378122 388226
rect 378178 388170 378246 388226
rect 378302 388170 378398 388226
rect 377778 388102 378398 388170
rect 377778 388046 377874 388102
rect 377930 388046 377998 388102
rect 378054 388046 378122 388102
rect 378178 388046 378246 388102
rect 378302 388046 378398 388102
rect 377778 387978 378398 388046
rect 377778 387922 377874 387978
rect 377930 387922 377998 387978
rect 378054 387922 378122 387978
rect 378178 387922 378246 387978
rect 378302 387922 378398 387978
rect 377778 370350 378398 387922
rect 404778 597212 405398 598268
rect 404778 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 405398 597212
rect 404778 597088 405398 597156
rect 404778 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 405398 597088
rect 404778 596964 405398 597032
rect 404778 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 405398 596964
rect 404778 596840 405398 596908
rect 404778 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 405398 596840
rect 404778 580350 405398 596784
rect 404778 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 405398 580350
rect 404778 580226 405398 580294
rect 404778 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 405398 580226
rect 404778 580102 405398 580170
rect 404778 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 405398 580102
rect 404778 579978 405398 580046
rect 404778 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 405398 579978
rect 404778 562350 405398 579922
rect 404778 562294 404874 562350
rect 404930 562294 404998 562350
rect 405054 562294 405122 562350
rect 405178 562294 405246 562350
rect 405302 562294 405398 562350
rect 404778 562226 405398 562294
rect 404778 562170 404874 562226
rect 404930 562170 404998 562226
rect 405054 562170 405122 562226
rect 405178 562170 405246 562226
rect 405302 562170 405398 562226
rect 404778 562102 405398 562170
rect 404778 562046 404874 562102
rect 404930 562046 404998 562102
rect 405054 562046 405122 562102
rect 405178 562046 405246 562102
rect 405302 562046 405398 562102
rect 404778 561978 405398 562046
rect 404778 561922 404874 561978
rect 404930 561922 404998 561978
rect 405054 561922 405122 561978
rect 405178 561922 405246 561978
rect 405302 561922 405398 561978
rect 404778 544350 405398 561922
rect 404778 544294 404874 544350
rect 404930 544294 404998 544350
rect 405054 544294 405122 544350
rect 405178 544294 405246 544350
rect 405302 544294 405398 544350
rect 404778 544226 405398 544294
rect 404778 544170 404874 544226
rect 404930 544170 404998 544226
rect 405054 544170 405122 544226
rect 405178 544170 405246 544226
rect 405302 544170 405398 544226
rect 404778 544102 405398 544170
rect 404778 544046 404874 544102
rect 404930 544046 404998 544102
rect 405054 544046 405122 544102
rect 405178 544046 405246 544102
rect 405302 544046 405398 544102
rect 404778 543978 405398 544046
rect 404778 543922 404874 543978
rect 404930 543922 404998 543978
rect 405054 543922 405122 543978
rect 405178 543922 405246 543978
rect 405302 543922 405398 543978
rect 404778 526350 405398 543922
rect 404778 526294 404874 526350
rect 404930 526294 404998 526350
rect 405054 526294 405122 526350
rect 405178 526294 405246 526350
rect 405302 526294 405398 526350
rect 404778 526226 405398 526294
rect 404778 526170 404874 526226
rect 404930 526170 404998 526226
rect 405054 526170 405122 526226
rect 405178 526170 405246 526226
rect 405302 526170 405398 526226
rect 404778 526102 405398 526170
rect 404778 526046 404874 526102
rect 404930 526046 404998 526102
rect 405054 526046 405122 526102
rect 405178 526046 405246 526102
rect 405302 526046 405398 526102
rect 404778 525978 405398 526046
rect 404778 525922 404874 525978
rect 404930 525922 404998 525978
rect 405054 525922 405122 525978
rect 405178 525922 405246 525978
rect 405302 525922 405398 525978
rect 404778 508350 405398 525922
rect 404778 508294 404874 508350
rect 404930 508294 404998 508350
rect 405054 508294 405122 508350
rect 405178 508294 405246 508350
rect 405302 508294 405398 508350
rect 404778 508226 405398 508294
rect 404778 508170 404874 508226
rect 404930 508170 404998 508226
rect 405054 508170 405122 508226
rect 405178 508170 405246 508226
rect 405302 508170 405398 508226
rect 404778 508102 405398 508170
rect 404778 508046 404874 508102
rect 404930 508046 404998 508102
rect 405054 508046 405122 508102
rect 405178 508046 405246 508102
rect 405302 508046 405398 508102
rect 404778 507978 405398 508046
rect 404778 507922 404874 507978
rect 404930 507922 404998 507978
rect 405054 507922 405122 507978
rect 405178 507922 405246 507978
rect 405302 507922 405398 507978
rect 404778 490350 405398 507922
rect 404778 490294 404874 490350
rect 404930 490294 404998 490350
rect 405054 490294 405122 490350
rect 405178 490294 405246 490350
rect 405302 490294 405398 490350
rect 404778 490226 405398 490294
rect 404778 490170 404874 490226
rect 404930 490170 404998 490226
rect 405054 490170 405122 490226
rect 405178 490170 405246 490226
rect 405302 490170 405398 490226
rect 404778 490102 405398 490170
rect 404778 490046 404874 490102
rect 404930 490046 404998 490102
rect 405054 490046 405122 490102
rect 405178 490046 405246 490102
rect 405302 490046 405398 490102
rect 404778 489978 405398 490046
rect 404778 489922 404874 489978
rect 404930 489922 404998 489978
rect 405054 489922 405122 489978
rect 405178 489922 405246 489978
rect 405302 489922 405398 489978
rect 404778 472350 405398 489922
rect 404778 472294 404874 472350
rect 404930 472294 404998 472350
rect 405054 472294 405122 472350
rect 405178 472294 405246 472350
rect 405302 472294 405398 472350
rect 404778 472226 405398 472294
rect 404778 472170 404874 472226
rect 404930 472170 404998 472226
rect 405054 472170 405122 472226
rect 405178 472170 405246 472226
rect 405302 472170 405398 472226
rect 404778 472102 405398 472170
rect 404778 472046 404874 472102
rect 404930 472046 404998 472102
rect 405054 472046 405122 472102
rect 405178 472046 405246 472102
rect 405302 472046 405398 472102
rect 404778 471978 405398 472046
rect 404778 471922 404874 471978
rect 404930 471922 404998 471978
rect 405054 471922 405122 471978
rect 405178 471922 405246 471978
rect 405302 471922 405398 471978
rect 404778 454350 405398 471922
rect 404778 454294 404874 454350
rect 404930 454294 404998 454350
rect 405054 454294 405122 454350
rect 405178 454294 405246 454350
rect 405302 454294 405398 454350
rect 404778 454226 405398 454294
rect 404778 454170 404874 454226
rect 404930 454170 404998 454226
rect 405054 454170 405122 454226
rect 405178 454170 405246 454226
rect 405302 454170 405398 454226
rect 404778 454102 405398 454170
rect 404778 454046 404874 454102
rect 404930 454046 404998 454102
rect 405054 454046 405122 454102
rect 405178 454046 405246 454102
rect 405302 454046 405398 454102
rect 404778 453978 405398 454046
rect 404778 453922 404874 453978
rect 404930 453922 404998 453978
rect 405054 453922 405122 453978
rect 405178 453922 405246 453978
rect 405302 453922 405398 453978
rect 404778 436350 405398 453922
rect 404778 436294 404874 436350
rect 404930 436294 404998 436350
rect 405054 436294 405122 436350
rect 405178 436294 405246 436350
rect 405302 436294 405398 436350
rect 404778 436226 405398 436294
rect 404778 436170 404874 436226
rect 404930 436170 404998 436226
rect 405054 436170 405122 436226
rect 405178 436170 405246 436226
rect 405302 436170 405398 436226
rect 404778 436102 405398 436170
rect 404778 436046 404874 436102
rect 404930 436046 404998 436102
rect 405054 436046 405122 436102
rect 405178 436046 405246 436102
rect 405302 436046 405398 436102
rect 404778 435978 405398 436046
rect 404778 435922 404874 435978
rect 404930 435922 404998 435978
rect 405054 435922 405122 435978
rect 405178 435922 405246 435978
rect 405302 435922 405398 435978
rect 404778 418350 405398 435922
rect 404778 418294 404874 418350
rect 404930 418294 404998 418350
rect 405054 418294 405122 418350
rect 405178 418294 405246 418350
rect 405302 418294 405398 418350
rect 404778 418226 405398 418294
rect 404778 418170 404874 418226
rect 404930 418170 404998 418226
rect 405054 418170 405122 418226
rect 405178 418170 405246 418226
rect 405302 418170 405398 418226
rect 404778 418102 405398 418170
rect 404778 418046 404874 418102
rect 404930 418046 404998 418102
rect 405054 418046 405122 418102
rect 405178 418046 405246 418102
rect 405302 418046 405398 418102
rect 404778 417978 405398 418046
rect 404778 417922 404874 417978
rect 404930 417922 404998 417978
rect 405054 417922 405122 417978
rect 405178 417922 405246 417978
rect 405302 417922 405398 417978
rect 404778 400350 405398 417922
rect 404778 400294 404874 400350
rect 404930 400294 404998 400350
rect 405054 400294 405122 400350
rect 405178 400294 405246 400350
rect 405302 400294 405398 400350
rect 404778 400226 405398 400294
rect 404778 400170 404874 400226
rect 404930 400170 404998 400226
rect 405054 400170 405122 400226
rect 405178 400170 405246 400226
rect 405302 400170 405398 400226
rect 404778 400102 405398 400170
rect 404778 400046 404874 400102
rect 404930 400046 404998 400102
rect 405054 400046 405122 400102
rect 405178 400046 405246 400102
rect 405302 400046 405398 400102
rect 404778 399978 405398 400046
rect 404778 399922 404874 399978
rect 404930 399922 404998 399978
rect 405054 399922 405122 399978
rect 405178 399922 405246 399978
rect 405302 399922 405398 399978
rect 404778 382350 405398 399922
rect 404778 382294 404874 382350
rect 404930 382294 404998 382350
rect 405054 382294 405122 382350
rect 405178 382294 405246 382350
rect 405302 382294 405398 382350
rect 404778 382226 405398 382294
rect 404778 382170 404874 382226
rect 404930 382170 404998 382226
rect 405054 382170 405122 382226
rect 405178 382170 405246 382226
rect 405302 382170 405398 382226
rect 404778 382102 405398 382170
rect 404778 382046 404874 382102
rect 404930 382046 404998 382102
rect 405054 382046 405122 382102
rect 405178 382046 405246 382102
rect 405302 382046 405398 382102
rect 404778 381978 405398 382046
rect 404778 381922 404874 381978
rect 404930 381922 404998 381978
rect 405054 381922 405122 381978
rect 405178 381922 405246 381978
rect 405302 381922 405398 381978
rect 377778 370294 377874 370350
rect 377930 370294 377998 370350
rect 378054 370294 378122 370350
rect 378178 370294 378246 370350
rect 378302 370294 378398 370350
rect 377778 370226 378398 370294
rect 377778 370170 377874 370226
rect 377930 370170 377998 370226
rect 378054 370170 378122 370226
rect 378178 370170 378246 370226
rect 378302 370170 378398 370226
rect 377778 370102 378398 370170
rect 377778 370046 377874 370102
rect 377930 370046 377998 370102
rect 378054 370046 378122 370102
rect 378178 370046 378246 370102
rect 378302 370046 378398 370102
rect 377778 369978 378398 370046
rect 377778 369922 377874 369978
rect 377930 369922 377998 369978
rect 378054 369922 378122 369978
rect 378178 369922 378246 369978
rect 378302 369922 378398 369978
rect 377778 352350 378398 369922
rect 377778 352294 377874 352350
rect 377930 352294 377998 352350
rect 378054 352294 378122 352350
rect 378178 352294 378246 352350
rect 378302 352294 378398 352350
rect 377778 352226 378398 352294
rect 377778 352170 377874 352226
rect 377930 352170 377998 352226
rect 378054 352170 378122 352226
rect 378178 352170 378246 352226
rect 378302 352170 378398 352226
rect 377778 352102 378398 352170
rect 377778 352046 377874 352102
rect 377930 352046 377998 352102
rect 378054 352046 378122 352102
rect 378178 352046 378246 352102
rect 378302 352046 378398 352102
rect 377778 351978 378398 352046
rect 377778 351922 377874 351978
rect 377930 351922 377998 351978
rect 378054 351922 378122 351978
rect 378178 351922 378246 351978
rect 378302 351922 378398 351978
rect 377778 334350 378398 351922
rect 377778 334294 377874 334350
rect 377930 334294 377998 334350
rect 378054 334294 378122 334350
rect 378178 334294 378246 334350
rect 378302 334294 378398 334350
rect 377778 334226 378398 334294
rect 377778 334170 377874 334226
rect 377930 334170 377998 334226
rect 378054 334170 378122 334226
rect 378178 334170 378246 334226
rect 378302 334170 378398 334226
rect 377778 334102 378398 334170
rect 377778 334046 377874 334102
rect 377930 334046 377998 334102
rect 378054 334046 378122 334102
rect 378178 334046 378246 334102
rect 378302 334046 378398 334102
rect 377778 333978 378398 334046
rect 377778 333922 377874 333978
rect 377930 333922 377998 333978
rect 378054 333922 378122 333978
rect 378178 333922 378246 333978
rect 378302 333922 378398 333978
rect 377580 324884 377636 324894
rect 376124 324772 376180 324782
rect 374058 310294 374154 310350
rect 374210 310294 374278 310350
rect 374334 310294 374402 310350
rect 374458 310294 374526 310350
rect 374582 310294 374678 310350
rect 374058 310226 374678 310294
rect 374058 310170 374154 310226
rect 374210 310170 374278 310226
rect 374334 310170 374402 310226
rect 374458 310170 374526 310226
rect 374582 310170 374678 310226
rect 374058 310102 374678 310170
rect 374058 310046 374154 310102
rect 374210 310046 374278 310102
rect 374334 310046 374402 310102
rect 374458 310046 374526 310102
rect 374582 310046 374678 310102
rect 374058 309978 374678 310046
rect 374058 309922 374154 309978
rect 374210 309922 374278 309978
rect 374334 309922 374402 309978
rect 374458 309922 374526 309978
rect 374582 309922 374678 309978
rect 373884 308084 373940 308094
rect 373884 298564 373940 308028
rect 373884 298498 373940 298508
rect 373772 295698 373828 295708
rect 373772 294644 373828 294654
rect 372876 293860 372932 293870
rect 372092 292404 372148 292414
rect 372092 277172 372148 292348
rect 372092 277106 372148 277116
rect 372428 289044 372484 289054
rect 372428 273812 372484 288988
rect 372428 273746 372484 273756
rect 372652 275716 372708 275726
rect 370972 271348 371028 271358
rect 370860 270658 370916 270668
rect 370748 266308 370804 266318
rect 370748 231252 370804 266252
rect 370748 231186 370804 231196
rect 370636 224354 370692 224364
rect 370636 224084 370692 224094
rect 370636 216580 370692 224028
rect 370636 216514 370692 216524
rect 370412 199042 370468 199052
rect 370524 215236 370580 215246
rect 370188 192322 370244 192332
rect 370076 184706 370132 184716
rect 214448 184350 214768 184384
rect 214448 184294 214518 184350
rect 214574 184294 214642 184350
rect 214698 184294 214768 184350
rect 214448 184226 214768 184294
rect 214448 184170 214518 184226
rect 214574 184170 214642 184226
rect 214698 184170 214768 184226
rect 214448 184102 214768 184170
rect 214448 184046 214518 184102
rect 214574 184046 214642 184102
rect 214698 184046 214768 184102
rect 214448 183978 214768 184046
rect 214448 183922 214518 183978
rect 214574 183922 214642 183978
rect 214698 183922 214768 183978
rect 214448 183888 214768 183922
rect 245168 184350 245488 184384
rect 245168 184294 245238 184350
rect 245294 184294 245362 184350
rect 245418 184294 245488 184350
rect 245168 184226 245488 184294
rect 245168 184170 245238 184226
rect 245294 184170 245362 184226
rect 245418 184170 245488 184226
rect 245168 184102 245488 184170
rect 245168 184046 245238 184102
rect 245294 184046 245362 184102
rect 245418 184046 245488 184102
rect 245168 183978 245488 184046
rect 245168 183922 245238 183978
rect 245294 183922 245362 183978
rect 245418 183922 245488 183978
rect 245168 183888 245488 183922
rect 275888 184350 276208 184384
rect 275888 184294 275958 184350
rect 276014 184294 276082 184350
rect 276138 184294 276208 184350
rect 275888 184226 276208 184294
rect 275888 184170 275958 184226
rect 276014 184170 276082 184226
rect 276138 184170 276208 184226
rect 275888 184102 276208 184170
rect 275888 184046 275958 184102
rect 276014 184046 276082 184102
rect 276138 184046 276208 184102
rect 275888 183978 276208 184046
rect 275888 183922 275958 183978
rect 276014 183922 276082 183978
rect 276138 183922 276208 183978
rect 275888 183888 276208 183922
rect 306608 184350 306928 184384
rect 306608 184294 306678 184350
rect 306734 184294 306802 184350
rect 306858 184294 306928 184350
rect 306608 184226 306928 184294
rect 306608 184170 306678 184226
rect 306734 184170 306802 184226
rect 306858 184170 306928 184226
rect 306608 184102 306928 184170
rect 306608 184046 306678 184102
rect 306734 184046 306802 184102
rect 306858 184046 306928 184102
rect 306608 183978 306928 184046
rect 306608 183922 306678 183978
rect 306734 183922 306802 183978
rect 306858 183922 306928 183978
rect 306608 183888 306928 183922
rect 337328 184350 337648 184384
rect 337328 184294 337398 184350
rect 337454 184294 337522 184350
rect 337578 184294 337648 184350
rect 337328 184226 337648 184294
rect 337328 184170 337398 184226
rect 337454 184170 337522 184226
rect 337578 184170 337648 184226
rect 337328 184102 337648 184170
rect 337328 184046 337398 184102
rect 337454 184046 337522 184102
rect 337578 184046 337648 184102
rect 337328 183978 337648 184046
rect 337328 183922 337398 183978
rect 337454 183922 337522 183978
rect 337578 183922 337648 183978
rect 337328 183888 337648 183922
rect 368048 184350 368368 184384
rect 368048 184294 368118 184350
rect 368174 184294 368242 184350
rect 368298 184294 368368 184350
rect 368048 184226 368368 184294
rect 368048 184170 368118 184226
rect 368174 184170 368242 184226
rect 368298 184170 368368 184226
rect 368048 184102 368368 184170
rect 368048 184046 368118 184102
rect 368174 184046 368242 184102
rect 368298 184046 368368 184102
rect 368048 183978 368368 184046
rect 368048 183922 368118 183978
rect 368174 183922 368242 183978
rect 368298 183922 368368 183978
rect 368048 183888 368368 183922
rect 370188 176708 370244 176718
rect 229808 172350 230128 172384
rect 229808 172294 229878 172350
rect 229934 172294 230002 172350
rect 230058 172294 230128 172350
rect 229808 172226 230128 172294
rect 229808 172170 229878 172226
rect 229934 172170 230002 172226
rect 230058 172170 230128 172226
rect 229808 172102 230128 172170
rect 229808 172046 229878 172102
rect 229934 172046 230002 172102
rect 230058 172046 230128 172102
rect 229808 171978 230128 172046
rect 229808 171922 229878 171978
rect 229934 171922 230002 171978
rect 230058 171922 230128 171978
rect 229808 171888 230128 171922
rect 260528 172350 260848 172384
rect 260528 172294 260598 172350
rect 260654 172294 260722 172350
rect 260778 172294 260848 172350
rect 260528 172226 260848 172294
rect 260528 172170 260598 172226
rect 260654 172170 260722 172226
rect 260778 172170 260848 172226
rect 260528 172102 260848 172170
rect 260528 172046 260598 172102
rect 260654 172046 260722 172102
rect 260778 172046 260848 172102
rect 260528 171978 260848 172046
rect 260528 171922 260598 171978
rect 260654 171922 260722 171978
rect 260778 171922 260848 171978
rect 260528 171888 260848 171922
rect 291248 172350 291568 172384
rect 291248 172294 291318 172350
rect 291374 172294 291442 172350
rect 291498 172294 291568 172350
rect 291248 172226 291568 172294
rect 291248 172170 291318 172226
rect 291374 172170 291442 172226
rect 291498 172170 291568 172226
rect 291248 172102 291568 172170
rect 291248 172046 291318 172102
rect 291374 172046 291442 172102
rect 291498 172046 291568 172102
rect 291248 171978 291568 172046
rect 291248 171922 291318 171978
rect 291374 171922 291442 171978
rect 291498 171922 291568 171978
rect 291248 171888 291568 171922
rect 321968 172350 322288 172384
rect 321968 172294 322038 172350
rect 322094 172294 322162 172350
rect 322218 172294 322288 172350
rect 321968 172226 322288 172294
rect 321968 172170 322038 172226
rect 322094 172170 322162 172226
rect 322218 172170 322288 172226
rect 321968 172102 322288 172170
rect 321968 172046 322038 172102
rect 322094 172046 322162 172102
rect 322218 172046 322288 172102
rect 321968 171978 322288 172046
rect 321968 171922 322038 171978
rect 322094 171922 322162 171978
rect 322218 171922 322288 171978
rect 321968 171888 322288 171922
rect 352688 172350 353008 172384
rect 352688 172294 352758 172350
rect 352814 172294 352882 172350
rect 352938 172294 353008 172350
rect 352688 172226 353008 172294
rect 352688 172170 352758 172226
rect 352814 172170 352882 172226
rect 352938 172170 353008 172226
rect 352688 172102 353008 172170
rect 352688 172046 352758 172102
rect 352814 172046 352882 172102
rect 352938 172046 353008 172102
rect 352688 171978 353008 172046
rect 352688 171922 352758 171978
rect 352814 171922 352882 171978
rect 352938 171922 353008 171978
rect 352688 171888 353008 171922
rect 370076 169204 370132 169214
rect 214448 166350 214768 166384
rect 214448 166294 214518 166350
rect 214574 166294 214642 166350
rect 214698 166294 214768 166350
rect 214448 166226 214768 166294
rect 214448 166170 214518 166226
rect 214574 166170 214642 166226
rect 214698 166170 214768 166226
rect 214448 166102 214768 166170
rect 214448 166046 214518 166102
rect 214574 166046 214642 166102
rect 214698 166046 214768 166102
rect 214448 165978 214768 166046
rect 214448 165922 214518 165978
rect 214574 165922 214642 165978
rect 214698 165922 214768 165978
rect 214448 165888 214768 165922
rect 245168 166350 245488 166384
rect 245168 166294 245238 166350
rect 245294 166294 245362 166350
rect 245418 166294 245488 166350
rect 245168 166226 245488 166294
rect 245168 166170 245238 166226
rect 245294 166170 245362 166226
rect 245418 166170 245488 166226
rect 245168 166102 245488 166170
rect 245168 166046 245238 166102
rect 245294 166046 245362 166102
rect 245418 166046 245488 166102
rect 245168 165978 245488 166046
rect 245168 165922 245238 165978
rect 245294 165922 245362 165978
rect 245418 165922 245488 165978
rect 245168 165888 245488 165922
rect 275888 166350 276208 166384
rect 275888 166294 275958 166350
rect 276014 166294 276082 166350
rect 276138 166294 276208 166350
rect 275888 166226 276208 166294
rect 275888 166170 275958 166226
rect 276014 166170 276082 166226
rect 276138 166170 276208 166226
rect 275888 166102 276208 166170
rect 275888 166046 275958 166102
rect 276014 166046 276082 166102
rect 276138 166046 276208 166102
rect 275888 165978 276208 166046
rect 275888 165922 275958 165978
rect 276014 165922 276082 165978
rect 276138 165922 276208 165978
rect 275888 165888 276208 165922
rect 306608 166350 306928 166384
rect 306608 166294 306678 166350
rect 306734 166294 306802 166350
rect 306858 166294 306928 166350
rect 306608 166226 306928 166294
rect 306608 166170 306678 166226
rect 306734 166170 306802 166226
rect 306858 166170 306928 166226
rect 306608 166102 306928 166170
rect 306608 166046 306678 166102
rect 306734 166046 306802 166102
rect 306858 166046 306928 166102
rect 306608 165978 306928 166046
rect 306608 165922 306678 165978
rect 306734 165922 306802 165978
rect 306858 165922 306928 165978
rect 306608 165888 306928 165922
rect 337328 166350 337648 166384
rect 337328 166294 337398 166350
rect 337454 166294 337522 166350
rect 337578 166294 337648 166350
rect 337328 166226 337648 166294
rect 337328 166170 337398 166226
rect 337454 166170 337522 166226
rect 337578 166170 337648 166226
rect 337328 166102 337648 166170
rect 337328 166046 337398 166102
rect 337454 166046 337522 166102
rect 337578 166046 337648 166102
rect 337328 165978 337648 166046
rect 337328 165922 337398 165978
rect 337454 165922 337522 165978
rect 337578 165922 337648 165978
rect 337328 165888 337648 165922
rect 368048 166350 368368 166384
rect 368048 166294 368118 166350
rect 368174 166294 368242 166350
rect 368298 166294 368368 166350
rect 368048 166226 368368 166294
rect 368048 166170 368118 166226
rect 368174 166170 368242 166226
rect 368298 166170 368368 166226
rect 368048 166102 368368 166170
rect 368048 166046 368118 166102
rect 368174 166046 368242 166102
rect 368298 166046 368368 166102
rect 368048 165978 368368 166046
rect 368048 165922 368118 165978
rect 368174 165922 368242 165978
rect 368298 165922 368368 165978
rect 368048 165888 368368 165922
rect 210588 161298 210644 161308
rect 210364 161074 210420 161084
rect 229808 154350 230128 154384
rect 229808 154294 229878 154350
rect 229934 154294 230002 154350
rect 230058 154294 230128 154350
rect 229808 154226 230128 154294
rect 229808 154170 229878 154226
rect 229934 154170 230002 154226
rect 230058 154170 230128 154226
rect 229808 154102 230128 154170
rect 229808 154046 229878 154102
rect 229934 154046 230002 154102
rect 230058 154046 230128 154102
rect 229808 153978 230128 154046
rect 229808 153922 229878 153978
rect 229934 153922 230002 153978
rect 230058 153922 230128 153978
rect 229808 153888 230128 153922
rect 260528 154350 260848 154384
rect 260528 154294 260598 154350
rect 260654 154294 260722 154350
rect 260778 154294 260848 154350
rect 260528 154226 260848 154294
rect 260528 154170 260598 154226
rect 260654 154170 260722 154226
rect 260778 154170 260848 154226
rect 260528 154102 260848 154170
rect 260528 154046 260598 154102
rect 260654 154046 260722 154102
rect 260778 154046 260848 154102
rect 260528 153978 260848 154046
rect 260528 153922 260598 153978
rect 260654 153922 260722 153978
rect 260778 153922 260848 153978
rect 260528 153888 260848 153922
rect 291248 154350 291568 154384
rect 291248 154294 291318 154350
rect 291374 154294 291442 154350
rect 291498 154294 291568 154350
rect 291248 154226 291568 154294
rect 291248 154170 291318 154226
rect 291374 154170 291442 154226
rect 291498 154170 291568 154226
rect 291248 154102 291568 154170
rect 291248 154046 291318 154102
rect 291374 154046 291442 154102
rect 291498 154046 291568 154102
rect 291248 153978 291568 154046
rect 291248 153922 291318 153978
rect 291374 153922 291442 153978
rect 291498 153922 291568 153978
rect 291248 153888 291568 153922
rect 321968 154350 322288 154384
rect 321968 154294 322038 154350
rect 322094 154294 322162 154350
rect 322218 154294 322288 154350
rect 321968 154226 322288 154294
rect 321968 154170 322038 154226
rect 322094 154170 322162 154226
rect 322218 154170 322288 154226
rect 321968 154102 322288 154170
rect 321968 154046 322038 154102
rect 322094 154046 322162 154102
rect 322218 154046 322288 154102
rect 321968 153978 322288 154046
rect 321968 153922 322038 153978
rect 322094 153922 322162 153978
rect 322218 153922 322288 153978
rect 321968 153888 322288 153922
rect 352688 154350 353008 154384
rect 352688 154294 352758 154350
rect 352814 154294 352882 154350
rect 352938 154294 353008 154350
rect 352688 154226 353008 154294
rect 352688 154170 352758 154226
rect 352814 154170 352882 154226
rect 352938 154170 353008 154226
rect 352688 154102 353008 154170
rect 352688 154046 352758 154102
rect 352814 154046 352882 154102
rect 352938 154046 353008 154102
rect 352688 153978 353008 154046
rect 352688 153922 352758 153978
rect 352814 153922 352882 153978
rect 352938 153922 353008 153978
rect 352688 153888 353008 153922
rect 214448 148350 214768 148384
rect 214448 148294 214518 148350
rect 214574 148294 214642 148350
rect 214698 148294 214768 148350
rect 214448 148226 214768 148294
rect 214448 148170 214518 148226
rect 214574 148170 214642 148226
rect 214698 148170 214768 148226
rect 214448 148102 214768 148170
rect 214448 148046 214518 148102
rect 214574 148046 214642 148102
rect 214698 148046 214768 148102
rect 214448 147978 214768 148046
rect 214448 147922 214518 147978
rect 214574 147922 214642 147978
rect 214698 147922 214768 147978
rect 214448 147888 214768 147922
rect 245168 148350 245488 148384
rect 245168 148294 245238 148350
rect 245294 148294 245362 148350
rect 245418 148294 245488 148350
rect 245168 148226 245488 148294
rect 245168 148170 245238 148226
rect 245294 148170 245362 148226
rect 245418 148170 245488 148226
rect 245168 148102 245488 148170
rect 245168 148046 245238 148102
rect 245294 148046 245362 148102
rect 245418 148046 245488 148102
rect 245168 147978 245488 148046
rect 245168 147922 245238 147978
rect 245294 147922 245362 147978
rect 245418 147922 245488 147978
rect 245168 147888 245488 147922
rect 275888 148350 276208 148384
rect 275888 148294 275958 148350
rect 276014 148294 276082 148350
rect 276138 148294 276208 148350
rect 275888 148226 276208 148294
rect 275888 148170 275958 148226
rect 276014 148170 276082 148226
rect 276138 148170 276208 148226
rect 275888 148102 276208 148170
rect 275888 148046 275958 148102
rect 276014 148046 276082 148102
rect 276138 148046 276208 148102
rect 275888 147978 276208 148046
rect 275888 147922 275958 147978
rect 276014 147922 276082 147978
rect 276138 147922 276208 147978
rect 275888 147888 276208 147922
rect 306608 148350 306928 148384
rect 306608 148294 306678 148350
rect 306734 148294 306802 148350
rect 306858 148294 306928 148350
rect 306608 148226 306928 148294
rect 306608 148170 306678 148226
rect 306734 148170 306802 148226
rect 306858 148170 306928 148226
rect 306608 148102 306928 148170
rect 306608 148046 306678 148102
rect 306734 148046 306802 148102
rect 306858 148046 306928 148102
rect 306608 147978 306928 148046
rect 306608 147922 306678 147978
rect 306734 147922 306802 147978
rect 306858 147922 306928 147978
rect 306608 147888 306928 147922
rect 337328 148350 337648 148384
rect 337328 148294 337398 148350
rect 337454 148294 337522 148350
rect 337578 148294 337648 148350
rect 337328 148226 337648 148294
rect 337328 148170 337398 148226
rect 337454 148170 337522 148226
rect 337578 148170 337648 148226
rect 337328 148102 337648 148170
rect 337328 148046 337398 148102
rect 337454 148046 337522 148102
rect 337578 148046 337648 148102
rect 337328 147978 337648 148046
rect 337328 147922 337398 147978
rect 337454 147922 337522 147978
rect 337578 147922 337648 147978
rect 337328 147888 337648 147922
rect 368048 148350 368368 148384
rect 368048 148294 368118 148350
rect 368174 148294 368242 148350
rect 368298 148294 368368 148350
rect 368048 148226 368368 148294
rect 368048 148170 368118 148226
rect 368174 148170 368242 148226
rect 368298 148170 368368 148226
rect 368048 148102 368368 148170
rect 368048 148046 368118 148102
rect 368174 148046 368242 148102
rect 368298 148046 368368 148102
rect 368048 147978 368368 148046
rect 368048 147922 368118 147978
rect 368174 147922 368242 147978
rect 368298 147922 368368 147978
rect 368048 147888 368368 147922
rect 229808 136350 230128 136384
rect 229808 136294 229878 136350
rect 229934 136294 230002 136350
rect 230058 136294 230128 136350
rect 229808 136226 230128 136294
rect 229808 136170 229878 136226
rect 229934 136170 230002 136226
rect 230058 136170 230128 136226
rect 229808 136102 230128 136170
rect 229808 136046 229878 136102
rect 229934 136046 230002 136102
rect 230058 136046 230128 136102
rect 229808 135978 230128 136046
rect 229808 135922 229878 135978
rect 229934 135922 230002 135978
rect 230058 135922 230128 135978
rect 229808 135888 230128 135922
rect 260528 136350 260848 136384
rect 260528 136294 260598 136350
rect 260654 136294 260722 136350
rect 260778 136294 260848 136350
rect 260528 136226 260848 136294
rect 260528 136170 260598 136226
rect 260654 136170 260722 136226
rect 260778 136170 260848 136226
rect 260528 136102 260848 136170
rect 260528 136046 260598 136102
rect 260654 136046 260722 136102
rect 260778 136046 260848 136102
rect 260528 135978 260848 136046
rect 260528 135922 260598 135978
rect 260654 135922 260722 135978
rect 260778 135922 260848 135978
rect 260528 135888 260848 135922
rect 291248 136350 291568 136384
rect 291248 136294 291318 136350
rect 291374 136294 291442 136350
rect 291498 136294 291568 136350
rect 291248 136226 291568 136294
rect 291248 136170 291318 136226
rect 291374 136170 291442 136226
rect 291498 136170 291568 136226
rect 291248 136102 291568 136170
rect 291248 136046 291318 136102
rect 291374 136046 291442 136102
rect 291498 136046 291568 136102
rect 291248 135978 291568 136046
rect 291248 135922 291318 135978
rect 291374 135922 291442 135978
rect 291498 135922 291568 135978
rect 291248 135888 291568 135922
rect 321968 136350 322288 136384
rect 321968 136294 322038 136350
rect 322094 136294 322162 136350
rect 322218 136294 322288 136350
rect 321968 136226 322288 136294
rect 321968 136170 322038 136226
rect 322094 136170 322162 136226
rect 322218 136170 322288 136226
rect 321968 136102 322288 136170
rect 321968 136046 322038 136102
rect 322094 136046 322162 136102
rect 322218 136046 322288 136102
rect 321968 135978 322288 136046
rect 321968 135922 322038 135978
rect 322094 135922 322162 135978
rect 322218 135922 322288 135978
rect 321968 135888 322288 135922
rect 352688 136350 353008 136384
rect 352688 136294 352758 136350
rect 352814 136294 352882 136350
rect 352938 136294 353008 136350
rect 352688 136226 353008 136294
rect 352688 136170 352758 136226
rect 352814 136170 352882 136226
rect 352938 136170 353008 136226
rect 352688 136102 353008 136170
rect 352688 136046 352758 136102
rect 352814 136046 352882 136102
rect 352938 136046 353008 136102
rect 352688 135978 353008 136046
rect 352688 135922 352758 135978
rect 352814 135922 352882 135978
rect 352938 135922 353008 135978
rect 352688 135888 353008 135922
rect 209692 133746 209748 133756
rect 214448 130350 214768 130384
rect 214448 130294 214518 130350
rect 214574 130294 214642 130350
rect 214698 130294 214768 130350
rect 214448 130226 214768 130294
rect 214448 130170 214518 130226
rect 214574 130170 214642 130226
rect 214698 130170 214768 130226
rect 214448 130102 214768 130170
rect 214448 130046 214518 130102
rect 214574 130046 214642 130102
rect 214698 130046 214768 130102
rect 214448 129978 214768 130046
rect 214448 129922 214518 129978
rect 214574 129922 214642 129978
rect 214698 129922 214768 129978
rect 214448 129888 214768 129922
rect 245168 130350 245488 130384
rect 245168 130294 245238 130350
rect 245294 130294 245362 130350
rect 245418 130294 245488 130350
rect 245168 130226 245488 130294
rect 245168 130170 245238 130226
rect 245294 130170 245362 130226
rect 245418 130170 245488 130226
rect 245168 130102 245488 130170
rect 245168 130046 245238 130102
rect 245294 130046 245362 130102
rect 245418 130046 245488 130102
rect 245168 129978 245488 130046
rect 245168 129922 245238 129978
rect 245294 129922 245362 129978
rect 245418 129922 245488 129978
rect 245168 129888 245488 129922
rect 275888 130350 276208 130384
rect 275888 130294 275958 130350
rect 276014 130294 276082 130350
rect 276138 130294 276208 130350
rect 275888 130226 276208 130294
rect 275888 130170 275958 130226
rect 276014 130170 276082 130226
rect 276138 130170 276208 130226
rect 275888 130102 276208 130170
rect 275888 130046 275958 130102
rect 276014 130046 276082 130102
rect 276138 130046 276208 130102
rect 275888 129978 276208 130046
rect 275888 129922 275958 129978
rect 276014 129922 276082 129978
rect 276138 129922 276208 129978
rect 275888 129888 276208 129922
rect 306608 130350 306928 130384
rect 306608 130294 306678 130350
rect 306734 130294 306802 130350
rect 306858 130294 306928 130350
rect 306608 130226 306928 130294
rect 306608 130170 306678 130226
rect 306734 130170 306802 130226
rect 306858 130170 306928 130226
rect 306608 130102 306928 130170
rect 306608 130046 306678 130102
rect 306734 130046 306802 130102
rect 306858 130046 306928 130102
rect 306608 129978 306928 130046
rect 306608 129922 306678 129978
rect 306734 129922 306802 129978
rect 306858 129922 306928 129978
rect 306608 129888 306928 129922
rect 337328 130350 337648 130384
rect 337328 130294 337398 130350
rect 337454 130294 337522 130350
rect 337578 130294 337648 130350
rect 337328 130226 337648 130294
rect 337328 130170 337398 130226
rect 337454 130170 337522 130226
rect 337578 130170 337648 130226
rect 337328 130102 337648 130170
rect 337328 130046 337398 130102
rect 337454 130046 337522 130102
rect 337578 130046 337648 130102
rect 337328 129978 337648 130046
rect 337328 129922 337398 129978
rect 337454 129922 337522 129978
rect 337578 129922 337648 129978
rect 337328 129888 337648 129922
rect 368048 130350 368368 130384
rect 368048 130294 368118 130350
rect 368174 130294 368242 130350
rect 368298 130294 368368 130350
rect 368048 130226 368368 130294
rect 368048 130170 368118 130226
rect 368174 130170 368242 130226
rect 368298 130170 368368 130226
rect 368048 130102 368368 130170
rect 368048 130046 368118 130102
rect 368174 130046 368242 130102
rect 368298 130046 368368 130102
rect 368048 129978 368368 130046
rect 368048 129922 368118 129978
rect 368174 129922 368242 129978
rect 368298 129922 368368 129978
rect 368048 129888 368368 129922
rect 209468 128370 209524 128380
rect 209244 122994 209300 123004
rect 229808 118350 230128 118384
rect 229808 118294 229878 118350
rect 229934 118294 230002 118350
rect 230058 118294 230128 118350
rect 229808 118226 230128 118294
rect 229808 118170 229878 118226
rect 229934 118170 230002 118226
rect 230058 118170 230128 118226
rect 229808 118102 230128 118170
rect 229808 118046 229878 118102
rect 229934 118046 230002 118102
rect 230058 118046 230128 118102
rect 229808 117978 230128 118046
rect 229808 117922 229878 117978
rect 229934 117922 230002 117978
rect 230058 117922 230128 117978
rect 229808 117888 230128 117922
rect 260528 118350 260848 118384
rect 260528 118294 260598 118350
rect 260654 118294 260722 118350
rect 260778 118294 260848 118350
rect 260528 118226 260848 118294
rect 260528 118170 260598 118226
rect 260654 118170 260722 118226
rect 260778 118170 260848 118226
rect 260528 118102 260848 118170
rect 260528 118046 260598 118102
rect 260654 118046 260722 118102
rect 260778 118046 260848 118102
rect 260528 117978 260848 118046
rect 260528 117922 260598 117978
rect 260654 117922 260722 117978
rect 260778 117922 260848 117978
rect 260528 117888 260848 117922
rect 291248 118350 291568 118384
rect 291248 118294 291318 118350
rect 291374 118294 291442 118350
rect 291498 118294 291568 118350
rect 291248 118226 291568 118294
rect 291248 118170 291318 118226
rect 291374 118170 291442 118226
rect 291498 118170 291568 118226
rect 291248 118102 291568 118170
rect 291248 118046 291318 118102
rect 291374 118046 291442 118102
rect 291498 118046 291568 118102
rect 291248 117978 291568 118046
rect 291248 117922 291318 117978
rect 291374 117922 291442 117978
rect 291498 117922 291568 117978
rect 291248 117888 291568 117922
rect 321968 118350 322288 118384
rect 321968 118294 322038 118350
rect 322094 118294 322162 118350
rect 322218 118294 322288 118350
rect 321968 118226 322288 118294
rect 321968 118170 322038 118226
rect 322094 118170 322162 118226
rect 322218 118170 322288 118226
rect 321968 118102 322288 118170
rect 321968 118046 322038 118102
rect 322094 118046 322162 118102
rect 322218 118046 322288 118102
rect 321968 117978 322288 118046
rect 321968 117922 322038 117978
rect 322094 117922 322162 117978
rect 322218 117922 322288 117978
rect 321968 117888 322288 117922
rect 352688 118350 353008 118384
rect 352688 118294 352758 118350
rect 352814 118294 352882 118350
rect 352938 118294 353008 118350
rect 352688 118226 353008 118294
rect 352688 118170 352758 118226
rect 352814 118170 352882 118226
rect 352938 118170 353008 118226
rect 352688 118102 353008 118170
rect 352688 118046 352758 118102
rect 352814 118046 352882 118102
rect 352938 118046 353008 118102
rect 352688 117978 353008 118046
rect 352688 117922 352758 117978
rect 352814 117922 352882 117978
rect 352938 117922 353008 117978
rect 352688 117888 353008 117922
rect 214448 112350 214768 112384
rect 214448 112294 214518 112350
rect 214574 112294 214642 112350
rect 214698 112294 214768 112350
rect 214448 112226 214768 112294
rect 214448 112170 214518 112226
rect 214574 112170 214642 112226
rect 214698 112170 214768 112226
rect 214448 112102 214768 112170
rect 214448 112046 214518 112102
rect 214574 112046 214642 112102
rect 214698 112046 214768 112102
rect 214448 111978 214768 112046
rect 214448 111922 214518 111978
rect 214574 111922 214642 111978
rect 214698 111922 214768 111978
rect 214448 111888 214768 111922
rect 245168 112350 245488 112384
rect 245168 112294 245238 112350
rect 245294 112294 245362 112350
rect 245418 112294 245488 112350
rect 245168 112226 245488 112294
rect 245168 112170 245238 112226
rect 245294 112170 245362 112226
rect 245418 112170 245488 112226
rect 245168 112102 245488 112170
rect 245168 112046 245238 112102
rect 245294 112046 245362 112102
rect 245418 112046 245488 112102
rect 245168 111978 245488 112046
rect 245168 111922 245238 111978
rect 245294 111922 245362 111978
rect 245418 111922 245488 111978
rect 245168 111888 245488 111922
rect 275888 112350 276208 112384
rect 275888 112294 275958 112350
rect 276014 112294 276082 112350
rect 276138 112294 276208 112350
rect 275888 112226 276208 112294
rect 275888 112170 275958 112226
rect 276014 112170 276082 112226
rect 276138 112170 276208 112226
rect 275888 112102 276208 112170
rect 275888 112046 275958 112102
rect 276014 112046 276082 112102
rect 276138 112046 276208 112102
rect 275888 111978 276208 112046
rect 275888 111922 275958 111978
rect 276014 111922 276082 111978
rect 276138 111922 276208 111978
rect 275888 111888 276208 111922
rect 306608 112350 306928 112384
rect 306608 112294 306678 112350
rect 306734 112294 306802 112350
rect 306858 112294 306928 112350
rect 306608 112226 306928 112294
rect 306608 112170 306678 112226
rect 306734 112170 306802 112226
rect 306858 112170 306928 112226
rect 306608 112102 306928 112170
rect 306608 112046 306678 112102
rect 306734 112046 306802 112102
rect 306858 112046 306928 112102
rect 306608 111978 306928 112046
rect 306608 111922 306678 111978
rect 306734 111922 306802 111978
rect 306858 111922 306928 111978
rect 306608 111888 306928 111922
rect 337328 112350 337648 112384
rect 337328 112294 337398 112350
rect 337454 112294 337522 112350
rect 337578 112294 337648 112350
rect 337328 112226 337648 112294
rect 337328 112170 337398 112226
rect 337454 112170 337522 112226
rect 337578 112170 337648 112226
rect 337328 112102 337648 112170
rect 337328 112046 337398 112102
rect 337454 112046 337522 112102
rect 337578 112046 337648 112102
rect 337328 111978 337648 112046
rect 337328 111922 337398 111978
rect 337454 111922 337522 111978
rect 337578 111922 337648 111978
rect 337328 111888 337648 111922
rect 368048 112350 368368 112384
rect 368048 112294 368118 112350
rect 368174 112294 368242 112350
rect 368298 112294 368368 112350
rect 368048 112226 368368 112294
rect 368048 112170 368118 112226
rect 368174 112170 368242 112226
rect 368298 112170 368368 112226
rect 368048 112102 368368 112170
rect 368048 112046 368118 112102
rect 368174 112046 368242 112102
rect 368298 112046 368368 112102
rect 368048 111978 368368 112046
rect 368048 111922 368118 111978
rect 368174 111922 368242 111978
rect 368298 111922 368368 111978
rect 368048 111888 368368 111922
rect 209132 104178 209188 104188
rect 229808 100350 230128 100384
rect 229808 100294 229878 100350
rect 229934 100294 230002 100350
rect 230058 100294 230128 100350
rect 229808 100226 230128 100294
rect 229808 100170 229878 100226
rect 229934 100170 230002 100226
rect 230058 100170 230128 100226
rect 229808 100102 230128 100170
rect 229808 100046 229878 100102
rect 229934 100046 230002 100102
rect 230058 100046 230128 100102
rect 229808 99978 230128 100046
rect 229808 99922 229878 99978
rect 229934 99922 230002 99978
rect 230058 99922 230128 99978
rect 229808 99888 230128 99922
rect 260528 100350 260848 100384
rect 260528 100294 260598 100350
rect 260654 100294 260722 100350
rect 260778 100294 260848 100350
rect 260528 100226 260848 100294
rect 260528 100170 260598 100226
rect 260654 100170 260722 100226
rect 260778 100170 260848 100226
rect 260528 100102 260848 100170
rect 260528 100046 260598 100102
rect 260654 100046 260722 100102
rect 260778 100046 260848 100102
rect 260528 99978 260848 100046
rect 260528 99922 260598 99978
rect 260654 99922 260722 99978
rect 260778 99922 260848 99978
rect 260528 99888 260848 99922
rect 291248 100350 291568 100384
rect 291248 100294 291318 100350
rect 291374 100294 291442 100350
rect 291498 100294 291568 100350
rect 291248 100226 291568 100294
rect 291248 100170 291318 100226
rect 291374 100170 291442 100226
rect 291498 100170 291568 100226
rect 291248 100102 291568 100170
rect 291248 100046 291318 100102
rect 291374 100046 291442 100102
rect 291498 100046 291568 100102
rect 291248 99978 291568 100046
rect 291248 99922 291318 99978
rect 291374 99922 291442 99978
rect 291498 99922 291568 99978
rect 291248 99888 291568 99922
rect 321968 100350 322288 100384
rect 321968 100294 322038 100350
rect 322094 100294 322162 100350
rect 322218 100294 322288 100350
rect 321968 100226 322288 100294
rect 321968 100170 322038 100226
rect 322094 100170 322162 100226
rect 322218 100170 322288 100226
rect 321968 100102 322288 100170
rect 321968 100046 322038 100102
rect 322094 100046 322162 100102
rect 322218 100046 322288 100102
rect 321968 99978 322288 100046
rect 321968 99922 322038 99978
rect 322094 99922 322162 99978
rect 322218 99922 322288 99978
rect 321968 99888 322288 99922
rect 352688 100350 353008 100384
rect 352688 100294 352758 100350
rect 352814 100294 352882 100350
rect 352938 100294 353008 100350
rect 352688 100226 353008 100294
rect 352688 100170 352758 100226
rect 352814 100170 352882 100226
rect 352938 100170 353008 100226
rect 352688 100102 353008 100170
rect 352688 100046 352758 100102
rect 352814 100046 352882 100102
rect 352938 100046 353008 100102
rect 352688 99978 353008 100046
rect 352688 99922 352758 99978
rect 352814 99922 352882 99978
rect 352938 99922 353008 99978
rect 352688 99888 353008 99922
rect 214448 94350 214768 94384
rect 214448 94294 214518 94350
rect 214574 94294 214642 94350
rect 214698 94294 214768 94350
rect 214448 94226 214768 94294
rect 214448 94170 214518 94226
rect 214574 94170 214642 94226
rect 214698 94170 214768 94226
rect 214448 94102 214768 94170
rect 214448 94046 214518 94102
rect 214574 94046 214642 94102
rect 214698 94046 214768 94102
rect 214448 93978 214768 94046
rect 214448 93922 214518 93978
rect 214574 93922 214642 93978
rect 214698 93922 214768 93978
rect 214448 93888 214768 93922
rect 245168 94350 245488 94384
rect 245168 94294 245238 94350
rect 245294 94294 245362 94350
rect 245418 94294 245488 94350
rect 245168 94226 245488 94294
rect 245168 94170 245238 94226
rect 245294 94170 245362 94226
rect 245418 94170 245488 94226
rect 245168 94102 245488 94170
rect 245168 94046 245238 94102
rect 245294 94046 245362 94102
rect 245418 94046 245488 94102
rect 245168 93978 245488 94046
rect 245168 93922 245238 93978
rect 245294 93922 245362 93978
rect 245418 93922 245488 93978
rect 245168 93888 245488 93922
rect 275888 94350 276208 94384
rect 275888 94294 275958 94350
rect 276014 94294 276082 94350
rect 276138 94294 276208 94350
rect 275888 94226 276208 94294
rect 275888 94170 275958 94226
rect 276014 94170 276082 94226
rect 276138 94170 276208 94226
rect 275888 94102 276208 94170
rect 275888 94046 275958 94102
rect 276014 94046 276082 94102
rect 276138 94046 276208 94102
rect 275888 93978 276208 94046
rect 275888 93922 275958 93978
rect 276014 93922 276082 93978
rect 276138 93922 276208 93978
rect 275888 93888 276208 93922
rect 306608 94350 306928 94384
rect 306608 94294 306678 94350
rect 306734 94294 306802 94350
rect 306858 94294 306928 94350
rect 306608 94226 306928 94294
rect 306608 94170 306678 94226
rect 306734 94170 306802 94226
rect 306858 94170 306928 94226
rect 306608 94102 306928 94170
rect 306608 94046 306678 94102
rect 306734 94046 306802 94102
rect 306858 94046 306928 94102
rect 306608 93978 306928 94046
rect 306608 93922 306678 93978
rect 306734 93922 306802 93978
rect 306858 93922 306928 93978
rect 306608 93888 306928 93922
rect 337328 94350 337648 94384
rect 337328 94294 337398 94350
rect 337454 94294 337522 94350
rect 337578 94294 337648 94350
rect 337328 94226 337648 94294
rect 337328 94170 337398 94226
rect 337454 94170 337522 94226
rect 337578 94170 337648 94226
rect 337328 94102 337648 94170
rect 337328 94046 337398 94102
rect 337454 94046 337522 94102
rect 337578 94046 337648 94102
rect 337328 93978 337648 94046
rect 337328 93922 337398 93978
rect 337454 93922 337522 93978
rect 337578 93922 337648 93978
rect 337328 93888 337648 93922
rect 368048 94350 368368 94384
rect 368048 94294 368118 94350
rect 368174 94294 368242 94350
rect 368298 94294 368368 94350
rect 368048 94226 368368 94294
rect 368048 94170 368118 94226
rect 368174 94170 368242 94226
rect 368298 94170 368368 94226
rect 368048 94102 368368 94170
rect 368048 94046 368118 94102
rect 368174 94046 368242 94102
rect 368298 94046 368368 94102
rect 368048 93978 368368 94046
rect 368048 93922 368118 93978
rect 368174 93922 368242 93978
rect 368298 93922 368368 93978
rect 368048 93888 368368 93922
rect 229808 82350 230128 82384
rect 229808 82294 229878 82350
rect 229934 82294 230002 82350
rect 230058 82294 230128 82350
rect 229808 82226 230128 82294
rect 229808 82170 229878 82226
rect 229934 82170 230002 82226
rect 230058 82170 230128 82226
rect 229808 82102 230128 82170
rect 229808 82046 229878 82102
rect 229934 82046 230002 82102
rect 230058 82046 230128 82102
rect 229808 81978 230128 82046
rect 229808 81922 229878 81978
rect 229934 81922 230002 81978
rect 230058 81922 230128 81978
rect 229808 81888 230128 81922
rect 260528 82350 260848 82384
rect 260528 82294 260598 82350
rect 260654 82294 260722 82350
rect 260778 82294 260848 82350
rect 260528 82226 260848 82294
rect 260528 82170 260598 82226
rect 260654 82170 260722 82226
rect 260778 82170 260848 82226
rect 260528 82102 260848 82170
rect 260528 82046 260598 82102
rect 260654 82046 260722 82102
rect 260778 82046 260848 82102
rect 260528 81978 260848 82046
rect 260528 81922 260598 81978
rect 260654 81922 260722 81978
rect 260778 81922 260848 81978
rect 260528 81888 260848 81922
rect 291248 82350 291568 82384
rect 291248 82294 291318 82350
rect 291374 82294 291442 82350
rect 291498 82294 291568 82350
rect 291248 82226 291568 82294
rect 291248 82170 291318 82226
rect 291374 82170 291442 82226
rect 291498 82170 291568 82226
rect 291248 82102 291568 82170
rect 291248 82046 291318 82102
rect 291374 82046 291442 82102
rect 291498 82046 291568 82102
rect 291248 81978 291568 82046
rect 291248 81922 291318 81978
rect 291374 81922 291442 81978
rect 291498 81922 291568 81978
rect 291248 81888 291568 81922
rect 321968 82350 322288 82384
rect 321968 82294 322038 82350
rect 322094 82294 322162 82350
rect 322218 82294 322288 82350
rect 321968 82226 322288 82294
rect 321968 82170 322038 82226
rect 322094 82170 322162 82226
rect 322218 82170 322288 82226
rect 321968 82102 322288 82170
rect 321968 82046 322038 82102
rect 322094 82046 322162 82102
rect 322218 82046 322288 82102
rect 321968 81978 322288 82046
rect 321968 81922 322038 81978
rect 322094 81922 322162 81978
rect 322218 81922 322288 81978
rect 321968 81888 322288 81922
rect 352688 82350 353008 82384
rect 352688 82294 352758 82350
rect 352814 82294 352882 82350
rect 352938 82294 353008 82350
rect 352688 82226 353008 82294
rect 352688 82170 352758 82226
rect 352814 82170 352882 82226
rect 352938 82170 353008 82226
rect 352688 82102 353008 82170
rect 352688 82046 352758 82102
rect 352814 82046 352882 82102
rect 352938 82046 353008 82102
rect 352688 81978 353008 82046
rect 352688 81922 352758 81978
rect 352814 81922 352882 81978
rect 352938 81922 353008 81978
rect 352688 81888 353008 81922
rect 370076 78708 370132 169148
rect 370188 88340 370244 176652
rect 370524 127652 370580 215180
rect 370748 209972 370804 209982
rect 370524 126028 370580 127596
rect 370188 88274 370244 88284
rect 370300 125972 370580 126028
rect 370636 170660 370692 170670
rect 370300 115444 370356 125972
rect 370076 78642 370132 78652
rect 214448 76350 214768 76384
rect 214448 76294 214518 76350
rect 214574 76294 214642 76350
rect 214698 76294 214768 76350
rect 214448 76226 214768 76294
rect 214448 76170 214518 76226
rect 214574 76170 214642 76226
rect 214698 76170 214768 76226
rect 214448 76102 214768 76170
rect 214448 76046 214518 76102
rect 214574 76046 214642 76102
rect 214698 76046 214768 76102
rect 214448 75978 214768 76046
rect 214448 75922 214518 75978
rect 214574 75922 214642 75978
rect 214698 75922 214768 75978
rect 214448 75888 214768 75922
rect 245168 76350 245488 76384
rect 245168 76294 245238 76350
rect 245294 76294 245362 76350
rect 245418 76294 245488 76350
rect 245168 76226 245488 76294
rect 245168 76170 245238 76226
rect 245294 76170 245362 76226
rect 245418 76170 245488 76226
rect 245168 76102 245488 76170
rect 245168 76046 245238 76102
rect 245294 76046 245362 76102
rect 245418 76046 245488 76102
rect 245168 75978 245488 76046
rect 245168 75922 245238 75978
rect 245294 75922 245362 75978
rect 245418 75922 245488 75978
rect 245168 75888 245488 75922
rect 275888 76350 276208 76384
rect 275888 76294 275958 76350
rect 276014 76294 276082 76350
rect 276138 76294 276208 76350
rect 275888 76226 276208 76294
rect 275888 76170 275958 76226
rect 276014 76170 276082 76226
rect 276138 76170 276208 76226
rect 275888 76102 276208 76170
rect 275888 76046 275958 76102
rect 276014 76046 276082 76102
rect 276138 76046 276208 76102
rect 275888 75978 276208 76046
rect 275888 75922 275958 75978
rect 276014 75922 276082 75978
rect 276138 75922 276208 75978
rect 275888 75888 276208 75922
rect 306608 76350 306928 76384
rect 306608 76294 306678 76350
rect 306734 76294 306802 76350
rect 306858 76294 306928 76350
rect 306608 76226 306928 76294
rect 306608 76170 306678 76226
rect 306734 76170 306802 76226
rect 306858 76170 306928 76226
rect 306608 76102 306928 76170
rect 306608 76046 306678 76102
rect 306734 76046 306802 76102
rect 306858 76046 306928 76102
rect 306608 75978 306928 76046
rect 306608 75922 306678 75978
rect 306734 75922 306802 75978
rect 306858 75922 306928 75978
rect 306608 75888 306928 75922
rect 337328 76350 337648 76384
rect 337328 76294 337398 76350
rect 337454 76294 337522 76350
rect 337578 76294 337648 76350
rect 337328 76226 337648 76294
rect 337328 76170 337398 76226
rect 337454 76170 337522 76226
rect 337578 76170 337648 76226
rect 337328 76102 337648 76170
rect 337328 76046 337398 76102
rect 337454 76046 337522 76102
rect 337578 76046 337648 76102
rect 337328 75978 337648 76046
rect 337328 75922 337398 75978
rect 337454 75922 337522 75978
rect 337578 75922 337648 75978
rect 337328 75888 337648 75922
rect 368048 76350 368368 76384
rect 368048 76294 368118 76350
rect 368174 76294 368242 76350
rect 368298 76294 368368 76350
rect 368048 76226 368368 76294
rect 368048 76170 368118 76226
rect 368174 76170 368242 76226
rect 368298 76170 368368 76226
rect 368048 76102 368368 76170
rect 368048 76046 368118 76102
rect 368174 76046 368242 76102
rect 368298 76046 368368 76102
rect 368048 75978 368368 76046
rect 368048 75922 368118 75978
rect 368174 75922 368242 75978
rect 368298 75922 368368 75978
rect 368048 75888 368368 75922
rect 370300 72660 370356 115388
rect 370636 99092 370692 170604
rect 370748 127204 370804 209916
rect 370860 205268 370916 270602
rect 370972 209098 371028 271292
rect 372540 269668 372596 269678
rect 372428 268212 372484 268222
rect 372092 258804 372148 258814
rect 370972 209032 371028 209042
rect 371084 248836 371140 248846
rect 370860 205202 370916 205212
rect 371084 183428 371140 248780
rect 371196 237860 371252 237870
rect 371196 234836 371252 237804
rect 371196 234770 371252 234780
rect 371756 231028 371812 231038
rect 371084 183362 371140 183372
rect 371196 229236 371252 229246
rect 370748 127138 370804 127148
rect 370860 182756 370916 182766
rect 370636 99026 370692 99036
rect 370860 95508 370916 182700
rect 371196 181412 371252 229180
rect 371644 228564 371700 228574
rect 371644 199220 371700 228508
rect 371644 199154 371700 199164
rect 371420 196084 371476 196094
rect 370860 95442 370916 95452
rect 371084 179396 371140 179406
rect 370300 72594 370356 72604
rect 370412 94164 370468 94174
rect 229808 64350 230128 64384
rect 229808 64294 229878 64350
rect 229934 64294 230002 64350
rect 230058 64294 230128 64350
rect 229808 64226 230128 64294
rect 229808 64170 229878 64226
rect 229934 64170 230002 64226
rect 230058 64170 230128 64226
rect 229808 64102 230128 64170
rect 229808 64046 229878 64102
rect 229934 64046 230002 64102
rect 230058 64046 230128 64102
rect 229808 63978 230128 64046
rect 229808 63922 229878 63978
rect 229934 63922 230002 63978
rect 230058 63922 230128 63978
rect 229808 63888 230128 63922
rect 260528 64350 260848 64384
rect 260528 64294 260598 64350
rect 260654 64294 260722 64350
rect 260778 64294 260848 64350
rect 260528 64226 260848 64294
rect 260528 64170 260598 64226
rect 260654 64170 260722 64226
rect 260778 64170 260848 64226
rect 260528 64102 260848 64170
rect 260528 64046 260598 64102
rect 260654 64046 260722 64102
rect 260778 64046 260848 64102
rect 260528 63978 260848 64046
rect 260528 63922 260598 63978
rect 260654 63922 260722 63978
rect 260778 63922 260848 63978
rect 260528 63888 260848 63922
rect 291248 64350 291568 64384
rect 291248 64294 291318 64350
rect 291374 64294 291442 64350
rect 291498 64294 291568 64350
rect 291248 64226 291568 64294
rect 291248 64170 291318 64226
rect 291374 64170 291442 64226
rect 291498 64170 291568 64226
rect 291248 64102 291568 64170
rect 291248 64046 291318 64102
rect 291374 64046 291442 64102
rect 291498 64046 291568 64102
rect 291248 63978 291568 64046
rect 291248 63922 291318 63978
rect 291374 63922 291442 63978
rect 291498 63922 291568 63978
rect 291248 63888 291568 63922
rect 321968 64350 322288 64384
rect 321968 64294 322038 64350
rect 322094 64294 322162 64350
rect 322218 64294 322288 64350
rect 321968 64226 322288 64294
rect 321968 64170 322038 64226
rect 322094 64170 322162 64226
rect 322218 64170 322288 64226
rect 321968 64102 322288 64170
rect 321968 64046 322038 64102
rect 322094 64046 322162 64102
rect 322218 64046 322288 64102
rect 321968 63978 322288 64046
rect 321968 63922 322038 63978
rect 322094 63922 322162 63978
rect 322218 63922 322288 63978
rect 321968 63888 322288 63922
rect 352688 64350 353008 64384
rect 352688 64294 352758 64350
rect 352814 64294 352882 64350
rect 352938 64294 353008 64350
rect 352688 64226 353008 64294
rect 352688 64170 352758 64226
rect 352814 64170 352882 64226
rect 352938 64170 353008 64226
rect 352688 64102 353008 64170
rect 352688 64046 352758 64102
rect 352814 64046 352882 64102
rect 352938 64046 353008 64102
rect 352688 63978 353008 64046
rect 352688 63922 352758 63978
rect 352814 63922 352882 63978
rect 352938 63922 353008 63978
rect 352688 63888 353008 63922
rect 214448 58350 214768 58384
rect 214448 58294 214518 58350
rect 214574 58294 214642 58350
rect 214698 58294 214768 58350
rect 214448 58226 214768 58294
rect 214448 58170 214518 58226
rect 214574 58170 214642 58226
rect 214698 58170 214768 58226
rect 214448 58102 214768 58170
rect 214448 58046 214518 58102
rect 214574 58046 214642 58102
rect 214698 58046 214768 58102
rect 214448 57978 214768 58046
rect 214448 57922 214518 57978
rect 214574 57922 214642 57978
rect 214698 57922 214768 57978
rect 214448 57888 214768 57922
rect 245168 58350 245488 58384
rect 245168 58294 245238 58350
rect 245294 58294 245362 58350
rect 245418 58294 245488 58350
rect 245168 58226 245488 58294
rect 245168 58170 245238 58226
rect 245294 58170 245362 58226
rect 245418 58170 245488 58226
rect 245168 58102 245488 58170
rect 245168 58046 245238 58102
rect 245294 58046 245362 58102
rect 245418 58046 245488 58102
rect 245168 57978 245488 58046
rect 245168 57922 245238 57978
rect 245294 57922 245362 57978
rect 245418 57922 245488 57978
rect 245168 57888 245488 57922
rect 275888 58350 276208 58384
rect 275888 58294 275958 58350
rect 276014 58294 276082 58350
rect 276138 58294 276208 58350
rect 275888 58226 276208 58294
rect 275888 58170 275958 58226
rect 276014 58170 276082 58226
rect 276138 58170 276208 58226
rect 275888 58102 276208 58170
rect 275888 58046 275958 58102
rect 276014 58046 276082 58102
rect 276138 58046 276208 58102
rect 275888 57978 276208 58046
rect 275888 57922 275958 57978
rect 276014 57922 276082 57978
rect 276138 57922 276208 57978
rect 275888 57888 276208 57922
rect 306608 58350 306928 58384
rect 306608 58294 306678 58350
rect 306734 58294 306802 58350
rect 306858 58294 306928 58350
rect 306608 58226 306928 58294
rect 306608 58170 306678 58226
rect 306734 58170 306802 58226
rect 306858 58170 306928 58226
rect 306608 58102 306928 58170
rect 306608 58046 306678 58102
rect 306734 58046 306802 58102
rect 306858 58046 306928 58102
rect 306608 57978 306928 58046
rect 306608 57922 306678 57978
rect 306734 57922 306802 57978
rect 306858 57922 306928 57978
rect 306608 57888 306928 57922
rect 337328 58350 337648 58384
rect 337328 58294 337398 58350
rect 337454 58294 337522 58350
rect 337578 58294 337648 58350
rect 337328 58226 337648 58294
rect 337328 58170 337398 58226
rect 337454 58170 337522 58226
rect 337578 58170 337648 58226
rect 337328 58102 337648 58170
rect 337328 58046 337398 58102
rect 337454 58046 337522 58102
rect 337578 58046 337648 58102
rect 337328 57978 337648 58046
rect 337328 57922 337398 57978
rect 337454 57922 337522 57978
rect 337578 57922 337648 57978
rect 337328 57888 337648 57922
rect 368048 58350 368368 58384
rect 368048 58294 368118 58350
rect 368174 58294 368242 58350
rect 368298 58294 368368 58350
rect 368048 58226 368368 58294
rect 368048 58170 368118 58226
rect 368174 58170 368242 58226
rect 368298 58170 368368 58226
rect 368048 58102 368368 58170
rect 368048 58046 368118 58102
rect 368174 58046 368242 58102
rect 368298 58046 368368 58102
rect 368048 57978 368368 58046
rect 368048 57922 368118 57978
rect 368174 57922 368242 57978
rect 368298 57922 368368 57978
rect 368048 57888 368368 57922
rect 209916 57876 209972 57886
rect 209916 56998 209972 57820
rect 209916 56932 209972 56942
rect 370412 56998 370468 94108
rect 370860 88340 370916 88350
rect 370860 87444 370916 88284
rect 370860 87378 370916 87388
rect 371084 86100 371140 179340
rect 371084 86034 371140 86044
rect 371196 85428 371252 181356
rect 371308 187124 371364 187134
rect 371308 163044 371364 187068
rect 371420 174692 371476 196028
rect 371420 174626 371476 174636
rect 371756 170660 371812 230972
rect 371980 222964 372036 222974
rect 371980 195748 372036 222908
rect 372092 219828 372148 258748
rect 372092 219762 372148 219772
rect 372204 236852 372260 236862
rect 371980 195682 372036 195692
rect 372092 199444 372148 199454
rect 371756 170594 371812 170604
rect 371868 173684 371924 173694
rect 371308 162978 371364 162988
rect 371868 123620 371924 173628
rect 371868 123554 371924 123564
rect 371980 163604 372036 163614
rect 371980 93492 372036 163548
rect 371980 93426 372036 93436
rect 371196 85362 371252 85372
rect 371308 86100 371364 86110
rect 208124 47730 208180 47740
rect 193458 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 194078 46350
rect 193458 46226 194078 46294
rect 193458 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 194078 46226
rect 193458 46102 194078 46170
rect 193458 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 194078 46102
rect 193458 45978 194078 46046
rect 193458 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 194078 45978
rect 193458 28350 194078 45922
rect 193458 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 194078 28350
rect 193458 28226 194078 28294
rect 193458 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 194078 28226
rect 193458 28102 194078 28170
rect 193458 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 194078 28102
rect 193458 27978 194078 28046
rect 193458 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 194078 27978
rect 193458 10350 194078 27922
rect 220458 40350 221078 56794
rect 220458 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 221078 40350
rect 220458 40226 221078 40294
rect 220458 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 221078 40226
rect 220458 40102 221078 40170
rect 220458 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 221078 40102
rect 220458 39978 221078 40046
rect 220458 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 221078 39978
rect 215140 22350 215460 22384
rect 215140 22294 215210 22350
rect 215266 22294 215334 22350
rect 215390 22294 215460 22350
rect 215140 22226 215460 22294
rect 215140 22170 215210 22226
rect 215266 22170 215334 22226
rect 215390 22170 215460 22226
rect 215140 22102 215460 22170
rect 215140 22046 215210 22102
rect 215266 22046 215334 22102
rect 215390 22046 215460 22102
rect 215140 21978 215460 22046
rect 215140 21922 215210 21978
rect 215266 21922 215334 21978
rect 215390 21922 215460 21978
rect 215140 21888 215460 21922
rect 220458 22350 221078 39922
rect 220458 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 221078 22350
rect 220458 22226 221078 22294
rect 220458 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 221078 22226
rect 220458 22102 221078 22170
rect 220458 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 221078 22102
rect 220458 21978 221078 22046
rect 220458 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 221078 21978
rect 193458 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 194078 10350
rect 193458 10226 194078 10294
rect 193458 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 194078 10226
rect 193458 10102 194078 10170
rect 193458 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 194078 10102
rect 193458 9978 194078 10046
rect 193458 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 194078 9978
rect 193458 -1120 194078 9922
rect 193458 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 194078 -1120
rect 193458 -1244 194078 -1176
rect 193458 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 194078 -1244
rect 193458 -1368 194078 -1300
rect 193458 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 194078 -1368
rect 193458 -1492 194078 -1424
rect 193458 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 194078 -1492
rect 193458 -1644 194078 -1548
rect 220458 4350 221078 21922
rect 220458 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 221078 4350
rect 220458 4226 221078 4294
rect 220458 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 221078 4226
rect 220458 4102 221078 4170
rect 220458 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 221078 4102
rect 220458 3978 221078 4046
rect 220458 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 221078 3978
rect 220458 -160 221078 3922
rect 220458 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 221078 -160
rect 220458 -284 221078 -216
rect 220458 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 221078 -284
rect 220458 -408 221078 -340
rect 220458 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 221078 -408
rect 220458 -532 221078 -464
rect 220458 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 221078 -532
rect 220458 -1644 221078 -588
rect 224178 46350 224798 56794
rect 224178 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 224798 46350
rect 224178 46226 224798 46294
rect 224178 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 224798 46226
rect 224178 46102 224798 46170
rect 224178 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 224798 46102
rect 224178 45978 224798 46046
rect 224178 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 224798 45978
rect 224178 28350 224798 45922
rect 224178 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 224798 28350
rect 224178 28226 224798 28294
rect 224178 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 224798 28226
rect 224178 28102 224798 28170
rect 224178 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 224798 28102
rect 224178 27978 224798 28046
rect 224178 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 224798 27978
rect 224178 10350 224798 27922
rect 224178 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 224798 10350
rect 224178 10226 224798 10294
rect 224178 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 224798 10226
rect 224178 10102 224798 10170
rect 224178 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 224798 10102
rect 224178 9978 224798 10046
rect 224178 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 224798 9978
rect 224178 -1120 224798 9922
rect 224178 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 224798 -1120
rect 224178 -1244 224798 -1176
rect 224178 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 224798 -1244
rect 224178 -1368 224798 -1300
rect 224178 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 224798 -1368
rect 224178 -1492 224798 -1424
rect 224178 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 224798 -1492
rect 224178 -1644 224798 -1548
rect 251178 40350 251798 56794
rect 251178 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 251798 40350
rect 251178 40226 251798 40294
rect 251178 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 251798 40226
rect 251178 40102 251798 40170
rect 251178 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 251798 40102
rect 251178 39978 251798 40046
rect 251178 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 251798 39978
rect 251178 22350 251798 39922
rect 251178 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 251798 22350
rect 251178 22226 251798 22294
rect 251178 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 251798 22226
rect 251178 22102 251798 22170
rect 251178 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 251798 22102
rect 251178 21978 251798 22046
rect 251178 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 251798 21978
rect 251178 4350 251798 21922
rect 251178 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 251798 4350
rect 251178 4226 251798 4294
rect 251178 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 251798 4226
rect 251178 4102 251798 4170
rect 251178 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 251798 4102
rect 251178 3978 251798 4046
rect 251178 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 251798 3978
rect 251178 -160 251798 3922
rect 251178 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 251798 -160
rect 251178 -284 251798 -216
rect 251178 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 251798 -284
rect 251178 -408 251798 -340
rect 251178 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 251798 -408
rect 251178 -532 251798 -464
rect 251178 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 251798 -532
rect 251178 -1644 251798 -588
rect 254898 46350 255518 56794
rect 254898 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 255518 46350
rect 254898 46226 255518 46294
rect 254898 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 255518 46226
rect 254898 46102 255518 46170
rect 254898 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 255518 46102
rect 254898 45978 255518 46046
rect 254898 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 255518 45978
rect 254898 28350 255518 45922
rect 281898 40350 282518 56794
rect 281898 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 282518 40350
rect 281898 40226 282518 40294
rect 281898 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 282518 40226
rect 281898 40102 282518 40170
rect 281898 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 282518 40102
rect 281898 39978 282518 40046
rect 281898 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 282518 39978
rect 254898 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 255518 28350
rect 254898 28226 255518 28294
rect 254898 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 255518 28226
rect 254898 28102 255518 28170
rect 254898 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 255518 28102
rect 254898 27978 255518 28046
rect 254898 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 255518 27978
rect 254898 10350 255518 27922
rect 279792 28350 280112 28384
rect 279792 28294 279862 28350
rect 279918 28294 279986 28350
rect 280042 28294 280112 28350
rect 279792 28226 280112 28294
rect 279792 28170 279862 28226
rect 279918 28170 279986 28226
rect 280042 28170 280112 28226
rect 279792 28102 280112 28170
rect 279792 28046 279862 28102
rect 279918 28046 279986 28102
rect 280042 28046 280112 28102
rect 279792 27978 280112 28046
rect 279792 27922 279862 27978
rect 279918 27922 279986 27978
rect 280042 27922 280112 27978
rect 279792 27888 280112 27922
rect 281898 22350 282518 39922
rect 281898 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 282518 22350
rect 281898 22226 282518 22294
rect 281898 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 282518 22226
rect 281898 22102 282518 22170
rect 281898 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 282518 22102
rect 281898 21978 282518 22046
rect 281898 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 282518 21978
rect 254898 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 255518 10350
rect 254898 10226 255518 10294
rect 254898 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 255518 10226
rect 254898 10102 255518 10170
rect 254898 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 255518 10102
rect 254898 9978 255518 10046
rect 254898 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 255518 9978
rect 254898 -1120 255518 9922
rect 279792 10350 280112 10384
rect 279792 10294 279862 10350
rect 279918 10294 279986 10350
rect 280042 10294 280112 10350
rect 279792 10226 280112 10294
rect 279792 10170 279862 10226
rect 279918 10170 279986 10226
rect 280042 10170 280112 10226
rect 279792 10102 280112 10170
rect 279792 10046 279862 10102
rect 279918 10046 279986 10102
rect 280042 10046 280112 10102
rect 279792 9978 280112 10046
rect 279792 9922 279862 9978
rect 279918 9922 279986 9978
rect 280042 9922 280112 9978
rect 279792 9888 280112 9922
rect 254898 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 255518 -1120
rect 254898 -1244 255518 -1176
rect 254898 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 255518 -1244
rect 254898 -1368 255518 -1300
rect 254898 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 255518 -1368
rect 254898 -1492 255518 -1424
rect 254898 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 255518 -1492
rect 254898 -1644 255518 -1548
rect 281898 4350 282518 21922
rect 281898 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 282518 4350
rect 281898 4226 282518 4294
rect 281898 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 282518 4226
rect 281898 4102 282518 4170
rect 281898 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 282518 4102
rect 281898 3978 282518 4046
rect 281898 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 282518 3978
rect 281898 -160 282518 3922
rect 281898 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 282518 -160
rect 281898 -284 282518 -216
rect 281898 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 282518 -284
rect 281898 -408 282518 -340
rect 281898 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 282518 -408
rect 281898 -532 282518 -464
rect 281898 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 282518 -532
rect 281898 -1644 282518 -588
rect 285618 46350 286238 56794
rect 285618 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 286238 46350
rect 285618 46226 286238 46294
rect 285618 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 286238 46226
rect 285618 46102 286238 46170
rect 285618 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 286238 46102
rect 285618 45978 286238 46046
rect 285618 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 286238 45978
rect 285618 28350 286238 45922
rect 285618 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 286238 28350
rect 285618 28226 286238 28294
rect 285618 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 286238 28226
rect 285618 28102 286238 28170
rect 285618 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 286238 28102
rect 285618 27978 286238 28046
rect 285618 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 286238 27978
rect 285618 10350 286238 27922
rect 285618 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 286238 10350
rect 285618 10226 286238 10294
rect 285618 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 286238 10226
rect 285618 10102 286238 10170
rect 285618 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 286238 10102
rect 285618 9978 286238 10046
rect 285618 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 286238 9978
rect 285618 -1120 286238 9922
rect 285618 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 286238 -1120
rect 285618 -1244 286238 -1176
rect 285618 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 286238 -1244
rect 285618 -1368 286238 -1300
rect 285618 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 286238 -1368
rect 285618 -1492 286238 -1424
rect 285618 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 286238 -1492
rect 285618 -1644 286238 -1548
rect 312618 40350 313238 56794
rect 312618 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 313238 40350
rect 312618 40226 313238 40294
rect 312618 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 313238 40226
rect 312618 40102 313238 40170
rect 312618 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 313238 40102
rect 312618 39978 313238 40046
rect 312618 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 313238 39978
rect 312618 22350 313238 39922
rect 312618 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 313238 22350
rect 312618 22226 313238 22294
rect 312618 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 313238 22226
rect 312618 22102 313238 22170
rect 312618 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 313238 22102
rect 312618 21978 313238 22046
rect 312618 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 313238 21978
rect 312618 4350 313238 21922
rect 312618 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 313238 4350
rect 312618 4226 313238 4294
rect 312618 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 313238 4226
rect 312618 4102 313238 4170
rect 312618 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 313238 4102
rect 312618 3978 313238 4046
rect 312618 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 313238 3978
rect 312618 -160 313238 3922
rect 312618 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 313238 -160
rect 312618 -284 313238 -216
rect 312618 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 313238 -284
rect 312618 -408 313238 -340
rect 312618 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 313238 -408
rect 312618 -532 313238 -464
rect 312618 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 313238 -532
rect 312618 -1644 313238 -588
rect 316338 46350 316958 56794
rect 316338 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 316958 46350
rect 316338 46226 316958 46294
rect 316338 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 316958 46226
rect 316338 46102 316958 46170
rect 316338 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 316958 46102
rect 316338 45978 316958 46046
rect 316338 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 316958 45978
rect 316338 28350 316958 45922
rect 316338 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 316958 28350
rect 316338 28226 316958 28294
rect 316338 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 316958 28226
rect 316338 28102 316958 28170
rect 316338 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 316958 28102
rect 316338 27978 316958 28046
rect 316338 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 316958 27978
rect 316338 10350 316958 27922
rect 316338 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 316958 10350
rect 316338 10226 316958 10294
rect 316338 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 316958 10226
rect 316338 10102 316958 10170
rect 316338 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 316958 10102
rect 316338 9978 316958 10046
rect 316338 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 316958 9978
rect 316338 -1120 316958 9922
rect 316338 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 316958 -1120
rect 316338 -1244 316958 -1176
rect 316338 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 316958 -1244
rect 316338 -1368 316958 -1300
rect 316338 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 316958 -1368
rect 316338 -1492 316958 -1424
rect 316338 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 316958 -1492
rect 316338 -1644 316958 -1548
rect 343338 40350 343958 56794
rect 343338 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 343958 40350
rect 343338 40226 343958 40294
rect 343338 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 343958 40226
rect 343338 40102 343958 40170
rect 343338 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 343958 40102
rect 343338 39978 343958 40046
rect 343338 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 343958 39978
rect 343338 22350 343958 39922
rect 347058 46350 347678 56794
rect 370412 51604 370468 56942
rect 371308 56084 371364 86044
rect 372092 83412 372148 199388
rect 372204 182756 372260 236796
rect 372204 182690 372260 182700
rect 372316 232596 372372 232606
rect 372316 176708 372372 232540
rect 372428 210898 372484 268156
rect 372540 232596 372596 269612
rect 372540 232530 372596 232540
rect 372652 229236 372708 275660
rect 372652 229170 372708 229180
rect 372764 268436 372820 268446
rect 372428 210832 372484 210842
rect 372540 218708 372596 218718
rect 372316 176642 372372 176652
rect 372428 177380 372484 177390
rect 372204 164724 372260 164734
rect 372204 92820 372260 164668
rect 372204 92754 372260 92764
rect 372316 134372 372372 134382
rect 372316 113204 372372 134316
rect 372092 83346 372148 83356
rect 372316 69972 372372 113148
rect 372316 69906 372372 69916
rect 372428 96180 372484 177324
rect 372540 134372 372596 218652
rect 372764 209278 372820 268380
rect 372876 217558 372932 293804
rect 373660 290164 373716 290174
rect 373324 284564 373380 284574
rect 373324 277060 373380 284508
rect 373324 276994 373380 277004
rect 373436 282324 373492 282334
rect 373436 275156 373492 282268
rect 373436 275090 373492 275100
rect 373548 276724 373604 276734
rect 373324 273364 373380 273374
rect 373324 266420 373380 273308
rect 373548 266756 373604 276668
rect 373660 275492 373716 290108
rect 373772 276948 373828 294588
rect 374058 292350 374678 309922
rect 375452 322868 375508 322878
rect 375452 309204 375508 322812
rect 375452 309138 375508 309148
rect 376012 316708 376068 316718
rect 374058 292294 374154 292350
rect 374210 292294 374278 292350
rect 374334 292294 374402 292350
rect 374458 292294 374526 292350
rect 374582 292294 374678 292350
rect 374058 292226 374678 292294
rect 374058 292170 374154 292226
rect 374210 292170 374278 292226
rect 374334 292170 374402 292226
rect 374458 292170 374526 292226
rect 374582 292170 374678 292226
rect 374058 292102 374678 292170
rect 374058 292046 374154 292102
rect 374210 292046 374278 292102
rect 374334 292046 374402 292102
rect 374458 292046 374526 292102
rect 374582 292046 374678 292102
rect 374058 291978 374678 292046
rect 374058 291922 374154 291978
rect 374210 291922 374278 291978
rect 374334 291922 374402 291978
rect 374458 291922 374526 291978
rect 374582 291922 374678 291978
rect 373772 276882 373828 276892
rect 373884 287924 373940 287934
rect 373660 275426 373716 275436
rect 373884 273700 373940 287868
rect 373884 273634 373940 273644
rect 374058 274350 374678 291922
rect 375452 293524 375508 293534
rect 374892 281204 374948 281214
rect 374780 280084 374836 280094
rect 374780 276612 374836 280028
rect 374780 276546 374836 276556
rect 374892 275380 374948 281148
rect 374892 275314 374948 275324
rect 375004 278964 375060 278974
rect 374058 274294 374154 274350
rect 374210 274294 374278 274350
rect 374334 274294 374402 274350
rect 374458 274294 374526 274350
rect 374582 274294 374678 274350
rect 374058 274226 374678 274294
rect 374058 274170 374154 274226
rect 374210 274170 374278 274226
rect 374334 274170 374402 274226
rect 374458 274170 374526 274226
rect 374582 274170 374678 274226
rect 374058 274102 374678 274170
rect 374058 274046 374154 274102
rect 374210 274046 374278 274102
rect 374334 274046 374402 274102
rect 374458 274046 374526 274102
rect 374582 274046 374678 274102
rect 374058 273978 374678 274046
rect 374058 273922 374154 273978
rect 374210 273922 374278 273978
rect 374334 273922 374402 273978
rect 374458 273922 374526 273978
rect 374582 273922 374678 273978
rect 373548 266690 373604 266700
rect 373324 266354 373380 266364
rect 373884 265188 373940 265198
rect 373436 263956 373492 263966
rect 373324 250964 373380 250974
rect 372988 249844 373044 249854
rect 372988 242004 373044 249788
rect 372988 241938 373044 241948
rect 373324 238644 373380 250908
rect 373436 246932 373492 263900
rect 373436 246866 373492 246876
rect 373660 263844 373716 263854
rect 373660 242788 373716 263788
rect 373772 262948 373828 262958
rect 373772 248836 373828 262892
rect 373884 261044 373940 265132
rect 373884 260978 373940 260988
rect 373772 248770 373828 248780
rect 374058 256350 374678 273922
rect 375004 273140 375060 278908
rect 375452 276836 375508 293468
rect 375676 291284 375732 291294
rect 375452 276770 375508 276780
rect 375564 283444 375620 283454
rect 375004 273074 375060 273084
rect 375116 275604 375172 275614
rect 374058 256294 374154 256350
rect 374210 256294 374278 256350
rect 374334 256294 374402 256350
rect 374458 256294 374526 256350
rect 374582 256294 374678 256350
rect 374058 256226 374678 256294
rect 374058 256170 374154 256226
rect 374210 256170 374278 256226
rect 374334 256170 374402 256226
rect 374458 256170 374526 256226
rect 374582 256170 374678 256226
rect 374058 256102 374678 256170
rect 374058 256046 374154 256102
rect 374210 256046 374278 256102
rect 374334 256046 374402 256102
rect 374458 256046 374526 256102
rect 374582 256046 374678 256102
rect 374058 255978 374678 256046
rect 374058 255922 374154 255978
rect 374210 255922 374278 255978
rect 374334 255922 374402 255978
rect 374458 255922 374526 255978
rect 374582 255922 374678 255978
rect 373660 242722 373716 242732
rect 373772 245364 373828 245374
rect 373772 242578 373828 245308
rect 373436 242522 373828 242578
rect 373884 244244 373940 244254
rect 373436 240884 373492 242522
rect 373884 242398 373940 244188
rect 373436 240818 373492 240828
rect 373660 242342 373940 242398
rect 373660 240598 373716 242342
rect 373884 242116 373940 242126
rect 373660 240542 373828 240598
rect 373660 240324 373716 240334
rect 373324 238578 373380 238588
rect 373548 238868 373604 238878
rect 373436 233492 373492 233502
rect 373436 231868 373492 233436
rect 372876 217492 372932 217502
rect 373324 231812 373492 231868
rect 373212 216580 373268 216590
rect 372764 209212 372820 209222
rect 373100 216244 373156 216254
rect 373100 200900 373156 216188
rect 373212 202468 373268 216524
rect 373324 215124 373380 231812
rect 373324 215058 373380 215068
rect 373436 229012 373492 229022
rect 373436 211652 373492 228956
rect 373548 215236 373604 238812
rect 373660 236852 373716 240268
rect 373660 235844 373716 236796
rect 373660 235778 373716 235788
rect 373772 234612 373828 240542
rect 373772 234546 373828 234556
rect 373884 233940 373940 242060
rect 373884 233874 373940 233884
rect 374058 238350 374678 255922
rect 374058 238294 374154 238350
rect 374210 238294 374278 238350
rect 374334 238294 374402 238350
rect 374458 238294 374526 238350
rect 374582 238294 374678 238350
rect 374058 238226 374678 238294
rect 374058 238170 374154 238226
rect 374210 238170 374278 238226
rect 374334 238170 374402 238226
rect 374458 238170 374526 238226
rect 374582 238170 374678 238226
rect 374058 238102 374678 238170
rect 374058 238046 374154 238102
rect 374210 238046 374278 238102
rect 374334 238046 374402 238102
rect 374458 238046 374526 238102
rect 374582 238046 374678 238102
rect 374058 237978 374678 238046
rect 374058 237922 374154 237978
rect 374210 237922 374278 237978
rect 374334 237922 374402 237978
rect 374458 237922 374526 237978
rect 374582 237922 374678 237978
rect 373548 215170 373604 215180
rect 373660 233044 373716 233054
rect 373660 214318 373716 232988
rect 373772 225092 373828 225102
rect 373772 216838 373828 225036
rect 374058 220350 374678 237922
rect 375004 270900 375060 270910
rect 374058 220294 374154 220350
rect 374210 220294 374278 220350
rect 374334 220294 374402 220350
rect 374458 220294 374526 220350
rect 374582 220294 374678 220350
rect 374058 220226 374678 220294
rect 374058 220170 374154 220226
rect 374210 220170 374278 220226
rect 374334 220170 374402 220226
rect 374458 220170 374526 220226
rect 374582 220170 374678 220226
rect 374058 220102 374678 220170
rect 374058 220046 374154 220102
rect 374210 220046 374278 220102
rect 374334 220046 374402 220102
rect 374458 220046 374526 220102
rect 374582 220046 374678 220102
rect 374058 219978 374678 220046
rect 374058 219922 374154 219978
rect 374210 219922 374278 219978
rect 374334 219922 374402 219978
rect 374458 219922 374526 219978
rect 374582 219922 374678 219978
rect 373884 218484 373940 218496
rect 373884 218392 373940 218402
rect 373772 216782 373940 216838
rect 373660 214252 373716 214262
rect 373772 216658 373828 216668
rect 373436 211586 373492 211596
rect 373212 202402 373268 202412
rect 373660 210644 373716 210654
rect 373548 201572 373604 201582
rect 373100 200834 373156 200844
rect 373324 201460 373380 201470
rect 373100 189028 373156 189038
rect 372764 184100 372820 184110
rect 372540 134306 372596 134316
rect 372652 173124 372708 173134
rect 372428 61684 372484 96124
rect 372540 116564 372596 116574
rect 372540 74676 372596 116508
rect 372652 85652 372708 173068
rect 372764 94108 372820 184044
rect 373100 182644 373156 188972
rect 373100 182578 373156 182588
rect 372876 182084 372932 182094
rect 372876 94500 372932 182028
rect 373324 179396 373380 201404
rect 373324 179330 373380 179340
rect 373436 187858 373492 187868
rect 373324 155428 373380 155438
rect 373324 128548 373380 155372
rect 373436 155204 373492 187802
rect 373548 174020 373604 201516
rect 373660 195972 373716 210588
rect 373660 195906 373716 195916
rect 373772 195418 373828 216602
rect 373884 214564 373940 216782
rect 373884 214498 373940 214508
rect 373884 214004 373940 214014
rect 373884 213418 373940 213948
rect 373884 213352 373940 213362
rect 373884 212884 373940 212894
rect 373884 211978 373940 212828
rect 373884 211912 373940 211922
rect 373884 211764 373940 211774
rect 373884 195860 373940 211708
rect 373884 195794 373940 195804
rect 374058 202350 374678 219922
rect 374058 202294 374154 202350
rect 374210 202294 374278 202350
rect 374334 202294 374402 202350
rect 374458 202294 374526 202350
rect 374582 202294 374678 202350
rect 374058 202226 374678 202294
rect 374058 202170 374154 202226
rect 374210 202170 374278 202226
rect 374334 202170 374402 202226
rect 374458 202170 374526 202226
rect 374582 202170 374678 202226
rect 374058 202102 374678 202170
rect 374058 202046 374154 202102
rect 374210 202046 374278 202102
rect 374334 202046 374402 202102
rect 374458 202046 374526 202102
rect 374582 202046 374678 202102
rect 374058 201978 374678 202046
rect 374058 201922 374154 201978
rect 374210 201922 374278 201978
rect 374334 201922 374402 201978
rect 374458 201922 374526 201978
rect 374582 201922 374678 201978
rect 373660 195362 373828 195418
rect 373660 194404 373716 195362
rect 373660 194338 373716 194348
rect 373772 194964 373828 194974
rect 373660 191828 373716 191838
rect 373660 183764 373716 191772
rect 373772 189364 373828 194908
rect 373772 189298 373828 189308
rect 373884 194740 373940 194750
rect 373884 188244 373940 194684
rect 373884 188178 373940 188188
rect 373884 186004 373940 186014
rect 373884 184978 373940 185948
rect 373884 184912 373940 184922
rect 373660 183698 373716 183708
rect 374058 184350 374678 201922
rect 374058 184294 374154 184350
rect 374210 184294 374278 184350
rect 374334 184294 374402 184350
rect 374458 184294 374526 184350
rect 374582 184294 374678 184350
rect 374058 184226 374678 184294
rect 374058 184170 374154 184226
rect 374210 184170 374278 184226
rect 374334 184170 374402 184226
rect 374458 184170 374526 184226
rect 374582 184170 374678 184226
rect 374058 184102 374678 184170
rect 374058 184046 374154 184102
rect 374210 184046 374278 184102
rect 374334 184046 374402 184102
rect 374458 184046 374526 184102
rect 374582 184046 374678 184102
rect 374058 183978 374678 184046
rect 374058 183922 374154 183978
rect 374210 183922 374278 183978
rect 374334 183922 374402 183978
rect 374458 183922 374526 183978
rect 374582 183922 374678 183978
rect 373884 183428 373940 183438
rect 373660 180404 373716 180414
rect 373660 176372 373716 180348
rect 373660 176306 373716 176316
rect 373772 179284 373828 179294
rect 373548 173124 373604 173964
rect 373548 173058 373604 173068
rect 373660 174916 373716 174926
rect 373436 155138 373492 155148
rect 373548 162484 373604 162494
rect 373324 128482 373380 128492
rect 373548 126868 373604 162428
rect 373660 133588 373716 174860
rect 373772 135828 373828 179228
rect 373772 135762 373828 135772
rect 373660 133522 373716 133532
rect 373548 126802 373604 126812
rect 373884 126028 373940 183372
rect 373772 125972 373940 126028
rect 374058 166350 374678 183922
rect 374892 226548 374948 226558
rect 374892 171332 374948 226492
rect 375004 213238 375060 270844
rect 375116 266532 375172 275548
rect 375564 275268 375620 283388
rect 375676 276724 375732 291228
rect 375676 276658 375732 276668
rect 375564 275202 375620 275212
rect 375788 274820 375844 274830
rect 375116 266466 375172 266476
rect 375228 274484 375284 274494
rect 375228 264628 375284 274428
rect 375228 264562 375284 264572
rect 375452 268858 375508 268868
rect 375004 213172 375060 213182
rect 375116 236404 375172 236414
rect 374892 169764 374948 171276
rect 375116 169988 375172 236348
rect 375452 233492 375508 268802
rect 375676 268548 375732 268558
rect 375452 233426 375508 233436
rect 375564 238756 375620 238766
rect 375340 231252 375396 231262
rect 375228 225204 375284 225214
rect 375228 206388 375284 225148
rect 375228 206322 375284 206332
rect 375228 188038 375284 188048
rect 375228 186564 375284 187982
rect 375228 186498 375284 186508
rect 375340 184100 375396 231196
rect 375452 213332 375508 213342
rect 375452 205044 375508 213276
rect 375452 204978 375508 204988
rect 375340 184034 375396 184044
rect 375452 198324 375508 198334
rect 375116 169922 375172 169932
rect 375340 172564 375396 172574
rect 374892 169698 374948 169708
rect 374058 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 374678 166350
rect 374058 166226 374678 166294
rect 374058 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 374678 166226
rect 374058 166102 374678 166170
rect 374058 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 374678 166102
rect 374058 165978 374678 166046
rect 374058 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 374678 165978
rect 374058 148350 374678 165922
rect 374058 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 374678 148350
rect 374058 148226 374678 148294
rect 374058 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 374678 148226
rect 374058 148102 374678 148170
rect 374058 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 374678 148102
rect 374058 147978 374678 148046
rect 374058 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 374678 147978
rect 374058 130350 374678 147922
rect 375340 133498 375396 172508
rect 375340 133432 375396 133442
rect 374058 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 374678 130350
rect 374058 130226 374678 130294
rect 374058 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 374678 130226
rect 374058 130102 374678 130170
rect 374058 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 374678 130102
rect 374058 129978 374678 130046
rect 374058 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 374678 129978
rect 373548 114996 373604 115006
rect 373548 114324 373604 114940
rect 372876 94434 372932 94444
rect 373100 99092 373156 99102
rect 373100 97524 373156 99036
rect 372988 94276 373044 94286
rect 372988 94108 373044 94220
rect 372764 94052 373044 94108
rect 372876 93828 372932 93838
rect 372876 87444 372932 93772
rect 372876 87378 372932 87388
rect 372652 85586 372708 85596
rect 372988 85204 373044 94052
rect 373100 89684 373156 97468
rect 373548 95732 373604 114268
rect 373548 95666 373604 95676
rect 373772 98196 373828 125972
rect 373884 120898 373940 120908
rect 373884 119924 373940 120842
rect 373884 119858 373940 119868
rect 373100 89618 373156 89628
rect 373772 86324 373828 98140
rect 373772 86258 373828 86268
rect 374058 112350 374678 129922
rect 374058 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 374678 112350
rect 374058 112226 374678 112294
rect 374058 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 374678 112226
rect 374058 112102 374678 112170
rect 374058 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 374678 112102
rect 374058 111978 374678 112046
rect 374058 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 374678 111978
rect 374058 94350 374678 111922
rect 374058 94294 374154 94350
rect 374210 94294 374278 94350
rect 374334 94294 374402 94350
rect 374458 94294 374526 94350
rect 374582 94294 374678 94350
rect 374058 94226 374678 94294
rect 374058 94170 374154 94226
rect 374210 94170 374278 94226
rect 374334 94170 374402 94226
rect 374458 94170 374526 94226
rect 374582 94170 374678 94226
rect 374058 94102 374678 94170
rect 374058 94046 374154 94102
rect 374210 94046 374278 94102
rect 374334 94046 374402 94102
rect 374458 94046 374526 94102
rect 374582 94046 374678 94102
rect 374058 93978 374678 94046
rect 374058 93922 374154 93978
rect 374210 93922 374278 93978
rect 374334 93922 374402 93978
rect 374458 93922 374526 93978
rect 374582 93922 374678 93978
rect 372988 85138 373044 85148
rect 372540 74610 372596 74620
rect 374058 76350 374678 93922
rect 375228 129332 375284 129342
rect 375228 90804 375284 129276
rect 375340 129220 375396 129230
rect 375340 112084 375396 129164
rect 375340 111076 375396 112028
rect 375340 111010 375396 111020
rect 375228 90738 375284 90748
rect 374058 76294 374154 76350
rect 374210 76294 374278 76350
rect 374334 76294 374402 76350
rect 374458 76294 374526 76350
rect 374582 76294 374678 76350
rect 374058 76226 374678 76294
rect 374058 76170 374154 76226
rect 374210 76170 374278 76226
rect 374334 76170 374402 76226
rect 374458 76170 374526 76226
rect 374582 76170 374678 76226
rect 374058 76102 374678 76170
rect 374058 76046 374154 76102
rect 374210 76046 374278 76102
rect 374334 76046 374402 76102
rect 374458 76046 374526 76102
rect 374582 76046 374678 76102
rect 374058 75978 374678 76046
rect 374058 75922 374154 75978
rect 374210 75922 374278 75978
rect 374334 75922 374402 75978
rect 374458 75922 374526 75978
rect 374582 75922 374678 75978
rect 372428 61618 372484 61628
rect 371308 56018 371364 56028
rect 374058 58350 374678 75922
rect 374058 58294 374154 58350
rect 374210 58294 374278 58350
rect 374334 58294 374402 58350
rect 374458 58294 374526 58350
rect 374582 58294 374678 58350
rect 374058 58226 374678 58294
rect 374058 58170 374154 58226
rect 374210 58170 374278 58226
rect 374334 58170 374402 58226
rect 374458 58170 374526 58226
rect 374582 58170 374678 58226
rect 374058 58102 374678 58170
rect 374058 58046 374154 58102
rect 374210 58046 374278 58102
rect 374334 58046 374402 58102
rect 374458 58046 374526 58102
rect 374582 58046 374678 58102
rect 374058 57978 374678 58046
rect 374058 57922 374154 57978
rect 374210 57922 374278 57978
rect 374334 57922 374402 57978
rect 374458 57922 374526 57978
rect 374582 57922 374678 57978
rect 370412 51538 370468 51548
rect 347058 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 347678 46350
rect 347058 46226 347678 46294
rect 347058 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 347678 46226
rect 347058 46102 347678 46170
rect 347058 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 347678 46102
rect 347058 45978 347678 46046
rect 347058 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 347678 45978
rect 347058 28350 347678 45922
rect 347058 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 347678 28350
rect 347058 28226 347678 28294
rect 347058 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 347678 28226
rect 347058 28102 347678 28170
rect 347058 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 347678 28102
rect 347058 27978 347678 28046
rect 347058 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 347678 27978
rect 343338 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 343958 22350
rect 343338 22226 343958 22294
rect 343338 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 343958 22226
rect 343338 22102 343958 22170
rect 343338 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 343958 22102
rect 343338 21978 343958 22046
rect 343338 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 343958 21978
rect 343338 4350 343958 21922
rect 344444 22350 344764 22384
rect 344444 22294 344514 22350
rect 344570 22294 344638 22350
rect 344694 22294 344764 22350
rect 344444 22226 344764 22294
rect 344444 22170 344514 22226
rect 344570 22170 344638 22226
rect 344694 22170 344764 22226
rect 344444 22102 344764 22170
rect 344444 22046 344514 22102
rect 344570 22046 344638 22102
rect 344694 22046 344764 22102
rect 344444 21978 344764 22046
rect 344444 21922 344514 21978
rect 344570 21922 344638 21978
rect 344694 21922 344764 21978
rect 344444 21888 344764 21922
rect 343338 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 343958 4350
rect 343338 4226 343958 4294
rect 343338 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 343958 4226
rect 343338 4102 343958 4170
rect 343338 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 343958 4102
rect 343338 3978 343958 4046
rect 343338 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 343958 3978
rect 343338 -160 343958 3922
rect 343338 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 343958 -160
rect 343338 -284 343958 -216
rect 343338 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 343958 -284
rect 343338 -408 343958 -340
rect 343338 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 343958 -408
rect 343338 -532 343958 -464
rect 343338 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 343958 -532
rect 343338 -1644 343958 -588
rect 347058 10350 347678 27922
rect 347058 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 347678 10350
rect 347058 10226 347678 10294
rect 347058 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 347678 10226
rect 347058 10102 347678 10170
rect 347058 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 347678 10102
rect 347058 9978 347678 10046
rect 347058 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 347678 9978
rect 347058 -1120 347678 9922
rect 347058 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 347678 -1120
rect 347058 -1244 347678 -1176
rect 347058 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 347678 -1244
rect 347058 -1368 347678 -1300
rect 347058 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 347678 -1368
rect 347058 -1492 347678 -1424
rect 347058 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 347678 -1492
rect 347058 -1644 347678 -1548
rect 374058 40350 374678 57922
rect 374780 87444 374836 87454
rect 374780 57204 374836 87388
rect 375452 81396 375508 198268
rect 375564 174692 375620 238700
rect 375676 212158 375732 268492
rect 375788 227220 375844 274764
rect 375788 227154 375844 227164
rect 376012 225316 376068 316652
rect 376012 225250 376068 225260
rect 376124 225204 376180 324716
rect 377468 316036 377524 316046
rect 376796 315364 376852 315374
rect 376236 303268 376292 303278
rect 376236 248052 376292 303212
rect 376460 301924 376516 301934
rect 376460 300244 376516 301868
rect 376460 300178 376516 300188
rect 376236 246932 376292 247996
rect 376460 252084 376516 252094
rect 376460 247380 376516 252028
rect 376460 247314 376516 247324
rect 376236 246866 376292 246876
rect 376460 246484 376516 246494
rect 376460 244692 376516 246428
rect 376460 244626 376516 244636
rect 376236 243124 376292 243134
rect 376236 235956 376292 243068
rect 376236 235890 376292 235900
rect 376124 225118 376180 225148
rect 375676 212092 375732 212102
rect 375788 225062 376180 225118
rect 375788 177380 375844 225062
rect 376124 224532 376180 224542
rect 376124 217018 376180 224476
rect 376796 224532 376852 315308
rect 377356 310660 377412 310670
rect 377244 302484 377300 302494
rect 377244 299908 377300 302428
rect 377244 299842 377300 299852
rect 377244 285124 377300 285134
rect 377132 260398 377188 260408
rect 377132 255892 377188 260342
rect 377132 255826 377188 255836
rect 377132 254324 377188 254334
rect 377132 229908 377188 254268
rect 377132 229842 377188 229852
rect 376796 224466 376852 224476
rect 377244 220108 377300 285068
rect 377356 221172 377412 310604
rect 377468 225988 377524 315980
rect 377580 315924 377636 324828
rect 377580 315858 377636 315868
rect 377778 316350 378398 333922
rect 387212 374724 387268 374734
rect 380268 327796 380324 327806
rect 379708 326004 379764 326014
rect 379036 323092 379092 323102
rect 377778 316294 377874 316350
rect 377930 316294 377998 316350
rect 378054 316294 378122 316350
rect 378178 316294 378246 316350
rect 378302 316294 378398 316350
rect 377778 316226 378398 316294
rect 377778 316170 377874 316226
rect 377930 316170 377998 316226
rect 378054 316170 378122 316226
rect 378178 316170 378246 316226
rect 378302 316170 378398 316226
rect 377778 316102 378398 316170
rect 377778 316046 377874 316102
rect 377930 316046 377998 316102
rect 378054 316046 378122 316102
rect 378178 316046 378246 316102
rect 378302 316046 378398 316102
rect 377778 315978 378398 316046
rect 377778 315922 377874 315978
rect 377930 315922 377998 315978
rect 378054 315922 378122 315978
rect 378178 315922 378246 315978
rect 378302 315922 378398 315978
rect 377778 298350 378398 315922
rect 378812 322980 378868 322990
rect 378812 311444 378868 322924
rect 379036 313684 379092 323036
rect 379036 313618 379092 313628
rect 378812 311378 378868 311388
rect 377778 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 378398 298350
rect 377778 298226 378398 298294
rect 377778 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 378398 298226
rect 377778 298102 378398 298170
rect 377778 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 378398 298102
rect 377778 297978 378398 298046
rect 377778 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 378398 297978
rect 377778 280350 378398 297922
rect 377778 280294 377874 280350
rect 377930 280294 377998 280350
rect 378054 280294 378122 280350
rect 378178 280294 378246 280350
rect 378302 280294 378398 280350
rect 377778 280226 378398 280294
rect 377778 280170 377874 280226
rect 377930 280170 377998 280226
rect 378054 280170 378122 280226
rect 378178 280170 378246 280226
rect 378302 280170 378398 280226
rect 377778 280102 378398 280170
rect 377778 280046 377874 280102
rect 377930 280046 377998 280102
rect 378054 280046 378122 280102
rect 378178 280046 378246 280102
rect 378302 280046 378398 280102
rect 377778 279978 378398 280046
rect 377778 279922 377874 279978
rect 377930 279922 377998 279978
rect 378054 279922 378122 279978
rect 378178 279922 378246 279978
rect 378302 279922 378398 279978
rect 377778 262350 378398 279922
rect 379372 291172 379428 291182
rect 377778 262294 377874 262350
rect 377930 262294 377998 262350
rect 378054 262294 378122 262350
rect 378178 262294 378246 262350
rect 378302 262294 378398 262350
rect 377778 262226 378398 262294
rect 377778 262170 377874 262226
rect 377930 262170 377998 262226
rect 378054 262170 378122 262226
rect 378178 262170 378246 262226
rect 378302 262170 378398 262226
rect 377778 262102 378398 262170
rect 377778 262046 377874 262102
rect 377930 262046 377998 262102
rect 378054 262046 378122 262102
rect 378178 262046 378246 262102
rect 378302 262046 378398 262102
rect 377778 261978 378398 262046
rect 377778 261922 377874 261978
rect 377930 261922 377998 261978
rect 378054 261922 378122 261978
rect 378178 261922 378246 261978
rect 378302 261922 378398 261978
rect 377580 261658 377636 261668
rect 377580 256116 377636 261602
rect 377580 256050 377636 256060
rect 377580 255892 377636 255902
rect 377580 250068 377636 255836
rect 377580 250002 377636 250012
rect 377778 244350 378398 261922
rect 377778 244294 377874 244350
rect 377930 244294 377998 244350
rect 378054 244294 378122 244350
rect 378178 244294 378246 244350
rect 378302 244294 378398 244350
rect 377778 244226 378398 244294
rect 377778 244170 377874 244226
rect 377930 244170 377998 244226
rect 378054 244170 378122 244226
rect 378178 244170 378246 244226
rect 378302 244170 378398 244226
rect 377778 244102 378398 244170
rect 377778 244046 377874 244102
rect 377930 244046 377998 244102
rect 378054 244046 378122 244102
rect 378178 244046 378246 244102
rect 378302 244046 378398 244102
rect 377778 243978 378398 244046
rect 377778 243922 377874 243978
rect 377930 243922 377998 243978
rect 378054 243922 378122 243978
rect 378178 243922 378246 243978
rect 378302 243922 378398 243978
rect 377468 225922 377524 225932
rect 377580 227220 377636 227230
rect 377356 221106 377412 221116
rect 377244 220052 377524 220108
rect 376124 216952 376180 216962
rect 375900 215796 375956 215806
rect 375900 178052 375956 215740
rect 375900 177986 375956 177996
rect 376124 213332 376180 213342
rect 375788 177314 375844 177324
rect 375564 174626 375620 174636
rect 375900 177044 375956 177054
rect 375452 81330 375508 81340
rect 375564 168084 375620 168094
rect 375564 76692 375620 168028
rect 375676 166964 375732 166974
rect 375676 88116 375732 166908
rect 375788 165844 375844 165854
rect 375788 92148 375844 165788
rect 375900 126980 375956 176988
rect 375900 126914 375956 126924
rect 376012 169764 376068 169774
rect 375788 92082 375844 92092
rect 375900 111076 375956 111086
rect 375676 88050 375732 88060
rect 375564 76626 375620 76636
rect 375900 69300 375956 111020
rect 376012 94836 376068 169708
rect 376124 130228 376180 213276
rect 377468 203028 377524 220052
rect 377468 202356 377524 202972
rect 377468 202290 377524 202300
rect 377468 201684 377524 201694
rect 377468 178724 377524 201628
rect 377468 178658 377524 178668
rect 376124 129220 376180 130172
rect 376124 129154 376180 129164
rect 376236 178052 376292 178062
rect 376124 105778 376180 105788
rect 376124 104244 376180 105722
rect 376124 104178 376180 104188
rect 376012 88564 376068 94780
rect 376124 91558 376180 91568
rect 376124 90804 376180 91502
rect 376124 90738 376180 90748
rect 376012 88498 376068 88508
rect 376236 76020 376292 177996
rect 377468 176036 377524 176046
rect 377356 156358 377412 156368
rect 376348 152740 376404 152750
rect 376348 151844 376404 152684
rect 376348 142324 376404 151788
rect 377132 152740 377188 152750
rect 377132 152404 377188 152684
rect 377132 145796 377188 152348
rect 377132 145730 377188 145740
rect 377244 151172 377300 151182
rect 377244 143444 377300 151116
rect 377244 143378 377300 143388
rect 376348 142258 376404 142268
rect 377356 134820 377412 156302
rect 377356 134596 377412 134764
rect 377356 134530 377412 134540
rect 376908 133678 376964 133688
rect 376908 132692 376964 133622
rect 376908 132626 376964 132636
rect 377468 114268 377524 175980
rect 377356 114212 377524 114268
rect 377580 175364 377636 227164
rect 376236 75718 376292 75964
rect 376460 87220 376516 87230
rect 376236 75662 376404 75718
rect 375900 69234 375956 69244
rect 374780 57138 374836 57148
rect 376348 54964 376404 75662
rect 376460 72212 376516 87164
rect 377356 84756 377412 114212
rect 377580 102508 377636 175308
rect 377468 102452 377636 102508
rect 377778 226350 378398 243922
rect 378812 267238 378868 267248
rect 378588 242676 378644 242686
rect 377778 226294 377874 226350
rect 377930 226294 377998 226350
rect 378054 226294 378122 226350
rect 378178 226294 378246 226350
rect 378302 226294 378398 226350
rect 377778 226226 378398 226294
rect 377778 226170 377874 226226
rect 377930 226170 377998 226226
rect 378054 226170 378122 226226
rect 378178 226170 378246 226226
rect 378302 226170 378398 226226
rect 377778 226102 378398 226170
rect 377778 226046 377874 226102
rect 377930 226046 377998 226102
rect 378054 226046 378122 226102
rect 378178 226046 378246 226102
rect 378302 226046 378398 226102
rect 377778 225978 378398 226046
rect 377778 225922 377874 225978
rect 377930 225922 377998 225978
rect 378054 225922 378122 225978
rect 378178 225922 378246 225978
rect 378302 225922 378398 225978
rect 377778 208350 378398 225922
rect 377778 208294 377874 208350
rect 377930 208294 377998 208350
rect 378054 208294 378122 208350
rect 378178 208294 378246 208350
rect 378302 208294 378398 208350
rect 377778 208226 378398 208294
rect 377778 208170 377874 208226
rect 377930 208170 377998 208226
rect 378054 208170 378122 208226
rect 378178 208170 378246 208226
rect 378302 208170 378398 208226
rect 377778 208102 378398 208170
rect 377778 208046 377874 208102
rect 377930 208046 377998 208102
rect 378054 208046 378122 208102
rect 378178 208046 378246 208102
rect 378302 208046 378398 208102
rect 377778 207978 378398 208046
rect 377778 207922 377874 207978
rect 377930 207922 377998 207978
rect 378054 207922 378122 207978
rect 378178 207922 378246 207978
rect 378302 207922 378398 207978
rect 377778 190350 378398 207922
rect 378476 229348 378532 229358
rect 378476 202580 378532 229292
rect 378476 202514 378532 202524
rect 377778 190294 377874 190350
rect 377930 190294 377998 190350
rect 378054 190294 378122 190350
rect 378178 190294 378246 190350
rect 378302 190294 378398 190350
rect 377778 190226 378398 190294
rect 377778 190170 377874 190226
rect 377930 190170 377998 190226
rect 378054 190170 378122 190226
rect 378178 190170 378246 190226
rect 378302 190170 378398 190226
rect 377778 190102 378398 190170
rect 377778 190046 377874 190102
rect 377930 190046 377998 190102
rect 378054 190046 378122 190102
rect 378178 190046 378246 190102
rect 378302 190046 378398 190102
rect 377778 189978 378398 190046
rect 377778 189922 377874 189978
rect 377930 189922 377998 189978
rect 378054 189922 378122 189978
rect 378178 189922 378246 189978
rect 378302 189922 378398 189978
rect 377778 172350 378398 189922
rect 377778 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 378398 172350
rect 377778 172226 378398 172294
rect 377778 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 378398 172226
rect 377778 172102 378398 172170
rect 377778 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 378398 172102
rect 377778 171978 378398 172046
rect 377778 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 378398 171978
rect 377778 154350 378398 171922
rect 377778 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 378398 154350
rect 377778 154226 378398 154294
rect 377778 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 378398 154226
rect 377778 154102 378398 154170
rect 377778 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 378398 154102
rect 377778 153978 378398 154046
rect 377778 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 378398 153978
rect 377778 136350 378398 153922
rect 377778 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 378398 136350
rect 377778 136226 378398 136294
rect 377778 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 378398 136226
rect 377778 136102 378398 136170
rect 377778 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 378398 136102
rect 377778 135978 378398 136046
rect 377778 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 378398 135978
rect 377778 118350 378398 135922
rect 378588 131796 378644 242620
rect 378700 219604 378756 219614
rect 378700 214138 378756 219548
rect 378700 214072 378756 214082
rect 378812 159572 378868 267182
rect 379260 264964 379316 264974
rect 379148 264852 379204 264862
rect 378924 237748 378980 237758
rect 378924 211078 378980 237692
rect 379148 231028 379204 264796
rect 379148 230962 379204 230972
rect 379260 226548 379316 264908
rect 379260 226482 379316 226492
rect 379260 215578 379316 215588
rect 379260 215484 379316 215516
rect 378924 211012 378980 211022
rect 379372 206276 379428 291116
rect 379484 264538 379540 264548
rect 379484 237860 379540 264482
rect 379484 237794 379540 237804
rect 379596 261298 379652 261308
rect 379484 217198 379540 217208
rect 379484 217140 379540 217142
rect 379484 217074 379540 217084
rect 379484 216478 379540 216488
rect 379484 215796 379540 216422
rect 379484 215730 379540 215740
rect 379484 215460 379540 215470
rect 379484 215398 379540 215404
rect 379484 215332 379540 215342
rect 379372 206210 379428 206220
rect 378812 159506 378868 159516
rect 378924 194628 378980 194638
rect 378588 131730 378644 131740
rect 378700 154532 378756 154542
rect 377778 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 378398 118350
rect 377778 118226 378398 118294
rect 377778 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 378398 118226
rect 377778 118102 378398 118170
rect 377778 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 378398 118102
rect 377778 117978 378398 118046
rect 377778 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 378398 117978
rect 377468 96598 377524 102452
rect 377580 102004 377636 102014
rect 377580 101638 377636 101948
rect 377580 101572 377636 101582
rect 377778 100350 378398 117922
rect 377778 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 378398 100350
rect 377778 100226 378398 100294
rect 377778 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 378398 100226
rect 377778 100102 378398 100170
rect 377778 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 378398 100102
rect 377778 99978 378398 100046
rect 377778 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 378398 99978
rect 377468 96542 377636 96598
rect 377356 84690 377412 84700
rect 377580 79380 377636 96542
rect 377580 78988 377636 79324
rect 376460 72146 376516 72156
rect 377132 78932 377636 78988
rect 377778 82350 378398 99922
rect 377778 82294 377874 82350
rect 377930 82294 377998 82350
rect 378054 82294 378122 82350
rect 378178 82294 378246 82350
rect 378302 82294 378398 82350
rect 377778 82226 378398 82294
rect 377778 82170 377874 82226
rect 377930 82170 377998 82226
rect 378054 82170 378122 82226
rect 378178 82170 378246 82226
rect 378302 82170 378398 82226
rect 377778 82102 378398 82170
rect 377778 82046 377874 82102
rect 377930 82046 377998 82102
rect 378054 82046 378122 82102
rect 378178 82046 378246 82102
rect 378302 82046 378398 82102
rect 377778 81978 378398 82046
rect 377778 81922 377874 81978
rect 377930 81922 377998 81978
rect 378054 81922 378122 81978
rect 378178 81922 378246 81978
rect 378302 81922 378398 81978
rect 376348 54898 376404 54908
rect 377132 53844 377188 78932
rect 377580 71764 377636 71774
rect 377580 71398 377636 71708
rect 377580 71332 377636 71342
rect 377580 65044 377636 65054
rect 377580 64918 377636 64988
rect 377580 64852 377636 64862
rect 377580 64738 377636 64748
rect 377580 63924 377636 64682
rect 377580 63858 377636 63868
rect 377778 64350 378398 81922
rect 378588 74278 378644 74288
rect 378588 74116 378644 74222
rect 378588 74050 378644 74060
rect 377778 64294 377874 64350
rect 377930 64294 377998 64350
rect 378054 64294 378122 64350
rect 378178 64294 378246 64350
rect 378302 64294 378398 64350
rect 377778 64226 378398 64294
rect 377778 64170 377874 64226
rect 377930 64170 377998 64226
rect 378054 64170 378122 64226
rect 378178 64170 378246 64226
rect 378302 64170 378398 64226
rect 377778 64102 378398 64170
rect 377778 64046 377874 64102
rect 377930 64046 377998 64102
rect 378054 64046 378122 64102
rect 378178 64046 378246 64102
rect 378302 64046 378398 64102
rect 377778 63978 378398 64046
rect 377778 63922 377874 63978
rect 377930 63922 377998 63978
rect 378054 63922 378122 63978
rect 378178 63922 378246 63978
rect 378302 63922 378398 63978
rect 377580 62938 377636 62948
rect 377580 62804 377636 62882
rect 377580 62738 377636 62748
rect 377132 53778 377188 53788
rect 376236 52164 376292 52176
rect 376236 52072 376292 52082
rect 374058 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 374678 40350
rect 374058 40226 374678 40294
rect 374058 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 374678 40226
rect 374058 40102 374678 40170
rect 374058 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 374678 40102
rect 374058 39978 374678 40046
rect 374058 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 374678 39978
rect 374058 22350 374678 39922
rect 374058 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 374678 22350
rect 374058 22226 374678 22294
rect 374058 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 374678 22226
rect 374058 22102 374678 22170
rect 374058 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 374678 22102
rect 374058 21978 374678 22046
rect 374058 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 374678 21978
rect 374058 4350 374678 21922
rect 374058 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 374678 4350
rect 374058 4226 374678 4294
rect 374058 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 374678 4226
rect 374058 4102 374678 4170
rect 374058 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 374678 4102
rect 374058 3978 374678 4046
rect 374058 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 374678 3978
rect 374058 -160 374678 3922
rect 374058 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 374678 -160
rect 374058 -284 374678 -216
rect 374058 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 374678 -284
rect 374058 -408 374678 -340
rect 374058 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 374678 -408
rect 374058 -532 374678 -464
rect 374058 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 374678 -532
rect 374058 -1644 374678 -588
rect 377778 46350 378398 63922
rect 377778 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 378398 46350
rect 377778 46226 378398 46294
rect 377778 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 378398 46226
rect 377778 46102 378398 46170
rect 377778 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 378398 46102
rect 377778 45978 378398 46046
rect 377778 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 378398 45978
rect 377778 28350 378398 45922
rect 378700 42868 378756 154476
rect 378924 152740 378980 194572
rect 379148 192612 379204 192622
rect 378924 152674 378980 152684
rect 379036 155764 379092 155774
rect 378812 142324 378868 142334
rect 378812 90748 378868 142268
rect 379036 137396 379092 155708
rect 379148 151284 379204 192556
rect 379148 148484 379204 151228
rect 379372 182278 379428 182288
rect 379372 151172 379428 182222
rect 379596 159908 379652 261242
rect 379708 221732 379764 325948
rect 379932 268138 379988 268148
rect 379708 221666 379764 221676
rect 379820 267958 379876 267968
rect 379708 217924 379764 217934
rect 379708 217738 379764 217868
rect 379708 217672 379764 217682
rect 379708 217364 379764 217374
rect 379708 212518 379764 217308
rect 379708 212452 379764 212462
rect 379708 209188 379764 209198
rect 379708 182084 379764 209132
rect 379708 182018 379764 182028
rect 379820 162596 379876 267902
rect 379932 249620 379988 268082
rect 380156 267652 380212 267662
rect 379932 249554 379988 249564
rect 380044 266644 380100 266654
rect 380044 249418 380100 266588
rect 379932 249362 380100 249418
rect 379932 238588 379988 249362
rect 380044 241858 380100 241868
rect 380044 241780 380100 241802
rect 380044 241714 380100 241724
rect 379932 238532 380100 238588
rect 379820 162530 379876 162540
rect 379932 236964 379988 236974
rect 379596 159842 379652 159852
rect 379820 156548 379876 156558
rect 379372 151106 379428 151116
rect 379596 152852 379652 152862
rect 379596 151138 379652 152796
rect 379596 151072 379652 151082
rect 379372 150500 379428 150510
rect 379148 148418 379204 148428
rect 379260 149156 379316 149166
rect 379036 137330 379092 137340
rect 379260 133700 379316 149100
rect 379260 133634 379316 133644
rect 378812 90692 378980 90748
rect 378812 81844 378868 81854
rect 378812 81658 378868 81788
rect 378812 81592 378868 81602
rect 378812 80836 378868 80846
rect 378812 80758 378868 80780
rect 378812 80692 378868 80702
rect 378812 80578 378868 80588
rect 378812 79604 378868 80522
rect 378812 79538 378868 79548
rect 378812 78484 378868 78494
rect 378812 78418 378868 78428
rect 378812 78352 378868 78362
rect 378812 78058 378868 78068
rect 378812 77364 378868 78002
rect 378812 77298 378868 77308
rect 378812 72884 378868 72894
rect 378812 72772 378868 72782
rect 378924 55468 378980 90692
rect 378812 55412 378980 55468
rect 378812 45556 378868 55412
rect 379372 47908 379428 150444
rect 379596 148484 379652 148494
rect 379596 137060 379652 148428
rect 379596 136994 379652 137004
rect 379708 143444 379764 143454
rect 379596 116340 379652 116350
rect 379596 115858 379652 116284
rect 379596 102508 379652 115802
rect 379484 102452 379652 102508
rect 379484 77364 379540 102452
rect 379484 77298 379540 77308
rect 379596 76618 379652 76628
rect 379596 76244 379652 76562
rect 379596 76178 379652 76188
rect 379596 75124 379652 75134
rect 379596 74098 379652 75068
rect 379596 74032 379652 74042
rect 379372 47842 379428 47852
rect 378812 45490 378868 45500
rect 379708 43678 379764 143388
rect 379708 43612 379764 43622
rect 378700 42802 378756 42812
rect 379820 40292 379876 156492
rect 379932 132356 379988 236908
rect 380044 159236 380100 238532
rect 380156 161924 380212 267596
rect 380268 223188 380324 327740
rect 380268 215218 380324 223132
rect 380380 324548 380436 324558
rect 380380 228564 380436 324492
rect 384448 310350 384768 310384
rect 384448 310294 384518 310350
rect 384574 310294 384642 310350
rect 384698 310294 384768 310350
rect 384448 310226 384768 310294
rect 384448 310170 384518 310226
rect 384574 310170 384642 310226
rect 384698 310170 384768 310226
rect 384448 310102 384768 310170
rect 384448 310046 384518 310102
rect 384574 310046 384642 310102
rect 384698 310046 384768 310102
rect 384448 309978 384768 310046
rect 384448 309922 384518 309978
rect 384574 309922 384642 309978
rect 384698 309922 384768 309978
rect 384448 309888 384768 309922
rect 384448 292350 384768 292384
rect 384448 292294 384518 292350
rect 384574 292294 384642 292350
rect 384698 292294 384768 292350
rect 384448 292226 384768 292294
rect 384448 292170 384518 292226
rect 384574 292170 384642 292226
rect 384698 292170 384768 292226
rect 384448 292102 384768 292170
rect 384448 292046 384518 292102
rect 384574 292046 384642 292102
rect 384698 292046 384768 292102
rect 384448 291978 384768 292046
rect 384448 291922 384518 291978
rect 384574 291922 384642 291978
rect 384698 291922 384768 291978
rect 384448 291888 384768 291922
rect 380380 216838 380436 228508
rect 380380 216772 380436 216782
rect 380492 289156 380548 289166
rect 380268 215152 380324 215162
rect 380380 216478 380436 216544
rect 380268 213668 380324 213678
rect 380268 213598 380324 213612
rect 380268 213532 380324 213542
rect 380268 213220 380324 213230
rect 380268 211798 380324 213164
rect 380268 211732 380324 211742
rect 380268 209278 380324 209288
rect 380268 205828 380324 209222
rect 380380 209188 380436 216412
rect 380380 209122 380436 209132
rect 380268 203924 380324 205772
rect 380492 204148 380548 289100
rect 380604 286138 380660 286142
rect 380716 286138 380772 286148
rect 380604 286132 380716 286138
rect 380660 286082 380716 286132
rect 380604 286066 380660 286076
rect 380716 286072 380772 286082
rect 385420 272132 385476 272142
rect 383852 272020 383908 272030
rect 381500 268100 381556 268110
rect 380604 263732 380660 263742
rect 380604 231868 380660 263676
rect 381500 241858 381556 268044
rect 383852 260398 383908 271964
rect 385420 270658 385476 272076
rect 387212 272132 387268 374668
rect 404778 364350 405398 381922
rect 404778 364294 404874 364350
rect 404930 364294 404998 364350
rect 405054 364294 405122 364350
rect 405178 364294 405246 364350
rect 405302 364294 405398 364350
rect 404778 364226 405398 364294
rect 404778 364170 404874 364226
rect 404930 364170 404998 364226
rect 405054 364170 405122 364226
rect 405178 364170 405246 364226
rect 405302 364170 405398 364226
rect 404778 364102 405398 364170
rect 404778 364046 404874 364102
rect 404930 364046 404998 364102
rect 405054 364046 405122 364102
rect 405178 364046 405246 364102
rect 405302 364046 405398 364102
rect 404778 363978 405398 364046
rect 404778 363922 404874 363978
rect 404930 363922 404998 363978
rect 405054 363922 405122 363978
rect 405178 363922 405246 363978
rect 405302 363922 405398 363978
rect 404778 346350 405398 363922
rect 404778 346294 404874 346350
rect 404930 346294 404998 346350
rect 405054 346294 405122 346350
rect 405178 346294 405246 346350
rect 405302 346294 405398 346350
rect 404778 346226 405398 346294
rect 404778 346170 404874 346226
rect 404930 346170 404998 346226
rect 405054 346170 405122 346226
rect 405178 346170 405246 346226
rect 405302 346170 405398 346226
rect 404778 346102 405398 346170
rect 404778 346046 404874 346102
rect 404930 346046 404998 346102
rect 405054 346046 405122 346102
rect 405178 346046 405246 346102
rect 405302 346046 405398 346102
rect 404778 345978 405398 346046
rect 404778 345922 404874 345978
rect 404930 345922 404998 345978
rect 405054 345922 405122 345978
rect 405178 345922 405246 345978
rect 405302 345922 405398 345978
rect 404778 328350 405398 345922
rect 404778 328294 404874 328350
rect 404930 328294 404998 328350
rect 405054 328294 405122 328350
rect 405178 328294 405246 328350
rect 405302 328294 405398 328350
rect 404778 328226 405398 328294
rect 404778 328170 404874 328226
rect 404930 328170 404998 328226
rect 405054 328170 405122 328226
rect 405178 328170 405246 328226
rect 405302 328170 405398 328226
rect 404778 328102 405398 328170
rect 404778 328046 404874 328102
rect 404930 328046 404998 328102
rect 405054 328046 405122 328102
rect 405178 328046 405246 328102
rect 405302 328046 405398 328102
rect 404778 327978 405398 328046
rect 404778 327922 404874 327978
rect 404930 327922 404998 327978
rect 405054 327922 405122 327978
rect 405178 327922 405246 327978
rect 405302 327922 405398 327978
rect 399808 316350 400128 316384
rect 399808 316294 399878 316350
rect 399934 316294 400002 316350
rect 400058 316294 400128 316350
rect 399808 316226 400128 316294
rect 399808 316170 399878 316226
rect 399934 316170 400002 316226
rect 400058 316170 400128 316226
rect 399808 316102 400128 316170
rect 399808 316046 399878 316102
rect 399934 316046 400002 316102
rect 400058 316046 400128 316102
rect 399808 315978 400128 316046
rect 399808 315922 399878 315978
rect 399934 315922 400002 315978
rect 400058 315922 400128 315978
rect 399808 315888 400128 315922
rect 404778 311926 405398 327922
rect 408498 598172 409118 598268
rect 408498 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 409118 598172
rect 408498 598048 409118 598116
rect 408498 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 409118 598048
rect 408498 597924 409118 597992
rect 408498 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 409118 597924
rect 408498 597800 409118 597868
rect 408498 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 409118 597800
rect 408498 586350 409118 597744
rect 408498 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 409118 586350
rect 408498 586226 409118 586294
rect 408498 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 409118 586226
rect 408498 586102 409118 586170
rect 408498 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 409118 586102
rect 408498 585978 409118 586046
rect 408498 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 409118 585978
rect 408498 568350 409118 585922
rect 408498 568294 408594 568350
rect 408650 568294 408718 568350
rect 408774 568294 408842 568350
rect 408898 568294 408966 568350
rect 409022 568294 409118 568350
rect 408498 568226 409118 568294
rect 408498 568170 408594 568226
rect 408650 568170 408718 568226
rect 408774 568170 408842 568226
rect 408898 568170 408966 568226
rect 409022 568170 409118 568226
rect 408498 568102 409118 568170
rect 408498 568046 408594 568102
rect 408650 568046 408718 568102
rect 408774 568046 408842 568102
rect 408898 568046 408966 568102
rect 409022 568046 409118 568102
rect 408498 567978 409118 568046
rect 408498 567922 408594 567978
rect 408650 567922 408718 567978
rect 408774 567922 408842 567978
rect 408898 567922 408966 567978
rect 409022 567922 409118 567978
rect 408498 550350 409118 567922
rect 408498 550294 408594 550350
rect 408650 550294 408718 550350
rect 408774 550294 408842 550350
rect 408898 550294 408966 550350
rect 409022 550294 409118 550350
rect 408498 550226 409118 550294
rect 408498 550170 408594 550226
rect 408650 550170 408718 550226
rect 408774 550170 408842 550226
rect 408898 550170 408966 550226
rect 409022 550170 409118 550226
rect 408498 550102 409118 550170
rect 408498 550046 408594 550102
rect 408650 550046 408718 550102
rect 408774 550046 408842 550102
rect 408898 550046 408966 550102
rect 409022 550046 409118 550102
rect 408498 549978 409118 550046
rect 408498 549922 408594 549978
rect 408650 549922 408718 549978
rect 408774 549922 408842 549978
rect 408898 549922 408966 549978
rect 409022 549922 409118 549978
rect 408498 532350 409118 549922
rect 408498 532294 408594 532350
rect 408650 532294 408718 532350
rect 408774 532294 408842 532350
rect 408898 532294 408966 532350
rect 409022 532294 409118 532350
rect 408498 532226 409118 532294
rect 408498 532170 408594 532226
rect 408650 532170 408718 532226
rect 408774 532170 408842 532226
rect 408898 532170 408966 532226
rect 409022 532170 409118 532226
rect 408498 532102 409118 532170
rect 408498 532046 408594 532102
rect 408650 532046 408718 532102
rect 408774 532046 408842 532102
rect 408898 532046 408966 532102
rect 409022 532046 409118 532102
rect 408498 531978 409118 532046
rect 408498 531922 408594 531978
rect 408650 531922 408718 531978
rect 408774 531922 408842 531978
rect 408898 531922 408966 531978
rect 409022 531922 409118 531978
rect 408498 514350 409118 531922
rect 408498 514294 408594 514350
rect 408650 514294 408718 514350
rect 408774 514294 408842 514350
rect 408898 514294 408966 514350
rect 409022 514294 409118 514350
rect 408498 514226 409118 514294
rect 408498 514170 408594 514226
rect 408650 514170 408718 514226
rect 408774 514170 408842 514226
rect 408898 514170 408966 514226
rect 409022 514170 409118 514226
rect 408498 514102 409118 514170
rect 408498 514046 408594 514102
rect 408650 514046 408718 514102
rect 408774 514046 408842 514102
rect 408898 514046 408966 514102
rect 409022 514046 409118 514102
rect 408498 513978 409118 514046
rect 408498 513922 408594 513978
rect 408650 513922 408718 513978
rect 408774 513922 408842 513978
rect 408898 513922 408966 513978
rect 409022 513922 409118 513978
rect 408498 496350 409118 513922
rect 408498 496294 408594 496350
rect 408650 496294 408718 496350
rect 408774 496294 408842 496350
rect 408898 496294 408966 496350
rect 409022 496294 409118 496350
rect 408498 496226 409118 496294
rect 408498 496170 408594 496226
rect 408650 496170 408718 496226
rect 408774 496170 408842 496226
rect 408898 496170 408966 496226
rect 409022 496170 409118 496226
rect 408498 496102 409118 496170
rect 408498 496046 408594 496102
rect 408650 496046 408718 496102
rect 408774 496046 408842 496102
rect 408898 496046 408966 496102
rect 409022 496046 409118 496102
rect 408498 495978 409118 496046
rect 408498 495922 408594 495978
rect 408650 495922 408718 495978
rect 408774 495922 408842 495978
rect 408898 495922 408966 495978
rect 409022 495922 409118 495978
rect 408498 478350 409118 495922
rect 408498 478294 408594 478350
rect 408650 478294 408718 478350
rect 408774 478294 408842 478350
rect 408898 478294 408966 478350
rect 409022 478294 409118 478350
rect 408498 478226 409118 478294
rect 408498 478170 408594 478226
rect 408650 478170 408718 478226
rect 408774 478170 408842 478226
rect 408898 478170 408966 478226
rect 409022 478170 409118 478226
rect 408498 478102 409118 478170
rect 408498 478046 408594 478102
rect 408650 478046 408718 478102
rect 408774 478046 408842 478102
rect 408898 478046 408966 478102
rect 409022 478046 409118 478102
rect 408498 477978 409118 478046
rect 408498 477922 408594 477978
rect 408650 477922 408718 477978
rect 408774 477922 408842 477978
rect 408898 477922 408966 477978
rect 409022 477922 409118 477978
rect 408498 460350 409118 477922
rect 408498 460294 408594 460350
rect 408650 460294 408718 460350
rect 408774 460294 408842 460350
rect 408898 460294 408966 460350
rect 409022 460294 409118 460350
rect 408498 460226 409118 460294
rect 408498 460170 408594 460226
rect 408650 460170 408718 460226
rect 408774 460170 408842 460226
rect 408898 460170 408966 460226
rect 409022 460170 409118 460226
rect 408498 460102 409118 460170
rect 408498 460046 408594 460102
rect 408650 460046 408718 460102
rect 408774 460046 408842 460102
rect 408898 460046 408966 460102
rect 409022 460046 409118 460102
rect 408498 459978 409118 460046
rect 408498 459922 408594 459978
rect 408650 459922 408718 459978
rect 408774 459922 408842 459978
rect 408898 459922 408966 459978
rect 409022 459922 409118 459978
rect 408498 442350 409118 459922
rect 408498 442294 408594 442350
rect 408650 442294 408718 442350
rect 408774 442294 408842 442350
rect 408898 442294 408966 442350
rect 409022 442294 409118 442350
rect 408498 442226 409118 442294
rect 408498 442170 408594 442226
rect 408650 442170 408718 442226
rect 408774 442170 408842 442226
rect 408898 442170 408966 442226
rect 409022 442170 409118 442226
rect 408498 442102 409118 442170
rect 408498 442046 408594 442102
rect 408650 442046 408718 442102
rect 408774 442046 408842 442102
rect 408898 442046 408966 442102
rect 409022 442046 409118 442102
rect 408498 441978 409118 442046
rect 408498 441922 408594 441978
rect 408650 441922 408718 441978
rect 408774 441922 408842 441978
rect 408898 441922 408966 441978
rect 409022 441922 409118 441978
rect 408498 424350 409118 441922
rect 408498 424294 408594 424350
rect 408650 424294 408718 424350
rect 408774 424294 408842 424350
rect 408898 424294 408966 424350
rect 409022 424294 409118 424350
rect 408498 424226 409118 424294
rect 408498 424170 408594 424226
rect 408650 424170 408718 424226
rect 408774 424170 408842 424226
rect 408898 424170 408966 424226
rect 409022 424170 409118 424226
rect 408498 424102 409118 424170
rect 408498 424046 408594 424102
rect 408650 424046 408718 424102
rect 408774 424046 408842 424102
rect 408898 424046 408966 424102
rect 409022 424046 409118 424102
rect 408498 423978 409118 424046
rect 408498 423922 408594 423978
rect 408650 423922 408718 423978
rect 408774 423922 408842 423978
rect 408898 423922 408966 423978
rect 409022 423922 409118 423978
rect 408498 406350 409118 423922
rect 408498 406294 408594 406350
rect 408650 406294 408718 406350
rect 408774 406294 408842 406350
rect 408898 406294 408966 406350
rect 409022 406294 409118 406350
rect 408498 406226 409118 406294
rect 408498 406170 408594 406226
rect 408650 406170 408718 406226
rect 408774 406170 408842 406226
rect 408898 406170 408966 406226
rect 409022 406170 409118 406226
rect 408498 406102 409118 406170
rect 408498 406046 408594 406102
rect 408650 406046 408718 406102
rect 408774 406046 408842 406102
rect 408898 406046 408966 406102
rect 409022 406046 409118 406102
rect 408498 405978 409118 406046
rect 408498 405922 408594 405978
rect 408650 405922 408718 405978
rect 408774 405922 408842 405978
rect 408898 405922 408966 405978
rect 409022 405922 409118 405978
rect 408498 388350 409118 405922
rect 408498 388294 408594 388350
rect 408650 388294 408718 388350
rect 408774 388294 408842 388350
rect 408898 388294 408966 388350
rect 409022 388294 409118 388350
rect 408498 388226 409118 388294
rect 408498 388170 408594 388226
rect 408650 388170 408718 388226
rect 408774 388170 408842 388226
rect 408898 388170 408966 388226
rect 409022 388170 409118 388226
rect 408498 388102 409118 388170
rect 408498 388046 408594 388102
rect 408650 388046 408718 388102
rect 408774 388046 408842 388102
rect 408898 388046 408966 388102
rect 409022 388046 409118 388102
rect 408498 387978 409118 388046
rect 408498 387922 408594 387978
rect 408650 387922 408718 387978
rect 408774 387922 408842 387978
rect 408898 387922 408966 387978
rect 409022 387922 409118 387978
rect 408498 370350 409118 387922
rect 408498 370294 408594 370350
rect 408650 370294 408718 370350
rect 408774 370294 408842 370350
rect 408898 370294 408966 370350
rect 409022 370294 409118 370350
rect 408498 370226 409118 370294
rect 408498 370170 408594 370226
rect 408650 370170 408718 370226
rect 408774 370170 408842 370226
rect 408898 370170 408966 370226
rect 409022 370170 409118 370226
rect 408498 370102 409118 370170
rect 408498 370046 408594 370102
rect 408650 370046 408718 370102
rect 408774 370046 408842 370102
rect 408898 370046 408966 370102
rect 409022 370046 409118 370102
rect 408498 369978 409118 370046
rect 408498 369922 408594 369978
rect 408650 369922 408718 369978
rect 408774 369922 408842 369978
rect 408898 369922 408966 369978
rect 409022 369922 409118 369978
rect 408498 352350 409118 369922
rect 408498 352294 408594 352350
rect 408650 352294 408718 352350
rect 408774 352294 408842 352350
rect 408898 352294 408966 352350
rect 409022 352294 409118 352350
rect 408498 352226 409118 352294
rect 408498 352170 408594 352226
rect 408650 352170 408718 352226
rect 408774 352170 408842 352226
rect 408898 352170 408966 352226
rect 409022 352170 409118 352226
rect 408498 352102 409118 352170
rect 408498 352046 408594 352102
rect 408650 352046 408718 352102
rect 408774 352046 408842 352102
rect 408898 352046 408966 352102
rect 409022 352046 409118 352102
rect 408498 351978 409118 352046
rect 408498 351922 408594 351978
rect 408650 351922 408718 351978
rect 408774 351922 408842 351978
rect 408898 351922 408966 351978
rect 409022 351922 409118 351978
rect 408498 334350 409118 351922
rect 408498 334294 408594 334350
rect 408650 334294 408718 334350
rect 408774 334294 408842 334350
rect 408898 334294 408966 334350
rect 409022 334294 409118 334350
rect 408498 334226 409118 334294
rect 408498 334170 408594 334226
rect 408650 334170 408718 334226
rect 408774 334170 408842 334226
rect 408898 334170 408966 334226
rect 409022 334170 409118 334226
rect 408498 334102 409118 334170
rect 408498 334046 408594 334102
rect 408650 334046 408718 334102
rect 408774 334046 408842 334102
rect 408898 334046 408966 334102
rect 409022 334046 409118 334102
rect 408498 333978 409118 334046
rect 408498 333922 408594 333978
rect 408650 333922 408718 333978
rect 408774 333922 408842 333978
rect 408898 333922 408966 333978
rect 409022 333922 409118 333978
rect 408498 316350 409118 333922
rect 435498 597212 436118 598268
rect 435498 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 436118 597212
rect 435498 597088 436118 597156
rect 435498 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 436118 597088
rect 435498 596964 436118 597032
rect 435498 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 436118 596964
rect 435498 596840 436118 596908
rect 435498 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 436118 596840
rect 435498 580350 436118 596784
rect 435498 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 436118 580350
rect 435498 580226 436118 580294
rect 435498 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 436118 580226
rect 435498 580102 436118 580170
rect 435498 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 436118 580102
rect 435498 579978 436118 580046
rect 435498 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 436118 579978
rect 435498 562350 436118 579922
rect 435498 562294 435594 562350
rect 435650 562294 435718 562350
rect 435774 562294 435842 562350
rect 435898 562294 435966 562350
rect 436022 562294 436118 562350
rect 435498 562226 436118 562294
rect 435498 562170 435594 562226
rect 435650 562170 435718 562226
rect 435774 562170 435842 562226
rect 435898 562170 435966 562226
rect 436022 562170 436118 562226
rect 435498 562102 436118 562170
rect 435498 562046 435594 562102
rect 435650 562046 435718 562102
rect 435774 562046 435842 562102
rect 435898 562046 435966 562102
rect 436022 562046 436118 562102
rect 435498 561978 436118 562046
rect 435498 561922 435594 561978
rect 435650 561922 435718 561978
rect 435774 561922 435842 561978
rect 435898 561922 435966 561978
rect 436022 561922 436118 561978
rect 435498 544350 436118 561922
rect 435498 544294 435594 544350
rect 435650 544294 435718 544350
rect 435774 544294 435842 544350
rect 435898 544294 435966 544350
rect 436022 544294 436118 544350
rect 435498 544226 436118 544294
rect 435498 544170 435594 544226
rect 435650 544170 435718 544226
rect 435774 544170 435842 544226
rect 435898 544170 435966 544226
rect 436022 544170 436118 544226
rect 435498 544102 436118 544170
rect 435498 544046 435594 544102
rect 435650 544046 435718 544102
rect 435774 544046 435842 544102
rect 435898 544046 435966 544102
rect 436022 544046 436118 544102
rect 435498 543978 436118 544046
rect 435498 543922 435594 543978
rect 435650 543922 435718 543978
rect 435774 543922 435842 543978
rect 435898 543922 435966 543978
rect 436022 543922 436118 543978
rect 435498 526350 436118 543922
rect 435498 526294 435594 526350
rect 435650 526294 435718 526350
rect 435774 526294 435842 526350
rect 435898 526294 435966 526350
rect 436022 526294 436118 526350
rect 435498 526226 436118 526294
rect 435498 526170 435594 526226
rect 435650 526170 435718 526226
rect 435774 526170 435842 526226
rect 435898 526170 435966 526226
rect 436022 526170 436118 526226
rect 435498 526102 436118 526170
rect 435498 526046 435594 526102
rect 435650 526046 435718 526102
rect 435774 526046 435842 526102
rect 435898 526046 435966 526102
rect 436022 526046 436118 526102
rect 435498 525978 436118 526046
rect 435498 525922 435594 525978
rect 435650 525922 435718 525978
rect 435774 525922 435842 525978
rect 435898 525922 435966 525978
rect 436022 525922 436118 525978
rect 435498 508350 436118 525922
rect 435498 508294 435594 508350
rect 435650 508294 435718 508350
rect 435774 508294 435842 508350
rect 435898 508294 435966 508350
rect 436022 508294 436118 508350
rect 435498 508226 436118 508294
rect 435498 508170 435594 508226
rect 435650 508170 435718 508226
rect 435774 508170 435842 508226
rect 435898 508170 435966 508226
rect 436022 508170 436118 508226
rect 435498 508102 436118 508170
rect 435498 508046 435594 508102
rect 435650 508046 435718 508102
rect 435774 508046 435842 508102
rect 435898 508046 435966 508102
rect 436022 508046 436118 508102
rect 435498 507978 436118 508046
rect 435498 507922 435594 507978
rect 435650 507922 435718 507978
rect 435774 507922 435842 507978
rect 435898 507922 435966 507978
rect 436022 507922 436118 507978
rect 435498 490350 436118 507922
rect 435498 490294 435594 490350
rect 435650 490294 435718 490350
rect 435774 490294 435842 490350
rect 435898 490294 435966 490350
rect 436022 490294 436118 490350
rect 435498 490226 436118 490294
rect 435498 490170 435594 490226
rect 435650 490170 435718 490226
rect 435774 490170 435842 490226
rect 435898 490170 435966 490226
rect 436022 490170 436118 490226
rect 435498 490102 436118 490170
rect 435498 490046 435594 490102
rect 435650 490046 435718 490102
rect 435774 490046 435842 490102
rect 435898 490046 435966 490102
rect 436022 490046 436118 490102
rect 435498 489978 436118 490046
rect 435498 489922 435594 489978
rect 435650 489922 435718 489978
rect 435774 489922 435842 489978
rect 435898 489922 435966 489978
rect 436022 489922 436118 489978
rect 435498 472350 436118 489922
rect 435498 472294 435594 472350
rect 435650 472294 435718 472350
rect 435774 472294 435842 472350
rect 435898 472294 435966 472350
rect 436022 472294 436118 472350
rect 435498 472226 436118 472294
rect 435498 472170 435594 472226
rect 435650 472170 435718 472226
rect 435774 472170 435842 472226
rect 435898 472170 435966 472226
rect 436022 472170 436118 472226
rect 435498 472102 436118 472170
rect 435498 472046 435594 472102
rect 435650 472046 435718 472102
rect 435774 472046 435842 472102
rect 435898 472046 435966 472102
rect 436022 472046 436118 472102
rect 435498 471978 436118 472046
rect 435498 471922 435594 471978
rect 435650 471922 435718 471978
rect 435774 471922 435842 471978
rect 435898 471922 435966 471978
rect 436022 471922 436118 471978
rect 435498 454350 436118 471922
rect 435498 454294 435594 454350
rect 435650 454294 435718 454350
rect 435774 454294 435842 454350
rect 435898 454294 435966 454350
rect 436022 454294 436118 454350
rect 435498 454226 436118 454294
rect 435498 454170 435594 454226
rect 435650 454170 435718 454226
rect 435774 454170 435842 454226
rect 435898 454170 435966 454226
rect 436022 454170 436118 454226
rect 435498 454102 436118 454170
rect 435498 454046 435594 454102
rect 435650 454046 435718 454102
rect 435774 454046 435842 454102
rect 435898 454046 435966 454102
rect 436022 454046 436118 454102
rect 435498 453978 436118 454046
rect 435498 453922 435594 453978
rect 435650 453922 435718 453978
rect 435774 453922 435842 453978
rect 435898 453922 435966 453978
rect 436022 453922 436118 453978
rect 435498 436350 436118 453922
rect 435498 436294 435594 436350
rect 435650 436294 435718 436350
rect 435774 436294 435842 436350
rect 435898 436294 435966 436350
rect 436022 436294 436118 436350
rect 435498 436226 436118 436294
rect 435498 436170 435594 436226
rect 435650 436170 435718 436226
rect 435774 436170 435842 436226
rect 435898 436170 435966 436226
rect 436022 436170 436118 436226
rect 435498 436102 436118 436170
rect 435498 436046 435594 436102
rect 435650 436046 435718 436102
rect 435774 436046 435842 436102
rect 435898 436046 435966 436102
rect 436022 436046 436118 436102
rect 435498 435978 436118 436046
rect 435498 435922 435594 435978
rect 435650 435922 435718 435978
rect 435774 435922 435842 435978
rect 435898 435922 435966 435978
rect 436022 435922 436118 435978
rect 435498 418350 436118 435922
rect 435498 418294 435594 418350
rect 435650 418294 435718 418350
rect 435774 418294 435842 418350
rect 435898 418294 435966 418350
rect 436022 418294 436118 418350
rect 435498 418226 436118 418294
rect 435498 418170 435594 418226
rect 435650 418170 435718 418226
rect 435774 418170 435842 418226
rect 435898 418170 435966 418226
rect 436022 418170 436118 418226
rect 435498 418102 436118 418170
rect 435498 418046 435594 418102
rect 435650 418046 435718 418102
rect 435774 418046 435842 418102
rect 435898 418046 435966 418102
rect 436022 418046 436118 418102
rect 435498 417978 436118 418046
rect 435498 417922 435594 417978
rect 435650 417922 435718 417978
rect 435774 417922 435842 417978
rect 435898 417922 435966 417978
rect 436022 417922 436118 417978
rect 435498 400350 436118 417922
rect 435498 400294 435594 400350
rect 435650 400294 435718 400350
rect 435774 400294 435842 400350
rect 435898 400294 435966 400350
rect 436022 400294 436118 400350
rect 435498 400226 436118 400294
rect 435498 400170 435594 400226
rect 435650 400170 435718 400226
rect 435774 400170 435842 400226
rect 435898 400170 435966 400226
rect 436022 400170 436118 400226
rect 435498 400102 436118 400170
rect 435498 400046 435594 400102
rect 435650 400046 435718 400102
rect 435774 400046 435842 400102
rect 435898 400046 435966 400102
rect 436022 400046 436118 400102
rect 435498 399978 436118 400046
rect 435498 399922 435594 399978
rect 435650 399922 435718 399978
rect 435774 399922 435842 399978
rect 435898 399922 435966 399978
rect 436022 399922 436118 399978
rect 435498 382350 436118 399922
rect 435498 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 436118 382350
rect 435498 382226 436118 382294
rect 435498 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 436118 382226
rect 435498 382102 436118 382170
rect 435498 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 436118 382102
rect 435498 381978 436118 382046
rect 435498 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 436118 381978
rect 435498 364350 436118 381922
rect 435498 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 436118 364350
rect 435498 364226 436118 364294
rect 435498 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 436118 364226
rect 435498 364102 436118 364170
rect 435498 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 436118 364102
rect 435498 363978 436118 364046
rect 435498 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 436118 363978
rect 435498 346350 436118 363922
rect 435498 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 436118 346350
rect 435498 346226 436118 346294
rect 435498 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 436118 346226
rect 435498 346102 436118 346170
rect 435498 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 436118 346102
rect 435498 345978 436118 346046
rect 435498 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 436118 345978
rect 435498 328350 436118 345922
rect 435498 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 436118 328350
rect 435498 328226 436118 328294
rect 435498 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 436118 328226
rect 423948 328132 424004 328142
rect 420140 327908 420196 327918
rect 420028 327796 420084 327806
rect 410732 324996 410788 325006
rect 410732 324436 410788 324940
rect 410732 324370 410788 324380
rect 411404 324436 411572 324478
rect 411460 324422 411572 324436
rect 411404 324370 411460 324380
rect 408498 316294 408594 316350
rect 408650 316294 408718 316350
rect 408774 316294 408842 316350
rect 408898 316294 408966 316350
rect 409022 316294 409118 316350
rect 408498 316226 409118 316294
rect 408498 316170 408594 316226
rect 408650 316170 408718 316226
rect 408774 316170 408842 316226
rect 408898 316170 408966 316226
rect 409022 316170 409118 316226
rect 408498 316102 409118 316170
rect 408498 316046 408594 316102
rect 408650 316046 408718 316102
rect 408774 316046 408842 316102
rect 408898 316046 408966 316102
rect 409022 316046 409118 316102
rect 408498 315978 409118 316046
rect 408498 315922 408594 315978
rect 408650 315922 408718 315978
rect 408774 315922 408842 315978
rect 408898 315922 408966 315978
rect 409022 315922 409118 315978
rect 408498 311926 409118 315922
rect 411516 312598 411572 324422
rect 418348 324436 418404 324446
rect 418348 314188 418404 324380
rect 418796 324436 418852 324446
rect 418348 314132 418516 314188
rect 411516 312532 411572 312542
rect 415168 310350 415488 310384
rect 415168 310294 415238 310350
rect 415294 310294 415362 310350
rect 415418 310294 415488 310350
rect 415168 310226 415488 310294
rect 415168 310170 415238 310226
rect 415294 310170 415362 310226
rect 415418 310170 415488 310226
rect 415168 310102 415488 310170
rect 415168 310046 415238 310102
rect 415294 310046 415362 310102
rect 415418 310046 415488 310102
rect 415168 309978 415488 310046
rect 415168 309922 415238 309978
rect 415294 309922 415362 309978
rect 415418 309922 415488 309978
rect 415168 309888 415488 309922
rect 399808 298350 400128 298384
rect 399808 298294 399878 298350
rect 399934 298294 400002 298350
rect 400058 298294 400128 298350
rect 399808 298226 400128 298294
rect 399808 298170 399878 298226
rect 399934 298170 400002 298226
rect 400058 298170 400128 298226
rect 399808 298102 400128 298170
rect 399808 298046 399878 298102
rect 399934 298046 400002 298102
rect 400058 298046 400128 298102
rect 399808 297978 400128 298046
rect 399808 297922 399878 297978
rect 399934 297922 400002 297978
rect 400058 297922 400128 297978
rect 399808 297888 400128 297922
rect 415168 292350 415488 292384
rect 415168 292294 415238 292350
rect 415294 292294 415362 292350
rect 415418 292294 415488 292350
rect 415168 292226 415488 292294
rect 415168 292170 415238 292226
rect 415294 292170 415362 292226
rect 415418 292170 415488 292226
rect 415168 292102 415488 292170
rect 415168 292046 415238 292102
rect 415294 292046 415362 292102
rect 415418 292046 415488 292102
rect 415168 291978 415488 292046
rect 415168 291922 415238 291978
rect 415294 291922 415362 291978
rect 415418 291922 415488 291978
rect 415168 291888 415488 291922
rect 387212 272066 387268 272076
rect 387324 286138 387380 286148
rect 387324 271348 387380 286082
rect 399808 280350 400128 280384
rect 399808 280294 399878 280350
rect 399934 280294 400002 280350
rect 400058 280294 400128 280350
rect 399808 280226 400128 280294
rect 399808 280170 399878 280226
rect 399934 280170 400002 280226
rect 400058 280170 400128 280226
rect 399808 280102 400128 280170
rect 399808 280046 399878 280102
rect 399934 280046 400002 280102
rect 400058 280046 400128 280102
rect 399808 279978 400128 280046
rect 399808 279922 399878 279978
rect 399934 279922 400002 279978
rect 400058 279922 400128 279978
rect 399808 279888 400128 279922
rect 404012 272244 404068 272254
rect 387324 271282 387380 271292
rect 387436 271908 387492 271918
rect 385420 270592 385476 270602
rect 387436 261658 387492 271852
rect 388108 271124 388164 271134
rect 387996 270452 388052 270462
rect 387996 268858 388052 270396
rect 387996 268792 388052 268802
rect 388108 261716 388164 271068
rect 388108 261650 388164 261660
rect 403564 265748 403620 265758
rect 403564 264292 403620 265692
rect 404012 265076 404068 272188
rect 404012 265010 404068 265020
rect 387436 261592 387492 261602
rect 403564 261298 403620 264236
rect 406252 264292 406308 264302
rect 406252 263396 406308 264236
rect 406252 263330 406308 263340
rect 406924 264292 406980 264302
rect 406924 263396 406980 264236
rect 406924 263330 406980 263340
rect 408498 262350 409118 275930
rect 416332 271684 416388 271694
rect 408498 262294 408594 262350
rect 408650 262294 408718 262350
rect 408774 262294 408842 262350
rect 408898 262294 408966 262350
rect 409022 262294 409118 262350
rect 408498 262226 409118 262294
rect 408498 262170 408594 262226
rect 408650 262170 408718 262226
rect 408774 262170 408842 262226
rect 408898 262170 408966 262226
rect 409022 262170 409118 262226
rect 408498 262102 409118 262170
rect 408498 262046 408594 262102
rect 408650 262046 408718 262102
rect 408774 262046 408842 262102
rect 408898 262046 408966 262102
rect 409022 262046 409118 262102
rect 408498 261978 409118 262046
rect 408498 261922 408594 261978
rect 408650 261922 408718 261978
rect 408774 261922 408842 261978
rect 408898 261922 408966 261978
rect 409022 261922 409118 261978
rect 408498 261638 409118 261922
rect 409948 271236 410004 271246
rect 409948 261604 410004 271180
rect 410060 271124 410116 271134
rect 410060 263060 410116 271068
rect 411628 271124 411684 271134
rect 410956 265748 411012 265758
rect 410956 264292 411012 265692
rect 410956 263732 411012 264236
rect 410956 263666 411012 263676
rect 411628 263620 411684 271068
rect 413308 271124 413364 271134
rect 411628 263554 411684 263564
rect 411740 268996 411796 269006
rect 411740 263396 411796 268940
rect 413308 264538 413364 271068
rect 413308 264472 413364 264482
rect 414988 271124 415044 271134
rect 411740 263330 411796 263340
rect 413644 264292 413700 264302
rect 413644 263172 413700 264236
rect 414988 263508 415044 271068
rect 416332 268138 416388 271628
rect 416332 268072 416388 268082
rect 418348 271124 418404 271134
rect 414988 263442 415044 263452
rect 413644 263106 413700 263116
rect 410060 262994 410116 263004
rect 418348 263060 418404 271068
rect 418460 270340 418516 314132
rect 418460 270274 418516 270284
rect 418572 312598 418628 312608
rect 418572 267204 418628 312542
rect 418796 268996 418852 324380
rect 418796 268930 418852 268940
rect 419916 272020 419972 272030
rect 419916 267316 419972 271964
rect 420028 269892 420084 327740
rect 420140 271236 420196 327852
rect 423388 324996 423444 325006
rect 421260 324436 421540 324478
rect 421316 324422 421540 324436
rect 421260 324370 421316 324380
rect 420140 271170 420196 271180
rect 420028 269826 420084 269836
rect 421484 268772 421540 324422
rect 422044 324436 422100 324446
rect 422044 270340 422100 324380
rect 422604 324436 422660 324446
rect 422604 273364 422660 324380
rect 422604 273298 422660 273308
rect 423388 272020 423444 324940
rect 423948 273252 424004 328076
rect 435498 328102 436118 328170
rect 435498 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 436118 328102
rect 431788 328020 431844 328030
rect 426860 327796 426916 327806
rect 426748 327684 426804 327694
rect 424172 324436 424228 324446
rect 424172 278908 424228 324380
rect 425068 324436 425124 324446
rect 424172 278852 424676 278908
rect 423948 273186 424004 273196
rect 423388 271954 423444 271964
rect 422044 270274 422100 270284
rect 421484 268706 421540 268716
rect 424620 267958 424676 278852
rect 425068 271684 425124 324380
rect 425068 271618 425124 271628
rect 426188 324436 426244 324446
rect 424620 267876 424676 267902
rect 424620 267810 424676 267820
rect 419916 267250 419972 267260
rect 418572 267138 418628 267148
rect 420364 267238 420420 267248
rect 420364 267138 420420 267148
rect 426188 263732 426244 324380
rect 426412 324436 426468 324446
rect 426412 323428 426468 324380
rect 426412 323362 426468 323372
rect 426748 268100 426804 327628
rect 426748 268034 426804 268044
rect 426860 267764 426916 327740
rect 426860 267698 426916 267708
rect 428428 326228 428484 326238
rect 428428 267428 428484 326172
rect 430528 316350 430848 316384
rect 430528 316294 430598 316350
rect 430654 316294 430722 316350
rect 430778 316294 430848 316350
rect 430528 316226 430848 316294
rect 430528 316170 430598 316226
rect 430654 316170 430722 316226
rect 430778 316170 430848 316226
rect 430528 316102 430848 316170
rect 430528 316046 430598 316102
rect 430654 316046 430722 316102
rect 430778 316046 430848 316102
rect 430528 315978 430848 316046
rect 430528 315922 430598 315978
rect 430654 315922 430722 315978
rect 430778 315922 430848 315978
rect 430528 315888 430848 315922
rect 430528 298350 430848 298384
rect 430528 298294 430598 298350
rect 430654 298294 430722 298350
rect 430778 298294 430848 298350
rect 430528 298226 430848 298294
rect 430528 298170 430598 298226
rect 430654 298170 430722 298226
rect 430778 298170 430848 298226
rect 430528 298102 430848 298170
rect 430528 298046 430598 298102
rect 430654 298046 430722 298102
rect 430778 298046 430848 298102
rect 430528 297978 430848 298046
rect 430528 297922 430598 297978
rect 430654 297922 430722 297978
rect 430778 297922 430848 297978
rect 430528 297888 430848 297922
rect 430528 280350 430848 280384
rect 430528 280294 430598 280350
rect 430654 280294 430722 280350
rect 430778 280294 430848 280350
rect 430528 280226 430848 280294
rect 430528 280170 430598 280226
rect 430654 280170 430722 280226
rect 430778 280170 430848 280226
rect 430528 280102 430848 280170
rect 430528 280046 430598 280102
rect 430654 280046 430722 280102
rect 430778 280046 430848 280102
rect 430528 279978 430848 280046
rect 430528 279922 430598 279978
rect 430654 279922 430722 279978
rect 430778 279922 430848 279978
rect 430528 279888 430848 279922
rect 431788 271796 431844 327964
rect 435498 327978 436118 328046
rect 435498 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 436118 327978
rect 433468 326116 433524 326126
rect 431788 271730 431844 271740
rect 432124 324548 432180 324558
rect 431788 271572 431844 271582
rect 428428 267362 428484 267372
rect 430108 271460 430164 271470
rect 426188 263666 426244 263676
rect 418348 262994 418404 263004
rect 409948 261538 410004 261548
rect 403564 261232 403620 261242
rect 383852 260332 383908 260342
rect 384448 256350 384768 256384
rect 384448 256294 384518 256350
rect 384574 256294 384642 256350
rect 384698 256294 384768 256350
rect 384448 256226 384768 256294
rect 384448 256170 384518 256226
rect 384574 256170 384642 256226
rect 384698 256170 384768 256226
rect 384448 256102 384768 256170
rect 384448 256046 384518 256102
rect 384574 256046 384642 256102
rect 384698 256046 384768 256102
rect 384448 255978 384768 256046
rect 384448 255922 384518 255978
rect 384574 255922 384642 255978
rect 384698 255922 384768 255978
rect 384448 255888 384768 255922
rect 415168 256350 415488 256384
rect 415168 256294 415238 256350
rect 415294 256294 415362 256350
rect 415418 256294 415488 256350
rect 415168 256226 415488 256294
rect 415168 256170 415238 256226
rect 415294 256170 415362 256226
rect 415418 256170 415488 256226
rect 415168 256102 415488 256170
rect 415168 256046 415238 256102
rect 415294 256046 415362 256102
rect 415418 256046 415488 256102
rect 415168 255978 415488 256046
rect 415168 255922 415238 255978
rect 415294 255922 415362 255978
rect 415418 255922 415488 255978
rect 415168 255888 415488 255922
rect 399808 244350 400128 244384
rect 399808 244294 399878 244350
rect 399934 244294 400002 244350
rect 400058 244294 400128 244350
rect 399808 244226 400128 244294
rect 399808 244170 399878 244226
rect 399934 244170 400002 244226
rect 400058 244170 400128 244226
rect 399808 244102 400128 244170
rect 399808 244046 399878 244102
rect 399934 244046 400002 244102
rect 400058 244046 400128 244102
rect 399808 243978 400128 244046
rect 399808 243922 399878 243978
rect 399934 243922 400002 243978
rect 400058 243922 400128 243978
rect 399808 243888 400128 243922
rect 381500 241792 381556 241802
rect 384448 238350 384768 238384
rect 384448 238294 384518 238350
rect 384574 238294 384642 238350
rect 384698 238294 384768 238350
rect 384448 238226 384768 238294
rect 384448 238170 384518 238226
rect 384574 238170 384642 238226
rect 384698 238170 384768 238226
rect 384448 238102 384768 238170
rect 384448 238046 384518 238102
rect 384574 238046 384642 238102
rect 384698 238046 384768 238102
rect 384448 237978 384768 238046
rect 384448 237922 384518 237978
rect 384574 237922 384642 237978
rect 384698 237922 384768 237978
rect 384448 237888 384768 237922
rect 415168 238350 415488 238384
rect 415168 238294 415238 238350
rect 415294 238294 415362 238350
rect 415418 238294 415488 238350
rect 415168 238226 415488 238294
rect 415168 238170 415238 238226
rect 415294 238170 415362 238226
rect 415418 238170 415488 238226
rect 415168 238102 415488 238170
rect 415168 238046 415238 238102
rect 415294 238046 415362 238102
rect 415418 238046 415488 238102
rect 415168 237978 415488 238046
rect 415168 237922 415238 237978
rect 415294 237922 415362 237978
rect 415418 237922 415488 237978
rect 415168 237888 415488 237922
rect 380604 231812 380884 231868
rect 380604 220500 380660 220510
rect 380604 220108 380660 220444
rect 380604 220052 380772 220108
rect 380716 215068 380772 220052
rect 380492 204082 380548 204092
rect 380604 215012 380772 215068
rect 380268 203858 380324 203868
rect 380604 203308 380660 215012
rect 380828 203308 380884 231812
rect 399808 226350 400128 226384
rect 399808 226294 399878 226350
rect 399934 226294 400002 226350
rect 400058 226294 400128 226350
rect 399808 226226 400128 226294
rect 399808 226170 399878 226226
rect 399934 226170 400002 226226
rect 400058 226170 400128 226226
rect 399808 226102 400128 226170
rect 399808 226046 399878 226102
rect 399934 226046 400002 226102
rect 400058 226046 400128 226102
rect 399808 225978 400128 226046
rect 399808 225922 399878 225978
rect 399934 225922 400002 225978
rect 400058 225922 400128 225978
rect 399808 225888 400128 225922
rect 384448 220350 384768 220384
rect 384448 220294 384518 220350
rect 384574 220294 384642 220350
rect 384698 220294 384768 220350
rect 384448 220226 384768 220294
rect 384448 220170 384518 220226
rect 384574 220170 384642 220226
rect 384698 220170 384768 220226
rect 384448 220102 384768 220170
rect 384448 220046 384518 220102
rect 384574 220046 384642 220102
rect 384698 220046 384768 220102
rect 384448 219978 384768 220046
rect 384448 219922 384518 219978
rect 384574 219922 384642 219978
rect 384698 219922 384768 219978
rect 384448 219888 384768 219922
rect 415168 220350 415488 220384
rect 415168 220294 415238 220350
rect 415294 220294 415362 220350
rect 415418 220294 415488 220350
rect 415168 220226 415488 220294
rect 415168 220170 415238 220226
rect 415294 220170 415362 220226
rect 415418 220170 415488 220226
rect 415168 220102 415488 220170
rect 415168 220046 415238 220102
rect 415294 220046 415362 220102
rect 415418 220046 415488 220102
rect 415168 219978 415488 220046
rect 415168 219922 415238 219978
rect 415294 219922 415362 219978
rect 415418 219922 415488 219978
rect 415168 219888 415488 219922
rect 381388 218458 381444 218468
rect 381388 215938 381444 218402
rect 383852 217738 383908 217748
rect 381724 217018 381780 217028
rect 381388 215872 381444 215882
rect 381500 216838 381556 216848
rect 381164 209098 381220 209108
rect 381164 205492 381220 209042
rect 381164 205426 381220 205436
rect 380156 161858 380212 161868
rect 380268 203252 380660 203308
rect 380716 203252 380884 203308
rect 380044 159170 380100 159180
rect 380044 145796 380100 145806
rect 380044 135156 380100 145740
rect 380044 135090 380100 135100
rect 379932 132290 379988 132300
rect 380268 133812 380324 203252
rect 380492 198324 380548 198334
rect 380380 166628 380436 166638
rect 380380 166534 380436 166562
rect 380380 158116 380436 158126
rect 380380 134932 380436 158060
rect 380380 134866 380436 134876
rect 380492 134148 380548 198268
rect 380716 196588 380772 203252
rect 380604 196532 380772 196588
rect 381276 199668 381332 199678
rect 380604 154756 380660 196532
rect 380604 151060 380660 154700
rect 380604 150994 380660 151004
rect 380604 149878 380660 149888
rect 380604 149762 380660 149772
rect 380604 145124 380660 145134
rect 380604 145018 380660 145068
rect 380604 144952 380660 144962
rect 380492 134082 380548 134092
rect 380604 141204 380660 141214
rect 380268 126028 380324 133756
rect 380268 125972 380436 126028
rect 380156 117684 380212 117694
rect 380156 117478 380212 117628
rect 380156 75348 380212 117422
rect 380380 114996 380436 125972
rect 380380 114930 380436 114940
rect 380156 75282 380212 75292
rect 379932 72118 379988 72128
rect 379932 66164 379988 72062
rect 379932 65604 379988 66108
rect 379932 65538 379988 65548
rect 380604 44996 380660 141148
rect 381276 134372 381332 199612
rect 381500 149878 381556 216782
rect 381612 215218 381668 215228
rect 381612 156358 381668 215162
rect 381724 195188 381780 216962
rect 382060 215578 382116 215588
rect 381836 215398 381892 215408
rect 381836 205716 381892 215342
rect 381836 205650 381892 205660
rect 381948 213598 382004 213608
rect 381724 195122 381780 195132
rect 381612 156292 381668 156302
rect 381724 166618 381780 166628
rect 381500 149812 381556 149822
rect 381276 134306 381332 134316
rect 381612 134820 381668 134830
rect 381388 132692 381444 132702
rect 381388 128884 381444 132636
rect 381388 128818 381444 128828
rect 381500 132468 381556 132478
rect 381500 126028 381556 132412
rect 381388 125972 381556 126028
rect 381388 72118 381444 125972
rect 381612 78988 381668 134764
rect 381724 127988 381780 166562
rect 381724 127922 381780 127932
rect 381836 132692 381892 132702
rect 381388 72052 381444 72062
rect 381500 78932 381668 78988
rect 381500 74278 381556 78932
rect 381388 71398 381444 71408
rect 381388 45780 381444 71342
rect 381388 45714 381444 45724
rect 381500 45556 381556 74222
rect 381836 72838 381892 132636
rect 381948 125972 382004 213542
rect 382060 205716 382116 215522
rect 382060 199948 382116 205660
rect 382508 213238 382564 213248
rect 382508 203308 382564 213182
rect 383404 211798 383460 211808
rect 383068 207284 383124 207294
rect 382508 203252 382676 203308
rect 382396 203028 382452 203038
rect 382060 199892 382228 199948
rect 382172 135716 382228 199892
rect 382172 135650 382228 135660
rect 382284 145018 382340 145028
rect 381948 124516 382004 125916
rect 381948 124450 382004 124460
rect 382284 124068 382340 144962
rect 382396 136052 382452 202972
rect 382620 161308 382676 203196
rect 383068 197876 383124 207228
rect 383404 205716 383460 211742
rect 383404 205650 383460 205660
rect 383068 197810 383124 197820
rect 383180 205492 383236 205502
rect 382956 196420 383012 196430
rect 382620 161252 382788 161308
rect 382508 151138 382564 151148
rect 382508 137956 382564 151082
rect 382508 137890 382564 137900
rect 382396 135986 382452 135996
rect 382732 134820 382788 161252
rect 382956 135828 383012 196364
rect 382956 135762 383012 135772
rect 383068 137956 383124 137966
rect 382732 134754 382788 134764
rect 383068 130340 383124 137900
rect 383068 130274 383124 130284
rect 383180 132580 383236 205436
rect 383628 203252 383684 203262
rect 383628 135716 383684 203196
rect 383852 201348 383908 217682
rect 383852 201282 383908 201292
rect 384076 217558 384132 217568
rect 384076 202020 384132 217502
rect 395724 214318 395780 214328
rect 386764 212158 386820 212168
rect 386092 210898 386148 210908
rect 385308 206276 385364 206286
rect 385308 205492 385364 206220
rect 385532 206276 385588 206286
rect 385532 205716 385588 206220
rect 385532 205650 385588 205660
rect 385308 205426 385364 205436
rect 386092 205268 386148 210842
rect 386092 205202 386148 205212
rect 386764 205268 386820 212102
rect 392252 211978 392308 211988
rect 386764 205202 386820 205212
rect 389452 211078 389508 211088
rect 389452 205268 389508 211022
rect 389452 205202 389508 205212
rect 384076 187858 384132 201964
rect 384636 202580 384804 202618
rect 384636 202562 384748 202580
rect 384636 202020 384692 202562
rect 384748 202514 384804 202524
rect 390572 202580 391076 202618
rect 390628 202562 391020 202580
rect 390572 202514 390628 202524
rect 391020 202514 391076 202524
rect 384636 201954 384692 201964
rect 384748 201460 384804 201470
rect 384748 199892 384804 201404
rect 392252 201124 392308 211922
rect 392252 201058 392308 201068
rect 395612 205268 395668 205278
rect 384748 199826 384804 199836
rect 389788 198118 389844 198138
rect 389788 198034 389844 198044
rect 384076 187792 384132 187802
rect 384448 184350 384768 184384
rect 384448 184294 384518 184350
rect 384574 184294 384642 184350
rect 384698 184294 384768 184350
rect 384448 184226 384768 184294
rect 384448 184170 384518 184226
rect 384574 184170 384642 184226
rect 384698 184170 384768 184226
rect 384448 184102 384768 184170
rect 384448 184046 384518 184102
rect 384574 184046 384642 184102
rect 384698 184046 384768 184102
rect 384448 183978 384768 184046
rect 384448 183922 384518 183978
rect 384574 183922 384642 183978
rect 384698 183922 384768 183978
rect 384448 183888 384768 183922
rect 395612 182278 395668 205212
rect 395724 197988 395780 214262
rect 399808 208393 400128 208446
rect 399808 208337 399836 208393
rect 399892 208337 399940 208393
rect 399996 208337 400044 208393
rect 400100 208337 400128 208393
rect 399808 208289 400128 208337
rect 399808 208233 399836 208289
rect 399892 208233 399940 208289
rect 399996 208233 400044 208289
rect 400100 208233 400128 208289
rect 399808 208185 400128 208233
rect 399808 208129 399836 208185
rect 399892 208129 399940 208185
rect 399996 208129 400044 208185
rect 400100 208129 400128 208185
rect 399808 208076 400128 208129
rect 399532 207172 399588 207182
rect 399532 205156 399588 207116
rect 399532 205090 399588 205100
rect 403340 206164 403396 206174
rect 403340 205156 403396 206108
rect 403340 205090 403396 205100
rect 402220 204058 402276 204068
rect 402220 203924 402276 204002
rect 402220 203858 402276 203868
rect 404778 202350 405398 215898
rect 408498 208350 409118 215898
rect 408498 208294 408594 208350
rect 408650 208294 408718 208350
rect 408774 208294 408842 208350
rect 408898 208294 408966 208350
rect 409022 208294 409118 208350
rect 408498 208226 409118 208294
rect 408498 208170 408594 208226
rect 408650 208170 408718 208226
rect 408774 208170 408842 208226
rect 408898 208170 408966 208226
rect 409022 208170 409118 208226
rect 408498 208102 409118 208170
rect 408498 208046 408594 208102
rect 408650 208046 408718 208102
rect 408774 208046 408842 208102
rect 408898 208046 408966 208102
rect 409022 208046 409118 208102
rect 408498 207978 409118 208046
rect 408498 207922 408594 207978
rect 408650 207922 408718 207978
rect 408774 207922 408842 207978
rect 408898 207922 408966 207978
rect 409022 207922 409118 207978
rect 407596 205828 407652 205838
rect 407596 205044 407652 205772
rect 407596 204978 407652 204988
rect 404778 202294 404874 202350
rect 404930 202294 404998 202350
rect 405054 202294 405122 202350
rect 405178 202294 405246 202350
rect 405302 202294 405398 202350
rect 404778 202226 405398 202294
rect 404778 202170 404874 202226
rect 404930 202170 404998 202226
rect 405054 202170 405122 202226
rect 405178 202170 405246 202226
rect 405302 202170 405398 202226
rect 404778 202102 405398 202170
rect 404778 202046 404874 202102
rect 404930 202046 404998 202102
rect 405054 202046 405122 202102
rect 405178 202046 405246 202102
rect 405302 202046 405398 202102
rect 404778 201978 405398 202046
rect 404778 201922 404874 201978
rect 404930 201922 404998 201978
rect 405054 201922 405122 201978
rect 405178 201922 405246 201978
rect 405302 201922 405398 201978
rect 395724 197922 395780 197932
rect 397292 201908 397348 201918
rect 397292 192612 397348 201852
rect 397292 192546 397348 192556
rect 399808 190350 400128 190384
rect 399808 190294 399878 190350
rect 399934 190294 400002 190350
rect 400058 190294 400128 190350
rect 399808 190226 400128 190294
rect 399808 190170 399878 190226
rect 399934 190170 400002 190226
rect 400058 190170 400128 190226
rect 399808 190102 400128 190170
rect 399808 190046 399878 190102
rect 399934 190046 400002 190102
rect 400058 190046 400128 190102
rect 399808 189978 400128 190046
rect 399808 189922 399878 189978
rect 399934 189922 400002 189978
rect 400058 189922 400128 189978
rect 399808 189888 400128 189922
rect 404778 184386 405398 201922
rect 404778 184330 404874 184386
rect 404930 184330 404998 184386
rect 405054 184330 405122 184386
rect 405178 184330 405246 184386
rect 405302 184330 405398 184386
rect 404778 184262 405398 184330
rect 404778 184206 404874 184262
rect 404930 184206 404998 184262
rect 405054 184206 405122 184262
rect 405178 184206 405246 184262
rect 405302 184206 405398 184262
rect 404778 184138 405398 184206
rect 404778 184082 404874 184138
rect 404930 184082 404998 184138
rect 405054 184082 405122 184138
rect 405178 184082 405246 184138
rect 405302 184082 405398 184138
rect 404778 184022 405398 184082
rect 408498 190350 409118 207922
rect 418348 213418 418404 213428
rect 410956 207396 411012 207406
rect 410956 205156 411012 207340
rect 417004 206052 417060 206062
rect 410956 205090 411012 205100
rect 414988 205492 415044 205502
rect 414988 205044 415044 205436
rect 417004 205492 417060 205996
rect 417004 205426 417060 205436
rect 414988 204978 415044 204988
rect 418348 198212 418404 213362
rect 418348 198146 418404 198156
rect 430108 198118 430164 271404
rect 430528 244350 430848 244384
rect 430528 244294 430598 244350
rect 430654 244294 430722 244350
rect 430778 244294 430848 244350
rect 430528 244226 430848 244294
rect 430528 244170 430598 244226
rect 430654 244170 430722 244226
rect 430778 244170 430848 244226
rect 430528 244102 430848 244170
rect 430528 244046 430598 244102
rect 430654 244046 430722 244102
rect 430778 244046 430848 244102
rect 430528 243978 430848 244046
rect 430528 243922 430598 243978
rect 430654 243922 430722 243978
rect 430778 243922 430848 243978
rect 430528 243888 430848 243922
rect 431004 242758 431060 242768
rect 430528 226350 430848 226384
rect 430528 226294 430598 226350
rect 430654 226294 430722 226350
rect 430778 226294 430848 226350
rect 430528 226226 430848 226294
rect 430528 226170 430598 226226
rect 430654 226170 430722 226226
rect 430778 226170 430848 226226
rect 430528 226102 430848 226170
rect 430528 226046 430598 226102
rect 430654 226046 430722 226102
rect 430778 226046 430848 226102
rect 430528 225978 430848 226046
rect 430528 225922 430598 225978
rect 430654 225922 430722 225978
rect 430778 225922 430848 225978
rect 430528 225888 430848 225922
rect 430528 208393 430848 208446
rect 430528 208337 430556 208393
rect 430612 208337 430660 208393
rect 430716 208337 430764 208393
rect 430820 208337 430848 208393
rect 430528 208289 430848 208337
rect 430528 208233 430556 208289
rect 430612 208233 430660 208289
rect 430716 208233 430764 208289
rect 430820 208233 430848 208289
rect 430528 208185 430848 208233
rect 430528 208129 430556 208185
rect 430612 208129 430660 208185
rect 430716 208129 430764 208185
rect 430820 208129 430848 208185
rect 430528 208076 430848 208129
rect 430108 198052 430164 198062
rect 423724 194852 423780 194862
rect 423332 194740 423388 194750
rect 423724 194698 423780 194796
rect 423388 194684 423780 194698
rect 423332 194642 423780 194684
rect 408498 190294 408594 190350
rect 408650 190294 408718 190350
rect 408774 190294 408842 190350
rect 408898 190294 408966 190350
rect 409022 190294 409118 190350
rect 408498 190226 409118 190294
rect 408498 190170 408594 190226
rect 408650 190170 408718 190226
rect 408774 190170 408842 190226
rect 408898 190170 408966 190226
rect 409022 190170 409118 190226
rect 408498 190102 409118 190170
rect 408498 190046 408594 190102
rect 408650 190046 408718 190102
rect 408774 190046 408842 190102
rect 408898 190046 408966 190102
rect 409022 190046 409118 190102
rect 408498 189978 409118 190046
rect 408498 189922 408594 189978
rect 408650 189922 408718 189978
rect 408774 189922 408842 189978
rect 408898 189922 408966 189978
rect 409022 189922 409118 189978
rect 408498 184022 409118 189922
rect 430528 190350 430848 190384
rect 430528 190294 430598 190350
rect 430654 190294 430722 190350
rect 430778 190294 430848 190350
rect 430528 190226 430848 190294
rect 430528 190170 430598 190226
rect 430654 190170 430722 190226
rect 430778 190170 430848 190226
rect 430528 190102 430848 190170
rect 430528 190046 430598 190102
rect 430654 190046 430722 190102
rect 430778 190046 430848 190102
rect 430528 189978 430848 190046
rect 430528 189922 430598 189978
rect 430654 189922 430722 189978
rect 430778 189922 430848 189978
rect 430528 189888 430848 189922
rect 431004 188038 431060 242702
rect 431788 206612 431844 271516
rect 431788 205268 431844 206556
rect 431788 205202 431844 205212
rect 431900 271348 431956 271358
rect 431900 205156 431956 271292
rect 431900 205090 431956 205100
rect 431004 187972 431060 187982
rect 431788 204260 431844 204270
rect 415168 184350 415488 184384
rect 415168 184294 415238 184350
rect 415294 184294 415362 184350
rect 415418 184294 415488 184350
rect 415168 184226 415488 184294
rect 415168 184170 415238 184226
rect 415294 184170 415362 184226
rect 415418 184170 415488 184226
rect 415168 184102 415488 184170
rect 415168 184046 415238 184102
rect 415294 184046 415362 184102
rect 415418 184046 415488 184102
rect 415168 183978 415488 184046
rect 415168 183922 415238 183978
rect 415294 183922 415362 183978
rect 415418 183922 415488 183978
rect 415168 183888 415488 183922
rect 395612 182212 395668 182222
rect 399808 172350 400128 172384
rect 399808 172294 399878 172350
rect 399934 172294 400002 172350
rect 400058 172294 400128 172350
rect 399808 172226 400128 172294
rect 399808 172170 399878 172226
rect 399934 172170 400002 172226
rect 400058 172170 400128 172226
rect 399808 172102 400128 172170
rect 399808 172046 399878 172102
rect 399934 172046 400002 172102
rect 400058 172046 400128 172102
rect 399808 171978 400128 172046
rect 399808 171922 399878 171978
rect 399934 171922 400002 171978
rect 400058 171922 400128 171978
rect 399808 171888 400128 171922
rect 430528 172350 430848 172384
rect 430528 172294 430598 172350
rect 430654 172294 430722 172350
rect 430778 172294 430848 172350
rect 430528 172226 430848 172294
rect 430528 172170 430598 172226
rect 430654 172170 430722 172226
rect 430778 172170 430848 172226
rect 430528 172102 430848 172170
rect 430528 172046 430598 172102
rect 430654 172046 430722 172102
rect 430778 172046 430848 172102
rect 430528 171978 430848 172046
rect 430528 171922 430598 171978
rect 430654 171922 430722 171978
rect 430778 171922 430848 171978
rect 430528 171888 430848 171922
rect 384448 166350 384768 166384
rect 384448 166294 384518 166350
rect 384574 166294 384642 166350
rect 384698 166294 384768 166350
rect 384448 166226 384768 166294
rect 384448 166170 384518 166226
rect 384574 166170 384642 166226
rect 384698 166170 384768 166226
rect 384448 166102 384768 166170
rect 384448 166046 384518 166102
rect 384574 166046 384642 166102
rect 384698 166046 384768 166102
rect 384448 165978 384768 166046
rect 384448 165922 384518 165978
rect 384574 165922 384642 165978
rect 384698 165922 384768 165978
rect 384448 165888 384768 165922
rect 415168 166350 415488 166384
rect 415168 166294 415238 166350
rect 415294 166294 415362 166350
rect 415418 166294 415488 166350
rect 415168 166226 415488 166294
rect 415168 166170 415238 166226
rect 415294 166170 415362 166226
rect 415418 166170 415488 166226
rect 415168 166102 415488 166170
rect 415168 166046 415238 166102
rect 415294 166046 415362 166102
rect 415418 166046 415488 166102
rect 415168 165978 415488 166046
rect 415168 165922 415238 165978
rect 415294 165922 415362 165978
rect 415418 165922 415488 165978
rect 415168 165888 415488 165922
rect 399808 154350 400128 154384
rect 399808 154294 399878 154350
rect 399934 154294 400002 154350
rect 400058 154294 400128 154350
rect 399808 154226 400128 154294
rect 399808 154170 399878 154226
rect 399934 154170 400002 154226
rect 400058 154170 400128 154226
rect 399808 154102 400128 154170
rect 399808 154046 399878 154102
rect 399934 154046 400002 154102
rect 400058 154046 400128 154102
rect 399808 153978 400128 154046
rect 399808 153922 399878 153978
rect 399934 153922 400002 153978
rect 400058 153922 400128 153978
rect 399808 153888 400128 153922
rect 430528 154350 430848 154384
rect 430528 154294 430598 154350
rect 430654 154294 430722 154350
rect 430778 154294 430848 154350
rect 430528 154226 430848 154294
rect 430528 154170 430598 154226
rect 430654 154170 430722 154226
rect 430778 154170 430848 154226
rect 430528 154102 430848 154170
rect 430528 154046 430598 154102
rect 430654 154046 430722 154102
rect 430778 154046 430848 154102
rect 430528 153978 430848 154046
rect 430528 153922 430598 153978
rect 430654 153922 430722 153978
rect 430778 153922 430848 153978
rect 430528 153888 430848 153922
rect 384448 148350 384768 148384
rect 384448 148294 384518 148350
rect 384574 148294 384642 148350
rect 384698 148294 384768 148350
rect 384448 148226 384768 148294
rect 384448 148170 384518 148226
rect 384574 148170 384642 148226
rect 384698 148170 384768 148226
rect 384448 148102 384768 148170
rect 384448 148046 384518 148102
rect 384574 148046 384642 148102
rect 384698 148046 384768 148102
rect 384448 147978 384768 148046
rect 384448 147922 384518 147978
rect 384574 147922 384642 147978
rect 384698 147922 384768 147978
rect 384448 147888 384768 147922
rect 415168 148350 415488 148384
rect 415168 148294 415238 148350
rect 415294 148294 415362 148350
rect 415418 148294 415488 148350
rect 415168 148226 415488 148294
rect 415168 148170 415238 148226
rect 415294 148170 415362 148226
rect 415418 148170 415488 148226
rect 415168 148102 415488 148170
rect 415168 148046 415238 148102
rect 415294 148046 415362 148102
rect 415418 148046 415488 148102
rect 415168 147978 415488 148046
rect 415168 147922 415238 147978
rect 415294 147922 415362 147978
rect 415418 147922 415488 147978
rect 415168 147888 415488 147922
rect 396844 137396 396900 137406
rect 393932 137172 393988 137182
rect 383628 135650 383684 135660
rect 385420 136724 385476 136734
rect 385420 135716 385476 136668
rect 385420 135650 385476 135660
rect 387212 136612 387268 136622
rect 385532 135604 385588 135614
rect 384748 135268 384804 135278
rect 382284 124002 382340 124012
rect 383180 78988 383236 132524
rect 384524 132692 384580 132702
rect 384524 125524 384580 132636
rect 384748 128996 384804 135212
rect 385532 135268 385588 135548
rect 385532 135202 385588 135212
rect 385756 135604 385812 135614
rect 385756 135156 385812 135548
rect 385756 135090 385812 135100
rect 385532 134708 385588 134718
rect 384748 128930 384804 128940
rect 384972 132580 385028 132590
rect 384524 125458 384580 125468
rect 384448 112350 384768 112384
rect 384448 112294 384518 112350
rect 384574 112294 384642 112350
rect 384698 112294 384768 112350
rect 384448 112226 384768 112294
rect 384448 112170 384518 112226
rect 384574 112170 384642 112226
rect 384698 112170 384768 112226
rect 384448 112102 384768 112170
rect 384448 112046 384518 112102
rect 384574 112046 384642 112102
rect 384698 112046 384768 112102
rect 384448 111978 384768 112046
rect 384448 111922 384518 111978
rect 384574 111922 384642 111978
rect 384698 111922 384768 111978
rect 384448 111888 384768 111922
rect 384448 94350 384768 94384
rect 384448 94294 384518 94350
rect 384574 94294 384642 94350
rect 384698 94294 384768 94350
rect 384448 94226 384768 94294
rect 384448 94170 384518 94226
rect 384574 94170 384642 94226
rect 384698 94170 384768 94226
rect 384448 94102 384768 94170
rect 384448 94046 384518 94102
rect 384574 94046 384642 94102
rect 384698 94046 384768 94102
rect 384448 93978 384768 94046
rect 384448 93922 384518 93978
rect 384574 93922 384642 93978
rect 384698 93922 384768 93978
rect 384448 93888 384768 93922
rect 381836 55468 381892 72782
rect 381612 55412 381892 55468
rect 383068 78932 383236 78988
rect 383068 76618 383124 78932
rect 381612 45780 381668 55412
rect 381612 45714 381668 45724
rect 383068 45780 383124 76562
rect 384972 78418 385028 132524
rect 384448 76350 384768 76384
rect 384448 76294 384518 76350
rect 384574 76294 384642 76350
rect 384698 76294 384768 76350
rect 384448 76226 384768 76294
rect 384448 76170 384518 76226
rect 384574 76170 384642 76226
rect 384698 76170 384768 76226
rect 384448 76102 384768 76170
rect 384448 76046 384518 76102
rect 384574 76046 384642 76102
rect 384698 76046 384768 76102
rect 384448 75978 384768 76046
rect 384448 75922 384518 75978
rect 384574 75922 384642 75978
rect 384698 75922 384768 75978
rect 384448 75888 384768 75922
rect 383068 45714 383124 45724
rect 383852 74098 383908 74108
rect 381500 45490 381556 45500
rect 383852 45556 383908 74042
rect 384448 58350 384768 58384
rect 384448 58294 384518 58350
rect 384574 58294 384642 58350
rect 384698 58294 384768 58350
rect 384448 58226 384768 58294
rect 384448 58170 384518 58226
rect 384574 58170 384642 58226
rect 384698 58170 384768 58226
rect 384448 58102 384768 58170
rect 384448 58046 384518 58102
rect 384574 58046 384642 58102
rect 384698 58046 384768 58102
rect 384448 57978 384768 58046
rect 384448 57922 384518 57978
rect 384574 57922 384642 57978
rect 384698 57922 384768 57978
rect 384448 57888 384768 57922
rect 383852 45490 383908 45500
rect 384972 45556 385028 78362
rect 385532 45892 385588 134652
rect 385644 132580 385700 132590
rect 385644 80578 385700 132524
rect 386540 132580 386596 132590
rect 385644 80512 385700 80522
rect 386428 131684 386484 131694
rect 386428 80758 386484 131628
rect 385532 45826 385588 45836
rect 385644 78058 385700 78068
rect 385644 45780 385700 78002
rect 385644 45714 385700 45724
rect 384972 45490 385028 45500
rect 386428 45556 386484 80702
rect 386540 81658 386596 132524
rect 386540 78988 386596 81602
rect 386540 78932 387044 78988
rect 386428 45490 386484 45500
rect 386988 45556 387044 78932
rect 386988 45490 387044 45500
rect 380604 44930 380660 44940
rect 385756 44436 385812 44446
rect 385756 44212 385812 44380
rect 385756 44146 385812 44156
rect 387212 41748 387268 136556
rect 388108 135828 388164 135838
rect 388108 64738 388164 135772
rect 390572 132804 390628 132814
rect 390572 132356 390628 132748
rect 390572 132290 390628 132300
rect 390796 132356 390852 132366
rect 390796 131796 390852 132300
rect 390796 131730 390852 131740
rect 392252 131572 392308 131582
rect 388220 131460 388276 131470
rect 388220 67228 388276 131404
rect 389788 129220 389844 129230
rect 388332 128884 388388 128894
rect 388332 71398 388388 128828
rect 388332 71332 388388 71342
rect 388220 67172 388388 67228
rect 388108 45444 388164 64682
rect 388332 64918 388388 67172
rect 388332 45556 388388 64862
rect 389788 62938 389844 129164
rect 390012 128996 390068 129006
rect 389788 45780 389844 62882
rect 389788 45714 389844 45724
rect 389900 80578 389956 80588
rect 388332 45490 388388 45500
rect 388108 45378 388164 45388
rect 389900 45220 389956 80522
rect 390012 78058 390068 128940
rect 390012 77992 390068 78002
rect 390572 124068 390628 124078
rect 389900 45154 389956 45164
rect 390572 43428 390628 124012
rect 391468 100918 391524 100928
rect 391468 45556 391524 100862
rect 391468 45490 391524 45500
rect 392252 45220 392308 131516
rect 392476 128996 392532 129006
rect 392364 125412 392420 125422
rect 392364 105778 392420 125356
rect 392364 105712 392420 105722
rect 392476 100918 392532 128940
rect 392476 100852 392532 100862
rect 393148 125524 393204 125534
rect 393148 74098 393204 125468
rect 393148 74032 393204 74042
rect 393820 46004 393876 46014
rect 393820 45556 393876 45948
rect 393820 45490 393876 45500
rect 392252 45154 392308 45164
rect 390572 43362 390628 43372
rect 393932 43316 393988 137116
rect 396844 136164 396900 137340
rect 396844 136098 396900 136108
rect 397516 137284 397572 137294
rect 397516 136276 397572 137228
rect 395724 135940 395780 135950
rect 394044 133476 394100 133486
rect 394044 48020 394100 133420
rect 394044 47954 394100 47964
rect 394156 91558 394212 91568
rect 394156 43540 394212 91502
rect 394828 52138 394884 52148
rect 394828 47012 394884 52082
rect 394828 46946 394884 46956
rect 395724 45220 395780 135884
rect 397516 135716 397572 136220
rect 397516 135650 397572 135660
rect 408044 137284 408100 137294
rect 408044 136276 408100 137228
rect 398188 131124 398244 131134
rect 395724 45154 395780 45164
rect 395836 131012 395892 131022
rect 395836 43652 395892 130956
rect 395836 43586 395892 43596
rect 396396 116038 396452 116048
rect 394156 43474 394212 43484
rect 393932 43250 393988 43260
rect 396396 42980 396452 115982
rect 398188 116038 398244 131068
rect 408044 127092 408100 136220
rect 408156 137172 408212 137182
rect 408156 136164 408212 137116
rect 408156 128884 408212 136108
rect 408156 128818 408212 128828
rect 408498 136350 409118 136602
rect 408498 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 409118 136350
rect 408498 136226 409118 136294
rect 408498 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 409118 136226
rect 408498 136102 409118 136170
rect 408498 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 409118 136102
rect 408498 135978 409118 136046
rect 408498 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 409118 135978
rect 408044 127026 408100 127036
rect 399808 118350 400128 118384
rect 399808 118294 399878 118350
rect 399934 118294 400002 118350
rect 400058 118294 400128 118350
rect 399808 118226 400128 118294
rect 399808 118170 399878 118226
rect 399934 118170 400002 118226
rect 400058 118170 400128 118226
rect 399808 118102 400128 118170
rect 399808 118046 399878 118102
rect 399934 118046 400002 118102
rect 400058 118046 400128 118102
rect 399808 117978 400128 118046
rect 399808 117922 399878 117978
rect 399934 117922 400002 117978
rect 400058 117922 400128 117978
rect 399808 117888 400128 117922
rect 408498 118350 409118 135922
rect 431788 132132 431844 204204
rect 432124 204058 432180 324492
rect 433468 278908 433524 326060
rect 435498 310350 436118 327922
rect 439218 598172 439838 598268
rect 439218 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 439838 598172
rect 439218 598048 439838 598116
rect 439218 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 439838 598048
rect 439218 597924 439838 597992
rect 439218 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 439838 597924
rect 439218 597800 439838 597868
rect 439218 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 439838 597800
rect 439218 586350 439838 597744
rect 439218 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 439838 586350
rect 439218 586226 439838 586294
rect 439218 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 439838 586226
rect 439218 586102 439838 586170
rect 439218 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 439838 586102
rect 439218 585978 439838 586046
rect 439218 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 439838 585978
rect 439218 568350 439838 585922
rect 439218 568294 439314 568350
rect 439370 568294 439438 568350
rect 439494 568294 439562 568350
rect 439618 568294 439686 568350
rect 439742 568294 439838 568350
rect 439218 568226 439838 568294
rect 439218 568170 439314 568226
rect 439370 568170 439438 568226
rect 439494 568170 439562 568226
rect 439618 568170 439686 568226
rect 439742 568170 439838 568226
rect 439218 568102 439838 568170
rect 439218 568046 439314 568102
rect 439370 568046 439438 568102
rect 439494 568046 439562 568102
rect 439618 568046 439686 568102
rect 439742 568046 439838 568102
rect 439218 567978 439838 568046
rect 439218 567922 439314 567978
rect 439370 567922 439438 567978
rect 439494 567922 439562 567978
rect 439618 567922 439686 567978
rect 439742 567922 439838 567978
rect 439218 550350 439838 567922
rect 439218 550294 439314 550350
rect 439370 550294 439438 550350
rect 439494 550294 439562 550350
rect 439618 550294 439686 550350
rect 439742 550294 439838 550350
rect 439218 550226 439838 550294
rect 439218 550170 439314 550226
rect 439370 550170 439438 550226
rect 439494 550170 439562 550226
rect 439618 550170 439686 550226
rect 439742 550170 439838 550226
rect 439218 550102 439838 550170
rect 439218 550046 439314 550102
rect 439370 550046 439438 550102
rect 439494 550046 439562 550102
rect 439618 550046 439686 550102
rect 439742 550046 439838 550102
rect 439218 549978 439838 550046
rect 439218 549922 439314 549978
rect 439370 549922 439438 549978
rect 439494 549922 439562 549978
rect 439618 549922 439686 549978
rect 439742 549922 439838 549978
rect 439218 532350 439838 549922
rect 439218 532294 439314 532350
rect 439370 532294 439438 532350
rect 439494 532294 439562 532350
rect 439618 532294 439686 532350
rect 439742 532294 439838 532350
rect 439218 532226 439838 532294
rect 439218 532170 439314 532226
rect 439370 532170 439438 532226
rect 439494 532170 439562 532226
rect 439618 532170 439686 532226
rect 439742 532170 439838 532226
rect 439218 532102 439838 532170
rect 439218 532046 439314 532102
rect 439370 532046 439438 532102
rect 439494 532046 439562 532102
rect 439618 532046 439686 532102
rect 439742 532046 439838 532102
rect 439218 531978 439838 532046
rect 439218 531922 439314 531978
rect 439370 531922 439438 531978
rect 439494 531922 439562 531978
rect 439618 531922 439686 531978
rect 439742 531922 439838 531978
rect 439218 514350 439838 531922
rect 439218 514294 439314 514350
rect 439370 514294 439438 514350
rect 439494 514294 439562 514350
rect 439618 514294 439686 514350
rect 439742 514294 439838 514350
rect 439218 514226 439838 514294
rect 439218 514170 439314 514226
rect 439370 514170 439438 514226
rect 439494 514170 439562 514226
rect 439618 514170 439686 514226
rect 439742 514170 439838 514226
rect 439218 514102 439838 514170
rect 439218 514046 439314 514102
rect 439370 514046 439438 514102
rect 439494 514046 439562 514102
rect 439618 514046 439686 514102
rect 439742 514046 439838 514102
rect 439218 513978 439838 514046
rect 439218 513922 439314 513978
rect 439370 513922 439438 513978
rect 439494 513922 439562 513978
rect 439618 513922 439686 513978
rect 439742 513922 439838 513978
rect 439218 496350 439838 513922
rect 439218 496294 439314 496350
rect 439370 496294 439438 496350
rect 439494 496294 439562 496350
rect 439618 496294 439686 496350
rect 439742 496294 439838 496350
rect 439218 496226 439838 496294
rect 439218 496170 439314 496226
rect 439370 496170 439438 496226
rect 439494 496170 439562 496226
rect 439618 496170 439686 496226
rect 439742 496170 439838 496226
rect 439218 496102 439838 496170
rect 439218 496046 439314 496102
rect 439370 496046 439438 496102
rect 439494 496046 439562 496102
rect 439618 496046 439686 496102
rect 439742 496046 439838 496102
rect 439218 495978 439838 496046
rect 439218 495922 439314 495978
rect 439370 495922 439438 495978
rect 439494 495922 439562 495978
rect 439618 495922 439686 495978
rect 439742 495922 439838 495978
rect 439218 478350 439838 495922
rect 439218 478294 439314 478350
rect 439370 478294 439438 478350
rect 439494 478294 439562 478350
rect 439618 478294 439686 478350
rect 439742 478294 439838 478350
rect 439218 478226 439838 478294
rect 439218 478170 439314 478226
rect 439370 478170 439438 478226
rect 439494 478170 439562 478226
rect 439618 478170 439686 478226
rect 439742 478170 439838 478226
rect 439218 478102 439838 478170
rect 439218 478046 439314 478102
rect 439370 478046 439438 478102
rect 439494 478046 439562 478102
rect 439618 478046 439686 478102
rect 439742 478046 439838 478102
rect 439218 477978 439838 478046
rect 439218 477922 439314 477978
rect 439370 477922 439438 477978
rect 439494 477922 439562 477978
rect 439618 477922 439686 477978
rect 439742 477922 439838 477978
rect 439218 460350 439838 477922
rect 439218 460294 439314 460350
rect 439370 460294 439438 460350
rect 439494 460294 439562 460350
rect 439618 460294 439686 460350
rect 439742 460294 439838 460350
rect 439218 460226 439838 460294
rect 439218 460170 439314 460226
rect 439370 460170 439438 460226
rect 439494 460170 439562 460226
rect 439618 460170 439686 460226
rect 439742 460170 439838 460226
rect 439218 460102 439838 460170
rect 439218 460046 439314 460102
rect 439370 460046 439438 460102
rect 439494 460046 439562 460102
rect 439618 460046 439686 460102
rect 439742 460046 439838 460102
rect 439218 459978 439838 460046
rect 439218 459922 439314 459978
rect 439370 459922 439438 459978
rect 439494 459922 439562 459978
rect 439618 459922 439686 459978
rect 439742 459922 439838 459978
rect 439218 442350 439838 459922
rect 439218 442294 439314 442350
rect 439370 442294 439438 442350
rect 439494 442294 439562 442350
rect 439618 442294 439686 442350
rect 439742 442294 439838 442350
rect 439218 442226 439838 442294
rect 439218 442170 439314 442226
rect 439370 442170 439438 442226
rect 439494 442170 439562 442226
rect 439618 442170 439686 442226
rect 439742 442170 439838 442226
rect 439218 442102 439838 442170
rect 439218 442046 439314 442102
rect 439370 442046 439438 442102
rect 439494 442046 439562 442102
rect 439618 442046 439686 442102
rect 439742 442046 439838 442102
rect 439218 441978 439838 442046
rect 439218 441922 439314 441978
rect 439370 441922 439438 441978
rect 439494 441922 439562 441978
rect 439618 441922 439686 441978
rect 439742 441922 439838 441978
rect 439218 424350 439838 441922
rect 439218 424294 439314 424350
rect 439370 424294 439438 424350
rect 439494 424294 439562 424350
rect 439618 424294 439686 424350
rect 439742 424294 439838 424350
rect 439218 424226 439838 424294
rect 439218 424170 439314 424226
rect 439370 424170 439438 424226
rect 439494 424170 439562 424226
rect 439618 424170 439686 424226
rect 439742 424170 439838 424226
rect 439218 424102 439838 424170
rect 439218 424046 439314 424102
rect 439370 424046 439438 424102
rect 439494 424046 439562 424102
rect 439618 424046 439686 424102
rect 439742 424046 439838 424102
rect 439218 423978 439838 424046
rect 439218 423922 439314 423978
rect 439370 423922 439438 423978
rect 439494 423922 439562 423978
rect 439618 423922 439686 423978
rect 439742 423922 439838 423978
rect 439218 406350 439838 423922
rect 439218 406294 439314 406350
rect 439370 406294 439438 406350
rect 439494 406294 439562 406350
rect 439618 406294 439686 406350
rect 439742 406294 439838 406350
rect 439218 406226 439838 406294
rect 439218 406170 439314 406226
rect 439370 406170 439438 406226
rect 439494 406170 439562 406226
rect 439618 406170 439686 406226
rect 439742 406170 439838 406226
rect 439218 406102 439838 406170
rect 439218 406046 439314 406102
rect 439370 406046 439438 406102
rect 439494 406046 439562 406102
rect 439618 406046 439686 406102
rect 439742 406046 439838 406102
rect 439218 405978 439838 406046
rect 439218 405922 439314 405978
rect 439370 405922 439438 405978
rect 439494 405922 439562 405978
rect 439618 405922 439686 405978
rect 439742 405922 439838 405978
rect 439218 388350 439838 405922
rect 439218 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 439838 388350
rect 439218 388226 439838 388294
rect 439218 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 439838 388226
rect 439218 388102 439838 388170
rect 439218 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 439838 388102
rect 439218 387978 439838 388046
rect 439218 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 439838 387978
rect 439218 370350 439838 387922
rect 439218 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 439838 370350
rect 439218 370226 439838 370294
rect 439218 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 439838 370226
rect 439218 370102 439838 370170
rect 439218 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 439838 370102
rect 439218 369978 439838 370046
rect 439218 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 439838 369978
rect 439218 352350 439838 369922
rect 439218 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 439838 352350
rect 439218 352226 439838 352294
rect 439218 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 439838 352226
rect 439218 352102 439838 352170
rect 439218 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 439838 352102
rect 439218 351978 439838 352046
rect 439218 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 439838 351978
rect 439218 334350 439838 351922
rect 439218 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 439838 334350
rect 439218 334226 439838 334294
rect 439218 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 439838 334226
rect 439218 334102 439838 334170
rect 439218 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 439838 334102
rect 439218 333978 439838 334046
rect 439218 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 439838 333978
rect 435498 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 436118 310350
rect 435498 310226 436118 310294
rect 435498 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 436118 310226
rect 435498 310102 436118 310170
rect 435498 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 436118 310102
rect 435498 309978 436118 310046
rect 435498 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 436118 309978
rect 435498 292350 436118 309922
rect 435498 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 436118 292350
rect 435498 292226 436118 292294
rect 435498 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 436118 292226
rect 435498 292102 436118 292170
rect 435498 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 436118 292102
rect 435498 291978 436118 292046
rect 435498 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 436118 291978
rect 433468 278852 433636 278908
rect 432124 203992 432180 204002
rect 433468 264516 433524 264526
rect 431788 132066 431844 132076
rect 431900 201684 431956 201694
rect 431900 132020 431956 201628
rect 432012 199668 432068 199678
rect 432012 132244 432068 199612
rect 433468 192500 433524 264460
rect 433580 263060 433636 278852
rect 435498 274350 436118 291922
rect 435498 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 436118 274350
rect 435498 274226 436118 274294
rect 435498 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 436118 274226
rect 435498 274102 436118 274170
rect 435498 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 436118 274102
rect 435498 273978 436118 274046
rect 435498 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 436118 273978
rect 433580 262994 433636 263004
rect 434252 263732 434308 263742
rect 434252 240058 434308 263676
rect 433468 192434 433524 192444
rect 433580 202692 433636 202702
rect 433580 132356 433636 202636
rect 433692 202468 433748 202478
rect 433692 132692 433748 202412
rect 434252 197428 434308 240002
rect 434252 197362 434308 197372
rect 435498 256350 436118 273922
rect 435498 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 436118 256350
rect 435498 256226 436118 256294
rect 435498 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 436118 256226
rect 435498 256102 436118 256170
rect 435498 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 436118 256102
rect 435498 255978 436118 256046
rect 435498 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 436118 255978
rect 435498 238350 436118 255922
rect 436828 323428 436884 323438
rect 436828 242758 436884 323372
rect 436828 242692 436884 242702
rect 439218 316350 439838 333922
rect 466218 597212 466838 598268
rect 466218 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 466838 597212
rect 466218 597088 466838 597156
rect 466218 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 466838 597088
rect 466218 596964 466838 597032
rect 466218 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 466838 596964
rect 466218 596840 466838 596908
rect 466218 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 466838 596840
rect 466218 580350 466838 596784
rect 466218 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 466838 580350
rect 466218 580226 466838 580294
rect 466218 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 466838 580226
rect 466218 580102 466838 580170
rect 466218 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 466838 580102
rect 466218 579978 466838 580046
rect 466218 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 466838 579978
rect 466218 562350 466838 579922
rect 466218 562294 466314 562350
rect 466370 562294 466438 562350
rect 466494 562294 466562 562350
rect 466618 562294 466686 562350
rect 466742 562294 466838 562350
rect 466218 562226 466838 562294
rect 466218 562170 466314 562226
rect 466370 562170 466438 562226
rect 466494 562170 466562 562226
rect 466618 562170 466686 562226
rect 466742 562170 466838 562226
rect 466218 562102 466838 562170
rect 466218 562046 466314 562102
rect 466370 562046 466438 562102
rect 466494 562046 466562 562102
rect 466618 562046 466686 562102
rect 466742 562046 466838 562102
rect 466218 561978 466838 562046
rect 466218 561922 466314 561978
rect 466370 561922 466438 561978
rect 466494 561922 466562 561978
rect 466618 561922 466686 561978
rect 466742 561922 466838 561978
rect 466218 544350 466838 561922
rect 466218 544294 466314 544350
rect 466370 544294 466438 544350
rect 466494 544294 466562 544350
rect 466618 544294 466686 544350
rect 466742 544294 466838 544350
rect 466218 544226 466838 544294
rect 466218 544170 466314 544226
rect 466370 544170 466438 544226
rect 466494 544170 466562 544226
rect 466618 544170 466686 544226
rect 466742 544170 466838 544226
rect 466218 544102 466838 544170
rect 466218 544046 466314 544102
rect 466370 544046 466438 544102
rect 466494 544046 466562 544102
rect 466618 544046 466686 544102
rect 466742 544046 466838 544102
rect 466218 543978 466838 544046
rect 466218 543922 466314 543978
rect 466370 543922 466438 543978
rect 466494 543922 466562 543978
rect 466618 543922 466686 543978
rect 466742 543922 466838 543978
rect 466218 526350 466838 543922
rect 466218 526294 466314 526350
rect 466370 526294 466438 526350
rect 466494 526294 466562 526350
rect 466618 526294 466686 526350
rect 466742 526294 466838 526350
rect 466218 526226 466838 526294
rect 466218 526170 466314 526226
rect 466370 526170 466438 526226
rect 466494 526170 466562 526226
rect 466618 526170 466686 526226
rect 466742 526170 466838 526226
rect 466218 526102 466838 526170
rect 466218 526046 466314 526102
rect 466370 526046 466438 526102
rect 466494 526046 466562 526102
rect 466618 526046 466686 526102
rect 466742 526046 466838 526102
rect 466218 525978 466838 526046
rect 466218 525922 466314 525978
rect 466370 525922 466438 525978
rect 466494 525922 466562 525978
rect 466618 525922 466686 525978
rect 466742 525922 466838 525978
rect 466218 508350 466838 525922
rect 466218 508294 466314 508350
rect 466370 508294 466438 508350
rect 466494 508294 466562 508350
rect 466618 508294 466686 508350
rect 466742 508294 466838 508350
rect 466218 508226 466838 508294
rect 466218 508170 466314 508226
rect 466370 508170 466438 508226
rect 466494 508170 466562 508226
rect 466618 508170 466686 508226
rect 466742 508170 466838 508226
rect 466218 508102 466838 508170
rect 466218 508046 466314 508102
rect 466370 508046 466438 508102
rect 466494 508046 466562 508102
rect 466618 508046 466686 508102
rect 466742 508046 466838 508102
rect 466218 507978 466838 508046
rect 466218 507922 466314 507978
rect 466370 507922 466438 507978
rect 466494 507922 466562 507978
rect 466618 507922 466686 507978
rect 466742 507922 466838 507978
rect 466218 490350 466838 507922
rect 466218 490294 466314 490350
rect 466370 490294 466438 490350
rect 466494 490294 466562 490350
rect 466618 490294 466686 490350
rect 466742 490294 466838 490350
rect 466218 490226 466838 490294
rect 466218 490170 466314 490226
rect 466370 490170 466438 490226
rect 466494 490170 466562 490226
rect 466618 490170 466686 490226
rect 466742 490170 466838 490226
rect 466218 490102 466838 490170
rect 466218 490046 466314 490102
rect 466370 490046 466438 490102
rect 466494 490046 466562 490102
rect 466618 490046 466686 490102
rect 466742 490046 466838 490102
rect 466218 489978 466838 490046
rect 466218 489922 466314 489978
rect 466370 489922 466438 489978
rect 466494 489922 466562 489978
rect 466618 489922 466686 489978
rect 466742 489922 466838 489978
rect 466218 472350 466838 489922
rect 466218 472294 466314 472350
rect 466370 472294 466438 472350
rect 466494 472294 466562 472350
rect 466618 472294 466686 472350
rect 466742 472294 466838 472350
rect 466218 472226 466838 472294
rect 466218 472170 466314 472226
rect 466370 472170 466438 472226
rect 466494 472170 466562 472226
rect 466618 472170 466686 472226
rect 466742 472170 466838 472226
rect 466218 472102 466838 472170
rect 466218 472046 466314 472102
rect 466370 472046 466438 472102
rect 466494 472046 466562 472102
rect 466618 472046 466686 472102
rect 466742 472046 466838 472102
rect 466218 471978 466838 472046
rect 466218 471922 466314 471978
rect 466370 471922 466438 471978
rect 466494 471922 466562 471978
rect 466618 471922 466686 471978
rect 466742 471922 466838 471978
rect 466218 454350 466838 471922
rect 466218 454294 466314 454350
rect 466370 454294 466438 454350
rect 466494 454294 466562 454350
rect 466618 454294 466686 454350
rect 466742 454294 466838 454350
rect 466218 454226 466838 454294
rect 466218 454170 466314 454226
rect 466370 454170 466438 454226
rect 466494 454170 466562 454226
rect 466618 454170 466686 454226
rect 466742 454170 466838 454226
rect 466218 454102 466838 454170
rect 466218 454046 466314 454102
rect 466370 454046 466438 454102
rect 466494 454046 466562 454102
rect 466618 454046 466686 454102
rect 466742 454046 466838 454102
rect 466218 453978 466838 454046
rect 466218 453922 466314 453978
rect 466370 453922 466438 453978
rect 466494 453922 466562 453978
rect 466618 453922 466686 453978
rect 466742 453922 466838 453978
rect 466218 436350 466838 453922
rect 466218 436294 466314 436350
rect 466370 436294 466438 436350
rect 466494 436294 466562 436350
rect 466618 436294 466686 436350
rect 466742 436294 466838 436350
rect 466218 436226 466838 436294
rect 466218 436170 466314 436226
rect 466370 436170 466438 436226
rect 466494 436170 466562 436226
rect 466618 436170 466686 436226
rect 466742 436170 466838 436226
rect 466218 436102 466838 436170
rect 466218 436046 466314 436102
rect 466370 436046 466438 436102
rect 466494 436046 466562 436102
rect 466618 436046 466686 436102
rect 466742 436046 466838 436102
rect 466218 435978 466838 436046
rect 466218 435922 466314 435978
rect 466370 435922 466438 435978
rect 466494 435922 466562 435978
rect 466618 435922 466686 435978
rect 466742 435922 466838 435978
rect 466218 418350 466838 435922
rect 466218 418294 466314 418350
rect 466370 418294 466438 418350
rect 466494 418294 466562 418350
rect 466618 418294 466686 418350
rect 466742 418294 466838 418350
rect 466218 418226 466838 418294
rect 466218 418170 466314 418226
rect 466370 418170 466438 418226
rect 466494 418170 466562 418226
rect 466618 418170 466686 418226
rect 466742 418170 466838 418226
rect 466218 418102 466838 418170
rect 466218 418046 466314 418102
rect 466370 418046 466438 418102
rect 466494 418046 466562 418102
rect 466618 418046 466686 418102
rect 466742 418046 466838 418102
rect 466218 417978 466838 418046
rect 466218 417922 466314 417978
rect 466370 417922 466438 417978
rect 466494 417922 466562 417978
rect 466618 417922 466686 417978
rect 466742 417922 466838 417978
rect 466218 400350 466838 417922
rect 466218 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 466838 400350
rect 466218 400226 466838 400294
rect 466218 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 466838 400226
rect 466218 400102 466838 400170
rect 466218 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 466838 400102
rect 466218 399978 466838 400046
rect 466218 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 466838 399978
rect 466218 382350 466838 399922
rect 466218 382294 466314 382350
rect 466370 382294 466438 382350
rect 466494 382294 466562 382350
rect 466618 382294 466686 382350
rect 466742 382294 466838 382350
rect 466218 382226 466838 382294
rect 466218 382170 466314 382226
rect 466370 382170 466438 382226
rect 466494 382170 466562 382226
rect 466618 382170 466686 382226
rect 466742 382170 466838 382226
rect 466218 382102 466838 382170
rect 466218 382046 466314 382102
rect 466370 382046 466438 382102
rect 466494 382046 466562 382102
rect 466618 382046 466686 382102
rect 466742 382046 466838 382102
rect 466218 381978 466838 382046
rect 466218 381922 466314 381978
rect 466370 381922 466438 381978
rect 466494 381922 466562 381978
rect 466618 381922 466686 381978
rect 466742 381922 466838 381978
rect 466218 364350 466838 381922
rect 466218 364294 466314 364350
rect 466370 364294 466438 364350
rect 466494 364294 466562 364350
rect 466618 364294 466686 364350
rect 466742 364294 466838 364350
rect 466218 364226 466838 364294
rect 466218 364170 466314 364226
rect 466370 364170 466438 364226
rect 466494 364170 466562 364226
rect 466618 364170 466686 364226
rect 466742 364170 466838 364226
rect 466218 364102 466838 364170
rect 466218 364046 466314 364102
rect 466370 364046 466438 364102
rect 466494 364046 466562 364102
rect 466618 364046 466686 364102
rect 466742 364046 466838 364102
rect 466218 363978 466838 364046
rect 466218 363922 466314 363978
rect 466370 363922 466438 363978
rect 466494 363922 466562 363978
rect 466618 363922 466686 363978
rect 466742 363922 466838 363978
rect 466218 346350 466838 363922
rect 466218 346294 466314 346350
rect 466370 346294 466438 346350
rect 466494 346294 466562 346350
rect 466618 346294 466686 346350
rect 466742 346294 466838 346350
rect 466218 346226 466838 346294
rect 466218 346170 466314 346226
rect 466370 346170 466438 346226
rect 466494 346170 466562 346226
rect 466618 346170 466686 346226
rect 466742 346170 466838 346226
rect 466218 346102 466838 346170
rect 466218 346046 466314 346102
rect 466370 346046 466438 346102
rect 466494 346046 466562 346102
rect 466618 346046 466686 346102
rect 466742 346046 466838 346102
rect 466218 345978 466838 346046
rect 466218 345922 466314 345978
rect 466370 345922 466438 345978
rect 466494 345922 466562 345978
rect 466618 345922 466686 345978
rect 466742 345922 466838 345978
rect 466218 328350 466838 345922
rect 466218 328294 466314 328350
rect 466370 328294 466438 328350
rect 466494 328294 466562 328350
rect 466618 328294 466686 328350
rect 466742 328294 466838 328350
rect 466218 328226 466838 328294
rect 466218 328170 466314 328226
rect 466370 328170 466438 328226
rect 466494 328170 466562 328226
rect 466618 328170 466686 328226
rect 466742 328170 466838 328226
rect 466218 328102 466838 328170
rect 466218 328046 466314 328102
rect 466370 328046 466438 328102
rect 466494 328046 466562 328102
rect 466618 328046 466686 328102
rect 466742 328046 466838 328102
rect 466218 327978 466838 328046
rect 466218 327922 466314 327978
rect 466370 327922 466438 327978
rect 466494 327922 466562 327978
rect 466618 327922 466686 327978
rect 466742 327922 466838 327978
rect 442092 324884 442148 324894
rect 441868 324772 441924 324782
rect 440300 324660 440356 324670
rect 439218 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 439838 316350
rect 439218 316226 439838 316294
rect 439218 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 439838 316226
rect 439218 316102 439838 316170
rect 439218 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 439838 316102
rect 439218 315978 439838 316046
rect 439218 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 439838 315978
rect 439218 298350 439838 315922
rect 439218 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 439838 298350
rect 439218 298226 439838 298294
rect 439218 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 439838 298226
rect 439218 298102 439838 298170
rect 439218 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 439838 298102
rect 439218 297978 439838 298046
rect 439218 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 439838 297978
rect 439218 280350 439838 297922
rect 440188 322644 440244 322654
rect 440188 294532 440244 322588
rect 440300 301252 440356 324604
rect 440300 301186 440356 301196
rect 440412 322756 440468 322766
rect 440412 299908 440468 322700
rect 441868 312004 441924 324716
rect 441868 311938 441924 311948
rect 441980 322868 442036 322878
rect 440412 299842 440468 299852
rect 440524 310978 440580 310988
rect 440524 296548 440580 310922
rect 440860 305284 440916 305294
rect 440524 296482 440580 296492
rect 440636 297220 440692 297230
rect 440188 294466 440244 294476
rect 440524 293860 440580 293870
rect 440300 293188 440356 293198
rect 439218 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 439838 280350
rect 439218 280226 439838 280294
rect 439218 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 439838 280226
rect 439218 280102 439838 280170
rect 439218 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 439838 280102
rect 439218 279978 439838 280046
rect 439218 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 439838 279978
rect 439218 262350 439838 279922
rect 440188 292516 440244 292526
rect 440188 275156 440244 292460
rect 440300 277060 440356 293132
rect 440300 276994 440356 277004
rect 440188 275090 440244 275100
rect 440524 273700 440580 293804
rect 440636 276948 440692 297164
rect 440636 276882 440692 276892
rect 440748 290500 440804 290510
rect 440748 275492 440804 290444
rect 440748 275426 440804 275436
rect 440524 273634 440580 273644
rect 440412 268884 440468 268894
rect 439218 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 439838 262350
rect 439218 262226 439838 262294
rect 439218 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 439838 262226
rect 439218 262102 439838 262170
rect 439218 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 439838 262102
rect 439218 261978 439838 262046
rect 439218 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 439838 261978
rect 439218 244350 439838 261922
rect 439218 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 439838 244350
rect 439218 244226 439838 244294
rect 439218 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 439838 244226
rect 439218 244102 439838 244170
rect 439218 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 439838 244102
rect 439218 243978 439838 244046
rect 439218 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 439838 243978
rect 435498 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 436118 238350
rect 435498 238226 436118 238294
rect 435498 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 436118 238226
rect 435498 238102 436118 238170
rect 435498 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 436118 238102
rect 435498 237978 436118 238046
rect 435498 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 436118 237978
rect 435498 220350 436118 237922
rect 435498 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 436118 220350
rect 435498 220226 436118 220294
rect 435498 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 436118 220226
rect 435498 220102 436118 220170
rect 435498 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 436118 220102
rect 435498 219978 436118 220046
rect 435498 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 436118 219978
rect 435498 202350 436118 219922
rect 435498 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 436118 202350
rect 435498 202226 436118 202294
rect 435498 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 436118 202226
rect 435498 202102 436118 202170
rect 435498 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 436118 202102
rect 435498 201978 436118 202046
rect 435498 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 436118 201978
rect 433692 132626 433748 132636
rect 435498 184350 436118 201922
rect 439218 226350 439838 243922
rect 440300 266756 440356 266766
rect 440188 242758 440244 242768
rect 440188 242004 440244 242702
rect 440188 241938 440244 241948
rect 439964 240058 440020 240068
rect 439964 239876 440020 240002
rect 439964 239810 440020 239820
rect 440300 235956 440356 266700
rect 440412 240660 440468 268828
rect 440412 240594 440468 240604
rect 440524 266420 440580 266430
rect 440300 235890 440356 235900
rect 440524 231924 440580 266364
rect 440860 262948 440916 305228
rect 441980 303268 442036 322812
rect 441980 303202 442036 303212
rect 441084 302596 441140 302606
rect 440972 301924 441028 301934
rect 440972 266308 441028 301868
rect 441084 269668 441140 302540
rect 442092 298564 442148 324828
rect 442316 323092 442372 323102
rect 442204 322980 442260 322990
rect 442204 303940 442260 322924
rect 442204 303874 442260 303884
rect 442092 298498 442148 298508
rect 442204 300580 442260 300590
rect 441868 295876 441924 295886
rect 441868 277172 441924 295820
rect 441868 277106 441924 277116
rect 441980 291844 442036 291854
rect 441980 275380 442036 291788
rect 442092 289828 442148 289838
rect 442092 276612 442148 289772
rect 442204 276836 442260 300524
rect 442316 299236 442372 323036
rect 443548 312676 443604 312686
rect 442316 299170 442372 299180
rect 442540 307972 442596 307982
rect 442204 276770 442260 276780
rect 442316 295204 442372 295214
rect 442092 276546 442148 276556
rect 441980 275314 442036 275324
rect 442316 275268 442372 295148
rect 442428 291172 442484 291182
rect 442428 276724 442484 291116
rect 442428 276658 442484 276668
rect 442316 275202 442372 275212
rect 441084 269602 441140 269612
rect 442092 273140 442148 273150
rect 440972 266242 441028 266252
rect 441980 266532 442036 266542
rect 440860 262882 440916 262892
rect 440972 263284 441028 263294
rect 440972 235172 441028 263228
rect 440972 235106 441028 235116
rect 441868 235172 441924 235182
rect 440524 231858 440580 231868
rect 441868 229236 441924 235116
rect 441980 232596 442036 266476
rect 442092 236628 442148 273084
rect 442428 265188 442484 265198
rect 442316 265076 442372 265086
rect 442092 236562 442148 236572
rect 442204 264628 442260 264638
rect 442204 233268 442260 264572
rect 442316 237300 442372 265020
rect 442316 237234 442372 237244
rect 442204 233202 442260 233212
rect 441980 232530 442036 232540
rect 442428 229908 442484 265132
rect 442540 264964 442596 307916
rect 442540 264898 442596 264908
rect 442652 304612 442708 304622
rect 442652 264852 442708 304556
rect 442764 297892 442820 297902
rect 442764 273812 442820 297836
rect 442764 273746 442820 273756
rect 442652 264786 442708 264796
rect 442428 229842 442484 229852
rect 441868 229170 441924 229180
rect 439218 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 439838 226350
rect 439218 226226 439838 226294
rect 439218 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 439838 226226
rect 439218 226102 439838 226170
rect 439218 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 439838 226102
rect 439218 225978 439838 226046
rect 439218 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 439838 225978
rect 439218 208350 439838 225922
rect 443548 216658 443604 312620
rect 445228 311332 445284 311342
rect 443660 306628 443716 306638
rect 443660 274820 443716 306572
rect 443660 274754 443716 274764
rect 443548 216592 443604 216602
rect 445228 216478 445284 311276
rect 466218 310350 466838 327922
rect 466218 310294 466314 310350
rect 466370 310294 466438 310350
rect 466494 310294 466562 310350
rect 466618 310294 466686 310350
rect 466742 310294 466838 310350
rect 466218 310226 466838 310294
rect 466218 310170 466314 310226
rect 466370 310170 466438 310226
rect 466494 310170 466562 310226
rect 466618 310170 466686 310226
rect 466742 310170 466838 310226
rect 466218 310102 466838 310170
rect 466218 310046 466314 310102
rect 466370 310046 466438 310102
rect 466494 310046 466562 310102
rect 466618 310046 466686 310102
rect 466742 310046 466838 310102
rect 466218 309978 466838 310046
rect 466218 309922 466314 309978
rect 466370 309922 466438 309978
rect 466494 309922 466562 309978
rect 466618 309922 466686 309978
rect 466742 309922 466838 309978
rect 445340 308644 445396 308654
rect 445340 217378 445396 308588
rect 445340 217312 445396 217322
rect 466218 292350 466838 309922
rect 466218 292294 466314 292350
rect 466370 292294 466438 292350
rect 466494 292294 466562 292350
rect 466618 292294 466686 292350
rect 466742 292294 466838 292350
rect 466218 292226 466838 292294
rect 466218 292170 466314 292226
rect 466370 292170 466438 292226
rect 466494 292170 466562 292226
rect 466618 292170 466686 292226
rect 466742 292170 466838 292226
rect 466218 292102 466838 292170
rect 466218 292046 466314 292102
rect 466370 292046 466438 292102
rect 466494 292046 466562 292102
rect 466618 292046 466686 292102
rect 466742 292046 466838 292102
rect 466218 291978 466838 292046
rect 466218 291922 466314 291978
rect 466370 291922 466438 291978
rect 466494 291922 466562 291978
rect 466618 291922 466686 291978
rect 466742 291922 466838 291978
rect 466218 274350 466838 291922
rect 466218 274294 466314 274350
rect 466370 274294 466438 274350
rect 466494 274294 466562 274350
rect 466618 274294 466686 274350
rect 466742 274294 466838 274350
rect 466218 274226 466838 274294
rect 466218 274170 466314 274226
rect 466370 274170 466438 274226
rect 466494 274170 466562 274226
rect 466618 274170 466686 274226
rect 466742 274170 466838 274226
rect 466218 274102 466838 274170
rect 466218 274046 466314 274102
rect 466370 274046 466438 274102
rect 466494 274046 466562 274102
rect 466618 274046 466686 274102
rect 466742 274046 466838 274102
rect 466218 273978 466838 274046
rect 466218 273922 466314 273978
rect 466370 273922 466438 273978
rect 466494 273922 466562 273978
rect 466618 273922 466686 273978
rect 466742 273922 466838 273978
rect 466218 256350 466838 273922
rect 466218 256294 466314 256350
rect 466370 256294 466438 256350
rect 466494 256294 466562 256350
rect 466618 256294 466686 256350
rect 466742 256294 466838 256350
rect 466218 256226 466838 256294
rect 466218 256170 466314 256226
rect 466370 256170 466438 256226
rect 466494 256170 466562 256226
rect 466618 256170 466686 256226
rect 466742 256170 466838 256226
rect 466218 256102 466838 256170
rect 466218 256046 466314 256102
rect 466370 256046 466438 256102
rect 466494 256046 466562 256102
rect 466618 256046 466686 256102
rect 466742 256046 466838 256102
rect 466218 255978 466838 256046
rect 466218 255922 466314 255978
rect 466370 255922 466438 255978
rect 466494 255922 466562 255978
rect 466618 255922 466686 255978
rect 466742 255922 466838 255978
rect 466218 238350 466838 255922
rect 466218 238294 466314 238350
rect 466370 238294 466438 238350
rect 466494 238294 466562 238350
rect 466618 238294 466686 238350
rect 466742 238294 466838 238350
rect 466218 238226 466838 238294
rect 466218 238170 466314 238226
rect 466370 238170 466438 238226
rect 466494 238170 466562 238226
rect 466618 238170 466686 238226
rect 466742 238170 466838 238226
rect 466218 238102 466838 238170
rect 466218 238046 466314 238102
rect 466370 238046 466438 238102
rect 466494 238046 466562 238102
rect 466618 238046 466686 238102
rect 466742 238046 466838 238102
rect 466218 237978 466838 238046
rect 466218 237922 466314 237978
rect 466370 237922 466438 237978
rect 466494 237922 466562 237978
rect 466618 237922 466686 237978
rect 466742 237922 466838 237978
rect 466218 220350 466838 237922
rect 466218 220294 466314 220350
rect 466370 220294 466438 220350
rect 466494 220294 466562 220350
rect 466618 220294 466686 220350
rect 466742 220294 466838 220350
rect 466218 220226 466838 220294
rect 466218 220170 466314 220226
rect 466370 220170 466438 220226
rect 466494 220170 466562 220226
rect 466618 220170 466686 220226
rect 466742 220170 466838 220226
rect 466218 220102 466838 220170
rect 466218 220046 466314 220102
rect 466370 220046 466438 220102
rect 466494 220046 466562 220102
rect 466618 220046 466686 220102
rect 466742 220046 466838 220102
rect 466218 219978 466838 220046
rect 466218 219922 466314 219978
rect 466370 219922 466438 219978
rect 466494 219922 466562 219978
rect 466618 219922 466686 219978
rect 466742 219922 466838 219978
rect 445228 216412 445284 216422
rect 439218 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 439838 208350
rect 439218 208226 439838 208294
rect 439218 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 439838 208226
rect 439218 208102 439838 208170
rect 439218 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 439838 208102
rect 439218 207978 439838 208046
rect 439218 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 439838 207978
rect 435498 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 436118 184350
rect 435498 184226 436118 184294
rect 435498 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 436118 184226
rect 435498 184102 436118 184170
rect 435498 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 436118 184102
rect 435498 183978 436118 184046
rect 435498 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 436118 183978
rect 435498 166350 436118 183922
rect 435498 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 436118 166350
rect 435498 166226 436118 166294
rect 435498 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 436118 166226
rect 435498 166102 436118 166170
rect 435498 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 436118 166102
rect 435498 165978 436118 166046
rect 435498 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 436118 165978
rect 435498 148350 436118 165922
rect 435498 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 436118 148350
rect 435498 148226 436118 148294
rect 435498 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 436118 148226
rect 435498 148102 436118 148170
rect 435498 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 436118 148102
rect 435498 147978 436118 148046
rect 435498 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 436118 147978
rect 433580 132290 433636 132300
rect 432012 132178 432068 132188
rect 431900 131954 431956 131964
rect 435498 130350 436118 147922
rect 436828 199556 436884 199566
rect 436828 132468 436884 199500
rect 436828 132402 436884 132412
rect 439218 190350 439838 207922
rect 442092 215938 442148 215948
rect 441868 200788 441924 200798
rect 440300 195972 440356 195982
rect 439218 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 439838 190350
rect 439218 190226 439838 190294
rect 439218 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 439838 190226
rect 439218 190102 439838 190170
rect 439218 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 439838 190102
rect 439218 189978 439838 190046
rect 439218 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 439838 189978
rect 439218 172350 439838 189922
rect 439218 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 439838 172350
rect 439218 172226 439838 172294
rect 439218 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 439838 172226
rect 439218 172102 439838 172170
rect 439218 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 439838 172102
rect 439218 171978 439838 172046
rect 439218 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 439838 171978
rect 439218 154350 439838 171922
rect 439218 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 439838 154350
rect 439218 154226 439838 154294
rect 439218 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 439838 154226
rect 439218 154102 439838 154170
rect 439218 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 439838 154102
rect 439218 153978 439838 154046
rect 439218 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 439838 153978
rect 439218 136350 439838 153922
rect 439218 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 439838 136350
rect 439218 136226 439838 136294
rect 439218 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 439838 136226
rect 439218 136102 439838 136170
rect 439218 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 439838 136102
rect 439218 135978 439838 136046
rect 439218 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 439838 135978
rect 408498 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 409118 118350
rect 408498 118226 409118 118294
rect 408498 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 409118 118226
rect 408498 118102 409118 118170
rect 408498 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 409118 118102
rect 408498 117978 409118 118046
rect 408498 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 409118 117978
rect 408498 116310 409118 117922
rect 429212 130340 429268 130350
rect 429212 124292 429268 130284
rect 435498 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 436118 130350
rect 435498 130226 436118 130294
rect 435498 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 436118 130226
rect 435498 130102 436118 130170
rect 435498 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 436118 130102
rect 435498 129978 436118 130046
rect 435498 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 436118 129978
rect 433468 128884 433524 128894
rect 398188 115972 398244 115982
rect 415168 112350 415488 112384
rect 415168 112294 415238 112350
rect 415294 112294 415362 112350
rect 415418 112294 415488 112350
rect 415168 112226 415488 112294
rect 415168 112170 415238 112226
rect 415294 112170 415362 112226
rect 415418 112170 415488 112226
rect 415168 112102 415488 112170
rect 415168 112046 415238 112102
rect 415294 112046 415362 112102
rect 415418 112046 415488 112102
rect 415168 111978 415488 112046
rect 415168 111922 415238 111978
rect 415294 111922 415362 111978
rect 415418 111922 415488 111978
rect 415168 111888 415488 111922
rect 399808 100350 400128 100384
rect 399808 100294 399878 100350
rect 399934 100294 400002 100350
rect 400058 100294 400128 100350
rect 399808 100226 400128 100294
rect 399808 100170 399878 100226
rect 399934 100170 400002 100226
rect 400058 100170 400128 100226
rect 399808 100102 400128 100170
rect 399808 100046 399878 100102
rect 399934 100046 400002 100102
rect 400058 100046 400128 100102
rect 399808 99978 400128 100046
rect 399808 99922 399878 99978
rect 399934 99922 400002 99978
rect 400058 99922 400128 99978
rect 399808 99888 400128 99922
rect 415168 94350 415488 94384
rect 415168 94294 415238 94350
rect 415294 94294 415362 94350
rect 415418 94294 415488 94350
rect 415168 94226 415488 94294
rect 415168 94170 415238 94226
rect 415294 94170 415362 94226
rect 415418 94170 415488 94226
rect 415168 94102 415488 94170
rect 415168 94046 415238 94102
rect 415294 94046 415362 94102
rect 415418 94046 415488 94102
rect 415168 93978 415488 94046
rect 415168 93922 415238 93978
rect 415294 93922 415362 93978
rect 415418 93922 415488 93978
rect 415168 93888 415488 93922
rect 399808 82350 400128 82384
rect 399808 82294 399878 82350
rect 399934 82294 400002 82350
rect 400058 82294 400128 82350
rect 399808 82226 400128 82294
rect 399808 82170 399878 82226
rect 399934 82170 400002 82226
rect 400058 82170 400128 82226
rect 399808 82102 400128 82170
rect 399808 82046 399878 82102
rect 399934 82046 400002 82102
rect 400058 82046 400128 82102
rect 399808 81978 400128 82046
rect 399808 81922 399878 81978
rect 399934 81922 400002 81978
rect 400058 81922 400128 81978
rect 399808 81888 400128 81922
rect 415168 76350 415488 76384
rect 415168 76294 415238 76350
rect 415294 76294 415362 76350
rect 415418 76294 415488 76350
rect 415168 76226 415488 76294
rect 415168 76170 415238 76226
rect 415294 76170 415362 76226
rect 415418 76170 415488 76226
rect 415168 76102 415488 76170
rect 415168 76046 415238 76102
rect 415294 76046 415362 76102
rect 415418 76046 415488 76102
rect 415168 75978 415488 76046
rect 415168 75922 415238 75978
rect 415294 75922 415362 75978
rect 415418 75922 415488 75978
rect 415168 75888 415488 75922
rect 399808 64350 400128 64384
rect 399808 64294 399878 64350
rect 399934 64294 400002 64350
rect 400058 64294 400128 64350
rect 399808 64226 400128 64294
rect 399808 64170 399878 64226
rect 399934 64170 400002 64226
rect 400058 64170 400128 64226
rect 399808 64102 400128 64170
rect 399808 64046 399878 64102
rect 399934 64046 400002 64102
rect 400058 64046 400128 64102
rect 399808 63978 400128 64046
rect 399808 63922 399878 63978
rect 399934 63922 400002 63978
rect 400058 63922 400128 63978
rect 399808 63888 400128 63922
rect 415168 58350 415488 58384
rect 415168 58294 415238 58350
rect 415294 58294 415362 58350
rect 415418 58294 415488 58350
rect 415168 58226 415488 58294
rect 415168 58170 415238 58226
rect 415294 58170 415362 58226
rect 415418 58170 415488 58226
rect 415168 58102 415488 58170
rect 415168 58046 415238 58102
rect 415294 58046 415362 58102
rect 415418 58046 415488 58102
rect 415168 57978 415488 58046
rect 415168 57922 415238 57978
rect 415294 57922 415362 57978
rect 415418 57922 415488 57978
rect 415168 57888 415488 57922
rect 403564 48020 403620 48030
rect 396844 46340 396900 46350
rect 396844 45780 396900 46284
rect 396844 45714 396900 45724
rect 398188 46228 398244 46238
rect 398188 45780 398244 46172
rect 398188 45714 398244 45724
rect 403564 45780 403620 47964
rect 417676 47908 417732 47918
rect 403564 45714 403620 45724
rect 396396 42914 396452 42924
rect 387212 41682 387268 41692
rect 379820 40226 379876 40236
rect 404778 40350 405398 46266
rect 404778 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 405398 40350
rect 404778 40226 405398 40294
rect 377778 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 378398 28350
rect 377778 28226 378398 28294
rect 377778 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 378398 28226
rect 377778 28102 378398 28170
rect 377778 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 378398 28102
rect 377778 27978 378398 28046
rect 377778 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 378398 27978
rect 377778 10350 378398 27922
rect 377778 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 378398 10350
rect 377778 10226 378398 10294
rect 377778 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 378398 10226
rect 377778 10102 378398 10170
rect 377778 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 378398 10102
rect 377778 9978 378398 10046
rect 377778 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 378398 9978
rect 377778 -1120 378398 9922
rect 377778 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 378398 -1120
rect 377778 -1244 378398 -1176
rect 377778 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 378398 -1244
rect 377778 -1368 378398 -1300
rect 377778 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 378398 -1368
rect 377778 -1492 378398 -1424
rect 377778 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 378398 -1492
rect 377778 -1644 378398 -1548
rect 404778 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 405398 40226
rect 404778 40102 405398 40170
rect 404778 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 405398 40102
rect 404778 39978 405398 40046
rect 404778 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 405398 39978
rect 404778 22350 405398 39922
rect 408498 46198 409118 46266
rect 408498 46142 408594 46198
rect 408650 46142 408718 46198
rect 408774 46142 408842 46198
rect 408898 46142 408966 46198
rect 409022 46142 409118 46198
rect 408498 46074 409118 46142
rect 408498 46018 408594 46074
rect 408650 46018 408718 46074
rect 408774 46018 408842 46074
rect 408898 46018 408966 46074
rect 409022 46018 409118 46074
rect 408498 45950 409118 46018
rect 408498 45894 408594 45950
rect 408650 45894 408718 45950
rect 408774 45894 408842 45950
rect 408898 45894 408966 45950
rect 409022 45894 409118 45950
rect 408498 33828 409118 45894
rect 417676 45780 417732 47852
rect 417676 45714 417732 45724
rect 419692 43678 419748 43688
rect 419692 43584 419748 43596
rect 429212 43652 429268 124236
rect 431788 127092 431844 127102
rect 430528 118350 430848 118384
rect 430528 118294 430598 118350
rect 430654 118294 430722 118350
rect 430778 118294 430848 118350
rect 430528 118226 430848 118294
rect 430528 118170 430598 118226
rect 430654 118170 430722 118226
rect 430778 118170 430848 118226
rect 430528 118102 430848 118170
rect 430528 118046 430598 118102
rect 430654 118046 430722 118102
rect 430778 118046 430848 118102
rect 430528 117978 430848 118046
rect 430528 117922 430598 117978
rect 430654 117922 430722 117978
rect 430778 117922 430848 117978
rect 430528 117888 430848 117922
rect 430528 100350 430848 100384
rect 430528 100294 430598 100350
rect 430654 100294 430722 100350
rect 430778 100294 430848 100350
rect 430528 100226 430848 100294
rect 430528 100170 430598 100226
rect 430654 100170 430722 100226
rect 430778 100170 430848 100226
rect 430528 100102 430848 100170
rect 430528 100046 430598 100102
rect 430654 100046 430722 100102
rect 430778 100046 430848 100102
rect 430528 99978 430848 100046
rect 430528 99922 430598 99978
rect 430654 99922 430722 99978
rect 430778 99922 430848 99978
rect 430528 99888 430848 99922
rect 430528 82350 430848 82384
rect 430528 82294 430598 82350
rect 430654 82294 430722 82350
rect 430778 82294 430848 82350
rect 430528 82226 430848 82294
rect 430528 82170 430598 82226
rect 430654 82170 430722 82226
rect 430778 82170 430848 82226
rect 430528 82102 430848 82170
rect 430528 82046 430598 82102
rect 430654 82046 430722 82102
rect 430778 82046 430848 82102
rect 430528 81978 430848 82046
rect 430528 81922 430598 81978
rect 430654 81922 430722 81978
rect 430778 81922 430848 81978
rect 430528 81888 430848 81922
rect 430528 64350 430848 64384
rect 430528 64294 430598 64350
rect 430654 64294 430722 64350
rect 430778 64294 430848 64350
rect 430528 64226 430848 64294
rect 430528 64170 430598 64226
rect 430654 64170 430722 64226
rect 430778 64170 430848 64226
rect 430528 64102 430848 64170
rect 430528 64046 430598 64102
rect 430654 64046 430722 64102
rect 430778 64046 430848 64102
rect 430528 63978 430848 64046
rect 430528 63922 430598 63978
rect 430654 63922 430722 63978
rect 430778 63922 430848 63978
rect 430528 63888 430848 63922
rect 429212 43586 429268 43596
rect 431788 43540 431844 127036
rect 431788 43474 431844 43484
rect 433468 43204 433524 128828
rect 433468 43138 433524 43148
rect 435498 112350 436118 129922
rect 435498 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 436118 112350
rect 435498 112226 436118 112294
rect 435498 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 436118 112226
rect 435498 112102 436118 112170
rect 435498 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 436118 112102
rect 435498 111978 436118 112046
rect 435498 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 436118 111978
rect 435498 94350 436118 111922
rect 435498 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 436118 94350
rect 435498 94226 436118 94294
rect 435498 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 436118 94226
rect 435498 94102 436118 94170
rect 435498 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 436118 94102
rect 435498 93978 436118 94046
rect 435498 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 436118 93978
rect 435498 76350 436118 93922
rect 435498 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 436118 76350
rect 435498 76226 436118 76294
rect 435498 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 436118 76226
rect 435498 76102 436118 76170
rect 435498 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 436118 76102
rect 435498 75978 436118 76046
rect 435498 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 436118 75978
rect 435498 58350 436118 75922
rect 435498 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 436118 58350
rect 435498 58226 436118 58294
rect 435498 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 436118 58226
rect 435498 58102 436118 58170
rect 435498 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 436118 58102
rect 435498 57978 436118 58046
rect 435498 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 436118 57978
rect 435498 40350 436118 57922
rect 435498 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 436118 40350
rect 435498 40226 436118 40294
rect 435498 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 436118 40226
rect 435498 40102 436118 40170
rect 435498 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 436118 40102
rect 435498 39978 436118 40046
rect 435498 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 436118 39978
rect 409096 28350 409416 28384
rect 409096 28294 409166 28350
rect 409222 28294 409290 28350
rect 409346 28294 409416 28350
rect 409096 28226 409416 28294
rect 409096 28170 409166 28226
rect 409222 28170 409290 28226
rect 409346 28170 409416 28226
rect 409096 28102 409416 28170
rect 409096 28046 409166 28102
rect 409222 28046 409290 28102
rect 409346 28046 409416 28102
rect 409096 27978 409416 28046
rect 409096 27922 409166 27978
rect 409222 27922 409290 27978
rect 409346 27922 409416 27978
rect 409096 27888 409416 27922
rect 404778 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 405398 22350
rect 404778 22226 405398 22294
rect 404778 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 405398 22226
rect 404778 22102 405398 22170
rect 404778 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 405398 22102
rect 404778 21978 405398 22046
rect 404778 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 405398 21978
rect 404778 4350 405398 21922
rect 435498 22350 436118 39922
rect 435498 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 436118 22350
rect 435498 22226 436118 22294
rect 435498 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 436118 22226
rect 435498 22102 436118 22170
rect 435498 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 436118 22102
rect 435498 21978 436118 22046
rect 435498 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 436118 21978
rect 409096 10350 409416 10384
rect 409096 10294 409166 10350
rect 409222 10294 409290 10350
rect 409346 10294 409416 10350
rect 409096 10226 409416 10294
rect 409096 10170 409166 10226
rect 409222 10170 409290 10226
rect 409346 10170 409416 10226
rect 409096 10102 409416 10170
rect 409096 10046 409166 10102
rect 409222 10046 409290 10102
rect 409346 10046 409416 10102
rect 409096 9978 409416 10046
rect 409096 9922 409166 9978
rect 409222 9922 409290 9978
rect 409346 9922 409416 9978
rect 409096 9888 409416 9922
rect 404778 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 405398 4350
rect 404778 4226 405398 4294
rect 404778 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 405398 4226
rect 404778 4102 405398 4170
rect 404778 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 405398 4102
rect 404778 3978 405398 4046
rect 404778 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 405398 3978
rect 404778 -160 405398 3922
rect 404778 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 405398 -160
rect 404778 -284 405398 -216
rect 404778 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 405398 -284
rect 404778 -408 405398 -340
rect 404778 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 405398 -408
rect 404778 -532 405398 -464
rect 404778 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 405398 -532
rect 404778 -1644 405398 -588
rect 435498 4350 436118 21922
rect 435498 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 436118 4350
rect 435498 4226 436118 4294
rect 435498 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 436118 4226
rect 435498 4102 436118 4170
rect 435498 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 436118 4102
rect 435498 3978 436118 4046
rect 435498 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 436118 3978
rect 435498 -160 436118 3922
rect 439218 118350 439838 135922
rect 439218 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 439838 118350
rect 439218 118226 439838 118294
rect 439218 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 439838 118226
rect 439218 118102 439838 118170
rect 439218 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 439838 118102
rect 439218 117978 439838 118046
rect 439218 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 439838 117978
rect 439218 100350 439838 117922
rect 439218 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 439838 100350
rect 439218 100226 439838 100294
rect 439218 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 439838 100226
rect 439218 100102 439838 100170
rect 439218 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 439838 100102
rect 439218 99978 439838 100046
rect 439218 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 439838 99978
rect 439218 82350 439838 99922
rect 439218 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 439838 82350
rect 439218 82226 439838 82294
rect 439218 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 439838 82226
rect 439218 82102 439838 82170
rect 439218 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 439838 82102
rect 439218 81978 439838 82046
rect 440188 191828 440244 191838
rect 440188 82068 440244 191772
rect 440300 174020 440356 195916
rect 441868 178724 441924 200732
rect 441980 199108 442036 199118
rect 441980 193396 442036 199052
rect 441980 193330 442036 193340
rect 441868 178658 441924 178668
rect 441980 193258 442036 193268
rect 440300 173954 440356 173964
rect 441980 173348 442036 193202
rect 442092 179396 442148 215882
rect 442540 214138 442596 214148
rect 442204 205716 442260 205726
rect 442204 191828 442260 205660
rect 442204 191762 442260 191772
rect 442316 199220 442372 199230
rect 442092 179330 442148 179340
rect 442316 175364 442372 199164
rect 442428 194404 442484 194414
rect 442428 178052 442484 194348
rect 442428 177986 442484 177996
rect 442540 176708 442596 214082
rect 442540 176642 442596 176652
rect 442652 212518 442708 212528
rect 442316 175298 442372 175308
rect 442652 174692 442708 212462
rect 466218 202350 466838 219922
rect 466218 202294 466314 202350
rect 466370 202294 466438 202350
rect 466494 202294 466562 202350
rect 466618 202294 466686 202350
rect 466742 202294 466838 202350
rect 466218 202226 466838 202294
rect 466218 202170 466314 202226
rect 466370 202170 466438 202226
rect 466494 202170 466562 202226
rect 466618 202170 466686 202226
rect 466742 202170 466838 202226
rect 466218 202102 466838 202170
rect 466218 202046 466314 202102
rect 466370 202046 466438 202102
rect 466494 202046 466562 202102
rect 466618 202046 466686 202102
rect 466742 202046 466838 202102
rect 466218 201978 466838 202046
rect 466218 201922 466314 201978
rect 466370 201922 466438 201978
rect 466494 201922 466562 201978
rect 466618 201922 466686 201978
rect 466742 201922 466838 201978
rect 443772 200900 443828 200910
rect 442876 195748 442932 195758
rect 442764 192388 442820 192398
rect 442764 176036 442820 192332
rect 442764 175970 442820 175980
rect 442652 174626 442708 174636
rect 441980 173282 442036 173292
rect 442876 169988 442932 195692
rect 442876 169922 442932 169932
rect 443548 194740 443604 194750
rect 440636 163268 440692 163278
rect 440412 161924 440468 161934
rect 440412 161308 440468 161868
rect 440412 161252 440580 161308
rect 440300 135268 440356 135278
rect 440300 82740 440356 135212
rect 440300 82674 440356 82684
rect 440412 126868 440468 126878
rect 440188 82002 440244 82012
rect 439218 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 439838 81978
rect 439218 64350 439838 81922
rect 440412 79380 440468 126812
rect 440524 115858 440580 161252
rect 440636 120898 440692 163212
rect 442316 162932 442372 162942
rect 441868 158564 441924 158574
rect 441868 133678 441924 158508
rect 442316 149548 442372 162876
rect 441868 133612 441924 133622
rect 442092 149492 442372 149548
rect 441980 133498 442036 133508
rect 440636 120832 440692 120842
rect 441868 126980 441924 126990
rect 440524 115792 440580 115802
rect 440412 79314 440468 79324
rect 441868 76692 441924 126924
rect 441980 84084 442036 133442
rect 442092 117478 442148 149492
rect 442092 117412 442148 117422
rect 442204 123620 442260 123630
rect 441980 84018 442036 84028
rect 442204 80724 442260 123564
rect 443548 88788 443604 194684
rect 443660 184978 443716 184988
rect 443660 90804 443716 184922
rect 443772 169316 443828 200844
rect 445228 200564 445284 200574
rect 443884 195860 443940 195870
rect 443884 171332 443940 195804
rect 443884 171266 443940 171276
rect 443772 169250 443828 169260
rect 443772 133588 443828 133598
rect 443772 91476 443828 133532
rect 443772 91410 443828 91420
rect 443660 90738 443716 90748
rect 443548 88722 443604 88732
rect 442204 80658 442260 80668
rect 445228 80052 445284 200508
rect 450268 197204 450324 197214
rect 447020 194964 447076 194974
rect 446908 192724 446964 192734
rect 445340 191604 445396 191614
rect 445340 88116 445396 191548
rect 445340 88050 445396 88060
rect 446908 86100 446964 192668
rect 447020 90132 447076 194908
rect 447020 90066 447076 90076
rect 448588 193844 448644 193854
rect 446908 86034 446964 86044
rect 448588 85428 448644 193788
rect 450268 86772 450324 197148
rect 450268 86706 450324 86716
rect 466218 184350 466838 201922
rect 466218 184294 466314 184350
rect 466370 184294 466438 184350
rect 466494 184294 466562 184350
rect 466618 184294 466686 184350
rect 466742 184294 466838 184350
rect 466218 184226 466838 184294
rect 466218 184170 466314 184226
rect 466370 184170 466438 184226
rect 466494 184170 466562 184226
rect 466618 184170 466686 184226
rect 466742 184170 466838 184226
rect 466218 184102 466838 184170
rect 466218 184046 466314 184102
rect 466370 184046 466438 184102
rect 466494 184046 466562 184102
rect 466618 184046 466686 184102
rect 466742 184046 466838 184102
rect 466218 183978 466838 184046
rect 466218 183922 466314 183978
rect 466370 183922 466438 183978
rect 466494 183922 466562 183978
rect 466618 183922 466686 183978
rect 466742 183922 466838 183978
rect 466218 166350 466838 183922
rect 466218 166294 466314 166350
rect 466370 166294 466438 166350
rect 466494 166294 466562 166350
rect 466618 166294 466686 166350
rect 466742 166294 466838 166350
rect 466218 166226 466838 166294
rect 466218 166170 466314 166226
rect 466370 166170 466438 166226
rect 466494 166170 466562 166226
rect 466618 166170 466686 166226
rect 466742 166170 466838 166226
rect 466218 166102 466838 166170
rect 466218 166046 466314 166102
rect 466370 166046 466438 166102
rect 466494 166046 466562 166102
rect 466618 166046 466686 166102
rect 466742 166046 466838 166102
rect 466218 165978 466838 166046
rect 466218 165922 466314 165978
rect 466370 165922 466438 165978
rect 466494 165922 466562 165978
rect 466618 165922 466686 165978
rect 466742 165922 466838 165978
rect 466218 148350 466838 165922
rect 466218 148294 466314 148350
rect 466370 148294 466438 148350
rect 466494 148294 466562 148350
rect 466618 148294 466686 148350
rect 466742 148294 466838 148350
rect 466218 148226 466838 148294
rect 466218 148170 466314 148226
rect 466370 148170 466438 148226
rect 466494 148170 466562 148226
rect 466618 148170 466686 148226
rect 466742 148170 466838 148226
rect 466218 148102 466838 148170
rect 466218 148046 466314 148102
rect 466370 148046 466438 148102
rect 466494 148046 466562 148102
rect 466618 148046 466686 148102
rect 466742 148046 466838 148102
rect 466218 147978 466838 148046
rect 466218 147922 466314 147978
rect 466370 147922 466438 147978
rect 466494 147922 466562 147978
rect 466618 147922 466686 147978
rect 466742 147922 466838 147978
rect 466218 130350 466838 147922
rect 466218 130294 466314 130350
rect 466370 130294 466438 130350
rect 466494 130294 466562 130350
rect 466618 130294 466686 130350
rect 466742 130294 466838 130350
rect 466218 130226 466838 130294
rect 466218 130170 466314 130226
rect 466370 130170 466438 130226
rect 466494 130170 466562 130226
rect 466618 130170 466686 130226
rect 466742 130170 466838 130226
rect 466218 130102 466838 130170
rect 466218 130046 466314 130102
rect 466370 130046 466438 130102
rect 466494 130046 466562 130102
rect 466618 130046 466686 130102
rect 466742 130046 466838 130102
rect 466218 129978 466838 130046
rect 466218 129922 466314 129978
rect 466370 129922 466438 129978
rect 466494 129922 466562 129978
rect 466618 129922 466686 129978
rect 466742 129922 466838 129978
rect 466218 112350 466838 129922
rect 466218 112294 466314 112350
rect 466370 112294 466438 112350
rect 466494 112294 466562 112350
rect 466618 112294 466686 112350
rect 466742 112294 466838 112350
rect 466218 112226 466838 112294
rect 466218 112170 466314 112226
rect 466370 112170 466438 112226
rect 466494 112170 466562 112226
rect 466618 112170 466686 112226
rect 466742 112170 466838 112226
rect 466218 112102 466838 112170
rect 466218 112046 466314 112102
rect 466370 112046 466438 112102
rect 466494 112046 466562 112102
rect 466618 112046 466686 112102
rect 466742 112046 466838 112102
rect 466218 111978 466838 112046
rect 466218 111922 466314 111978
rect 466370 111922 466438 111978
rect 466494 111922 466562 111978
rect 466618 111922 466686 111978
rect 466742 111922 466838 111978
rect 466218 94350 466838 111922
rect 466218 94294 466314 94350
rect 466370 94294 466438 94350
rect 466494 94294 466562 94350
rect 466618 94294 466686 94350
rect 466742 94294 466838 94350
rect 466218 94226 466838 94294
rect 466218 94170 466314 94226
rect 466370 94170 466438 94226
rect 466494 94170 466562 94226
rect 466618 94170 466686 94226
rect 466742 94170 466838 94226
rect 466218 94102 466838 94170
rect 466218 94046 466314 94102
rect 466370 94046 466438 94102
rect 466494 94046 466562 94102
rect 466618 94046 466686 94102
rect 466742 94046 466838 94102
rect 466218 93978 466838 94046
rect 466218 93922 466314 93978
rect 466370 93922 466438 93978
rect 466494 93922 466562 93978
rect 466618 93922 466686 93978
rect 466742 93922 466838 93978
rect 448588 85362 448644 85372
rect 445228 79986 445284 79996
rect 441868 76626 441924 76636
rect 464448 76350 464768 76384
rect 464448 76294 464518 76350
rect 464574 76294 464642 76350
rect 464698 76294 464768 76350
rect 464448 76226 464768 76294
rect 464448 76170 464518 76226
rect 464574 76170 464642 76226
rect 464698 76170 464768 76226
rect 464448 76102 464768 76170
rect 464448 76046 464518 76102
rect 464574 76046 464642 76102
rect 464698 76046 464768 76102
rect 464448 75978 464768 76046
rect 464448 75922 464518 75978
rect 464574 75922 464642 75978
rect 464698 75922 464768 75978
rect 464448 75888 464768 75922
rect 466218 76350 466838 93922
rect 466218 76294 466314 76350
rect 466370 76294 466438 76350
rect 466494 76294 466562 76350
rect 466618 76294 466686 76350
rect 466742 76294 466838 76350
rect 466218 76226 466838 76294
rect 466218 76170 466314 76226
rect 466370 76170 466438 76226
rect 466494 76170 466562 76226
rect 466618 76170 466686 76226
rect 466742 76170 466838 76226
rect 466218 76102 466838 76170
rect 466218 76046 466314 76102
rect 466370 76046 466438 76102
rect 466494 76046 466562 76102
rect 466618 76046 466686 76102
rect 466742 76046 466838 76102
rect 466218 75978 466838 76046
rect 466218 75922 466314 75978
rect 466370 75922 466438 75978
rect 466494 75922 466562 75978
rect 466618 75922 466686 75978
rect 466742 75922 466838 75978
rect 439218 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 439838 64350
rect 439218 64226 439838 64294
rect 439218 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 439838 64226
rect 439218 64102 439838 64170
rect 439218 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 439838 64102
rect 439218 63978 439838 64046
rect 439218 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 439838 63978
rect 439218 46350 439838 63922
rect 464448 58350 464768 58384
rect 464448 58294 464518 58350
rect 464574 58294 464642 58350
rect 464698 58294 464768 58350
rect 464448 58226 464768 58294
rect 464448 58170 464518 58226
rect 464574 58170 464642 58226
rect 464698 58170 464768 58226
rect 464448 58102 464768 58170
rect 464448 58046 464518 58102
rect 464574 58046 464642 58102
rect 464698 58046 464768 58102
rect 464448 57978 464768 58046
rect 464448 57922 464518 57978
rect 464574 57922 464642 57978
rect 464698 57922 464768 57978
rect 464448 57888 464768 57922
rect 466218 58350 466838 75922
rect 466218 58294 466314 58350
rect 466370 58294 466438 58350
rect 466494 58294 466562 58350
rect 466618 58294 466686 58350
rect 466742 58294 466838 58350
rect 466218 58226 466838 58294
rect 466218 58170 466314 58226
rect 466370 58170 466438 58226
rect 466494 58170 466562 58226
rect 466618 58170 466686 58226
rect 466742 58170 466838 58226
rect 466218 58102 466838 58170
rect 466218 58046 466314 58102
rect 466370 58046 466438 58102
rect 466494 58046 466562 58102
rect 466618 58046 466686 58102
rect 466742 58046 466838 58102
rect 466218 57978 466838 58046
rect 466218 57922 466314 57978
rect 466370 57922 466438 57978
rect 466494 57922 466562 57978
rect 466618 57922 466686 57978
rect 466742 57922 466838 57978
rect 439218 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 439838 46350
rect 439218 46226 439838 46294
rect 439218 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 439838 46226
rect 439218 46102 439838 46170
rect 439218 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 439838 46102
rect 439218 45978 439838 46046
rect 439218 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 439838 45978
rect 439218 28350 439838 45922
rect 439218 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 439838 28350
rect 439218 28226 439838 28294
rect 439218 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 439838 28226
rect 439218 28102 439838 28170
rect 439218 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 439838 28102
rect 439218 27978 439838 28046
rect 439218 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 439838 27978
rect 439218 10350 439838 27922
rect 439218 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 439838 10350
rect 439218 10226 439838 10294
rect 439218 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 439838 10226
rect 439218 10102 439838 10170
rect 439218 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 439838 10102
rect 439218 9978 439838 10046
rect 439218 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 439838 9978
rect 436828 1876 436884 1886
rect 436828 196 436884 1820
rect 436828 130 436884 140
rect 435498 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 436118 -160
rect 435498 -284 436118 -216
rect 435498 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 436118 -284
rect 435498 -408 436118 -340
rect 435498 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 436118 -408
rect 435498 -532 436118 -464
rect 435498 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 436118 -532
rect 435498 -1644 436118 -588
rect 439218 -1120 439838 9922
rect 466218 40350 466838 57922
rect 466218 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 466838 40350
rect 466218 40226 466838 40294
rect 466218 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 466838 40226
rect 466218 40102 466838 40170
rect 466218 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 466838 40102
rect 466218 39978 466838 40046
rect 466218 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 466838 39978
rect 466218 22350 466838 39922
rect 466218 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 466838 22350
rect 466218 22226 466838 22294
rect 466218 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 466838 22226
rect 466218 22102 466838 22170
rect 466218 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 466838 22102
rect 466218 21978 466838 22046
rect 466218 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 466838 21978
rect 442988 5158 443044 5168
rect 442988 5058 443044 5068
rect 466218 4350 466838 21922
rect 466218 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 466838 4350
rect 466218 4226 466838 4294
rect 466218 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 466838 4226
rect 466218 4102 466838 4170
rect 466218 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 466838 4102
rect 466218 3978 466838 4046
rect 466218 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 466838 3978
rect 447692 3358 447748 3370
rect 447692 3266 447748 3276
rect 457100 2996 457156 3006
rect 457100 478 457156 2940
rect 457100 412 457156 422
rect 439218 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 439838 -1120
rect 439218 -1244 439838 -1176
rect 439218 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 439838 -1244
rect 439218 -1368 439838 -1300
rect 439218 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 439838 -1368
rect 439218 -1492 439838 -1424
rect 439218 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 439838 -1492
rect 439218 -1644 439838 -1548
rect 466218 -160 466838 3922
rect 466218 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 466838 -160
rect 466218 -284 466838 -216
rect 466218 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 466838 -284
rect 466218 -408 466838 -340
rect 466218 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 466838 -408
rect 466218 -532 466838 -464
rect 466218 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 466838 -532
rect 466218 -1644 466838 -588
rect 469938 598172 470558 598268
rect 469938 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 470558 598172
rect 469938 598048 470558 598116
rect 469938 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 470558 598048
rect 469938 597924 470558 597992
rect 469938 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 470558 597924
rect 469938 597800 470558 597868
rect 469938 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 470558 597800
rect 469938 586350 470558 597744
rect 469938 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 470558 586350
rect 469938 586226 470558 586294
rect 469938 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 470558 586226
rect 469938 586102 470558 586170
rect 469938 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 470558 586102
rect 469938 585978 470558 586046
rect 469938 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 470558 585978
rect 469938 568350 470558 585922
rect 469938 568294 470034 568350
rect 470090 568294 470158 568350
rect 470214 568294 470282 568350
rect 470338 568294 470406 568350
rect 470462 568294 470558 568350
rect 469938 568226 470558 568294
rect 469938 568170 470034 568226
rect 470090 568170 470158 568226
rect 470214 568170 470282 568226
rect 470338 568170 470406 568226
rect 470462 568170 470558 568226
rect 469938 568102 470558 568170
rect 469938 568046 470034 568102
rect 470090 568046 470158 568102
rect 470214 568046 470282 568102
rect 470338 568046 470406 568102
rect 470462 568046 470558 568102
rect 469938 567978 470558 568046
rect 469938 567922 470034 567978
rect 470090 567922 470158 567978
rect 470214 567922 470282 567978
rect 470338 567922 470406 567978
rect 470462 567922 470558 567978
rect 469938 550350 470558 567922
rect 469938 550294 470034 550350
rect 470090 550294 470158 550350
rect 470214 550294 470282 550350
rect 470338 550294 470406 550350
rect 470462 550294 470558 550350
rect 469938 550226 470558 550294
rect 469938 550170 470034 550226
rect 470090 550170 470158 550226
rect 470214 550170 470282 550226
rect 470338 550170 470406 550226
rect 470462 550170 470558 550226
rect 469938 550102 470558 550170
rect 469938 550046 470034 550102
rect 470090 550046 470158 550102
rect 470214 550046 470282 550102
rect 470338 550046 470406 550102
rect 470462 550046 470558 550102
rect 469938 549978 470558 550046
rect 469938 549922 470034 549978
rect 470090 549922 470158 549978
rect 470214 549922 470282 549978
rect 470338 549922 470406 549978
rect 470462 549922 470558 549978
rect 469938 532350 470558 549922
rect 469938 532294 470034 532350
rect 470090 532294 470158 532350
rect 470214 532294 470282 532350
rect 470338 532294 470406 532350
rect 470462 532294 470558 532350
rect 469938 532226 470558 532294
rect 469938 532170 470034 532226
rect 470090 532170 470158 532226
rect 470214 532170 470282 532226
rect 470338 532170 470406 532226
rect 470462 532170 470558 532226
rect 469938 532102 470558 532170
rect 469938 532046 470034 532102
rect 470090 532046 470158 532102
rect 470214 532046 470282 532102
rect 470338 532046 470406 532102
rect 470462 532046 470558 532102
rect 469938 531978 470558 532046
rect 469938 531922 470034 531978
rect 470090 531922 470158 531978
rect 470214 531922 470282 531978
rect 470338 531922 470406 531978
rect 470462 531922 470558 531978
rect 469938 514350 470558 531922
rect 469938 514294 470034 514350
rect 470090 514294 470158 514350
rect 470214 514294 470282 514350
rect 470338 514294 470406 514350
rect 470462 514294 470558 514350
rect 469938 514226 470558 514294
rect 469938 514170 470034 514226
rect 470090 514170 470158 514226
rect 470214 514170 470282 514226
rect 470338 514170 470406 514226
rect 470462 514170 470558 514226
rect 469938 514102 470558 514170
rect 469938 514046 470034 514102
rect 470090 514046 470158 514102
rect 470214 514046 470282 514102
rect 470338 514046 470406 514102
rect 470462 514046 470558 514102
rect 469938 513978 470558 514046
rect 469938 513922 470034 513978
rect 470090 513922 470158 513978
rect 470214 513922 470282 513978
rect 470338 513922 470406 513978
rect 470462 513922 470558 513978
rect 469938 496350 470558 513922
rect 469938 496294 470034 496350
rect 470090 496294 470158 496350
rect 470214 496294 470282 496350
rect 470338 496294 470406 496350
rect 470462 496294 470558 496350
rect 469938 496226 470558 496294
rect 469938 496170 470034 496226
rect 470090 496170 470158 496226
rect 470214 496170 470282 496226
rect 470338 496170 470406 496226
rect 470462 496170 470558 496226
rect 469938 496102 470558 496170
rect 469938 496046 470034 496102
rect 470090 496046 470158 496102
rect 470214 496046 470282 496102
rect 470338 496046 470406 496102
rect 470462 496046 470558 496102
rect 469938 495978 470558 496046
rect 469938 495922 470034 495978
rect 470090 495922 470158 495978
rect 470214 495922 470282 495978
rect 470338 495922 470406 495978
rect 470462 495922 470558 495978
rect 469938 478350 470558 495922
rect 469938 478294 470034 478350
rect 470090 478294 470158 478350
rect 470214 478294 470282 478350
rect 470338 478294 470406 478350
rect 470462 478294 470558 478350
rect 469938 478226 470558 478294
rect 469938 478170 470034 478226
rect 470090 478170 470158 478226
rect 470214 478170 470282 478226
rect 470338 478170 470406 478226
rect 470462 478170 470558 478226
rect 469938 478102 470558 478170
rect 469938 478046 470034 478102
rect 470090 478046 470158 478102
rect 470214 478046 470282 478102
rect 470338 478046 470406 478102
rect 470462 478046 470558 478102
rect 469938 477978 470558 478046
rect 469938 477922 470034 477978
rect 470090 477922 470158 477978
rect 470214 477922 470282 477978
rect 470338 477922 470406 477978
rect 470462 477922 470558 477978
rect 469938 460350 470558 477922
rect 469938 460294 470034 460350
rect 470090 460294 470158 460350
rect 470214 460294 470282 460350
rect 470338 460294 470406 460350
rect 470462 460294 470558 460350
rect 469938 460226 470558 460294
rect 469938 460170 470034 460226
rect 470090 460170 470158 460226
rect 470214 460170 470282 460226
rect 470338 460170 470406 460226
rect 470462 460170 470558 460226
rect 469938 460102 470558 460170
rect 469938 460046 470034 460102
rect 470090 460046 470158 460102
rect 470214 460046 470282 460102
rect 470338 460046 470406 460102
rect 470462 460046 470558 460102
rect 469938 459978 470558 460046
rect 469938 459922 470034 459978
rect 470090 459922 470158 459978
rect 470214 459922 470282 459978
rect 470338 459922 470406 459978
rect 470462 459922 470558 459978
rect 469938 442350 470558 459922
rect 469938 442294 470034 442350
rect 470090 442294 470158 442350
rect 470214 442294 470282 442350
rect 470338 442294 470406 442350
rect 470462 442294 470558 442350
rect 469938 442226 470558 442294
rect 469938 442170 470034 442226
rect 470090 442170 470158 442226
rect 470214 442170 470282 442226
rect 470338 442170 470406 442226
rect 470462 442170 470558 442226
rect 469938 442102 470558 442170
rect 469938 442046 470034 442102
rect 470090 442046 470158 442102
rect 470214 442046 470282 442102
rect 470338 442046 470406 442102
rect 470462 442046 470558 442102
rect 469938 441978 470558 442046
rect 469938 441922 470034 441978
rect 470090 441922 470158 441978
rect 470214 441922 470282 441978
rect 470338 441922 470406 441978
rect 470462 441922 470558 441978
rect 469938 424350 470558 441922
rect 469938 424294 470034 424350
rect 470090 424294 470158 424350
rect 470214 424294 470282 424350
rect 470338 424294 470406 424350
rect 470462 424294 470558 424350
rect 469938 424226 470558 424294
rect 469938 424170 470034 424226
rect 470090 424170 470158 424226
rect 470214 424170 470282 424226
rect 470338 424170 470406 424226
rect 470462 424170 470558 424226
rect 469938 424102 470558 424170
rect 469938 424046 470034 424102
rect 470090 424046 470158 424102
rect 470214 424046 470282 424102
rect 470338 424046 470406 424102
rect 470462 424046 470558 424102
rect 469938 423978 470558 424046
rect 469938 423922 470034 423978
rect 470090 423922 470158 423978
rect 470214 423922 470282 423978
rect 470338 423922 470406 423978
rect 470462 423922 470558 423978
rect 469938 406350 470558 423922
rect 469938 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 470558 406350
rect 469938 406226 470558 406294
rect 469938 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 470558 406226
rect 469938 406102 470558 406170
rect 469938 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 470558 406102
rect 469938 405978 470558 406046
rect 469938 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 470558 405978
rect 469938 388350 470558 405922
rect 469938 388294 470034 388350
rect 470090 388294 470158 388350
rect 470214 388294 470282 388350
rect 470338 388294 470406 388350
rect 470462 388294 470558 388350
rect 469938 388226 470558 388294
rect 469938 388170 470034 388226
rect 470090 388170 470158 388226
rect 470214 388170 470282 388226
rect 470338 388170 470406 388226
rect 470462 388170 470558 388226
rect 469938 388102 470558 388170
rect 469938 388046 470034 388102
rect 470090 388046 470158 388102
rect 470214 388046 470282 388102
rect 470338 388046 470406 388102
rect 470462 388046 470558 388102
rect 469938 387978 470558 388046
rect 469938 387922 470034 387978
rect 470090 387922 470158 387978
rect 470214 387922 470282 387978
rect 470338 387922 470406 387978
rect 470462 387922 470558 387978
rect 469938 370350 470558 387922
rect 469938 370294 470034 370350
rect 470090 370294 470158 370350
rect 470214 370294 470282 370350
rect 470338 370294 470406 370350
rect 470462 370294 470558 370350
rect 469938 370226 470558 370294
rect 469938 370170 470034 370226
rect 470090 370170 470158 370226
rect 470214 370170 470282 370226
rect 470338 370170 470406 370226
rect 470462 370170 470558 370226
rect 469938 370102 470558 370170
rect 469938 370046 470034 370102
rect 470090 370046 470158 370102
rect 470214 370046 470282 370102
rect 470338 370046 470406 370102
rect 470462 370046 470558 370102
rect 469938 369978 470558 370046
rect 469938 369922 470034 369978
rect 470090 369922 470158 369978
rect 470214 369922 470282 369978
rect 470338 369922 470406 369978
rect 470462 369922 470558 369978
rect 469938 352350 470558 369922
rect 469938 352294 470034 352350
rect 470090 352294 470158 352350
rect 470214 352294 470282 352350
rect 470338 352294 470406 352350
rect 470462 352294 470558 352350
rect 469938 352226 470558 352294
rect 469938 352170 470034 352226
rect 470090 352170 470158 352226
rect 470214 352170 470282 352226
rect 470338 352170 470406 352226
rect 470462 352170 470558 352226
rect 469938 352102 470558 352170
rect 469938 352046 470034 352102
rect 470090 352046 470158 352102
rect 470214 352046 470282 352102
rect 470338 352046 470406 352102
rect 470462 352046 470558 352102
rect 469938 351978 470558 352046
rect 469938 351922 470034 351978
rect 470090 351922 470158 351978
rect 470214 351922 470282 351978
rect 470338 351922 470406 351978
rect 470462 351922 470558 351978
rect 469938 334350 470558 351922
rect 469938 334294 470034 334350
rect 470090 334294 470158 334350
rect 470214 334294 470282 334350
rect 470338 334294 470406 334350
rect 470462 334294 470558 334350
rect 469938 334226 470558 334294
rect 469938 334170 470034 334226
rect 470090 334170 470158 334226
rect 470214 334170 470282 334226
rect 470338 334170 470406 334226
rect 470462 334170 470558 334226
rect 469938 334102 470558 334170
rect 469938 334046 470034 334102
rect 470090 334046 470158 334102
rect 470214 334046 470282 334102
rect 470338 334046 470406 334102
rect 470462 334046 470558 334102
rect 469938 333978 470558 334046
rect 469938 333922 470034 333978
rect 470090 333922 470158 333978
rect 470214 333922 470282 333978
rect 470338 333922 470406 333978
rect 470462 333922 470558 333978
rect 469938 316350 470558 333922
rect 469938 316294 470034 316350
rect 470090 316294 470158 316350
rect 470214 316294 470282 316350
rect 470338 316294 470406 316350
rect 470462 316294 470558 316350
rect 469938 316226 470558 316294
rect 469938 316170 470034 316226
rect 470090 316170 470158 316226
rect 470214 316170 470282 316226
rect 470338 316170 470406 316226
rect 470462 316170 470558 316226
rect 469938 316102 470558 316170
rect 469938 316046 470034 316102
rect 470090 316046 470158 316102
rect 470214 316046 470282 316102
rect 470338 316046 470406 316102
rect 470462 316046 470558 316102
rect 469938 315978 470558 316046
rect 469938 315922 470034 315978
rect 470090 315922 470158 315978
rect 470214 315922 470282 315978
rect 470338 315922 470406 315978
rect 470462 315922 470558 315978
rect 469938 298350 470558 315922
rect 469938 298294 470034 298350
rect 470090 298294 470158 298350
rect 470214 298294 470282 298350
rect 470338 298294 470406 298350
rect 470462 298294 470558 298350
rect 469938 298226 470558 298294
rect 469938 298170 470034 298226
rect 470090 298170 470158 298226
rect 470214 298170 470282 298226
rect 470338 298170 470406 298226
rect 470462 298170 470558 298226
rect 469938 298102 470558 298170
rect 469938 298046 470034 298102
rect 470090 298046 470158 298102
rect 470214 298046 470282 298102
rect 470338 298046 470406 298102
rect 470462 298046 470558 298102
rect 469938 297978 470558 298046
rect 469938 297922 470034 297978
rect 470090 297922 470158 297978
rect 470214 297922 470282 297978
rect 470338 297922 470406 297978
rect 470462 297922 470558 297978
rect 469938 280350 470558 297922
rect 469938 280294 470034 280350
rect 470090 280294 470158 280350
rect 470214 280294 470282 280350
rect 470338 280294 470406 280350
rect 470462 280294 470558 280350
rect 469938 280226 470558 280294
rect 469938 280170 470034 280226
rect 470090 280170 470158 280226
rect 470214 280170 470282 280226
rect 470338 280170 470406 280226
rect 470462 280170 470558 280226
rect 469938 280102 470558 280170
rect 469938 280046 470034 280102
rect 470090 280046 470158 280102
rect 470214 280046 470282 280102
rect 470338 280046 470406 280102
rect 470462 280046 470558 280102
rect 469938 279978 470558 280046
rect 469938 279922 470034 279978
rect 470090 279922 470158 279978
rect 470214 279922 470282 279978
rect 470338 279922 470406 279978
rect 470462 279922 470558 279978
rect 469938 262350 470558 279922
rect 469938 262294 470034 262350
rect 470090 262294 470158 262350
rect 470214 262294 470282 262350
rect 470338 262294 470406 262350
rect 470462 262294 470558 262350
rect 469938 262226 470558 262294
rect 469938 262170 470034 262226
rect 470090 262170 470158 262226
rect 470214 262170 470282 262226
rect 470338 262170 470406 262226
rect 470462 262170 470558 262226
rect 469938 262102 470558 262170
rect 469938 262046 470034 262102
rect 470090 262046 470158 262102
rect 470214 262046 470282 262102
rect 470338 262046 470406 262102
rect 470462 262046 470558 262102
rect 469938 261978 470558 262046
rect 469938 261922 470034 261978
rect 470090 261922 470158 261978
rect 470214 261922 470282 261978
rect 470338 261922 470406 261978
rect 470462 261922 470558 261978
rect 469938 244350 470558 261922
rect 469938 244294 470034 244350
rect 470090 244294 470158 244350
rect 470214 244294 470282 244350
rect 470338 244294 470406 244350
rect 470462 244294 470558 244350
rect 469938 244226 470558 244294
rect 469938 244170 470034 244226
rect 470090 244170 470158 244226
rect 470214 244170 470282 244226
rect 470338 244170 470406 244226
rect 470462 244170 470558 244226
rect 469938 244102 470558 244170
rect 469938 244046 470034 244102
rect 470090 244046 470158 244102
rect 470214 244046 470282 244102
rect 470338 244046 470406 244102
rect 470462 244046 470558 244102
rect 469938 243978 470558 244046
rect 469938 243922 470034 243978
rect 470090 243922 470158 243978
rect 470214 243922 470282 243978
rect 470338 243922 470406 243978
rect 470462 243922 470558 243978
rect 469938 226350 470558 243922
rect 469938 226294 470034 226350
rect 470090 226294 470158 226350
rect 470214 226294 470282 226350
rect 470338 226294 470406 226350
rect 470462 226294 470558 226350
rect 469938 226226 470558 226294
rect 469938 226170 470034 226226
rect 470090 226170 470158 226226
rect 470214 226170 470282 226226
rect 470338 226170 470406 226226
rect 470462 226170 470558 226226
rect 469938 226102 470558 226170
rect 469938 226046 470034 226102
rect 470090 226046 470158 226102
rect 470214 226046 470282 226102
rect 470338 226046 470406 226102
rect 470462 226046 470558 226102
rect 469938 225978 470558 226046
rect 469938 225922 470034 225978
rect 470090 225922 470158 225978
rect 470214 225922 470282 225978
rect 470338 225922 470406 225978
rect 470462 225922 470558 225978
rect 469938 208350 470558 225922
rect 469938 208294 470034 208350
rect 470090 208294 470158 208350
rect 470214 208294 470282 208350
rect 470338 208294 470406 208350
rect 470462 208294 470558 208350
rect 469938 208226 470558 208294
rect 469938 208170 470034 208226
rect 470090 208170 470158 208226
rect 470214 208170 470282 208226
rect 470338 208170 470406 208226
rect 470462 208170 470558 208226
rect 469938 208102 470558 208170
rect 469938 208046 470034 208102
rect 470090 208046 470158 208102
rect 470214 208046 470282 208102
rect 470338 208046 470406 208102
rect 470462 208046 470558 208102
rect 469938 207978 470558 208046
rect 469938 207922 470034 207978
rect 470090 207922 470158 207978
rect 470214 207922 470282 207978
rect 470338 207922 470406 207978
rect 470462 207922 470558 207978
rect 469938 190350 470558 207922
rect 469938 190294 470034 190350
rect 470090 190294 470158 190350
rect 470214 190294 470282 190350
rect 470338 190294 470406 190350
rect 470462 190294 470558 190350
rect 469938 190226 470558 190294
rect 469938 190170 470034 190226
rect 470090 190170 470158 190226
rect 470214 190170 470282 190226
rect 470338 190170 470406 190226
rect 470462 190170 470558 190226
rect 469938 190102 470558 190170
rect 469938 190046 470034 190102
rect 470090 190046 470158 190102
rect 470214 190046 470282 190102
rect 470338 190046 470406 190102
rect 470462 190046 470558 190102
rect 469938 189978 470558 190046
rect 469938 189922 470034 189978
rect 470090 189922 470158 189978
rect 470214 189922 470282 189978
rect 470338 189922 470406 189978
rect 470462 189922 470558 189978
rect 469938 172350 470558 189922
rect 469938 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 470558 172350
rect 469938 172226 470558 172294
rect 469938 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 470558 172226
rect 469938 172102 470558 172170
rect 469938 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 470558 172102
rect 469938 171978 470558 172046
rect 469938 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 470558 171978
rect 469938 154350 470558 171922
rect 469938 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 470558 154350
rect 469938 154226 470558 154294
rect 469938 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 470558 154226
rect 469938 154102 470558 154170
rect 469938 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 470558 154102
rect 469938 153978 470558 154046
rect 469938 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 470558 153978
rect 469938 136350 470558 153922
rect 469938 136294 470034 136350
rect 470090 136294 470158 136350
rect 470214 136294 470282 136350
rect 470338 136294 470406 136350
rect 470462 136294 470558 136350
rect 469938 136226 470558 136294
rect 469938 136170 470034 136226
rect 470090 136170 470158 136226
rect 470214 136170 470282 136226
rect 470338 136170 470406 136226
rect 470462 136170 470558 136226
rect 469938 136102 470558 136170
rect 469938 136046 470034 136102
rect 470090 136046 470158 136102
rect 470214 136046 470282 136102
rect 470338 136046 470406 136102
rect 470462 136046 470558 136102
rect 469938 135978 470558 136046
rect 469938 135922 470034 135978
rect 470090 135922 470158 135978
rect 470214 135922 470282 135978
rect 470338 135922 470406 135978
rect 470462 135922 470558 135978
rect 469938 118350 470558 135922
rect 469938 118294 470034 118350
rect 470090 118294 470158 118350
rect 470214 118294 470282 118350
rect 470338 118294 470406 118350
rect 470462 118294 470558 118350
rect 469938 118226 470558 118294
rect 469938 118170 470034 118226
rect 470090 118170 470158 118226
rect 470214 118170 470282 118226
rect 470338 118170 470406 118226
rect 470462 118170 470558 118226
rect 469938 118102 470558 118170
rect 469938 118046 470034 118102
rect 470090 118046 470158 118102
rect 470214 118046 470282 118102
rect 470338 118046 470406 118102
rect 470462 118046 470558 118102
rect 469938 117978 470558 118046
rect 469938 117922 470034 117978
rect 470090 117922 470158 117978
rect 470214 117922 470282 117978
rect 470338 117922 470406 117978
rect 470462 117922 470558 117978
rect 469938 100350 470558 117922
rect 469938 100294 470034 100350
rect 470090 100294 470158 100350
rect 470214 100294 470282 100350
rect 470338 100294 470406 100350
rect 470462 100294 470558 100350
rect 469938 100226 470558 100294
rect 469938 100170 470034 100226
rect 470090 100170 470158 100226
rect 470214 100170 470282 100226
rect 470338 100170 470406 100226
rect 470462 100170 470558 100226
rect 469938 100102 470558 100170
rect 469938 100046 470034 100102
rect 470090 100046 470158 100102
rect 470214 100046 470282 100102
rect 470338 100046 470406 100102
rect 470462 100046 470558 100102
rect 469938 99978 470558 100046
rect 469938 99922 470034 99978
rect 470090 99922 470158 99978
rect 470214 99922 470282 99978
rect 470338 99922 470406 99978
rect 470462 99922 470558 99978
rect 469938 82350 470558 99922
rect 496938 597212 497558 598268
rect 496938 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 497558 597212
rect 496938 597088 497558 597156
rect 496938 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 497558 597088
rect 496938 596964 497558 597032
rect 496938 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 497558 596964
rect 496938 596840 497558 596908
rect 496938 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 497558 596840
rect 496938 580350 497558 596784
rect 496938 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 497558 580350
rect 496938 580226 497558 580294
rect 496938 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 497558 580226
rect 496938 580102 497558 580170
rect 496938 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 497558 580102
rect 496938 579978 497558 580046
rect 496938 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 497558 579978
rect 496938 562350 497558 579922
rect 496938 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 497558 562350
rect 496938 562226 497558 562294
rect 496938 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 497558 562226
rect 496938 562102 497558 562170
rect 496938 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 497558 562102
rect 496938 561978 497558 562046
rect 496938 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 497558 561978
rect 496938 544350 497558 561922
rect 496938 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 497558 544350
rect 496938 544226 497558 544294
rect 496938 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 497558 544226
rect 496938 544102 497558 544170
rect 496938 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 497558 544102
rect 496938 543978 497558 544046
rect 496938 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 497558 543978
rect 496938 526350 497558 543922
rect 496938 526294 497034 526350
rect 497090 526294 497158 526350
rect 497214 526294 497282 526350
rect 497338 526294 497406 526350
rect 497462 526294 497558 526350
rect 496938 526226 497558 526294
rect 496938 526170 497034 526226
rect 497090 526170 497158 526226
rect 497214 526170 497282 526226
rect 497338 526170 497406 526226
rect 497462 526170 497558 526226
rect 496938 526102 497558 526170
rect 496938 526046 497034 526102
rect 497090 526046 497158 526102
rect 497214 526046 497282 526102
rect 497338 526046 497406 526102
rect 497462 526046 497558 526102
rect 496938 525978 497558 526046
rect 496938 525922 497034 525978
rect 497090 525922 497158 525978
rect 497214 525922 497282 525978
rect 497338 525922 497406 525978
rect 497462 525922 497558 525978
rect 496938 508350 497558 525922
rect 496938 508294 497034 508350
rect 497090 508294 497158 508350
rect 497214 508294 497282 508350
rect 497338 508294 497406 508350
rect 497462 508294 497558 508350
rect 496938 508226 497558 508294
rect 496938 508170 497034 508226
rect 497090 508170 497158 508226
rect 497214 508170 497282 508226
rect 497338 508170 497406 508226
rect 497462 508170 497558 508226
rect 496938 508102 497558 508170
rect 496938 508046 497034 508102
rect 497090 508046 497158 508102
rect 497214 508046 497282 508102
rect 497338 508046 497406 508102
rect 497462 508046 497558 508102
rect 496938 507978 497558 508046
rect 496938 507922 497034 507978
rect 497090 507922 497158 507978
rect 497214 507922 497282 507978
rect 497338 507922 497406 507978
rect 497462 507922 497558 507978
rect 496938 490350 497558 507922
rect 496938 490294 497034 490350
rect 497090 490294 497158 490350
rect 497214 490294 497282 490350
rect 497338 490294 497406 490350
rect 497462 490294 497558 490350
rect 496938 490226 497558 490294
rect 496938 490170 497034 490226
rect 497090 490170 497158 490226
rect 497214 490170 497282 490226
rect 497338 490170 497406 490226
rect 497462 490170 497558 490226
rect 496938 490102 497558 490170
rect 496938 490046 497034 490102
rect 497090 490046 497158 490102
rect 497214 490046 497282 490102
rect 497338 490046 497406 490102
rect 497462 490046 497558 490102
rect 496938 489978 497558 490046
rect 496938 489922 497034 489978
rect 497090 489922 497158 489978
rect 497214 489922 497282 489978
rect 497338 489922 497406 489978
rect 497462 489922 497558 489978
rect 496938 472350 497558 489922
rect 496938 472294 497034 472350
rect 497090 472294 497158 472350
rect 497214 472294 497282 472350
rect 497338 472294 497406 472350
rect 497462 472294 497558 472350
rect 496938 472226 497558 472294
rect 496938 472170 497034 472226
rect 497090 472170 497158 472226
rect 497214 472170 497282 472226
rect 497338 472170 497406 472226
rect 497462 472170 497558 472226
rect 496938 472102 497558 472170
rect 496938 472046 497034 472102
rect 497090 472046 497158 472102
rect 497214 472046 497282 472102
rect 497338 472046 497406 472102
rect 497462 472046 497558 472102
rect 496938 471978 497558 472046
rect 496938 471922 497034 471978
rect 497090 471922 497158 471978
rect 497214 471922 497282 471978
rect 497338 471922 497406 471978
rect 497462 471922 497558 471978
rect 496938 454350 497558 471922
rect 496938 454294 497034 454350
rect 497090 454294 497158 454350
rect 497214 454294 497282 454350
rect 497338 454294 497406 454350
rect 497462 454294 497558 454350
rect 496938 454226 497558 454294
rect 496938 454170 497034 454226
rect 497090 454170 497158 454226
rect 497214 454170 497282 454226
rect 497338 454170 497406 454226
rect 497462 454170 497558 454226
rect 496938 454102 497558 454170
rect 496938 454046 497034 454102
rect 497090 454046 497158 454102
rect 497214 454046 497282 454102
rect 497338 454046 497406 454102
rect 497462 454046 497558 454102
rect 496938 453978 497558 454046
rect 496938 453922 497034 453978
rect 497090 453922 497158 453978
rect 497214 453922 497282 453978
rect 497338 453922 497406 453978
rect 497462 453922 497558 453978
rect 496938 436350 497558 453922
rect 496938 436294 497034 436350
rect 497090 436294 497158 436350
rect 497214 436294 497282 436350
rect 497338 436294 497406 436350
rect 497462 436294 497558 436350
rect 496938 436226 497558 436294
rect 496938 436170 497034 436226
rect 497090 436170 497158 436226
rect 497214 436170 497282 436226
rect 497338 436170 497406 436226
rect 497462 436170 497558 436226
rect 496938 436102 497558 436170
rect 496938 436046 497034 436102
rect 497090 436046 497158 436102
rect 497214 436046 497282 436102
rect 497338 436046 497406 436102
rect 497462 436046 497558 436102
rect 496938 435978 497558 436046
rect 496938 435922 497034 435978
rect 497090 435922 497158 435978
rect 497214 435922 497282 435978
rect 497338 435922 497406 435978
rect 497462 435922 497558 435978
rect 496938 418350 497558 435922
rect 496938 418294 497034 418350
rect 497090 418294 497158 418350
rect 497214 418294 497282 418350
rect 497338 418294 497406 418350
rect 497462 418294 497558 418350
rect 496938 418226 497558 418294
rect 496938 418170 497034 418226
rect 497090 418170 497158 418226
rect 497214 418170 497282 418226
rect 497338 418170 497406 418226
rect 497462 418170 497558 418226
rect 496938 418102 497558 418170
rect 496938 418046 497034 418102
rect 497090 418046 497158 418102
rect 497214 418046 497282 418102
rect 497338 418046 497406 418102
rect 497462 418046 497558 418102
rect 496938 417978 497558 418046
rect 496938 417922 497034 417978
rect 497090 417922 497158 417978
rect 497214 417922 497282 417978
rect 497338 417922 497406 417978
rect 497462 417922 497558 417978
rect 496938 400350 497558 417922
rect 496938 400294 497034 400350
rect 497090 400294 497158 400350
rect 497214 400294 497282 400350
rect 497338 400294 497406 400350
rect 497462 400294 497558 400350
rect 496938 400226 497558 400294
rect 496938 400170 497034 400226
rect 497090 400170 497158 400226
rect 497214 400170 497282 400226
rect 497338 400170 497406 400226
rect 497462 400170 497558 400226
rect 496938 400102 497558 400170
rect 496938 400046 497034 400102
rect 497090 400046 497158 400102
rect 497214 400046 497282 400102
rect 497338 400046 497406 400102
rect 497462 400046 497558 400102
rect 496938 399978 497558 400046
rect 496938 399922 497034 399978
rect 497090 399922 497158 399978
rect 497214 399922 497282 399978
rect 497338 399922 497406 399978
rect 497462 399922 497558 399978
rect 496938 382350 497558 399922
rect 496938 382294 497034 382350
rect 497090 382294 497158 382350
rect 497214 382294 497282 382350
rect 497338 382294 497406 382350
rect 497462 382294 497558 382350
rect 496938 382226 497558 382294
rect 496938 382170 497034 382226
rect 497090 382170 497158 382226
rect 497214 382170 497282 382226
rect 497338 382170 497406 382226
rect 497462 382170 497558 382226
rect 496938 382102 497558 382170
rect 496938 382046 497034 382102
rect 497090 382046 497158 382102
rect 497214 382046 497282 382102
rect 497338 382046 497406 382102
rect 497462 382046 497558 382102
rect 496938 381978 497558 382046
rect 496938 381922 497034 381978
rect 497090 381922 497158 381978
rect 497214 381922 497282 381978
rect 497338 381922 497406 381978
rect 497462 381922 497558 381978
rect 496938 364350 497558 381922
rect 496938 364294 497034 364350
rect 497090 364294 497158 364350
rect 497214 364294 497282 364350
rect 497338 364294 497406 364350
rect 497462 364294 497558 364350
rect 496938 364226 497558 364294
rect 496938 364170 497034 364226
rect 497090 364170 497158 364226
rect 497214 364170 497282 364226
rect 497338 364170 497406 364226
rect 497462 364170 497558 364226
rect 496938 364102 497558 364170
rect 496938 364046 497034 364102
rect 497090 364046 497158 364102
rect 497214 364046 497282 364102
rect 497338 364046 497406 364102
rect 497462 364046 497558 364102
rect 496938 363978 497558 364046
rect 496938 363922 497034 363978
rect 497090 363922 497158 363978
rect 497214 363922 497282 363978
rect 497338 363922 497406 363978
rect 497462 363922 497558 363978
rect 496938 346350 497558 363922
rect 496938 346294 497034 346350
rect 497090 346294 497158 346350
rect 497214 346294 497282 346350
rect 497338 346294 497406 346350
rect 497462 346294 497558 346350
rect 496938 346226 497558 346294
rect 496938 346170 497034 346226
rect 497090 346170 497158 346226
rect 497214 346170 497282 346226
rect 497338 346170 497406 346226
rect 497462 346170 497558 346226
rect 496938 346102 497558 346170
rect 496938 346046 497034 346102
rect 497090 346046 497158 346102
rect 497214 346046 497282 346102
rect 497338 346046 497406 346102
rect 497462 346046 497558 346102
rect 496938 345978 497558 346046
rect 496938 345922 497034 345978
rect 497090 345922 497158 345978
rect 497214 345922 497282 345978
rect 497338 345922 497406 345978
rect 497462 345922 497558 345978
rect 496938 328350 497558 345922
rect 496938 328294 497034 328350
rect 497090 328294 497158 328350
rect 497214 328294 497282 328350
rect 497338 328294 497406 328350
rect 497462 328294 497558 328350
rect 496938 328226 497558 328294
rect 496938 328170 497034 328226
rect 497090 328170 497158 328226
rect 497214 328170 497282 328226
rect 497338 328170 497406 328226
rect 497462 328170 497558 328226
rect 496938 328102 497558 328170
rect 496938 328046 497034 328102
rect 497090 328046 497158 328102
rect 497214 328046 497282 328102
rect 497338 328046 497406 328102
rect 497462 328046 497558 328102
rect 496938 327978 497558 328046
rect 496938 327922 497034 327978
rect 497090 327922 497158 327978
rect 497214 327922 497282 327978
rect 497338 327922 497406 327978
rect 497462 327922 497558 327978
rect 496938 310350 497558 327922
rect 496938 310294 497034 310350
rect 497090 310294 497158 310350
rect 497214 310294 497282 310350
rect 497338 310294 497406 310350
rect 497462 310294 497558 310350
rect 496938 310226 497558 310294
rect 496938 310170 497034 310226
rect 497090 310170 497158 310226
rect 497214 310170 497282 310226
rect 497338 310170 497406 310226
rect 497462 310170 497558 310226
rect 496938 310102 497558 310170
rect 496938 310046 497034 310102
rect 497090 310046 497158 310102
rect 497214 310046 497282 310102
rect 497338 310046 497406 310102
rect 497462 310046 497558 310102
rect 496938 309978 497558 310046
rect 496938 309922 497034 309978
rect 497090 309922 497158 309978
rect 497214 309922 497282 309978
rect 497338 309922 497406 309978
rect 497462 309922 497558 309978
rect 496938 292350 497558 309922
rect 496938 292294 497034 292350
rect 497090 292294 497158 292350
rect 497214 292294 497282 292350
rect 497338 292294 497406 292350
rect 497462 292294 497558 292350
rect 496938 292226 497558 292294
rect 496938 292170 497034 292226
rect 497090 292170 497158 292226
rect 497214 292170 497282 292226
rect 497338 292170 497406 292226
rect 497462 292170 497558 292226
rect 496938 292102 497558 292170
rect 496938 292046 497034 292102
rect 497090 292046 497158 292102
rect 497214 292046 497282 292102
rect 497338 292046 497406 292102
rect 497462 292046 497558 292102
rect 496938 291978 497558 292046
rect 496938 291922 497034 291978
rect 497090 291922 497158 291978
rect 497214 291922 497282 291978
rect 497338 291922 497406 291978
rect 497462 291922 497558 291978
rect 496938 274350 497558 291922
rect 496938 274294 497034 274350
rect 497090 274294 497158 274350
rect 497214 274294 497282 274350
rect 497338 274294 497406 274350
rect 497462 274294 497558 274350
rect 496938 274226 497558 274294
rect 496938 274170 497034 274226
rect 497090 274170 497158 274226
rect 497214 274170 497282 274226
rect 497338 274170 497406 274226
rect 497462 274170 497558 274226
rect 496938 274102 497558 274170
rect 496938 274046 497034 274102
rect 497090 274046 497158 274102
rect 497214 274046 497282 274102
rect 497338 274046 497406 274102
rect 497462 274046 497558 274102
rect 496938 273978 497558 274046
rect 496938 273922 497034 273978
rect 497090 273922 497158 273978
rect 497214 273922 497282 273978
rect 497338 273922 497406 273978
rect 497462 273922 497558 273978
rect 496938 256350 497558 273922
rect 496938 256294 497034 256350
rect 497090 256294 497158 256350
rect 497214 256294 497282 256350
rect 497338 256294 497406 256350
rect 497462 256294 497558 256350
rect 496938 256226 497558 256294
rect 496938 256170 497034 256226
rect 497090 256170 497158 256226
rect 497214 256170 497282 256226
rect 497338 256170 497406 256226
rect 497462 256170 497558 256226
rect 496938 256102 497558 256170
rect 496938 256046 497034 256102
rect 497090 256046 497158 256102
rect 497214 256046 497282 256102
rect 497338 256046 497406 256102
rect 497462 256046 497558 256102
rect 496938 255978 497558 256046
rect 496938 255922 497034 255978
rect 497090 255922 497158 255978
rect 497214 255922 497282 255978
rect 497338 255922 497406 255978
rect 497462 255922 497558 255978
rect 496938 238350 497558 255922
rect 496938 238294 497034 238350
rect 497090 238294 497158 238350
rect 497214 238294 497282 238350
rect 497338 238294 497406 238350
rect 497462 238294 497558 238350
rect 496938 238226 497558 238294
rect 496938 238170 497034 238226
rect 497090 238170 497158 238226
rect 497214 238170 497282 238226
rect 497338 238170 497406 238226
rect 497462 238170 497558 238226
rect 496938 238102 497558 238170
rect 496938 238046 497034 238102
rect 497090 238046 497158 238102
rect 497214 238046 497282 238102
rect 497338 238046 497406 238102
rect 497462 238046 497558 238102
rect 496938 237978 497558 238046
rect 496938 237922 497034 237978
rect 497090 237922 497158 237978
rect 497214 237922 497282 237978
rect 497338 237922 497406 237978
rect 497462 237922 497558 237978
rect 496938 220350 497558 237922
rect 496938 220294 497034 220350
rect 497090 220294 497158 220350
rect 497214 220294 497282 220350
rect 497338 220294 497406 220350
rect 497462 220294 497558 220350
rect 496938 220226 497558 220294
rect 496938 220170 497034 220226
rect 497090 220170 497158 220226
rect 497214 220170 497282 220226
rect 497338 220170 497406 220226
rect 497462 220170 497558 220226
rect 496938 220102 497558 220170
rect 496938 220046 497034 220102
rect 497090 220046 497158 220102
rect 497214 220046 497282 220102
rect 497338 220046 497406 220102
rect 497462 220046 497558 220102
rect 496938 219978 497558 220046
rect 496938 219922 497034 219978
rect 497090 219922 497158 219978
rect 497214 219922 497282 219978
rect 497338 219922 497406 219978
rect 497462 219922 497558 219978
rect 496938 202350 497558 219922
rect 496938 202294 497034 202350
rect 497090 202294 497158 202350
rect 497214 202294 497282 202350
rect 497338 202294 497406 202350
rect 497462 202294 497558 202350
rect 496938 202226 497558 202294
rect 496938 202170 497034 202226
rect 497090 202170 497158 202226
rect 497214 202170 497282 202226
rect 497338 202170 497406 202226
rect 497462 202170 497558 202226
rect 496938 202102 497558 202170
rect 496938 202046 497034 202102
rect 497090 202046 497158 202102
rect 497214 202046 497282 202102
rect 497338 202046 497406 202102
rect 497462 202046 497558 202102
rect 496938 201978 497558 202046
rect 496938 201922 497034 201978
rect 497090 201922 497158 201978
rect 497214 201922 497282 201978
rect 497338 201922 497406 201978
rect 497462 201922 497558 201978
rect 496938 184350 497558 201922
rect 496938 184294 497034 184350
rect 497090 184294 497158 184350
rect 497214 184294 497282 184350
rect 497338 184294 497406 184350
rect 497462 184294 497558 184350
rect 496938 184226 497558 184294
rect 496938 184170 497034 184226
rect 497090 184170 497158 184226
rect 497214 184170 497282 184226
rect 497338 184170 497406 184226
rect 497462 184170 497558 184226
rect 496938 184102 497558 184170
rect 496938 184046 497034 184102
rect 497090 184046 497158 184102
rect 497214 184046 497282 184102
rect 497338 184046 497406 184102
rect 497462 184046 497558 184102
rect 496938 183978 497558 184046
rect 496938 183922 497034 183978
rect 497090 183922 497158 183978
rect 497214 183922 497282 183978
rect 497338 183922 497406 183978
rect 497462 183922 497558 183978
rect 496938 166350 497558 183922
rect 496938 166294 497034 166350
rect 497090 166294 497158 166350
rect 497214 166294 497282 166350
rect 497338 166294 497406 166350
rect 497462 166294 497558 166350
rect 496938 166226 497558 166294
rect 496938 166170 497034 166226
rect 497090 166170 497158 166226
rect 497214 166170 497282 166226
rect 497338 166170 497406 166226
rect 497462 166170 497558 166226
rect 496938 166102 497558 166170
rect 496938 166046 497034 166102
rect 497090 166046 497158 166102
rect 497214 166046 497282 166102
rect 497338 166046 497406 166102
rect 497462 166046 497558 166102
rect 496938 165978 497558 166046
rect 496938 165922 497034 165978
rect 497090 165922 497158 165978
rect 497214 165922 497282 165978
rect 497338 165922 497406 165978
rect 497462 165922 497558 165978
rect 496938 148350 497558 165922
rect 496938 148294 497034 148350
rect 497090 148294 497158 148350
rect 497214 148294 497282 148350
rect 497338 148294 497406 148350
rect 497462 148294 497558 148350
rect 496938 148226 497558 148294
rect 496938 148170 497034 148226
rect 497090 148170 497158 148226
rect 497214 148170 497282 148226
rect 497338 148170 497406 148226
rect 497462 148170 497558 148226
rect 496938 148102 497558 148170
rect 496938 148046 497034 148102
rect 497090 148046 497158 148102
rect 497214 148046 497282 148102
rect 497338 148046 497406 148102
rect 497462 148046 497558 148102
rect 496938 147978 497558 148046
rect 496938 147922 497034 147978
rect 497090 147922 497158 147978
rect 497214 147922 497282 147978
rect 497338 147922 497406 147978
rect 497462 147922 497558 147978
rect 496938 130350 497558 147922
rect 496938 130294 497034 130350
rect 497090 130294 497158 130350
rect 497214 130294 497282 130350
rect 497338 130294 497406 130350
rect 497462 130294 497558 130350
rect 496938 130226 497558 130294
rect 496938 130170 497034 130226
rect 497090 130170 497158 130226
rect 497214 130170 497282 130226
rect 497338 130170 497406 130226
rect 497462 130170 497558 130226
rect 496938 130102 497558 130170
rect 496938 130046 497034 130102
rect 497090 130046 497158 130102
rect 497214 130046 497282 130102
rect 497338 130046 497406 130102
rect 497462 130046 497558 130102
rect 496938 129978 497558 130046
rect 496938 129922 497034 129978
rect 497090 129922 497158 129978
rect 497214 129922 497282 129978
rect 497338 129922 497406 129978
rect 497462 129922 497558 129978
rect 496938 112350 497558 129922
rect 496938 112294 497034 112350
rect 497090 112294 497158 112350
rect 497214 112294 497282 112350
rect 497338 112294 497406 112350
rect 497462 112294 497558 112350
rect 496938 112226 497558 112294
rect 496938 112170 497034 112226
rect 497090 112170 497158 112226
rect 497214 112170 497282 112226
rect 497338 112170 497406 112226
rect 497462 112170 497558 112226
rect 496938 112102 497558 112170
rect 496938 112046 497034 112102
rect 497090 112046 497158 112102
rect 497214 112046 497282 112102
rect 497338 112046 497406 112102
rect 497462 112046 497558 112102
rect 496938 111978 497558 112046
rect 496938 111922 497034 111978
rect 497090 111922 497158 111978
rect 497214 111922 497282 111978
rect 497338 111922 497406 111978
rect 497462 111922 497558 111978
rect 496938 94350 497558 111922
rect 496938 94294 497034 94350
rect 497090 94294 497158 94350
rect 497214 94294 497282 94350
rect 497338 94294 497406 94350
rect 497462 94294 497558 94350
rect 496938 94226 497558 94294
rect 496938 94170 497034 94226
rect 497090 94170 497158 94226
rect 497214 94170 497282 94226
rect 497338 94170 497406 94226
rect 497462 94170 497558 94226
rect 496938 94102 497558 94170
rect 496938 94046 497034 94102
rect 497090 94046 497158 94102
rect 497214 94046 497282 94102
rect 497338 94046 497406 94102
rect 497462 94046 497558 94102
rect 496938 93978 497558 94046
rect 496938 93922 497034 93978
rect 497090 93922 497158 93978
rect 497214 93922 497282 93978
rect 497338 93922 497406 93978
rect 497462 93922 497558 93978
rect 469938 82294 470034 82350
rect 470090 82294 470158 82350
rect 470214 82294 470282 82350
rect 470338 82294 470406 82350
rect 470462 82294 470558 82350
rect 469938 82226 470558 82294
rect 469938 82170 470034 82226
rect 470090 82170 470158 82226
rect 470214 82170 470282 82226
rect 470338 82170 470406 82226
rect 470462 82170 470558 82226
rect 469938 82102 470558 82170
rect 469938 82046 470034 82102
rect 470090 82046 470158 82102
rect 470214 82046 470282 82102
rect 470338 82046 470406 82102
rect 470462 82046 470558 82102
rect 469938 81978 470558 82046
rect 469938 81922 470034 81978
rect 470090 81922 470158 81978
rect 470214 81922 470282 81978
rect 470338 81922 470406 81978
rect 470462 81922 470558 81978
rect 469938 64350 470558 81922
rect 479808 82350 480128 82384
rect 479808 82294 479878 82350
rect 479934 82294 480002 82350
rect 480058 82294 480128 82350
rect 479808 82226 480128 82294
rect 479808 82170 479878 82226
rect 479934 82170 480002 82226
rect 480058 82170 480128 82226
rect 479808 82102 480128 82170
rect 479808 82046 479878 82102
rect 479934 82046 480002 82102
rect 480058 82046 480128 82102
rect 479808 81978 480128 82046
rect 479808 81922 479878 81978
rect 479934 81922 480002 81978
rect 480058 81922 480128 81978
rect 479808 81888 480128 81922
rect 495168 76350 495488 76384
rect 495168 76294 495238 76350
rect 495294 76294 495362 76350
rect 495418 76294 495488 76350
rect 495168 76226 495488 76294
rect 495168 76170 495238 76226
rect 495294 76170 495362 76226
rect 495418 76170 495488 76226
rect 495168 76102 495488 76170
rect 495168 76046 495238 76102
rect 495294 76046 495362 76102
rect 495418 76046 495488 76102
rect 495168 75978 495488 76046
rect 495168 75922 495238 75978
rect 495294 75922 495362 75978
rect 495418 75922 495488 75978
rect 495168 75888 495488 75922
rect 496938 76350 497558 93922
rect 496938 76294 497034 76350
rect 497090 76294 497158 76350
rect 497214 76294 497282 76350
rect 497338 76294 497406 76350
rect 497462 76294 497558 76350
rect 496938 76226 497558 76294
rect 496938 76170 497034 76226
rect 497090 76170 497158 76226
rect 497214 76170 497282 76226
rect 497338 76170 497406 76226
rect 497462 76170 497558 76226
rect 496938 76102 497558 76170
rect 496938 76046 497034 76102
rect 497090 76046 497158 76102
rect 497214 76046 497282 76102
rect 497338 76046 497406 76102
rect 497462 76046 497558 76102
rect 496938 75978 497558 76046
rect 496938 75922 497034 75978
rect 497090 75922 497158 75978
rect 497214 75922 497282 75978
rect 497338 75922 497406 75978
rect 497462 75922 497558 75978
rect 469938 64294 470034 64350
rect 470090 64294 470158 64350
rect 470214 64294 470282 64350
rect 470338 64294 470406 64350
rect 470462 64294 470558 64350
rect 469938 64226 470558 64294
rect 469938 64170 470034 64226
rect 470090 64170 470158 64226
rect 470214 64170 470282 64226
rect 470338 64170 470406 64226
rect 470462 64170 470558 64226
rect 469938 64102 470558 64170
rect 469938 64046 470034 64102
rect 470090 64046 470158 64102
rect 470214 64046 470282 64102
rect 470338 64046 470406 64102
rect 470462 64046 470558 64102
rect 469938 63978 470558 64046
rect 469938 63922 470034 63978
rect 470090 63922 470158 63978
rect 470214 63922 470282 63978
rect 470338 63922 470406 63978
rect 470462 63922 470558 63978
rect 469938 46350 470558 63922
rect 479808 64350 480128 64384
rect 479808 64294 479878 64350
rect 479934 64294 480002 64350
rect 480058 64294 480128 64350
rect 479808 64226 480128 64294
rect 479808 64170 479878 64226
rect 479934 64170 480002 64226
rect 480058 64170 480128 64226
rect 479808 64102 480128 64170
rect 479808 64046 479878 64102
rect 479934 64046 480002 64102
rect 480058 64046 480128 64102
rect 479808 63978 480128 64046
rect 479808 63922 479878 63978
rect 479934 63922 480002 63978
rect 480058 63922 480128 63978
rect 479808 63888 480128 63922
rect 495168 58350 495488 58384
rect 495168 58294 495238 58350
rect 495294 58294 495362 58350
rect 495418 58294 495488 58350
rect 495168 58226 495488 58294
rect 495168 58170 495238 58226
rect 495294 58170 495362 58226
rect 495418 58170 495488 58226
rect 495168 58102 495488 58170
rect 495168 58046 495238 58102
rect 495294 58046 495362 58102
rect 495418 58046 495488 58102
rect 495168 57978 495488 58046
rect 495168 57922 495238 57978
rect 495294 57922 495362 57978
rect 495418 57922 495488 57978
rect 495168 57888 495488 57922
rect 496938 58350 497558 75922
rect 496938 58294 497034 58350
rect 497090 58294 497158 58350
rect 497214 58294 497282 58350
rect 497338 58294 497406 58350
rect 497462 58294 497558 58350
rect 496938 58226 497558 58294
rect 496938 58170 497034 58226
rect 497090 58170 497158 58226
rect 497214 58170 497282 58226
rect 497338 58170 497406 58226
rect 497462 58170 497558 58226
rect 496938 58102 497558 58170
rect 496938 58046 497034 58102
rect 497090 58046 497158 58102
rect 497214 58046 497282 58102
rect 497338 58046 497406 58102
rect 497462 58046 497558 58102
rect 496938 57978 497558 58046
rect 496938 57922 497034 57978
rect 497090 57922 497158 57978
rect 497214 57922 497282 57978
rect 497338 57922 497406 57978
rect 497462 57922 497558 57978
rect 469938 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 470558 46350
rect 469938 46226 470558 46294
rect 469938 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 470558 46226
rect 469938 46102 470558 46170
rect 469938 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 470558 46102
rect 469938 45978 470558 46046
rect 469938 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 470558 45978
rect 469938 28350 470558 45922
rect 469938 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 470558 28350
rect 469938 28226 470558 28294
rect 469938 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 470558 28226
rect 469938 28102 470558 28170
rect 469938 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 470558 28102
rect 469938 27978 470558 28046
rect 469938 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 470558 27978
rect 469938 10350 470558 27922
rect 496938 40350 497558 57922
rect 496938 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 497558 40350
rect 496938 40226 497558 40294
rect 496938 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 497558 40226
rect 496938 40102 497558 40170
rect 496938 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 497558 40102
rect 496938 39978 497558 40046
rect 496938 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 497558 39978
rect 473748 22350 474068 22384
rect 473748 22294 473818 22350
rect 473874 22294 473942 22350
rect 473998 22294 474068 22350
rect 473748 22226 474068 22294
rect 473748 22170 473818 22226
rect 473874 22170 473942 22226
rect 473998 22170 474068 22226
rect 473748 22102 474068 22170
rect 473748 22046 473818 22102
rect 473874 22046 473942 22102
rect 473998 22046 474068 22102
rect 473748 21978 474068 22046
rect 473748 21922 473818 21978
rect 473874 21922 473942 21978
rect 473998 21922 474068 21978
rect 473748 21888 474068 21922
rect 496938 22350 497558 39922
rect 496938 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 497558 22350
rect 496938 22226 497558 22294
rect 496938 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 497558 22226
rect 496938 22102 497558 22170
rect 496938 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 497558 22102
rect 496938 21978 497558 22046
rect 496938 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 497558 21978
rect 469938 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 470558 10350
rect 469938 10226 470558 10294
rect 469938 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 470558 10226
rect 469938 10102 470558 10170
rect 469938 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 470558 10102
rect 469938 9978 470558 10046
rect 469938 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 470558 9978
rect 469938 -1120 470558 9922
rect 475468 5338 475524 5348
rect 475468 3332 475524 5282
rect 494956 5158 495012 5168
rect 494956 3444 495012 5102
rect 494956 3378 495012 3388
rect 496938 4350 497558 21922
rect 500658 598172 501278 598268
rect 500658 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 501278 598172
rect 500658 598048 501278 598116
rect 500658 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 501278 598048
rect 500658 597924 501278 597992
rect 500658 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 501278 597924
rect 500658 597800 501278 597868
rect 500658 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 501278 597800
rect 500658 586350 501278 597744
rect 500658 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 501278 586350
rect 500658 586226 501278 586294
rect 500658 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 501278 586226
rect 500658 586102 501278 586170
rect 500658 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 501278 586102
rect 500658 585978 501278 586046
rect 500658 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 501278 585978
rect 500658 568350 501278 585922
rect 500658 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 501278 568350
rect 500658 568226 501278 568294
rect 500658 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 501278 568226
rect 500658 568102 501278 568170
rect 500658 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 501278 568102
rect 500658 567978 501278 568046
rect 500658 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 501278 567978
rect 500658 550350 501278 567922
rect 500658 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 501278 550350
rect 500658 550226 501278 550294
rect 500658 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 501278 550226
rect 500658 550102 501278 550170
rect 500658 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 501278 550102
rect 500658 549978 501278 550046
rect 500658 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 501278 549978
rect 500658 532350 501278 549922
rect 500658 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 501278 532350
rect 500658 532226 501278 532294
rect 500658 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 501278 532226
rect 500658 532102 501278 532170
rect 500658 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 501278 532102
rect 500658 531978 501278 532046
rect 500658 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 501278 531978
rect 500658 514350 501278 531922
rect 500658 514294 500754 514350
rect 500810 514294 500878 514350
rect 500934 514294 501002 514350
rect 501058 514294 501126 514350
rect 501182 514294 501278 514350
rect 500658 514226 501278 514294
rect 500658 514170 500754 514226
rect 500810 514170 500878 514226
rect 500934 514170 501002 514226
rect 501058 514170 501126 514226
rect 501182 514170 501278 514226
rect 500658 514102 501278 514170
rect 500658 514046 500754 514102
rect 500810 514046 500878 514102
rect 500934 514046 501002 514102
rect 501058 514046 501126 514102
rect 501182 514046 501278 514102
rect 500658 513978 501278 514046
rect 500658 513922 500754 513978
rect 500810 513922 500878 513978
rect 500934 513922 501002 513978
rect 501058 513922 501126 513978
rect 501182 513922 501278 513978
rect 500658 496350 501278 513922
rect 500658 496294 500754 496350
rect 500810 496294 500878 496350
rect 500934 496294 501002 496350
rect 501058 496294 501126 496350
rect 501182 496294 501278 496350
rect 500658 496226 501278 496294
rect 500658 496170 500754 496226
rect 500810 496170 500878 496226
rect 500934 496170 501002 496226
rect 501058 496170 501126 496226
rect 501182 496170 501278 496226
rect 500658 496102 501278 496170
rect 500658 496046 500754 496102
rect 500810 496046 500878 496102
rect 500934 496046 501002 496102
rect 501058 496046 501126 496102
rect 501182 496046 501278 496102
rect 500658 495978 501278 496046
rect 500658 495922 500754 495978
rect 500810 495922 500878 495978
rect 500934 495922 501002 495978
rect 501058 495922 501126 495978
rect 501182 495922 501278 495978
rect 500658 478350 501278 495922
rect 500658 478294 500754 478350
rect 500810 478294 500878 478350
rect 500934 478294 501002 478350
rect 501058 478294 501126 478350
rect 501182 478294 501278 478350
rect 500658 478226 501278 478294
rect 500658 478170 500754 478226
rect 500810 478170 500878 478226
rect 500934 478170 501002 478226
rect 501058 478170 501126 478226
rect 501182 478170 501278 478226
rect 500658 478102 501278 478170
rect 500658 478046 500754 478102
rect 500810 478046 500878 478102
rect 500934 478046 501002 478102
rect 501058 478046 501126 478102
rect 501182 478046 501278 478102
rect 500658 477978 501278 478046
rect 500658 477922 500754 477978
rect 500810 477922 500878 477978
rect 500934 477922 501002 477978
rect 501058 477922 501126 477978
rect 501182 477922 501278 477978
rect 500658 460350 501278 477922
rect 500658 460294 500754 460350
rect 500810 460294 500878 460350
rect 500934 460294 501002 460350
rect 501058 460294 501126 460350
rect 501182 460294 501278 460350
rect 500658 460226 501278 460294
rect 500658 460170 500754 460226
rect 500810 460170 500878 460226
rect 500934 460170 501002 460226
rect 501058 460170 501126 460226
rect 501182 460170 501278 460226
rect 500658 460102 501278 460170
rect 500658 460046 500754 460102
rect 500810 460046 500878 460102
rect 500934 460046 501002 460102
rect 501058 460046 501126 460102
rect 501182 460046 501278 460102
rect 500658 459978 501278 460046
rect 500658 459922 500754 459978
rect 500810 459922 500878 459978
rect 500934 459922 501002 459978
rect 501058 459922 501126 459978
rect 501182 459922 501278 459978
rect 500658 442350 501278 459922
rect 500658 442294 500754 442350
rect 500810 442294 500878 442350
rect 500934 442294 501002 442350
rect 501058 442294 501126 442350
rect 501182 442294 501278 442350
rect 500658 442226 501278 442294
rect 500658 442170 500754 442226
rect 500810 442170 500878 442226
rect 500934 442170 501002 442226
rect 501058 442170 501126 442226
rect 501182 442170 501278 442226
rect 500658 442102 501278 442170
rect 500658 442046 500754 442102
rect 500810 442046 500878 442102
rect 500934 442046 501002 442102
rect 501058 442046 501126 442102
rect 501182 442046 501278 442102
rect 500658 441978 501278 442046
rect 500658 441922 500754 441978
rect 500810 441922 500878 441978
rect 500934 441922 501002 441978
rect 501058 441922 501126 441978
rect 501182 441922 501278 441978
rect 500658 424350 501278 441922
rect 500658 424294 500754 424350
rect 500810 424294 500878 424350
rect 500934 424294 501002 424350
rect 501058 424294 501126 424350
rect 501182 424294 501278 424350
rect 500658 424226 501278 424294
rect 500658 424170 500754 424226
rect 500810 424170 500878 424226
rect 500934 424170 501002 424226
rect 501058 424170 501126 424226
rect 501182 424170 501278 424226
rect 500658 424102 501278 424170
rect 500658 424046 500754 424102
rect 500810 424046 500878 424102
rect 500934 424046 501002 424102
rect 501058 424046 501126 424102
rect 501182 424046 501278 424102
rect 500658 423978 501278 424046
rect 500658 423922 500754 423978
rect 500810 423922 500878 423978
rect 500934 423922 501002 423978
rect 501058 423922 501126 423978
rect 501182 423922 501278 423978
rect 500658 406350 501278 423922
rect 500658 406294 500754 406350
rect 500810 406294 500878 406350
rect 500934 406294 501002 406350
rect 501058 406294 501126 406350
rect 501182 406294 501278 406350
rect 500658 406226 501278 406294
rect 500658 406170 500754 406226
rect 500810 406170 500878 406226
rect 500934 406170 501002 406226
rect 501058 406170 501126 406226
rect 501182 406170 501278 406226
rect 500658 406102 501278 406170
rect 500658 406046 500754 406102
rect 500810 406046 500878 406102
rect 500934 406046 501002 406102
rect 501058 406046 501126 406102
rect 501182 406046 501278 406102
rect 500658 405978 501278 406046
rect 500658 405922 500754 405978
rect 500810 405922 500878 405978
rect 500934 405922 501002 405978
rect 501058 405922 501126 405978
rect 501182 405922 501278 405978
rect 500658 388350 501278 405922
rect 527658 597212 528278 598268
rect 527658 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 528278 597212
rect 527658 597088 528278 597156
rect 527658 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 528278 597088
rect 527658 596964 528278 597032
rect 527658 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 528278 596964
rect 527658 596840 528278 596908
rect 527658 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 528278 596840
rect 527658 580350 528278 596784
rect 527658 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 528278 580350
rect 527658 580226 528278 580294
rect 527658 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 528278 580226
rect 527658 580102 528278 580170
rect 527658 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 528278 580102
rect 527658 579978 528278 580046
rect 527658 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 528278 579978
rect 527658 562350 528278 579922
rect 527658 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 528278 562350
rect 527658 562226 528278 562294
rect 527658 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 528278 562226
rect 527658 562102 528278 562170
rect 527658 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 528278 562102
rect 527658 561978 528278 562046
rect 527658 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 528278 561978
rect 527658 544350 528278 561922
rect 527658 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 528278 544350
rect 527658 544226 528278 544294
rect 527658 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 528278 544226
rect 527658 544102 528278 544170
rect 527658 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 528278 544102
rect 527658 543978 528278 544046
rect 527658 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 528278 543978
rect 527658 526350 528278 543922
rect 527658 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 528278 526350
rect 527658 526226 528278 526294
rect 527658 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 528278 526226
rect 527658 526102 528278 526170
rect 527658 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 528278 526102
rect 527658 525978 528278 526046
rect 527658 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 528278 525978
rect 527658 508350 528278 525922
rect 527658 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 528278 508350
rect 527658 508226 528278 508294
rect 527658 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 528278 508226
rect 527658 508102 528278 508170
rect 527658 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 528278 508102
rect 527658 507978 528278 508046
rect 527658 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 528278 507978
rect 527658 490350 528278 507922
rect 527658 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 528278 490350
rect 527658 490226 528278 490294
rect 527658 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 528278 490226
rect 527658 490102 528278 490170
rect 527658 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 528278 490102
rect 527658 489978 528278 490046
rect 527658 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 528278 489978
rect 527658 472350 528278 489922
rect 527658 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 528278 472350
rect 527658 472226 528278 472294
rect 527658 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 528278 472226
rect 527658 472102 528278 472170
rect 527658 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 528278 472102
rect 527658 471978 528278 472046
rect 527658 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 528278 471978
rect 527658 454350 528278 471922
rect 527658 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 528278 454350
rect 527658 454226 528278 454294
rect 527658 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 528278 454226
rect 527658 454102 528278 454170
rect 527658 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 528278 454102
rect 527658 453978 528278 454046
rect 527658 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 528278 453978
rect 527658 436350 528278 453922
rect 527658 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 528278 436350
rect 527658 436226 528278 436294
rect 527658 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 528278 436226
rect 527658 436102 528278 436170
rect 527658 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 528278 436102
rect 527658 435978 528278 436046
rect 527658 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 528278 435978
rect 527658 418350 528278 435922
rect 527658 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 528278 418350
rect 527658 418226 528278 418294
rect 527658 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 528278 418226
rect 527658 418102 528278 418170
rect 527658 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 528278 418102
rect 527658 417978 528278 418046
rect 527658 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 528278 417978
rect 527658 400350 528278 417922
rect 527658 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 528278 400350
rect 527658 400226 528278 400294
rect 527658 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 528278 400226
rect 527658 400102 528278 400170
rect 527658 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 528278 400102
rect 527658 399978 528278 400046
rect 527658 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 528278 399978
rect 500658 388294 500754 388350
rect 500810 388294 500878 388350
rect 500934 388294 501002 388350
rect 501058 388294 501126 388350
rect 501182 388294 501278 388350
rect 500658 388226 501278 388294
rect 500658 388170 500754 388226
rect 500810 388170 500878 388226
rect 500934 388170 501002 388226
rect 501058 388170 501126 388226
rect 501182 388170 501278 388226
rect 500658 388102 501278 388170
rect 500658 388046 500754 388102
rect 500810 388046 500878 388102
rect 500934 388046 501002 388102
rect 501058 388046 501126 388102
rect 501182 388046 501278 388102
rect 500658 387978 501278 388046
rect 500658 387922 500754 387978
rect 500810 387922 500878 387978
rect 500934 387922 501002 387978
rect 501058 387922 501126 387978
rect 501182 387922 501278 387978
rect 500658 370350 501278 387922
rect 500658 370294 500754 370350
rect 500810 370294 500878 370350
rect 500934 370294 501002 370350
rect 501058 370294 501126 370350
rect 501182 370294 501278 370350
rect 500658 370226 501278 370294
rect 500658 370170 500754 370226
rect 500810 370170 500878 370226
rect 500934 370170 501002 370226
rect 501058 370170 501126 370226
rect 501182 370170 501278 370226
rect 500658 370102 501278 370170
rect 500658 370046 500754 370102
rect 500810 370046 500878 370102
rect 500934 370046 501002 370102
rect 501058 370046 501126 370102
rect 501182 370046 501278 370102
rect 500658 369978 501278 370046
rect 500658 369922 500754 369978
rect 500810 369922 500878 369978
rect 500934 369922 501002 369978
rect 501058 369922 501126 369978
rect 501182 369922 501278 369978
rect 500658 352350 501278 369922
rect 500658 352294 500754 352350
rect 500810 352294 500878 352350
rect 500934 352294 501002 352350
rect 501058 352294 501126 352350
rect 501182 352294 501278 352350
rect 500658 352226 501278 352294
rect 500658 352170 500754 352226
rect 500810 352170 500878 352226
rect 500934 352170 501002 352226
rect 501058 352170 501126 352226
rect 501182 352170 501278 352226
rect 500658 352102 501278 352170
rect 500658 352046 500754 352102
rect 500810 352046 500878 352102
rect 500934 352046 501002 352102
rect 501058 352046 501126 352102
rect 501182 352046 501278 352102
rect 500658 351978 501278 352046
rect 500658 351922 500754 351978
rect 500810 351922 500878 351978
rect 500934 351922 501002 351978
rect 501058 351922 501126 351978
rect 501182 351922 501278 351978
rect 500658 334350 501278 351922
rect 500658 334294 500754 334350
rect 500810 334294 500878 334350
rect 500934 334294 501002 334350
rect 501058 334294 501126 334350
rect 501182 334294 501278 334350
rect 500658 334226 501278 334294
rect 500658 334170 500754 334226
rect 500810 334170 500878 334226
rect 500934 334170 501002 334226
rect 501058 334170 501126 334226
rect 501182 334170 501278 334226
rect 500658 334102 501278 334170
rect 500658 334046 500754 334102
rect 500810 334046 500878 334102
rect 500934 334046 501002 334102
rect 501058 334046 501126 334102
rect 501182 334046 501278 334102
rect 500658 333978 501278 334046
rect 500658 333922 500754 333978
rect 500810 333922 500878 333978
rect 500934 333922 501002 333978
rect 501058 333922 501126 333978
rect 501182 333922 501278 333978
rect 500658 316350 501278 333922
rect 500658 316294 500754 316350
rect 500810 316294 500878 316350
rect 500934 316294 501002 316350
rect 501058 316294 501126 316350
rect 501182 316294 501278 316350
rect 500658 316226 501278 316294
rect 500658 316170 500754 316226
rect 500810 316170 500878 316226
rect 500934 316170 501002 316226
rect 501058 316170 501126 316226
rect 501182 316170 501278 316226
rect 500658 316102 501278 316170
rect 500658 316046 500754 316102
rect 500810 316046 500878 316102
rect 500934 316046 501002 316102
rect 501058 316046 501126 316102
rect 501182 316046 501278 316102
rect 500658 315978 501278 316046
rect 500658 315922 500754 315978
rect 500810 315922 500878 315978
rect 500934 315922 501002 315978
rect 501058 315922 501126 315978
rect 501182 315922 501278 315978
rect 500658 298350 501278 315922
rect 500658 298294 500754 298350
rect 500810 298294 500878 298350
rect 500934 298294 501002 298350
rect 501058 298294 501126 298350
rect 501182 298294 501278 298350
rect 500658 298226 501278 298294
rect 500658 298170 500754 298226
rect 500810 298170 500878 298226
rect 500934 298170 501002 298226
rect 501058 298170 501126 298226
rect 501182 298170 501278 298226
rect 500658 298102 501278 298170
rect 500658 298046 500754 298102
rect 500810 298046 500878 298102
rect 500934 298046 501002 298102
rect 501058 298046 501126 298102
rect 501182 298046 501278 298102
rect 500658 297978 501278 298046
rect 500658 297922 500754 297978
rect 500810 297922 500878 297978
rect 500934 297922 501002 297978
rect 501058 297922 501126 297978
rect 501182 297922 501278 297978
rect 500658 280350 501278 297922
rect 500658 280294 500754 280350
rect 500810 280294 500878 280350
rect 500934 280294 501002 280350
rect 501058 280294 501126 280350
rect 501182 280294 501278 280350
rect 500658 280226 501278 280294
rect 500658 280170 500754 280226
rect 500810 280170 500878 280226
rect 500934 280170 501002 280226
rect 501058 280170 501126 280226
rect 501182 280170 501278 280226
rect 500658 280102 501278 280170
rect 500658 280046 500754 280102
rect 500810 280046 500878 280102
rect 500934 280046 501002 280102
rect 501058 280046 501126 280102
rect 501182 280046 501278 280102
rect 500658 279978 501278 280046
rect 500658 279922 500754 279978
rect 500810 279922 500878 279978
rect 500934 279922 501002 279978
rect 501058 279922 501126 279978
rect 501182 279922 501278 279978
rect 500658 262350 501278 279922
rect 500658 262294 500754 262350
rect 500810 262294 500878 262350
rect 500934 262294 501002 262350
rect 501058 262294 501126 262350
rect 501182 262294 501278 262350
rect 500658 262226 501278 262294
rect 500658 262170 500754 262226
rect 500810 262170 500878 262226
rect 500934 262170 501002 262226
rect 501058 262170 501126 262226
rect 501182 262170 501278 262226
rect 500658 262102 501278 262170
rect 500658 262046 500754 262102
rect 500810 262046 500878 262102
rect 500934 262046 501002 262102
rect 501058 262046 501126 262102
rect 501182 262046 501278 262102
rect 500658 261978 501278 262046
rect 500658 261922 500754 261978
rect 500810 261922 500878 261978
rect 500934 261922 501002 261978
rect 501058 261922 501126 261978
rect 501182 261922 501278 261978
rect 500658 244350 501278 261922
rect 500658 244294 500754 244350
rect 500810 244294 500878 244350
rect 500934 244294 501002 244350
rect 501058 244294 501126 244350
rect 501182 244294 501278 244350
rect 500658 244226 501278 244294
rect 500658 244170 500754 244226
rect 500810 244170 500878 244226
rect 500934 244170 501002 244226
rect 501058 244170 501126 244226
rect 501182 244170 501278 244226
rect 500658 244102 501278 244170
rect 500658 244046 500754 244102
rect 500810 244046 500878 244102
rect 500934 244046 501002 244102
rect 501058 244046 501126 244102
rect 501182 244046 501278 244102
rect 500658 243978 501278 244046
rect 500658 243922 500754 243978
rect 500810 243922 500878 243978
rect 500934 243922 501002 243978
rect 501058 243922 501126 243978
rect 501182 243922 501278 243978
rect 500658 226350 501278 243922
rect 500658 226294 500754 226350
rect 500810 226294 500878 226350
rect 500934 226294 501002 226350
rect 501058 226294 501126 226350
rect 501182 226294 501278 226350
rect 500658 226226 501278 226294
rect 500658 226170 500754 226226
rect 500810 226170 500878 226226
rect 500934 226170 501002 226226
rect 501058 226170 501126 226226
rect 501182 226170 501278 226226
rect 500658 226102 501278 226170
rect 500658 226046 500754 226102
rect 500810 226046 500878 226102
rect 500934 226046 501002 226102
rect 501058 226046 501126 226102
rect 501182 226046 501278 226102
rect 500658 225978 501278 226046
rect 500658 225922 500754 225978
rect 500810 225922 500878 225978
rect 500934 225922 501002 225978
rect 501058 225922 501126 225978
rect 501182 225922 501278 225978
rect 500658 208350 501278 225922
rect 500658 208294 500754 208350
rect 500810 208294 500878 208350
rect 500934 208294 501002 208350
rect 501058 208294 501126 208350
rect 501182 208294 501278 208350
rect 500658 208226 501278 208294
rect 500658 208170 500754 208226
rect 500810 208170 500878 208226
rect 500934 208170 501002 208226
rect 501058 208170 501126 208226
rect 501182 208170 501278 208226
rect 500658 208102 501278 208170
rect 500658 208046 500754 208102
rect 500810 208046 500878 208102
rect 500934 208046 501002 208102
rect 501058 208046 501126 208102
rect 501182 208046 501278 208102
rect 500658 207978 501278 208046
rect 500658 207922 500754 207978
rect 500810 207922 500878 207978
rect 500934 207922 501002 207978
rect 501058 207922 501126 207978
rect 501182 207922 501278 207978
rect 500658 190350 501278 207922
rect 500658 190294 500754 190350
rect 500810 190294 500878 190350
rect 500934 190294 501002 190350
rect 501058 190294 501126 190350
rect 501182 190294 501278 190350
rect 500658 190226 501278 190294
rect 500658 190170 500754 190226
rect 500810 190170 500878 190226
rect 500934 190170 501002 190226
rect 501058 190170 501126 190226
rect 501182 190170 501278 190226
rect 500658 190102 501278 190170
rect 500658 190046 500754 190102
rect 500810 190046 500878 190102
rect 500934 190046 501002 190102
rect 501058 190046 501126 190102
rect 501182 190046 501278 190102
rect 500658 189978 501278 190046
rect 500658 189922 500754 189978
rect 500810 189922 500878 189978
rect 500934 189922 501002 189978
rect 501058 189922 501126 189978
rect 501182 189922 501278 189978
rect 500658 172350 501278 189922
rect 500658 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 501278 172350
rect 500658 172226 501278 172294
rect 500658 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 501278 172226
rect 500658 172102 501278 172170
rect 500658 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 501278 172102
rect 500658 171978 501278 172046
rect 500658 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 501278 171978
rect 500658 154350 501278 171922
rect 500658 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 501278 154350
rect 500658 154226 501278 154294
rect 500658 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 501278 154226
rect 500658 154102 501278 154170
rect 500658 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 501278 154102
rect 500658 153978 501278 154046
rect 500658 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 501278 153978
rect 500658 136350 501278 153922
rect 500658 136294 500754 136350
rect 500810 136294 500878 136350
rect 500934 136294 501002 136350
rect 501058 136294 501126 136350
rect 501182 136294 501278 136350
rect 500658 136226 501278 136294
rect 500658 136170 500754 136226
rect 500810 136170 500878 136226
rect 500934 136170 501002 136226
rect 501058 136170 501126 136226
rect 501182 136170 501278 136226
rect 500658 136102 501278 136170
rect 500658 136046 500754 136102
rect 500810 136046 500878 136102
rect 500934 136046 501002 136102
rect 501058 136046 501126 136102
rect 501182 136046 501278 136102
rect 500658 135978 501278 136046
rect 500658 135922 500754 135978
rect 500810 135922 500878 135978
rect 500934 135922 501002 135978
rect 501058 135922 501126 135978
rect 501182 135922 501278 135978
rect 500658 118350 501278 135922
rect 500658 118294 500754 118350
rect 500810 118294 500878 118350
rect 500934 118294 501002 118350
rect 501058 118294 501126 118350
rect 501182 118294 501278 118350
rect 500658 118226 501278 118294
rect 500658 118170 500754 118226
rect 500810 118170 500878 118226
rect 500934 118170 501002 118226
rect 501058 118170 501126 118226
rect 501182 118170 501278 118226
rect 500658 118102 501278 118170
rect 500658 118046 500754 118102
rect 500810 118046 500878 118102
rect 500934 118046 501002 118102
rect 501058 118046 501126 118102
rect 501182 118046 501278 118102
rect 500658 117978 501278 118046
rect 500658 117922 500754 117978
rect 500810 117922 500878 117978
rect 500934 117922 501002 117978
rect 501058 117922 501126 117978
rect 501182 117922 501278 117978
rect 500658 100350 501278 117922
rect 500658 100294 500754 100350
rect 500810 100294 500878 100350
rect 500934 100294 501002 100350
rect 501058 100294 501126 100350
rect 501182 100294 501278 100350
rect 500658 100226 501278 100294
rect 500658 100170 500754 100226
rect 500810 100170 500878 100226
rect 500934 100170 501002 100226
rect 501058 100170 501126 100226
rect 501182 100170 501278 100226
rect 500658 100102 501278 100170
rect 500658 100046 500754 100102
rect 500810 100046 500878 100102
rect 500934 100046 501002 100102
rect 501058 100046 501126 100102
rect 501182 100046 501278 100102
rect 500658 99978 501278 100046
rect 500658 99922 500754 99978
rect 500810 99922 500878 99978
rect 500934 99922 501002 99978
rect 501058 99922 501126 99978
rect 501182 99922 501278 99978
rect 500658 82350 501278 99922
rect 500658 82294 500754 82350
rect 500810 82294 500878 82350
rect 500934 82294 501002 82350
rect 501058 82294 501126 82350
rect 501182 82294 501278 82350
rect 500658 82226 501278 82294
rect 500658 82170 500754 82226
rect 500810 82170 500878 82226
rect 500934 82170 501002 82226
rect 501058 82170 501126 82226
rect 501182 82170 501278 82226
rect 500658 82102 501278 82170
rect 500658 82046 500754 82102
rect 500810 82046 500878 82102
rect 500934 82046 501002 82102
rect 501058 82046 501126 82102
rect 501182 82046 501278 82102
rect 500658 81978 501278 82046
rect 500658 81922 500754 81978
rect 500810 81922 500878 81978
rect 500934 81922 501002 81978
rect 501058 81922 501126 81978
rect 501182 81922 501278 81978
rect 500658 64350 501278 81922
rect 513212 390404 513268 390414
rect 513212 70644 513268 390348
rect 513212 70578 513268 70588
rect 527658 382350 528278 399922
rect 527658 382294 527754 382350
rect 527810 382294 527878 382350
rect 527934 382294 528002 382350
rect 528058 382294 528126 382350
rect 528182 382294 528278 382350
rect 527658 382226 528278 382294
rect 527658 382170 527754 382226
rect 527810 382170 527878 382226
rect 527934 382170 528002 382226
rect 528058 382170 528126 382226
rect 528182 382170 528278 382226
rect 527658 382102 528278 382170
rect 527658 382046 527754 382102
rect 527810 382046 527878 382102
rect 527934 382046 528002 382102
rect 528058 382046 528126 382102
rect 528182 382046 528278 382102
rect 527658 381978 528278 382046
rect 527658 381922 527754 381978
rect 527810 381922 527878 381978
rect 527934 381922 528002 381978
rect 528058 381922 528126 381978
rect 528182 381922 528278 381978
rect 527658 364350 528278 381922
rect 527658 364294 527754 364350
rect 527810 364294 527878 364350
rect 527934 364294 528002 364350
rect 528058 364294 528126 364350
rect 528182 364294 528278 364350
rect 527658 364226 528278 364294
rect 527658 364170 527754 364226
rect 527810 364170 527878 364226
rect 527934 364170 528002 364226
rect 528058 364170 528126 364226
rect 528182 364170 528278 364226
rect 527658 364102 528278 364170
rect 527658 364046 527754 364102
rect 527810 364046 527878 364102
rect 527934 364046 528002 364102
rect 528058 364046 528126 364102
rect 528182 364046 528278 364102
rect 527658 363978 528278 364046
rect 527658 363922 527754 363978
rect 527810 363922 527878 363978
rect 527934 363922 528002 363978
rect 528058 363922 528126 363978
rect 528182 363922 528278 363978
rect 527658 346350 528278 363922
rect 527658 346294 527754 346350
rect 527810 346294 527878 346350
rect 527934 346294 528002 346350
rect 528058 346294 528126 346350
rect 528182 346294 528278 346350
rect 527658 346226 528278 346294
rect 527658 346170 527754 346226
rect 527810 346170 527878 346226
rect 527934 346170 528002 346226
rect 528058 346170 528126 346226
rect 528182 346170 528278 346226
rect 527658 346102 528278 346170
rect 527658 346046 527754 346102
rect 527810 346046 527878 346102
rect 527934 346046 528002 346102
rect 528058 346046 528126 346102
rect 528182 346046 528278 346102
rect 527658 345978 528278 346046
rect 527658 345922 527754 345978
rect 527810 345922 527878 345978
rect 527934 345922 528002 345978
rect 528058 345922 528126 345978
rect 528182 345922 528278 345978
rect 527658 328350 528278 345922
rect 527658 328294 527754 328350
rect 527810 328294 527878 328350
rect 527934 328294 528002 328350
rect 528058 328294 528126 328350
rect 528182 328294 528278 328350
rect 527658 328226 528278 328294
rect 527658 328170 527754 328226
rect 527810 328170 527878 328226
rect 527934 328170 528002 328226
rect 528058 328170 528126 328226
rect 528182 328170 528278 328226
rect 527658 328102 528278 328170
rect 527658 328046 527754 328102
rect 527810 328046 527878 328102
rect 527934 328046 528002 328102
rect 528058 328046 528126 328102
rect 528182 328046 528278 328102
rect 527658 327978 528278 328046
rect 527658 327922 527754 327978
rect 527810 327922 527878 327978
rect 527934 327922 528002 327978
rect 528058 327922 528126 327978
rect 528182 327922 528278 327978
rect 527658 310350 528278 327922
rect 527658 310294 527754 310350
rect 527810 310294 527878 310350
rect 527934 310294 528002 310350
rect 528058 310294 528126 310350
rect 528182 310294 528278 310350
rect 527658 310226 528278 310294
rect 527658 310170 527754 310226
rect 527810 310170 527878 310226
rect 527934 310170 528002 310226
rect 528058 310170 528126 310226
rect 528182 310170 528278 310226
rect 527658 310102 528278 310170
rect 527658 310046 527754 310102
rect 527810 310046 527878 310102
rect 527934 310046 528002 310102
rect 528058 310046 528126 310102
rect 528182 310046 528278 310102
rect 527658 309978 528278 310046
rect 527658 309922 527754 309978
rect 527810 309922 527878 309978
rect 527934 309922 528002 309978
rect 528058 309922 528126 309978
rect 528182 309922 528278 309978
rect 527658 292350 528278 309922
rect 527658 292294 527754 292350
rect 527810 292294 527878 292350
rect 527934 292294 528002 292350
rect 528058 292294 528126 292350
rect 528182 292294 528278 292350
rect 527658 292226 528278 292294
rect 527658 292170 527754 292226
rect 527810 292170 527878 292226
rect 527934 292170 528002 292226
rect 528058 292170 528126 292226
rect 528182 292170 528278 292226
rect 527658 292102 528278 292170
rect 527658 292046 527754 292102
rect 527810 292046 527878 292102
rect 527934 292046 528002 292102
rect 528058 292046 528126 292102
rect 528182 292046 528278 292102
rect 527658 291978 528278 292046
rect 527658 291922 527754 291978
rect 527810 291922 527878 291978
rect 527934 291922 528002 291978
rect 528058 291922 528126 291978
rect 528182 291922 528278 291978
rect 527658 274350 528278 291922
rect 531378 598172 531998 598268
rect 531378 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 531998 598172
rect 531378 598048 531998 598116
rect 531378 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 531998 598048
rect 531378 597924 531998 597992
rect 531378 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 531998 597924
rect 531378 597800 531998 597868
rect 531378 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 531998 597800
rect 531378 586350 531998 597744
rect 531378 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 531998 586350
rect 531378 586226 531998 586294
rect 531378 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 531998 586226
rect 531378 586102 531998 586170
rect 531378 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 531998 586102
rect 531378 585978 531998 586046
rect 531378 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 531998 585978
rect 531378 568350 531998 585922
rect 531378 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 531998 568350
rect 531378 568226 531998 568294
rect 531378 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 531998 568226
rect 531378 568102 531998 568170
rect 531378 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 531998 568102
rect 531378 567978 531998 568046
rect 531378 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 531998 567978
rect 531378 550350 531998 567922
rect 531378 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 531998 550350
rect 531378 550226 531998 550294
rect 531378 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 531998 550226
rect 531378 550102 531998 550170
rect 531378 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 531998 550102
rect 531378 549978 531998 550046
rect 531378 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 531998 549978
rect 531378 532350 531998 549922
rect 531378 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 531998 532350
rect 531378 532226 531998 532294
rect 531378 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 531998 532226
rect 531378 532102 531998 532170
rect 531378 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 531998 532102
rect 531378 531978 531998 532046
rect 531378 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 531998 531978
rect 531378 514350 531998 531922
rect 531378 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 531998 514350
rect 531378 514226 531998 514294
rect 531378 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 531998 514226
rect 531378 514102 531998 514170
rect 531378 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 531998 514102
rect 531378 513978 531998 514046
rect 531378 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 531998 513978
rect 531378 496350 531998 513922
rect 531378 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 531998 496350
rect 531378 496226 531998 496294
rect 531378 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 531998 496226
rect 531378 496102 531998 496170
rect 531378 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 531998 496102
rect 531378 495978 531998 496046
rect 531378 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 531998 495978
rect 531378 478350 531998 495922
rect 531378 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 531998 478350
rect 531378 478226 531998 478294
rect 531378 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 531998 478226
rect 531378 478102 531998 478170
rect 531378 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 531998 478102
rect 531378 477978 531998 478046
rect 531378 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 531998 477978
rect 531378 460350 531998 477922
rect 531378 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 531998 460350
rect 531378 460226 531998 460294
rect 531378 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 531998 460226
rect 531378 460102 531998 460170
rect 531378 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 531998 460102
rect 531378 459978 531998 460046
rect 531378 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 531998 459978
rect 531378 442350 531998 459922
rect 531378 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 531998 442350
rect 531378 442226 531998 442294
rect 531378 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 531998 442226
rect 531378 442102 531998 442170
rect 531378 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 531998 442102
rect 531378 441978 531998 442046
rect 531378 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 531998 441978
rect 531378 424350 531998 441922
rect 531378 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 531998 424350
rect 531378 424226 531998 424294
rect 531378 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 531998 424226
rect 531378 424102 531998 424170
rect 531378 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 531998 424102
rect 531378 423978 531998 424046
rect 531378 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 531998 423978
rect 531378 406350 531998 423922
rect 531378 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 531998 406350
rect 531378 406226 531998 406294
rect 531378 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 531998 406226
rect 531378 406102 531998 406170
rect 531378 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 531998 406102
rect 531378 405978 531998 406046
rect 531378 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 531998 405978
rect 531378 388350 531998 405922
rect 531378 388294 531474 388350
rect 531530 388294 531598 388350
rect 531654 388294 531722 388350
rect 531778 388294 531846 388350
rect 531902 388294 531998 388350
rect 531378 388226 531998 388294
rect 531378 388170 531474 388226
rect 531530 388170 531598 388226
rect 531654 388170 531722 388226
rect 531778 388170 531846 388226
rect 531902 388170 531998 388226
rect 531378 388102 531998 388170
rect 531378 388046 531474 388102
rect 531530 388046 531598 388102
rect 531654 388046 531722 388102
rect 531778 388046 531846 388102
rect 531902 388046 531998 388102
rect 531378 387978 531998 388046
rect 531378 387922 531474 387978
rect 531530 387922 531598 387978
rect 531654 387922 531722 387978
rect 531778 387922 531846 387978
rect 531902 387922 531998 387978
rect 531378 370350 531998 387922
rect 531378 370294 531474 370350
rect 531530 370294 531598 370350
rect 531654 370294 531722 370350
rect 531778 370294 531846 370350
rect 531902 370294 531998 370350
rect 531378 370226 531998 370294
rect 531378 370170 531474 370226
rect 531530 370170 531598 370226
rect 531654 370170 531722 370226
rect 531778 370170 531846 370226
rect 531902 370170 531998 370226
rect 531378 370102 531998 370170
rect 531378 370046 531474 370102
rect 531530 370046 531598 370102
rect 531654 370046 531722 370102
rect 531778 370046 531846 370102
rect 531902 370046 531998 370102
rect 531378 369978 531998 370046
rect 531378 369922 531474 369978
rect 531530 369922 531598 369978
rect 531654 369922 531722 369978
rect 531778 369922 531846 369978
rect 531902 369922 531998 369978
rect 531378 352350 531998 369922
rect 531378 352294 531474 352350
rect 531530 352294 531598 352350
rect 531654 352294 531722 352350
rect 531778 352294 531846 352350
rect 531902 352294 531998 352350
rect 531378 352226 531998 352294
rect 531378 352170 531474 352226
rect 531530 352170 531598 352226
rect 531654 352170 531722 352226
rect 531778 352170 531846 352226
rect 531902 352170 531998 352226
rect 531378 352102 531998 352170
rect 531378 352046 531474 352102
rect 531530 352046 531598 352102
rect 531654 352046 531722 352102
rect 531778 352046 531846 352102
rect 531902 352046 531998 352102
rect 531378 351978 531998 352046
rect 531378 351922 531474 351978
rect 531530 351922 531598 351978
rect 531654 351922 531722 351978
rect 531778 351922 531846 351978
rect 531902 351922 531998 351978
rect 531378 334350 531998 351922
rect 531378 334294 531474 334350
rect 531530 334294 531598 334350
rect 531654 334294 531722 334350
rect 531778 334294 531846 334350
rect 531902 334294 531998 334350
rect 531378 334226 531998 334294
rect 531378 334170 531474 334226
rect 531530 334170 531598 334226
rect 531654 334170 531722 334226
rect 531778 334170 531846 334226
rect 531902 334170 531998 334226
rect 531378 334102 531998 334170
rect 531378 334046 531474 334102
rect 531530 334046 531598 334102
rect 531654 334046 531722 334102
rect 531778 334046 531846 334102
rect 531902 334046 531998 334102
rect 531378 333978 531998 334046
rect 531378 333922 531474 333978
rect 531530 333922 531598 333978
rect 531654 333922 531722 333978
rect 531778 333922 531846 333978
rect 531902 333922 531998 333978
rect 531378 316350 531998 333922
rect 531378 316294 531474 316350
rect 531530 316294 531598 316350
rect 531654 316294 531722 316350
rect 531778 316294 531846 316350
rect 531902 316294 531998 316350
rect 531378 316226 531998 316294
rect 531378 316170 531474 316226
rect 531530 316170 531598 316226
rect 531654 316170 531722 316226
rect 531778 316170 531846 316226
rect 531902 316170 531998 316226
rect 531378 316102 531998 316170
rect 531378 316046 531474 316102
rect 531530 316046 531598 316102
rect 531654 316046 531722 316102
rect 531778 316046 531846 316102
rect 531902 316046 531998 316102
rect 531378 315978 531998 316046
rect 531378 315922 531474 315978
rect 531530 315922 531598 315978
rect 531654 315922 531722 315978
rect 531778 315922 531846 315978
rect 531902 315922 531998 315978
rect 531378 298350 531998 315922
rect 558378 597212 558998 598268
rect 558378 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 558998 597212
rect 558378 597088 558998 597156
rect 558378 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 558998 597088
rect 558378 596964 558998 597032
rect 558378 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 558998 596964
rect 558378 596840 558998 596908
rect 558378 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 558998 596840
rect 558378 580350 558998 596784
rect 558378 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 558998 580350
rect 558378 580226 558998 580294
rect 558378 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 558998 580226
rect 558378 580102 558998 580170
rect 558378 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 558998 580102
rect 558378 579978 558998 580046
rect 558378 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 558998 579978
rect 558378 562350 558998 579922
rect 558378 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 558998 562350
rect 558378 562226 558998 562294
rect 558378 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 558998 562226
rect 558378 562102 558998 562170
rect 558378 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 558998 562102
rect 558378 561978 558998 562046
rect 558378 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 558998 561978
rect 558378 544350 558998 561922
rect 558378 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 558998 544350
rect 558378 544226 558998 544294
rect 558378 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 558998 544226
rect 558378 544102 558998 544170
rect 558378 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 558998 544102
rect 558378 543978 558998 544046
rect 558378 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 558998 543978
rect 558378 526350 558998 543922
rect 558378 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 558998 526350
rect 558378 526226 558998 526294
rect 558378 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 558998 526226
rect 558378 526102 558998 526170
rect 558378 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 558998 526102
rect 558378 525978 558998 526046
rect 558378 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 558998 525978
rect 558378 508350 558998 525922
rect 558378 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 558998 508350
rect 558378 508226 558998 508294
rect 558378 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 558998 508226
rect 558378 508102 558998 508170
rect 558378 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 558998 508102
rect 558378 507978 558998 508046
rect 558378 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 558998 507978
rect 558378 490350 558998 507922
rect 558378 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 558998 490350
rect 558378 490226 558998 490294
rect 558378 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 558998 490226
rect 558378 490102 558998 490170
rect 558378 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 558998 490102
rect 558378 489978 558998 490046
rect 558378 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 558998 489978
rect 558378 472350 558998 489922
rect 558378 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 558998 472350
rect 558378 472226 558998 472294
rect 558378 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 558998 472226
rect 558378 472102 558998 472170
rect 558378 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 558998 472102
rect 558378 471978 558998 472046
rect 558378 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 558998 471978
rect 558378 454350 558998 471922
rect 558378 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 558998 454350
rect 558378 454226 558998 454294
rect 558378 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 558998 454226
rect 558378 454102 558998 454170
rect 558378 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 558998 454102
rect 558378 453978 558998 454046
rect 558378 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 558998 453978
rect 558378 436350 558998 453922
rect 558378 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 558998 436350
rect 558378 436226 558998 436294
rect 558378 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 558998 436226
rect 558378 436102 558998 436170
rect 558378 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 558998 436102
rect 558378 435978 558998 436046
rect 558378 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 558998 435978
rect 558378 418350 558998 435922
rect 558378 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 558998 418350
rect 558378 418226 558998 418294
rect 558378 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 558998 418226
rect 558378 418102 558998 418170
rect 558378 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 558998 418102
rect 558378 417978 558998 418046
rect 558378 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 558998 417978
rect 558378 400350 558998 417922
rect 558378 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 558998 400350
rect 558378 400226 558998 400294
rect 558378 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 558998 400226
rect 558378 400102 558998 400170
rect 558378 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 558998 400102
rect 558378 399978 558998 400046
rect 558378 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 558998 399978
rect 558378 382350 558998 399922
rect 558378 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 558998 382350
rect 558378 382226 558998 382294
rect 558378 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 558998 382226
rect 558378 382102 558998 382170
rect 558378 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 558998 382102
rect 558378 381978 558998 382046
rect 558378 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 558998 381978
rect 558378 364350 558998 381922
rect 558378 364294 558474 364350
rect 558530 364294 558598 364350
rect 558654 364294 558722 364350
rect 558778 364294 558846 364350
rect 558902 364294 558998 364350
rect 558378 364226 558998 364294
rect 558378 364170 558474 364226
rect 558530 364170 558598 364226
rect 558654 364170 558722 364226
rect 558778 364170 558846 364226
rect 558902 364170 558998 364226
rect 558378 364102 558998 364170
rect 558378 364046 558474 364102
rect 558530 364046 558598 364102
rect 558654 364046 558722 364102
rect 558778 364046 558846 364102
rect 558902 364046 558998 364102
rect 558378 363978 558998 364046
rect 558378 363922 558474 363978
rect 558530 363922 558598 363978
rect 558654 363922 558722 363978
rect 558778 363922 558846 363978
rect 558902 363922 558998 363978
rect 558378 346350 558998 363922
rect 558378 346294 558474 346350
rect 558530 346294 558598 346350
rect 558654 346294 558722 346350
rect 558778 346294 558846 346350
rect 558902 346294 558998 346350
rect 558378 346226 558998 346294
rect 558378 346170 558474 346226
rect 558530 346170 558598 346226
rect 558654 346170 558722 346226
rect 558778 346170 558846 346226
rect 558902 346170 558998 346226
rect 558378 346102 558998 346170
rect 558378 346046 558474 346102
rect 558530 346046 558598 346102
rect 558654 346046 558722 346102
rect 558778 346046 558846 346102
rect 558902 346046 558998 346102
rect 558378 345978 558998 346046
rect 558378 345922 558474 345978
rect 558530 345922 558598 345978
rect 558654 345922 558722 345978
rect 558778 345922 558846 345978
rect 558902 345922 558998 345978
rect 558378 328350 558998 345922
rect 558378 328294 558474 328350
rect 558530 328294 558598 328350
rect 558654 328294 558722 328350
rect 558778 328294 558846 328350
rect 558902 328294 558998 328350
rect 558378 328226 558998 328294
rect 558378 328170 558474 328226
rect 558530 328170 558598 328226
rect 558654 328170 558722 328226
rect 558778 328170 558846 328226
rect 558902 328170 558998 328226
rect 558378 328102 558998 328170
rect 558378 328046 558474 328102
rect 558530 328046 558598 328102
rect 558654 328046 558722 328102
rect 558778 328046 558846 328102
rect 558902 328046 558998 328102
rect 558378 327978 558998 328046
rect 558378 327922 558474 327978
rect 558530 327922 558598 327978
rect 558654 327922 558722 327978
rect 558778 327922 558846 327978
rect 558902 327922 558998 327978
rect 531378 298294 531474 298350
rect 531530 298294 531598 298350
rect 531654 298294 531722 298350
rect 531778 298294 531846 298350
rect 531902 298294 531998 298350
rect 531378 298226 531998 298294
rect 531378 298170 531474 298226
rect 531530 298170 531598 298226
rect 531654 298170 531722 298226
rect 531778 298170 531846 298226
rect 531902 298170 531998 298226
rect 531378 298102 531998 298170
rect 531378 298046 531474 298102
rect 531530 298046 531598 298102
rect 531654 298046 531722 298102
rect 531778 298046 531846 298102
rect 531902 298046 531998 298102
rect 531378 297978 531998 298046
rect 531378 297922 531474 297978
rect 531530 297922 531598 297978
rect 531654 297922 531722 297978
rect 531778 297922 531846 297978
rect 531902 297922 531998 297978
rect 531378 280350 531998 297922
rect 531378 280294 531474 280350
rect 531530 280294 531598 280350
rect 531654 280294 531722 280350
rect 531778 280294 531846 280350
rect 531902 280294 531998 280350
rect 531378 280226 531998 280294
rect 531378 280170 531474 280226
rect 531530 280170 531598 280226
rect 531654 280170 531722 280226
rect 531778 280170 531846 280226
rect 531902 280170 531998 280226
rect 531378 280102 531998 280170
rect 531378 280046 531474 280102
rect 531530 280046 531598 280102
rect 531654 280046 531722 280102
rect 531778 280046 531846 280102
rect 531902 280046 531998 280102
rect 531378 279978 531998 280046
rect 531378 279922 531474 279978
rect 531530 279922 531598 279978
rect 531654 279922 531722 279978
rect 531778 279922 531846 279978
rect 531902 279922 531998 279978
rect 527658 274294 527754 274350
rect 527810 274294 527878 274350
rect 527934 274294 528002 274350
rect 528058 274294 528126 274350
rect 528182 274294 528278 274350
rect 527658 274226 528278 274294
rect 527658 274170 527754 274226
rect 527810 274170 527878 274226
rect 527934 274170 528002 274226
rect 528058 274170 528126 274226
rect 528182 274170 528278 274226
rect 527658 274102 528278 274170
rect 527658 274046 527754 274102
rect 527810 274046 527878 274102
rect 527934 274046 528002 274102
rect 528058 274046 528126 274102
rect 528182 274046 528278 274102
rect 527658 273978 528278 274046
rect 527658 273922 527754 273978
rect 527810 273922 527878 273978
rect 527934 273922 528002 273978
rect 528058 273922 528126 273978
rect 528182 273922 528278 273978
rect 527658 256350 528278 273922
rect 527658 256294 527754 256350
rect 527810 256294 527878 256350
rect 527934 256294 528002 256350
rect 528058 256294 528126 256350
rect 528182 256294 528278 256350
rect 527658 256226 528278 256294
rect 527658 256170 527754 256226
rect 527810 256170 527878 256226
rect 527934 256170 528002 256226
rect 528058 256170 528126 256226
rect 528182 256170 528278 256226
rect 527658 256102 528278 256170
rect 527658 256046 527754 256102
rect 527810 256046 527878 256102
rect 527934 256046 528002 256102
rect 528058 256046 528126 256102
rect 528182 256046 528278 256102
rect 527658 255978 528278 256046
rect 527658 255922 527754 255978
rect 527810 255922 527878 255978
rect 527934 255922 528002 255978
rect 528058 255922 528126 255978
rect 528182 255922 528278 255978
rect 527658 238350 528278 255922
rect 527658 238294 527754 238350
rect 527810 238294 527878 238350
rect 527934 238294 528002 238350
rect 528058 238294 528126 238350
rect 528182 238294 528278 238350
rect 527658 238226 528278 238294
rect 527658 238170 527754 238226
rect 527810 238170 527878 238226
rect 527934 238170 528002 238226
rect 528058 238170 528126 238226
rect 528182 238170 528278 238226
rect 527658 238102 528278 238170
rect 527658 238046 527754 238102
rect 527810 238046 527878 238102
rect 527934 238046 528002 238102
rect 528058 238046 528126 238102
rect 528182 238046 528278 238102
rect 527658 237978 528278 238046
rect 527658 237922 527754 237978
rect 527810 237922 527878 237978
rect 527934 237922 528002 237978
rect 528058 237922 528126 237978
rect 528182 237922 528278 237978
rect 527658 220350 528278 237922
rect 527658 220294 527754 220350
rect 527810 220294 527878 220350
rect 527934 220294 528002 220350
rect 528058 220294 528126 220350
rect 528182 220294 528278 220350
rect 527658 220226 528278 220294
rect 527658 220170 527754 220226
rect 527810 220170 527878 220226
rect 527934 220170 528002 220226
rect 528058 220170 528126 220226
rect 528182 220170 528278 220226
rect 527658 220102 528278 220170
rect 527658 220046 527754 220102
rect 527810 220046 527878 220102
rect 527934 220046 528002 220102
rect 528058 220046 528126 220102
rect 528182 220046 528278 220102
rect 527658 219978 528278 220046
rect 527658 219922 527754 219978
rect 527810 219922 527878 219978
rect 527934 219922 528002 219978
rect 528058 219922 528126 219978
rect 528182 219922 528278 219978
rect 527658 202350 528278 219922
rect 527658 202294 527754 202350
rect 527810 202294 527878 202350
rect 527934 202294 528002 202350
rect 528058 202294 528126 202350
rect 528182 202294 528278 202350
rect 527658 202226 528278 202294
rect 527658 202170 527754 202226
rect 527810 202170 527878 202226
rect 527934 202170 528002 202226
rect 528058 202170 528126 202226
rect 528182 202170 528278 202226
rect 527658 202102 528278 202170
rect 527658 202046 527754 202102
rect 527810 202046 527878 202102
rect 527934 202046 528002 202102
rect 528058 202046 528126 202102
rect 528182 202046 528278 202102
rect 527658 201978 528278 202046
rect 527658 201922 527754 201978
rect 527810 201922 527878 201978
rect 527934 201922 528002 201978
rect 528058 201922 528126 201978
rect 528182 201922 528278 201978
rect 527658 184350 528278 201922
rect 527658 184294 527754 184350
rect 527810 184294 527878 184350
rect 527934 184294 528002 184350
rect 528058 184294 528126 184350
rect 528182 184294 528278 184350
rect 527658 184226 528278 184294
rect 527658 184170 527754 184226
rect 527810 184170 527878 184226
rect 527934 184170 528002 184226
rect 528058 184170 528126 184226
rect 528182 184170 528278 184226
rect 527658 184102 528278 184170
rect 527658 184046 527754 184102
rect 527810 184046 527878 184102
rect 527934 184046 528002 184102
rect 528058 184046 528126 184102
rect 528182 184046 528278 184102
rect 527658 183978 528278 184046
rect 527658 183922 527754 183978
rect 527810 183922 527878 183978
rect 527934 183922 528002 183978
rect 528058 183922 528126 183978
rect 528182 183922 528278 183978
rect 527658 166350 528278 183922
rect 527658 166294 527754 166350
rect 527810 166294 527878 166350
rect 527934 166294 528002 166350
rect 528058 166294 528126 166350
rect 528182 166294 528278 166350
rect 527658 166226 528278 166294
rect 527658 166170 527754 166226
rect 527810 166170 527878 166226
rect 527934 166170 528002 166226
rect 528058 166170 528126 166226
rect 528182 166170 528278 166226
rect 527658 166102 528278 166170
rect 527658 166046 527754 166102
rect 527810 166046 527878 166102
rect 527934 166046 528002 166102
rect 528058 166046 528126 166102
rect 528182 166046 528278 166102
rect 527658 165978 528278 166046
rect 527658 165922 527754 165978
rect 527810 165922 527878 165978
rect 527934 165922 528002 165978
rect 528058 165922 528126 165978
rect 528182 165922 528278 165978
rect 527658 148350 528278 165922
rect 527658 148294 527754 148350
rect 527810 148294 527878 148350
rect 527934 148294 528002 148350
rect 528058 148294 528126 148350
rect 528182 148294 528278 148350
rect 527658 148226 528278 148294
rect 527658 148170 527754 148226
rect 527810 148170 527878 148226
rect 527934 148170 528002 148226
rect 528058 148170 528126 148226
rect 528182 148170 528278 148226
rect 527658 148102 528278 148170
rect 527658 148046 527754 148102
rect 527810 148046 527878 148102
rect 527934 148046 528002 148102
rect 528058 148046 528126 148102
rect 528182 148046 528278 148102
rect 527658 147978 528278 148046
rect 527658 147922 527754 147978
rect 527810 147922 527878 147978
rect 527934 147922 528002 147978
rect 528058 147922 528126 147978
rect 528182 147922 528278 147978
rect 527658 130350 528278 147922
rect 527658 130294 527754 130350
rect 527810 130294 527878 130350
rect 527934 130294 528002 130350
rect 528058 130294 528126 130350
rect 528182 130294 528278 130350
rect 527658 130226 528278 130294
rect 527658 130170 527754 130226
rect 527810 130170 527878 130226
rect 527934 130170 528002 130226
rect 528058 130170 528126 130226
rect 528182 130170 528278 130226
rect 527658 130102 528278 130170
rect 527658 130046 527754 130102
rect 527810 130046 527878 130102
rect 527934 130046 528002 130102
rect 528058 130046 528126 130102
rect 528182 130046 528278 130102
rect 527658 129978 528278 130046
rect 527658 129922 527754 129978
rect 527810 129922 527878 129978
rect 527934 129922 528002 129978
rect 528058 129922 528126 129978
rect 528182 129922 528278 129978
rect 527658 112350 528278 129922
rect 527658 112294 527754 112350
rect 527810 112294 527878 112350
rect 527934 112294 528002 112350
rect 528058 112294 528126 112350
rect 528182 112294 528278 112350
rect 527658 112226 528278 112294
rect 527658 112170 527754 112226
rect 527810 112170 527878 112226
rect 527934 112170 528002 112226
rect 528058 112170 528126 112226
rect 528182 112170 528278 112226
rect 527658 112102 528278 112170
rect 527658 112046 527754 112102
rect 527810 112046 527878 112102
rect 527934 112046 528002 112102
rect 528058 112046 528126 112102
rect 528182 112046 528278 112102
rect 527658 111978 528278 112046
rect 527658 111922 527754 111978
rect 527810 111922 527878 111978
rect 527934 111922 528002 111978
rect 528058 111922 528126 111978
rect 528182 111922 528278 111978
rect 527658 94350 528278 111922
rect 527658 94294 527754 94350
rect 527810 94294 527878 94350
rect 527934 94294 528002 94350
rect 528058 94294 528126 94350
rect 528182 94294 528278 94350
rect 527658 94226 528278 94294
rect 527658 94170 527754 94226
rect 527810 94170 527878 94226
rect 527934 94170 528002 94226
rect 528058 94170 528126 94226
rect 528182 94170 528278 94226
rect 527658 94102 528278 94170
rect 527658 94046 527754 94102
rect 527810 94046 527878 94102
rect 527934 94046 528002 94102
rect 528058 94046 528126 94102
rect 528182 94046 528278 94102
rect 527658 93978 528278 94046
rect 527658 93922 527754 93978
rect 527810 93922 527878 93978
rect 527934 93922 528002 93978
rect 528058 93922 528126 93978
rect 528182 93922 528278 93978
rect 527658 76350 528278 93922
rect 527658 76294 527754 76350
rect 527810 76294 527878 76350
rect 527934 76294 528002 76350
rect 528058 76294 528126 76350
rect 528182 76294 528278 76350
rect 527658 76226 528278 76294
rect 527658 76170 527754 76226
rect 527810 76170 527878 76226
rect 527934 76170 528002 76226
rect 528058 76170 528126 76226
rect 528182 76170 528278 76226
rect 527658 76102 528278 76170
rect 527658 76046 527754 76102
rect 527810 76046 527878 76102
rect 527934 76046 528002 76102
rect 528058 76046 528126 76102
rect 528182 76046 528278 76102
rect 527658 75978 528278 76046
rect 527658 75922 527754 75978
rect 527810 75922 527878 75978
rect 527934 75922 528002 75978
rect 528058 75922 528126 75978
rect 528182 75922 528278 75978
rect 500658 64294 500754 64350
rect 500810 64294 500878 64350
rect 500934 64294 501002 64350
rect 501058 64294 501126 64350
rect 501182 64294 501278 64350
rect 500658 64226 501278 64294
rect 500658 64170 500754 64226
rect 500810 64170 500878 64226
rect 500934 64170 501002 64226
rect 501058 64170 501126 64226
rect 501182 64170 501278 64226
rect 500658 64102 501278 64170
rect 500658 64046 500754 64102
rect 500810 64046 500878 64102
rect 500934 64046 501002 64102
rect 501058 64046 501126 64102
rect 501182 64046 501278 64102
rect 500658 63978 501278 64046
rect 500658 63922 500754 63978
rect 500810 63922 500878 63978
rect 500934 63922 501002 63978
rect 501058 63922 501126 63978
rect 501182 63922 501278 63978
rect 500658 46350 501278 63922
rect 500658 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 501278 46350
rect 500658 46226 501278 46294
rect 500658 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 501278 46226
rect 500658 46102 501278 46170
rect 500658 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 501278 46102
rect 500658 45978 501278 46046
rect 500658 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 501278 45978
rect 500658 28350 501278 45922
rect 500658 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 501278 28350
rect 500658 28226 501278 28294
rect 500658 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 501278 28226
rect 500658 28102 501278 28170
rect 500658 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 501278 28102
rect 500658 27978 501278 28046
rect 500658 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 501278 27978
rect 500658 10350 501278 27922
rect 500658 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 501278 10350
rect 500658 10226 501278 10294
rect 500658 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 501278 10226
rect 500658 10102 501278 10170
rect 500658 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 501278 10102
rect 500658 9978 501278 10046
rect 500658 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 501278 9978
rect 498988 5158 499044 5168
rect 498988 5058 499044 5068
rect 496938 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 497558 4350
rect 496938 4226 497558 4294
rect 496938 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 497558 4226
rect 496938 4102 497558 4170
rect 496938 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 497558 4102
rect 496938 3978 497558 4046
rect 496938 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 497558 3978
rect 475468 3266 475524 3276
rect 487676 1204 487732 1214
rect 487676 308 487732 1148
rect 487676 242 487732 252
rect 469938 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 470558 -1120
rect 469938 -1244 470558 -1176
rect 469938 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 470558 -1244
rect 469938 -1368 470558 -1300
rect 469938 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 470558 -1368
rect 469938 -1492 470558 -1424
rect 469938 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 470558 -1492
rect 469938 -1644 470558 -1548
rect 496938 -160 497558 3922
rect 498988 3444 499044 3454
rect 498988 3358 499044 3388
rect 498988 3292 499044 3302
rect 499436 3332 499492 3342
rect 499436 3178 499492 3276
rect 499436 3112 499492 3122
rect 496938 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 497558 -160
rect 496938 -284 497558 -216
rect 496938 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 497558 -284
rect 496938 -408 497558 -340
rect 496938 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 497558 -408
rect 496938 -532 497558 -464
rect 496938 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 497558 -532
rect 496938 -1644 497558 -588
rect 500658 -1120 501278 9922
rect 527658 58350 528278 75922
rect 530012 278068 530068 278078
rect 530012 68628 530068 278012
rect 530012 68562 530068 68572
rect 531378 262350 531998 279922
rect 531378 262294 531474 262350
rect 531530 262294 531598 262350
rect 531654 262294 531722 262350
rect 531778 262294 531846 262350
rect 531902 262294 531998 262350
rect 531378 262226 531998 262294
rect 531378 262170 531474 262226
rect 531530 262170 531598 262226
rect 531654 262170 531722 262226
rect 531778 262170 531846 262226
rect 531902 262170 531998 262226
rect 531378 262102 531998 262170
rect 531378 262046 531474 262102
rect 531530 262046 531598 262102
rect 531654 262046 531722 262102
rect 531778 262046 531846 262102
rect 531902 262046 531998 262102
rect 531378 261978 531998 262046
rect 531378 261922 531474 261978
rect 531530 261922 531598 261978
rect 531654 261922 531722 261978
rect 531778 261922 531846 261978
rect 531902 261922 531998 261978
rect 531378 244350 531998 261922
rect 531378 244294 531474 244350
rect 531530 244294 531598 244350
rect 531654 244294 531722 244350
rect 531778 244294 531846 244350
rect 531902 244294 531998 244350
rect 531378 244226 531998 244294
rect 531378 244170 531474 244226
rect 531530 244170 531598 244226
rect 531654 244170 531722 244226
rect 531778 244170 531846 244226
rect 531902 244170 531998 244226
rect 531378 244102 531998 244170
rect 531378 244046 531474 244102
rect 531530 244046 531598 244102
rect 531654 244046 531722 244102
rect 531778 244046 531846 244102
rect 531902 244046 531998 244102
rect 531378 243978 531998 244046
rect 531378 243922 531474 243978
rect 531530 243922 531598 243978
rect 531654 243922 531722 243978
rect 531778 243922 531846 243978
rect 531902 243922 531998 243978
rect 531378 226350 531998 243922
rect 531378 226294 531474 226350
rect 531530 226294 531598 226350
rect 531654 226294 531722 226350
rect 531778 226294 531846 226350
rect 531902 226294 531998 226350
rect 531378 226226 531998 226294
rect 531378 226170 531474 226226
rect 531530 226170 531598 226226
rect 531654 226170 531722 226226
rect 531778 226170 531846 226226
rect 531902 226170 531998 226226
rect 531378 226102 531998 226170
rect 531378 226046 531474 226102
rect 531530 226046 531598 226102
rect 531654 226046 531722 226102
rect 531778 226046 531846 226102
rect 531902 226046 531998 226102
rect 531378 225978 531998 226046
rect 531378 225922 531474 225978
rect 531530 225922 531598 225978
rect 531654 225922 531722 225978
rect 531778 225922 531846 225978
rect 531902 225922 531998 225978
rect 531378 208350 531998 225922
rect 531378 208294 531474 208350
rect 531530 208294 531598 208350
rect 531654 208294 531722 208350
rect 531778 208294 531846 208350
rect 531902 208294 531998 208350
rect 531378 208226 531998 208294
rect 531378 208170 531474 208226
rect 531530 208170 531598 208226
rect 531654 208170 531722 208226
rect 531778 208170 531846 208226
rect 531902 208170 531998 208226
rect 531378 208102 531998 208170
rect 531378 208046 531474 208102
rect 531530 208046 531598 208102
rect 531654 208046 531722 208102
rect 531778 208046 531846 208102
rect 531902 208046 531998 208102
rect 531378 207978 531998 208046
rect 531378 207922 531474 207978
rect 531530 207922 531598 207978
rect 531654 207922 531722 207978
rect 531778 207922 531846 207978
rect 531902 207922 531998 207978
rect 531378 190350 531998 207922
rect 531378 190294 531474 190350
rect 531530 190294 531598 190350
rect 531654 190294 531722 190350
rect 531778 190294 531846 190350
rect 531902 190294 531998 190350
rect 531378 190226 531998 190294
rect 531378 190170 531474 190226
rect 531530 190170 531598 190226
rect 531654 190170 531722 190226
rect 531778 190170 531846 190226
rect 531902 190170 531998 190226
rect 531378 190102 531998 190170
rect 531378 190046 531474 190102
rect 531530 190046 531598 190102
rect 531654 190046 531722 190102
rect 531778 190046 531846 190102
rect 531902 190046 531998 190102
rect 531378 189978 531998 190046
rect 531378 189922 531474 189978
rect 531530 189922 531598 189978
rect 531654 189922 531722 189978
rect 531778 189922 531846 189978
rect 531902 189922 531998 189978
rect 531378 172350 531998 189922
rect 531378 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 531998 172350
rect 531378 172226 531998 172294
rect 531378 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 531998 172226
rect 531378 172102 531998 172170
rect 531378 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 531998 172102
rect 531378 171978 531998 172046
rect 531378 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 531998 171978
rect 531378 154350 531998 171922
rect 531378 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 531998 154350
rect 531378 154226 531998 154294
rect 531378 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 531998 154226
rect 531378 154102 531998 154170
rect 531378 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 531998 154102
rect 531378 153978 531998 154046
rect 531378 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 531998 153978
rect 531378 136350 531998 153922
rect 531378 136294 531474 136350
rect 531530 136294 531598 136350
rect 531654 136294 531722 136350
rect 531778 136294 531846 136350
rect 531902 136294 531998 136350
rect 531378 136226 531998 136294
rect 531378 136170 531474 136226
rect 531530 136170 531598 136226
rect 531654 136170 531722 136226
rect 531778 136170 531846 136226
rect 531902 136170 531998 136226
rect 531378 136102 531998 136170
rect 531378 136046 531474 136102
rect 531530 136046 531598 136102
rect 531654 136046 531722 136102
rect 531778 136046 531846 136102
rect 531902 136046 531998 136102
rect 531378 135978 531998 136046
rect 531378 135922 531474 135978
rect 531530 135922 531598 135978
rect 531654 135922 531722 135978
rect 531778 135922 531846 135978
rect 531902 135922 531998 135978
rect 531378 118350 531998 135922
rect 531378 118294 531474 118350
rect 531530 118294 531598 118350
rect 531654 118294 531722 118350
rect 531778 118294 531846 118350
rect 531902 118294 531998 118350
rect 531378 118226 531998 118294
rect 531378 118170 531474 118226
rect 531530 118170 531598 118226
rect 531654 118170 531722 118226
rect 531778 118170 531846 118226
rect 531902 118170 531998 118226
rect 531378 118102 531998 118170
rect 531378 118046 531474 118102
rect 531530 118046 531598 118102
rect 531654 118046 531722 118102
rect 531778 118046 531846 118102
rect 531902 118046 531998 118102
rect 531378 117978 531998 118046
rect 531378 117922 531474 117978
rect 531530 117922 531598 117978
rect 531654 117922 531722 117978
rect 531778 117922 531846 117978
rect 531902 117922 531998 117978
rect 531378 100350 531998 117922
rect 531378 100294 531474 100350
rect 531530 100294 531598 100350
rect 531654 100294 531722 100350
rect 531778 100294 531846 100350
rect 531902 100294 531998 100350
rect 531378 100226 531998 100294
rect 531378 100170 531474 100226
rect 531530 100170 531598 100226
rect 531654 100170 531722 100226
rect 531778 100170 531846 100226
rect 531902 100170 531998 100226
rect 531378 100102 531998 100170
rect 531378 100046 531474 100102
rect 531530 100046 531598 100102
rect 531654 100046 531722 100102
rect 531778 100046 531846 100102
rect 531902 100046 531998 100102
rect 531378 99978 531998 100046
rect 531378 99922 531474 99978
rect 531530 99922 531598 99978
rect 531654 99922 531722 99978
rect 531778 99922 531846 99978
rect 531902 99922 531998 99978
rect 531378 82350 531998 99922
rect 531378 82294 531474 82350
rect 531530 82294 531598 82350
rect 531654 82294 531722 82350
rect 531778 82294 531846 82350
rect 531902 82294 531998 82350
rect 531378 82226 531998 82294
rect 531378 82170 531474 82226
rect 531530 82170 531598 82226
rect 531654 82170 531722 82226
rect 531778 82170 531846 82226
rect 531902 82170 531998 82226
rect 531378 82102 531998 82170
rect 531378 82046 531474 82102
rect 531530 82046 531598 82102
rect 531654 82046 531722 82102
rect 531778 82046 531846 82102
rect 531902 82046 531998 82102
rect 531378 81978 531998 82046
rect 531378 81922 531474 81978
rect 531530 81922 531598 81978
rect 531654 81922 531722 81978
rect 531778 81922 531846 81978
rect 531902 81922 531998 81978
rect 527658 58294 527754 58350
rect 527810 58294 527878 58350
rect 527934 58294 528002 58350
rect 528058 58294 528126 58350
rect 528182 58294 528278 58350
rect 527658 58226 528278 58294
rect 527658 58170 527754 58226
rect 527810 58170 527878 58226
rect 527934 58170 528002 58226
rect 528058 58170 528126 58226
rect 528182 58170 528278 58226
rect 527658 58102 528278 58170
rect 527658 58046 527754 58102
rect 527810 58046 527878 58102
rect 527934 58046 528002 58102
rect 528058 58046 528126 58102
rect 528182 58046 528278 58102
rect 527658 57978 528278 58046
rect 527658 57922 527754 57978
rect 527810 57922 527878 57978
rect 527934 57922 528002 57978
rect 528058 57922 528126 57978
rect 528182 57922 528278 57978
rect 527658 40350 528278 57922
rect 527658 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 528278 40350
rect 527658 40226 528278 40294
rect 527658 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 528278 40226
rect 527658 40102 528278 40170
rect 527658 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 528278 40102
rect 527658 39978 528278 40046
rect 527658 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 528278 39978
rect 527658 22350 528278 39922
rect 527658 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 528278 22350
rect 527658 22226 528278 22294
rect 527658 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 528278 22226
rect 527658 22102 528278 22170
rect 527658 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 528278 22102
rect 527658 21978 528278 22046
rect 527658 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 528278 21978
rect 527658 4350 528278 21922
rect 531378 64350 531998 81922
rect 531378 64294 531474 64350
rect 531530 64294 531598 64350
rect 531654 64294 531722 64350
rect 531778 64294 531846 64350
rect 531902 64294 531998 64350
rect 531378 64226 531998 64294
rect 531378 64170 531474 64226
rect 531530 64170 531598 64226
rect 531654 64170 531722 64226
rect 531778 64170 531846 64226
rect 531902 64170 531998 64226
rect 531378 64102 531998 64170
rect 531378 64046 531474 64102
rect 531530 64046 531598 64102
rect 531654 64046 531722 64102
rect 531778 64046 531846 64102
rect 531902 64046 531998 64102
rect 531378 63978 531998 64046
rect 531378 63922 531474 63978
rect 531530 63922 531598 63978
rect 531654 63922 531722 63978
rect 531778 63922 531846 63978
rect 531902 63922 531998 63978
rect 531378 46350 531998 63922
rect 531378 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 531998 46350
rect 531378 46226 531998 46294
rect 531378 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 531998 46226
rect 531378 46102 531998 46170
rect 531378 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 531998 46102
rect 531378 45978 531998 46046
rect 531378 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 531998 45978
rect 531378 28350 531998 45922
rect 543452 311108 543508 311118
rect 543452 32900 543508 311052
rect 558378 310350 558998 327922
rect 558378 310294 558474 310350
rect 558530 310294 558598 310350
rect 558654 310294 558722 310350
rect 558778 310294 558846 310350
rect 558902 310294 558998 310350
rect 558378 310226 558998 310294
rect 558378 310170 558474 310226
rect 558530 310170 558598 310226
rect 558654 310170 558722 310226
rect 558778 310170 558846 310226
rect 558902 310170 558998 310226
rect 558378 310102 558998 310170
rect 558378 310046 558474 310102
rect 558530 310046 558598 310102
rect 558654 310046 558722 310102
rect 558778 310046 558846 310102
rect 558902 310046 558998 310102
rect 558378 309978 558998 310046
rect 558378 309922 558474 309978
rect 558530 309922 558598 309978
rect 558654 309922 558722 309978
rect 558778 309922 558846 309978
rect 558902 309922 558998 309978
rect 558378 292350 558998 309922
rect 558378 292294 558474 292350
rect 558530 292294 558598 292350
rect 558654 292294 558722 292350
rect 558778 292294 558846 292350
rect 558902 292294 558998 292350
rect 558378 292226 558998 292294
rect 558378 292170 558474 292226
rect 558530 292170 558598 292226
rect 558654 292170 558722 292226
rect 558778 292170 558846 292226
rect 558902 292170 558998 292226
rect 558378 292102 558998 292170
rect 558378 292046 558474 292102
rect 558530 292046 558598 292102
rect 558654 292046 558722 292102
rect 558778 292046 558846 292102
rect 558902 292046 558998 292102
rect 558378 291978 558998 292046
rect 558378 291922 558474 291978
rect 558530 291922 558598 291978
rect 558654 291922 558722 291978
rect 558778 291922 558846 291978
rect 558902 291922 558998 291978
rect 558378 274350 558998 291922
rect 558378 274294 558474 274350
rect 558530 274294 558598 274350
rect 558654 274294 558722 274350
rect 558778 274294 558846 274350
rect 558902 274294 558998 274350
rect 558378 274226 558998 274294
rect 558378 274170 558474 274226
rect 558530 274170 558598 274226
rect 558654 274170 558722 274226
rect 558778 274170 558846 274226
rect 558902 274170 558998 274226
rect 558378 274102 558998 274170
rect 558378 274046 558474 274102
rect 558530 274046 558598 274102
rect 558654 274046 558722 274102
rect 558778 274046 558846 274102
rect 558902 274046 558998 274102
rect 558378 273978 558998 274046
rect 558378 273922 558474 273978
rect 558530 273922 558598 273978
rect 558654 273922 558722 273978
rect 558778 273922 558846 273978
rect 558902 273922 558998 273978
rect 550172 271460 550228 271470
rect 543452 32834 543508 32844
rect 543564 231924 543620 231934
rect 531378 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 531998 28350
rect 531378 28226 531998 28294
rect 531378 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 531998 28226
rect 531378 28102 531998 28170
rect 531378 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 531998 28102
rect 531378 27978 531998 28046
rect 531378 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 531998 27978
rect 531378 10350 531998 27922
rect 538400 28350 538720 28384
rect 538400 28294 538470 28350
rect 538526 28294 538594 28350
rect 538650 28294 538720 28350
rect 538400 28226 538720 28294
rect 538400 28170 538470 28226
rect 538526 28170 538594 28226
rect 538650 28170 538720 28226
rect 538400 28102 538720 28170
rect 538400 28046 538470 28102
rect 538526 28046 538594 28102
rect 538650 28046 538720 28102
rect 538400 27978 538720 28046
rect 538400 27922 538470 27978
rect 538526 27922 538594 27978
rect 538650 27922 538720 27978
rect 538400 27888 538720 27922
rect 543564 26180 543620 231868
rect 543564 26114 543620 26124
rect 543676 218596 543732 218606
rect 543676 25060 543732 218540
rect 548492 192164 548548 192174
rect 543676 24994 543732 25004
rect 543788 152516 543844 152526
rect 543788 19460 543844 152460
rect 543788 19394 543844 19404
rect 543900 139300 543956 139310
rect 543900 18340 543956 139244
rect 546812 112868 546868 112878
rect 545132 73220 545188 73230
rect 543900 18274 543956 18284
rect 544012 60004 544068 60014
rect 544012 11620 544068 59948
rect 544236 29428 544292 29438
rect 544236 27300 544292 29372
rect 544236 27234 544292 27244
rect 544348 24388 544404 24398
rect 544348 20580 544404 24332
rect 544348 20514 544404 20524
rect 545132 12740 545188 73164
rect 546812 16100 546868 112812
rect 548492 22820 548548 192108
rect 550172 29540 550228 271404
rect 555212 258244 555268 258254
rect 553532 178948 553588 178958
rect 551852 98308 551908 98318
rect 550172 29474 550228 29484
rect 550284 33684 550340 33694
rect 548492 22754 548548 22764
rect 546812 16034 546868 16044
rect 548492 19348 548548 19358
rect 545132 12674 545188 12684
rect 544012 11554 544068 11564
rect 544348 12628 544404 12638
rect 544348 10500 544404 12572
rect 544348 10434 544404 10444
rect 531378 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 531998 10350
rect 531378 10226 531998 10294
rect 531378 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 531998 10226
rect 531378 10102 531998 10170
rect 531378 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 531998 10102
rect 531378 9978 531998 10046
rect 531378 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 531998 9978
rect 527658 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 528278 4350
rect 527658 4226 528278 4294
rect 527658 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 528278 4226
rect 527658 4102 528278 4170
rect 527658 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 528278 4102
rect 527658 3978 528278 4046
rect 527658 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 528278 3978
rect 501676 3358 501732 3370
rect 501676 3266 501732 3276
rect 504140 2548 504196 2558
rect 504140 118 504196 2492
rect 510748 2548 510804 2558
rect 510748 298 510804 2492
rect 512092 756 512148 766
rect 512092 478 512148 700
rect 512092 412 512148 422
rect 510748 232 510804 242
rect 504140 52 504196 62
rect 500658 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 501278 -1120
rect 500658 -1244 501278 -1176
rect 500658 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 501278 -1244
rect 500658 -1368 501278 -1300
rect 500658 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 501278 -1368
rect 500658 -1492 501278 -1424
rect 500658 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 501278 -1492
rect 500658 -1644 501278 -1548
rect 527658 -160 528278 3922
rect 529228 5338 529284 5348
rect 529228 3444 529284 5282
rect 529228 3378 529284 3388
rect 527658 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 528278 -160
rect 527658 -284 528278 -216
rect 527658 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 528278 -284
rect 527658 -408 528278 -340
rect 527658 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 528278 -408
rect 527658 -532 528278 -464
rect 527658 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 528278 -532
rect 527658 -1644 528278 -588
rect 531378 -1120 531998 9922
rect 538400 10350 538720 10384
rect 538400 10294 538470 10350
rect 538526 10294 538594 10350
rect 538650 10294 538720 10350
rect 538400 10226 538720 10294
rect 538400 10170 538470 10226
rect 538526 10170 538594 10226
rect 538650 10170 538720 10226
rect 538400 10102 538720 10170
rect 538400 10046 538470 10102
rect 538526 10046 538594 10102
rect 538650 10046 538720 10102
rect 538400 9978 538720 10046
rect 538400 9922 538470 9978
rect 538526 9922 538594 9978
rect 538650 9922 538720 9978
rect 538400 9888 538720 9922
rect 548492 8260 548548 19292
rect 550284 9380 550340 33628
rect 551852 14980 551908 98252
rect 553532 21700 553588 178892
rect 555212 28420 555268 258188
rect 558378 256350 558998 273922
rect 558378 256294 558474 256350
rect 558530 256294 558598 256350
rect 558654 256294 558722 256350
rect 558778 256294 558846 256350
rect 558902 256294 558998 256350
rect 558378 256226 558998 256294
rect 558378 256170 558474 256226
rect 558530 256170 558598 256226
rect 558654 256170 558722 256226
rect 558778 256170 558846 256226
rect 558902 256170 558998 256226
rect 558378 256102 558998 256170
rect 558378 256046 558474 256102
rect 558530 256046 558598 256102
rect 558654 256046 558722 256102
rect 558778 256046 558846 256102
rect 558902 256046 558998 256102
rect 558378 255978 558998 256046
rect 558378 255922 558474 255978
rect 558530 255922 558598 255978
rect 558654 255922 558722 255978
rect 558778 255922 558846 255978
rect 558902 255922 558998 255978
rect 558378 238350 558998 255922
rect 558378 238294 558474 238350
rect 558530 238294 558598 238350
rect 558654 238294 558722 238350
rect 558778 238294 558846 238350
rect 558902 238294 558998 238350
rect 558378 238226 558998 238294
rect 558378 238170 558474 238226
rect 558530 238170 558598 238226
rect 558654 238170 558722 238226
rect 558778 238170 558846 238226
rect 558902 238170 558998 238226
rect 558378 238102 558998 238170
rect 558378 238046 558474 238102
rect 558530 238046 558598 238102
rect 558654 238046 558722 238102
rect 558778 238046 558846 238102
rect 558902 238046 558998 238102
rect 558378 237978 558998 238046
rect 558378 237922 558474 237978
rect 558530 237922 558598 237978
rect 558654 237922 558722 237978
rect 558778 237922 558846 237978
rect 558902 237922 558998 237978
rect 558378 220350 558998 237922
rect 558378 220294 558474 220350
rect 558530 220294 558598 220350
rect 558654 220294 558722 220350
rect 558778 220294 558846 220350
rect 558902 220294 558998 220350
rect 558378 220226 558998 220294
rect 558378 220170 558474 220226
rect 558530 220170 558598 220226
rect 558654 220170 558722 220226
rect 558778 220170 558846 220226
rect 558902 220170 558998 220226
rect 558378 220102 558998 220170
rect 558378 220046 558474 220102
rect 558530 220046 558598 220102
rect 558654 220046 558722 220102
rect 558778 220046 558846 220102
rect 558902 220046 558998 220102
rect 558378 219978 558998 220046
rect 558378 219922 558474 219978
rect 558530 219922 558598 219978
rect 558654 219922 558722 219978
rect 558778 219922 558846 219978
rect 558902 219922 558998 219978
rect 558378 202350 558998 219922
rect 562098 598172 562718 598268
rect 562098 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 562718 598172
rect 562098 598048 562718 598116
rect 562098 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 562718 598048
rect 562098 597924 562718 597992
rect 562098 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 562718 597924
rect 562098 597800 562718 597868
rect 562098 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 562718 597800
rect 562098 586350 562718 597744
rect 589098 597212 589718 598268
rect 589098 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 589718 597212
rect 589098 597088 589718 597156
rect 589098 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 589718 597088
rect 589098 596964 589718 597032
rect 589098 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 589718 596964
rect 589098 596840 589718 596908
rect 589098 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 589718 596840
rect 562098 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 562718 586350
rect 562098 586226 562718 586294
rect 562098 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 562718 586226
rect 562098 586102 562718 586170
rect 562098 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 562718 586102
rect 562098 585978 562718 586046
rect 562098 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 562718 585978
rect 562098 568350 562718 585922
rect 562098 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 562718 568350
rect 562098 568226 562718 568294
rect 562098 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 562718 568226
rect 562098 568102 562718 568170
rect 562098 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 562718 568102
rect 562098 567978 562718 568046
rect 562098 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 562718 567978
rect 562098 550350 562718 567922
rect 562098 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 562718 550350
rect 562098 550226 562718 550294
rect 562098 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 562718 550226
rect 562098 550102 562718 550170
rect 562098 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 562718 550102
rect 562098 549978 562718 550046
rect 562098 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 562718 549978
rect 562098 532350 562718 549922
rect 562098 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 562718 532350
rect 562098 532226 562718 532294
rect 562098 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 562718 532226
rect 562098 532102 562718 532170
rect 562098 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 562718 532102
rect 562098 531978 562718 532046
rect 562098 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 562718 531978
rect 562098 514350 562718 531922
rect 562098 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 562718 514350
rect 562098 514226 562718 514294
rect 562098 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 562718 514226
rect 562098 514102 562718 514170
rect 562098 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 562718 514102
rect 562098 513978 562718 514046
rect 562098 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 562718 513978
rect 562098 496350 562718 513922
rect 562098 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 562718 496350
rect 562098 496226 562718 496294
rect 562098 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 562718 496226
rect 562098 496102 562718 496170
rect 562098 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 562718 496102
rect 562098 495978 562718 496046
rect 562098 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 562718 495978
rect 562098 478350 562718 495922
rect 562098 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 562718 478350
rect 562098 478226 562718 478294
rect 562098 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 562718 478226
rect 562098 478102 562718 478170
rect 562098 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 562718 478102
rect 562098 477978 562718 478046
rect 562098 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 562718 477978
rect 562098 460350 562718 477922
rect 562098 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 562718 460350
rect 562098 460226 562718 460294
rect 562098 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 562718 460226
rect 562098 460102 562718 460170
rect 562098 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 562718 460102
rect 562098 459978 562718 460046
rect 562098 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 562718 459978
rect 562098 442350 562718 459922
rect 562098 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 562718 442350
rect 562098 442226 562718 442294
rect 562098 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 562718 442226
rect 562098 442102 562718 442170
rect 562098 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 562718 442102
rect 562098 441978 562718 442046
rect 562098 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 562718 441978
rect 562098 424350 562718 441922
rect 562098 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 562718 424350
rect 562098 424226 562718 424294
rect 562098 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 562718 424226
rect 562098 424102 562718 424170
rect 562098 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 562718 424102
rect 562098 423978 562718 424046
rect 562098 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 562718 423978
rect 562098 406350 562718 423922
rect 562098 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 562718 406350
rect 562098 406226 562718 406294
rect 562098 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 562718 406226
rect 562098 406102 562718 406170
rect 562098 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 562718 406102
rect 562098 405978 562718 406046
rect 562098 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 562718 405978
rect 562098 388350 562718 405922
rect 562098 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 562718 388350
rect 562098 388226 562718 388294
rect 562098 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 562718 388226
rect 562098 388102 562718 388170
rect 562098 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 562718 388102
rect 562098 387978 562718 388046
rect 562098 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 562718 387978
rect 562098 370350 562718 387922
rect 562098 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 562718 370350
rect 562098 370226 562718 370294
rect 562098 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 562718 370226
rect 562098 370102 562718 370170
rect 562098 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 562718 370102
rect 562098 369978 562718 370046
rect 562098 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 562718 369978
rect 562098 352350 562718 369922
rect 584668 590212 584724 590222
rect 584668 368758 584724 590156
rect 584668 368692 584724 368702
rect 589098 580350 589718 596784
rect 592818 598172 593438 598268
rect 592818 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 593438 598172
rect 592818 598048 593438 598116
rect 592818 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 593438 598048
rect 592818 597924 593438 597992
rect 592818 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 593438 597924
rect 592818 597800 593438 597868
rect 592818 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 593438 597800
rect 589098 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 589718 580350
rect 589098 580226 589718 580294
rect 589098 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 589718 580226
rect 589098 580102 589718 580170
rect 589098 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 589718 580102
rect 589098 579978 589718 580046
rect 589098 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 589718 579978
rect 589098 562350 589718 579922
rect 589098 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 589718 562350
rect 589098 562226 589718 562294
rect 589098 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 589718 562226
rect 589098 562102 589718 562170
rect 589098 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 589718 562102
rect 589098 561978 589718 562046
rect 589098 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 589718 561978
rect 589098 544350 589718 561922
rect 589098 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 589718 544350
rect 589098 544226 589718 544294
rect 589098 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 589718 544226
rect 589098 544102 589718 544170
rect 589098 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 589718 544102
rect 589098 543978 589718 544046
rect 589098 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 589718 543978
rect 589098 526350 589718 543922
rect 589098 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 589718 526350
rect 589098 526226 589718 526294
rect 589098 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 589718 526226
rect 589098 526102 589718 526170
rect 589098 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 589718 526102
rect 589098 525978 589718 526046
rect 589098 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 589718 525978
rect 589098 508350 589718 525922
rect 589098 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 589718 508350
rect 589098 508226 589718 508294
rect 589098 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 589718 508226
rect 589098 508102 589718 508170
rect 589098 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 589718 508102
rect 589098 507978 589718 508046
rect 589098 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 589718 507978
rect 589098 490350 589718 507922
rect 589098 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 589718 490350
rect 589098 490226 589718 490294
rect 589098 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 589718 490226
rect 589098 490102 589718 490170
rect 589098 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 589718 490102
rect 589098 489978 589718 490046
rect 589098 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 589718 489978
rect 589098 472350 589718 489922
rect 590492 588644 590548 588654
rect 590492 483028 590548 588588
rect 592818 586350 593438 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 592818 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 593438 586350
rect 592818 586226 593438 586294
rect 592818 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 593438 586226
rect 592818 586102 593438 586170
rect 592818 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 593438 586102
rect 592818 585978 593438 586046
rect 592818 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 593438 585978
rect 592818 568350 593438 585922
rect 592818 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 593438 568350
rect 592818 568226 593438 568294
rect 592818 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 593438 568226
rect 592818 568102 593438 568170
rect 592818 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 593438 568102
rect 592818 567978 593438 568046
rect 592818 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 593438 567978
rect 590604 562212 590660 562222
rect 590604 523348 590660 562156
rect 590604 523282 590660 523292
rect 592818 550350 593438 567922
rect 592818 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 593438 550350
rect 592818 550226 593438 550294
rect 592818 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 593438 550226
rect 592818 550102 593438 550170
rect 592818 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 593438 550102
rect 592818 549978 593438 550046
rect 592818 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 593438 549978
rect 592818 532350 593438 549922
rect 592818 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 593438 532350
rect 592818 532226 593438 532294
rect 592818 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 593438 532226
rect 592818 532102 593438 532170
rect 592818 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 593438 532102
rect 592818 531978 593438 532046
rect 592818 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 593438 531978
rect 590492 482962 590548 482972
rect 592818 514350 593438 531922
rect 592818 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 593438 514350
rect 592818 514226 593438 514294
rect 592818 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 593438 514226
rect 592818 514102 593438 514170
rect 592818 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 593438 514102
rect 592818 513978 593438 514046
rect 592818 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 593438 513978
rect 592818 496350 593438 513922
rect 592818 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 593438 496350
rect 592818 496226 593438 496294
rect 592818 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 593438 496226
rect 592818 496102 593438 496170
rect 592818 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 593438 496102
rect 592818 495978 593438 496046
rect 592818 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 593438 495978
rect 589098 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 589718 472350
rect 589098 472226 589718 472294
rect 589098 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 589718 472226
rect 589098 472102 589718 472170
rect 589098 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 589718 472102
rect 589098 471978 589718 472046
rect 589098 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 589718 471978
rect 589098 454350 589718 471922
rect 589098 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 589718 454350
rect 589098 454226 589718 454294
rect 589098 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 589718 454226
rect 589098 454102 589718 454170
rect 589098 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 589718 454102
rect 589098 453978 589718 454046
rect 589098 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 589718 453978
rect 589098 436350 589718 453922
rect 589098 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 589718 436350
rect 589098 436226 589718 436294
rect 589098 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 589718 436226
rect 589098 436102 589718 436170
rect 589098 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 589718 436102
rect 589098 435978 589718 436046
rect 589098 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 589718 435978
rect 589098 418350 589718 435922
rect 589098 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 589718 418350
rect 589098 418226 589718 418294
rect 589098 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 589718 418226
rect 589098 418102 589718 418170
rect 589098 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 589718 418102
rect 589098 417978 589718 418046
rect 589098 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 589718 417978
rect 589098 400350 589718 417922
rect 589098 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 589718 400350
rect 589098 400226 589718 400294
rect 589098 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 589718 400226
rect 589098 400102 589718 400170
rect 589098 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 589718 400102
rect 589098 399978 589718 400046
rect 589098 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 589718 399978
rect 589098 382350 589718 399922
rect 589098 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 589718 382350
rect 589098 382226 589718 382294
rect 589098 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 589718 382226
rect 589098 382102 589718 382170
rect 589098 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 589718 382102
rect 589098 381978 589718 382046
rect 589098 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 589718 381978
rect 562098 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 562718 352350
rect 562098 352226 562718 352294
rect 562098 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 562718 352226
rect 562098 352102 562718 352170
rect 562098 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 562718 352102
rect 562098 351978 562718 352046
rect 562098 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 562718 351978
rect 562098 334350 562718 351922
rect 562098 334294 562194 334350
rect 562250 334294 562318 334350
rect 562374 334294 562442 334350
rect 562498 334294 562566 334350
rect 562622 334294 562718 334350
rect 562098 334226 562718 334294
rect 562098 334170 562194 334226
rect 562250 334170 562318 334226
rect 562374 334170 562442 334226
rect 562498 334170 562566 334226
rect 562622 334170 562718 334226
rect 562098 334102 562718 334170
rect 562098 334046 562194 334102
rect 562250 334046 562318 334102
rect 562374 334046 562442 334102
rect 562498 334046 562566 334102
rect 562622 334046 562718 334102
rect 562098 333978 562718 334046
rect 562098 333922 562194 333978
rect 562250 333922 562318 333978
rect 562374 333922 562442 333978
rect 562498 333922 562566 333978
rect 562622 333922 562718 333978
rect 562098 316350 562718 333922
rect 562098 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 562718 316350
rect 562098 316226 562718 316294
rect 562098 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 562718 316226
rect 562098 316102 562718 316170
rect 562098 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 562718 316102
rect 562098 315978 562718 316046
rect 562098 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 562718 315978
rect 562098 298350 562718 315922
rect 562098 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 562718 298350
rect 562098 298226 562718 298294
rect 562098 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 562718 298226
rect 562098 298102 562718 298170
rect 562098 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 562718 298102
rect 562098 297978 562718 298046
rect 562098 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 562718 297978
rect 562098 280350 562718 297922
rect 589098 364350 589718 381922
rect 589098 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 589718 364350
rect 589098 364226 589718 364294
rect 589098 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 589718 364226
rect 589098 364102 589718 364170
rect 589098 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 589718 364102
rect 589098 363978 589718 364046
rect 592818 478350 593438 495922
rect 592818 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 593438 478350
rect 592818 478226 593438 478294
rect 592818 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 593438 478226
rect 592818 478102 593438 478170
rect 592818 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 593438 478102
rect 592818 477978 593438 478046
rect 592818 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 593438 477978
rect 592818 460350 593438 477922
rect 592818 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 593438 460350
rect 592818 460226 593438 460294
rect 592818 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 593438 460226
rect 592818 460102 593438 460170
rect 592818 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 593438 460102
rect 592818 459978 593438 460046
rect 592818 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 593438 459978
rect 592818 442350 593438 459922
rect 592818 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 593438 442350
rect 592818 442226 593438 442294
rect 592818 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 593438 442226
rect 592818 442102 593438 442170
rect 592818 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 593438 442102
rect 592818 441978 593438 442046
rect 592818 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 593438 441978
rect 592818 424350 593438 441922
rect 592818 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 593438 424350
rect 592818 424226 593438 424294
rect 592818 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 593438 424226
rect 592818 424102 593438 424170
rect 592818 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 593438 424102
rect 592818 423978 593438 424046
rect 592818 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 593438 423978
rect 592818 406350 593438 423922
rect 592818 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 593438 406350
rect 592818 406226 593438 406294
rect 592818 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 593438 406226
rect 592818 406102 593438 406170
rect 592818 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 593438 406102
rect 592818 405978 593438 406046
rect 592818 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 593438 405978
rect 592818 388350 593438 405922
rect 592818 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 593438 388350
rect 592818 388226 593438 388294
rect 592818 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 593438 388226
rect 592818 388102 593438 388170
rect 592818 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 593438 388102
rect 592818 387978 593438 388046
rect 592818 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 593438 387978
rect 592818 370350 593438 387922
rect 592818 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 593438 370350
rect 592818 370226 593438 370294
rect 592818 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 593438 370226
rect 592818 370102 593438 370170
rect 592818 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 593438 370102
rect 592818 369978 593438 370046
rect 592818 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 593438 369978
rect 589098 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 589718 363978
rect 589098 346350 589718 363922
rect 589098 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 589718 346350
rect 589098 346226 589718 346294
rect 589098 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 589718 346226
rect 589098 346102 589718 346170
rect 589098 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 589718 346102
rect 589098 345978 589718 346046
rect 589098 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 589718 345978
rect 589098 328350 589718 345922
rect 589098 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 589718 328350
rect 589098 328226 589718 328294
rect 589098 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 589718 328226
rect 589098 328102 589718 328170
rect 589098 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 589718 328102
rect 589098 327978 589718 328046
rect 589098 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 589718 327978
rect 589098 310350 589718 327922
rect 589098 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 589718 310350
rect 589098 310226 589718 310294
rect 589098 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 589718 310226
rect 589098 310102 589718 310170
rect 589098 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 589718 310102
rect 589098 309978 589718 310046
rect 589098 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 589718 309978
rect 562098 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 562718 280350
rect 562098 280226 562718 280294
rect 562098 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 562718 280226
rect 562098 280102 562718 280170
rect 562098 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 562718 280102
rect 562098 279978 562718 280046
rect 562098 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 562718 279978
rect 562098 262350 562718 279922
rect 562098 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 562718 262350
rect 562098 262226 562718 262294
rect 562098 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 562718 262226
rect 562098 262102 562718 262170
rect 562098 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 562718 262102
rect 562098 261978 562718 262046
rect 562098 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 562718 261978
rect 562098 244350 562718 261922
rect 562098 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 562718 244350
rect 562098 244226 562718 244294
rect 562098 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 562718 244226
rect 562098 244102 562718 244170
rect 562098 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 562718 244102
rect 562098 243978 562718 244046
rect 562098 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 562718 243978
rect 562098 226350 562718 243922
rect 562098 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 562718 226350
rect 562098 226226 562718 226294
rect 562098 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 562718 226226
rect 562098 226102 562718 226170
rect 562098 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 562718 226102
rect 562098 225978 562718 226046
rect 562098 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 562718 225978
rect 562098 208350 562718 225922
rect 562098 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 562718 208350
rect 562098 208226 562718 208294
rect 562098 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 562718 208226
rect 562098 208102 562718 208170
rect 562098 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 562718 208102
rect 562098 207978 562718 208046
rect 562098 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 562718 207978
rect 558378 202294 558474 202350
rect 558530 202294 558598 202350
rect 558654 202294 558722 202350
rect 558778 202294 558846 202350
rect 558902 202294 558998 202350
rect 558378 202226 558998 202294
rect 558378 202170 558474 202226
rect 558530 202170 558598 202226
rect 558654 202170 558722 202226
rect 558778 202170 558846 202226
rect 558902 202170 558998 202226
rect 558378 202102 558998 202170
rect 558378 202046 558474 202102
rect 558530 202046 558598 202102
rect 558654 202046 558722 202102
rect 558778 202046 558846 202102
rect 558902 202046 558998 202102
rect 558378 201978 558998 202046
rect 558378 201922 558474 201978
rect 558530 201922 558598 201978
rect 558654 201922 558722 201978
rect 558778 201922 558846 201978
rect 558902 201922 558998 201978
rect 558378 184350 558998 201922
rect 558378 184294 558474 184350
rect 558530 184294 558598 184350
rect 558654 184294 558722 184350
rect 558778 184294 558846 184350
rect 558902 184294 558998 184350
rect 558378 184226 558998 184294
rect 558378 184170 558474 184226
rect 558530 184170 558598 184226
rect 558654 184170 558722 184226
rect 558778 184170 558846 184226
rect 558902 184170 558998 184226
rect 558378 184102 558998 184170
rect 558378 184046 558474 184102
rect 558530 184046 558598 184102
rect 558654 184046 558722 184102
rect 558778 184046 558846 184102
rect 558902 184046 558998 184102
rect 558378 183978 558998 184046
rect 558378 183922 558474 183978
rect 558530 183922 558598 183978
rect 558654 183922 558722 183978
rect 558778 183922 558846 183978
rect 558902 183922 558998 183978
rect 558378 166350 558998 183922
rect 558378 166294 558474 166350
rect 558530 166294 558598 166350
rect 558654 166294 558722 166350
rect 558778 166294 558846 166350
rect 558902 166294 558998 166350
rect 558378 166226 558998 166294
rect 558378 166170 558474 166226
rect 558530 166170 558598 166226
rect 558654 166170 558722 166226
rect 558778 166170 558846 166226
rect 558902 166170 558998 166226
rect 558378 166102 558998 166170
rect 558378 166046 558474 166102
rect 558530 166046 558598 166102
rect 558654 166046 558722 166102
rect 558778 166046 558846 166102
rect 558902 166046 558998 166102
rect 558378 165978 558998 166046
rect 558378 165922 558474 165978
rect 558530 165922 558598 165978
rect 558654 165922 558722 165978
rect 558778 165922 558846 165978
rect 558902 165922 558998 165978
rect 558378 148350 558998 165922
rect 558378 148294 558474 148350
rect 558530 148294 558598 148350
rect 558654 148294 558722 148350
rect 558778 148294 558846 148350
rect 558902 148294 558998 148350
rect 558378 148226 558998 148294
rect 558378 148170 558474 148226
rect 558530 148170 558598 148226
rect 558654 148170 558722 148226
rect 558778 148170 558846 148226
rect 558902 148170 558998 148226
rect 558378 148102 558998 148170
rect 558378 148046 558474 148102
rect 558530 148046 558598 148102
rect 558654 148046 558722 148102
rect 558778 148046 558846 148102
rect 558902 148046 558998 148102
rect 558378 147978 558998 148046
rect 558378 147922 558474 147978
rect 558530 147922 558598 147978
rect 558654 147922 558722 147978
rect 558778 147922 558846 147978
rect 558902 147922 558998 147978
rect 558378 130350 558998 147922
rect 558378 130294 558474 130350
rect 558530 130294 558598 130350
rect 558654 130294 558722 130350
rect 558778 130294 558846 130350
rect 558902 130294 558998 130350
rect 558378 130226 558998 130294
rect 558378 130170 558474 130226
rect 558530 130170 558598 130226
rect 558654 130170 558722 130226
rect 558778 130170 558846 130226
rect 558902 130170 558998 130226
rect 558378 130102 558998 130170
rect 558378 130046 558474 130102
rect 558530 130046 558598 130102
rect 558654 130046 558722 130102
rect 558778 130046 558846 130102
rect 558902 130046 558998 130102
rect 558378 129978 558998 130046
rect 558378 129922 558474 129978
rect 558530 129922 558598 129978
rect 558654 129922 558722 129978
rect 558778 129922 558846 129978
rect 558902 129922 558998 129978
rect 558378 112350 558998 129922
rect 558378 112294 558474 112350
rect 558530 112294 558598 112350
rect 558654 112294 558722 112350
rect 558778 112294 558846 112350
rect 558902 112294 558998 112350
rect 558378 112226 558998 112294
rect 558378 112170 558474 112226
rect 558530 112170 558598 112226
rect 558654 112170 558722 112226
rect 558778 112170 558846 112226
rect 558902 112170 558998 112226
rect 558378 112102 558998 112170
rect 558378 112046 558474 112102
rect 558530 112046 558598 112102
rect 558654 112046 558722 112102
rect 558778 112046 558846 112102
rect 558902 112046 558998 112102
rect 558378 111978 558998 112046
rect 558378 111922 558474 111978
rect 558530 111922 558598 111978
rect 558654 111922 558722 111978
rect 558778 111922 558846 111978
rect 558902 111922 558998 111978
rect 558378 94350 558998 111922
rect 558378 94294 558474 94350
rect 558530 94294 558598 94350
rect 558654 94294 558722 94350
rect 558778 94294 558846 94350
rect 558902 94294 558998 94350
rect 558378 94226 558998 94294
rect 558378 94170 558474 94226
rect 558530 94170 558598 94226
rect 558654 94170 558722 94226
rect 558778 94170 558846 94226
rect 558902 94170 558998 94226
rect 558378 94102 558998 94170
rect 558378 94046 558474 94102
rect 558530 94046 558598 94102
rect 558654 94046 558722 94102
rect 558778 94046 558846 94102
rect 558902 94046 558998 94102
rect 558378 93978 558998 94046
rect 558378 93922 558474 93978
rect 558530 93922 558598 93978
rect 558654 93922 558722 93978
rect 558778 93922 558846 93978
rect 558902 93922 558998 93978
rect 555212 28354 555268 28364
rect 556892 86436 556948 86446
rect 553532 21634 553588 21644
rect 551852 14914 551908 14924
rect 556892 13860 556948 86380
rect 556892 13794 556948 13804
rect 558378 76350 558998 93922
rect 558378 76294 558474 76350
rect 558530 76294 558598 76350
rect 558654 76294 558722 76350
rect 558778 76294 558846 76350
rect 558902 76294 558998 76350
rect 558378 76226 558998 76294
rect 558378 76170 558474 76226
rect 558530 76170 558598 76226
rect 558654 76170 558722 76226
rect 558778 76170 558846 76226
rect 558902 76170 558998 76226
rect 558378 76102 558998 76170
rect 558378 76046 558474 76102
rect 558530 76046 558598 76102
rect 558654 76046 558722 76102
rect 558778 76046 558846 76102
rect 558902 76046 558998 76102
rect 558378 75978 558998 76046
rect 558378 75922 558474 75978
rect 558530 75922 558598 75978
rect 558654 75922 558722 75978
rect 558778 75922 558846 75978
rect 558902 75922 558998 75978
rect 558378 58350 558998 75922
rect 558378 58294 558474 58350
rect 558530 58294 558598 58350
rect 558654 58294 558722 58350
rect 558778 58294 558846 58350
rect 558902 58294 558998 58350
rect 558378 58226 558998 58294
rect 558378 58170 558474 58226
rect 558530 58170 558598 58226
rect 558654 58170 558722 58226
rect 558778 58170 558846 58226
rect 558902 58170 558998 58226
rect 558378 58102 558998 58170
rect 558378 58046 558474 58102
rect 558530 58046 558598 58102
rect 558654 58046 558722 58102
rect 558778 58046 558846 58102
rect 558902 58046 558998 58102
rect 558378 57978 558998 58046
rect 558378 57922 558474 57978
rect 558530 57922 558598 57978
rect 558654 57922 558722 57978
rect 558778 57922 558846 57978
rect 558902 57922 558998 57978
rect 558378 40350 558998 57922
rect 558378 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 558998 40350
rect 558378 40226 558998 40294
rect 558378 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 558998 40226
rect 558378 40102 558998 40170
rect 558378 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 558998 40102
rect 558378 39978 558998 40046
rect 558378 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 558998 39978
rect 558378 22350 558998 39922
rect 560252 205380 560308 205390
rect 560252 23940 560308 205324
rect 560252 23874 560308 23884
rect 562098 190350 562718 207922
rect 562098 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 562718 190350
rect 562098 190226 562718 190294
rect 562098 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 562718 190226
rect 562098 190102 562718 190170
rect 562098 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 562718 190102
rect 562098 189978 562718 190046
rect 562098 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 562718 189978
rect 562098 172350 562718 189922
rect 562098 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 562718 172350
rect 562098 172226 562718 172294
rect 562098 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 562718 172226
rect 562098 172102 562718 172170
rect 562098 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 562718 172102
rect 562098 171978 562718 172046
rect 562098 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 562718 171978
rect 562098 154350 562718 171922
rect 562098 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 562718 154350
rect 562098 154226 562718 154294
rect 562098 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 562718 154226
rect 562098 154102 562718 154170
rect 562098 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 562718 154102
rect 562098 153978 562718 154046
rect 562098 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 562718 153978
rect 562098 136350 562718 153922
rect 562098 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 562718 136350
rect 562098 136226 562718 136294
rect 562098 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 562718 136226
rect 562098 136102 562718 136170
rect 562098 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 562718 136102
rect 562098 135978 562718 136046
rect 562098 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 562718 135978
rect 562098 118350 562718 135922
rect 562098 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 562718 118350
rect 562098 118226 562718 118294
rect 562098 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 562718 118226
rect 562098 118102 562718 118170
rect 562098 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 562718 118102
rect 562098 117978 562718 118046
rect 562098 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 562718 117978
rect 562098 100350 562718 117922
rect 562098 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 562718 100350
rect 562098 100226 562718 100294
rect 562098 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 562718 100226
rect 562098 100102 562718 100170
rect 562098 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 562718 100102
rect 562098 99978 562718 100046
rect 562098 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 562718 99978
rect 562098 82350 562718 99922
rect 562098 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 562718 82350
rect 562098 82226 562718 82294
rect 562098 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 562718 82226
rect 562098 82102 562718 82170
rect 562098 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 562718 82102
rect 562098 81978 562718 82046
rect 562098 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 562718 81978
rect 562098 64350 562718 81922
rect 562098 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 562718 64350
rect 562098 64226 562718 64294
rect 562098 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 562718 64226
rect 562098 64102 562718 64170
rect 562098 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 562718 64102
rect 562098 63978 562718 64046
rect 562098 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 562718 63978
rect 562098 46350 562718 63922
rect 562098 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 562718 46350
rect 562098 46226 562718 46294
rect 562098 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 562718 46226
rect 562098 46102 562718 46170
rect 562098 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 562718 46102
rect 562098 45978 562718 46046
rect 562098 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 562718 45978
rect 562098 28350 562718 45922
rect 563612 296548 563668 296558
rect 563612 31780 563668 296492
rect 589098 292350 589718 309922
rect 590492 363972 590548 363982
rect 590156 297892 590212 297902
rect 590156 296548 590212 297836
rect 590156 296482 590212 296492
rect 589098 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 589718 292350
rect 589098 292226 589718 292294
rect 589098 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 589718 292226
rect 589098 292102 589718 292170
rect 589098 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 589718 292102
rect 589098 291978 589718 292046
rect 589098 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 589718 291978
rect 563612 31714 563668 31724
rect 565292 284676 565348 284686
rect 565292 30660 565348 284620
rect 589098 274350 589718 291922
rect 590492 278068 590548 363916
rect 590492 278002 590548 278012
rect 592818 352350 593438 369922
rect 592818 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 593438 352350
rect 592818 352226 593438 352294
rect 592818 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 593438 352226
rect 592818 352102 593438 352170
rect 592818 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 593438 352102
rect 592818 351978 593438 352046
rect 592818 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 593438 351978
rect 592818 334350 593438 351922
rect 592818 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 593438 334350
rect 592818 334226 593438 334294
rect 592818 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 593438 334226
rect 592818 334102 593438 334170
rect 592818 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 593438 334102
rect 592818 333978 593438 334046
rect 592818 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 593438 333978
rect 592818 316350 593438 333922
rect 592818 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 593438 316350
rect 592818 316226 593438 316294
rect 592818 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 593438 316226
rect 592818 316102 593438 316170
rect 592818 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 593438 316102
rect 592818 315978 593438 316046
rect 592818 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 593438 315978
rect 592818 298350 593438 315922
rect 592818 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 593438 298350
rect 592818 298226 593438 298294
rect 592818 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 593438 298226
rect 592818 298102 593438 298170
rect 592818 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 593438 298102
rect 592818 297978 593438 298046
rect 592818 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 593438 297978
rect 592818 280350 593438 297922
rect 592818 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 593438 280350
rect 592818 280226 593438 280294
rect 592818 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 593438 280226
rect 592818 280102 593438 280170
rect 592818 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 593438 280102
rect 592818 279978 593438 280046
rect 592818 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 593438 279978
rect 589098 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 589718 274350
rect 589098 274226 589718 274294
rect 589098 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 589718 274226
rect 589098 274102 589718 274170
rect 589098 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 589718 274102
rect 589098 273978 589718 274046
rect 589098 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 589718 273978
rect 589098 256350 589718 273922
rect 589098 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 589718 256350
rect 589098 256226 589718 256294
rect 589098 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 589718 256226
rect 589098 256102 589718 256170
rect 589098 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 589718 256102
rect 589098 255978 589718 256046
rect 589098 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 589718 255978
rect 587132 245028 587188 245038
rect 565292 30594 565348 30604
rect 572012 126084 572068 126094
rect 562098 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 562718 28350
rect 562098 28226 562718 28294
rect 562098 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 562718 28226
rect 562098 28102 562718 28170
rect 562098 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 562718 28102
rect 562098 27978 562718 28046
rect 562098 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 562718 27978
rect 558378 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 558998 22350
rect 558378 22226 558998 22294
rect 558378 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 558998 22226
rect 558378 22102 558998 22170
rect 558378 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 558998 22102
rect 558378 21978 558998 22046
rect 558378 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 558998 21978
rect 550284 9314 550340 9324
rect 548492 8194 548548 8204
rect 557788 5158 557844 5168
rect 557788 3444 557844 5102
rect 557788 3378 557844 3388
rect 558378 4350 558998 21922
rect 558378 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 558998 4350
rect 558378 4226 558998 4294
rect 558378 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 558998 4226
rect 558378 4102 558998 4170
rect 558378 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 558998 4102
rect 558378 3978 558998 4046
rect 558378 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 558998 3978
rect 531378 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 531998 -1120
rect 531378 -1244 531998 -1176
rect 531378 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 531998 -1244
rect 531378 -1368 531998 -1300
rect 531378 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 531998 -1368
rect 531378 -1492 531998 -1424
rect 531378 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 531998 -1492
rect 531378 -1644 531998 -1548
rect 558378 -160 558998 3922
rect 558378 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 558998 -160
rect 558378 -284 558998 -216
rect 558378 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 558998 -284
rect 558378 -408 558998 -340
rect 558378 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 558998 -408
rect 558378 -532 558998 -464
rect 558378 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 558998 -532
rect 558378 -1644 558998 -588
rect 562098 10350 562718 27922
rect 572012 17220 572068 126028
rect 587132 29428 587188 244972
rect 587132 29362 587188 29372
rect 589098 238350 589718 255922
rect 589098 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 589718 238350
rect 589098 238226 589718 238294
rect 589098 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 589718 238226
rect 589098 238102 589718 238170
rect 589098 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 589718 238102
rect 589098 237978 589718 238046
rect 589098 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 589718 237978
rect 589098 220350 589718 237922
rect 589098 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 589718 220350
rect 589098 220226 589718 220294
rect 589098 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 589718 220226
rect 589098 220102 589718 220170
rect 589098 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 589718 220102
rect 589098 219978 589718 220046
rect 589098 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 589718 219978
rect 589098 202350 589718 219922
rect 589098 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 589718 202350
rect 589098 202226 589718 202294
rect 589098 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 589718 202226
rect 589098 202102 589718 202170
rect 589098 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 589718 202102
rect 589098 201978 589718 202046
rect 589098 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 589718 201978
rect 589098 184350 589718 201922
rect 589098 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 589718 184350
rect 589098 184226 589718 184294
rect 589098 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 589718 184226
rect 589098 184102 589718 184170
rect 589098 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 589718 184102
rect 589098 183978 589718 184046
rect 589098 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 589718 183978
rect 589098 166350 589718 183922
rect 589098 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 589718 166350
rect 589098 166226 589718 166294
rect 589098 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 589718 166226
rect 589098 166102 589718 166170
rect 589098 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 589718 166102
rect 589098 165978 589718 166046
rect 589098 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 589718 165978
rect 589098 148350 589718 165922
rect 592818 262350 593438 279922
rect 592818 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 593438 262350
rect 592818 262226 593438 262294
rect 592818 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 593438 262226
rect 592818 262102 593438 262170
rect 592818 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 593438 262102
rect 592818 261978 593438 262046
rect 592818 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 593438 261978
rect 592818 244350 593438 261922
rect 592818 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 593438 244350
rect 592818 244226 593438 244294
rect 592818 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 593438 244226
rect 592818 244102 593438 244170
rect 592818 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 593438 244102
rect 592818 243978 593438 244046
rect 592818 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 593438 243978
rect 592818 226350 593438 243922
rect 592818 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 593438 226350
rect 592818 226226 593438 226294
rect 592818 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 593438 226226
rect 592818 226102 593438 226170
rect 592818 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 593438 226102
rect 592818 225978 593438 226046
rect 592818 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 593438 225978
rect 592818 208350 593438 225922
rect 592818 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 593438 208350
rect 592818 208226 593438 208294
rect 592818 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 593438 208226
rect 592818 208102 593438 208170
rect 592818 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 593438 208102
rect 592818 207978 593438 208046
rect 592818 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 593438 207978
rect 592818 190350 593438 207922
rect 592818 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 593438 190350
rect 592818 190226 593438 190294
rect 592818 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 593438 190226
rect 592818 190102 593438 190170
rect 592818 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 593438 190102
rect 592818 189978 593438 190046
rect 592818 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 593438 189978
rect 592818 172350 593438 189922
rect 592818 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 593438 172350
rect 592818 172226 593438 172294
rect 592818 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 593438 172226
rect 592818 172102 593438 172170
rect 592818 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 593438 172102
rect 592818 171978 593438 172046
rect 592818 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 593438 171978
rect 589098 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 589718 148350
rect 589098 148226 589718 148294
rect 589098 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 589718 148226
rect 589098 148102 589718 148170
rect 589098 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 589718 148102
rect 589098 147978 589718 148046
rect 589098 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 589718 147978
rect 589098 130350 589718 147922
rect 589098 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 589718 130350
rect 589098 130226 589718 130294
rect 589098 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 589718 130226
rect 589098 130102 589718 130170
rect 589098 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 589718 130102
rect 589098 129978 589718 130046
rect 589098 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 589718 129978
rect 589098 112350 589718 129922
rect 589098 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 589718 112350
rect 589098 112226 589718 112294
rect 589098 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 589718 112226
rect 589098 112102 589718 112170
rect 589098 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 589718 112102
rect 589098 111978 589718 112046
rect 589098 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 589718 111978
rect 589098 94350 589718 111922
rect 590492 165732 590548 165742
rect 590156 99652 590212 99662
rect 590156 98308 590212 99596
rect 590156 98242 590212 98252
rect 589098 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 589718 94350
rect 589098 94226 589718 94294
rect 589098 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 589718 94226
rect 589098 94102 589718 94170
rect 589098 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 589718 94102
rect 589098 93978 589718 94046
rect 589098 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 589718 93978
rect 589098 76350 589718 93922
rect 589098 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 589718 76350
rect 589098 76226 589718 76294
rect 589098 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 589718 76226
rect 589098 76102 589718 76170
rect 589098 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 589718 76102
rect 589098 75978 589718 76046
rect 589098 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 589718 75978
rect 589098 58350 589718 75922
rect 589098 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 589718 58350
rect 589098 58226 589718 58294
rect 589098 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 589718 58226
rect 589098 58102 589718 58170
rect 589098 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 589718 58102
rect 589098 57978 589718 58046
rect 589098 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 589718 57978
rect 589098 40350 589718 57922
rect 589098 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 589718 40350
rect 589098 40226 589718 40294
rect 589098 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 589718 40226
rect 589098 40102 589718 40170
rect 589098 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 589718 40102
rect 589098 39978 589718 40046
rect 589098 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 589718 39978
rect 572012 17154 572068 17164
rect 589098 22350 589718 39922
rect 590492 24388 590548 165676
rect 592818 154350 593438 171922
rect 592818 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 593438 154350
rect 592818 154226 593438 154294
rect 592818 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 593438 154226
rect 592818 154102 593438 154170
rect 592818 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 593438 154102
rect 592818 153978 593438 154046
rect 592818 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 593438 153978
rect 592818 136350 593438 153922
rect 592818 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 593438 136350
rect 592818 136226 593438 136294
rect 592818 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 593438 136226
rect 592818 136102 593438 136170
rect 592818 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 593438 136102
rect 592818 135978 593438 136046
rect 592818 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 593438 135978
rect 592818 118350 593438 135922
rect 592818 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 593438 118350
rect 592818 118226 593438 118294
rect 592818 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 593438 118226
rect 592818 118102 593438 118170
rect 592818 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 593438 118102
rect 592818 117978 593438 118046
rect 592818 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 593438 117978
rect 592818 100350 593438 117922
rect 592818 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 593438 100350
rect 592818 100226 593438 100294
rect 592818 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 593438 100226
rect 592818 100102 593438 100170
rect 592818 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 593438 100102
rect 592818 99978 593438 100046
rect 592818 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 593438 99978
rect 592818 82350 593438 99922
rect 592818 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 593438 82350
rect 592818 82226 593438 82294
rect 592818 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 593438 82226
rect 592818 82102 593438 82170
rect 592818 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 593438 82102
rect 592818 81978 593438 82046
rect 592818 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 593438 81978
rect 592818 64350 593438 81922
rect 592818 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 593438 64350
rect 592818 64226 593438 64294
rect 592818 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 593438 64226
rect 592818 64102 593438 64170
rect 592818 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 593438 64102
rect 592818 63978 593438 64046
rect 592818 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 593438 63978
rect 590492 24322 590548 24332
rect 590604 46788 590660 46798
rect 589098 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 589718 22350
rect 589098 22226 589718 22294
rect 589098 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 589718 22226
rect 589098 22102 589718 22170
rect 589098 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 589718 22102
rect 589098 21978 589718 22046
rect 589098 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 589718 21978
rect 562098 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 562718 10350
rect 562098 10226 562718 10294
rect 562098 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 562718 10226
rect 562098 10102 562718 10170
rect 562098 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 562718 10102
rect 562098 9978 562718 10046
rect 562098 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 562718 9978
rect 562098 -1120 562718 9922
rect 589098 4350 589718 21922
rect 590604 12628 590660 46732
rect 592818 46350 593438 63922
rect 592818 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 593438 46350
rect 592818 46226 593438 46294
rect 592818 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 593438 46226
rect 592818 46102 593438 46170
rect 592818 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 593438 46102
rect 592818 45978 593438 46046
rect 592818 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 593438 45978
rect 592818 28350 593438 45922
rect 592818 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 593438 28350
rect 592818 28226 593438 28294
rect 592818 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 593438 28226
rect 592818 28102 593438 28170
rect 592818 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 593438 28102
rect 592818 27978 593438 28046
rect 592818 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 593438 27978
rect 591276 20356 591332 20366
rect 591276 19348 591332 20300
rect 591276 19282 591332 19292
rect 590604 12562 590660 12572
rect 589098 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 589718 4350
rect 589098 4226 589718 4294
rect 589098 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 589718 4226
rect 589098 4102 589718 4170
rect 589098 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 589718 4102
rect 589098 3978 589718 4046
rect 589098 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 589718 3978
rect 565404 3444 565460 3454
rect 565404 3358 565460 3388
rect 565404 3292 565460 3302
rect 563500 3178 563556 3188
rect 563500 1764 563556 3122
rect 563500 1698 563556 1708
rect 569212 644 569268 654
rect 569212 118 569268 588
rect 571228 644 571284 654
rect 571228 298 571284 588
rect 571228 232 571284 242
rect 569212 52 569268 62
rect 562098 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 562718 -1120
rect 562098 -1244 562718 -1176
rect 562098 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 562718 -1244
rect 562098 -1368 562718 -1300
rect 562098 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 562718 -1368
rect 562098 -1492 562718 -1424
rect 562098 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 562718 -1492
rect 562098 -1644 562718 -1548
rect 589098 -160 589718 3922
rect 589098 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 589718 -160
rect 589098 -284 589718 -216
rect 589098 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 589718 -284
rect 589098 -408 589718 -340
rect 589098 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 589718 -408
rect 589098 -532 589718 -464
rect 589098 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 589718 -532
rect 589098 -1644 589718 -588
rect 592818 10350 593438 27922
rect 592818 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 593438 10350
rect 592818 10226 593438 10294
rect 592818 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 593438 10226
rect 592818 10102 593438 10170
rect 592818 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 593438 10102
rect 592818 9978 593438 10046
rect 592818 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 593438 9978
rect 592818 -1120 593438 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 592818 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 593438 -1120
rect 592818 -1244 593438 -1176
rect 592818 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 593438 -1244
rect 592818 -1368 593438 -1300
rect 592818 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 593438 -1368
rect 592818 -1492 593438 -1424
rect 592818 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 593438 -1492
rect 592818 -1644 593438 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect 5514 597156 5570 597212
rect 5638 597156 5694 597212
rect 5762 597156 5818 597212
rect 5886 597156 5942 597212
rect 5514 597032 5570 597088
rect 5638 597032 5694 597088
rect 5762 597032 5818 597088
rect 5886 597032 5942 597088
rect 5514 596908 5570 596964
rect 5638 596908 5694 596964
rect 5762 596908 5818 596964
rect 5886 596908 5942 596964
rect 5514 596784 5570 596840
rect 5638 596784 5694 596840
rect 5762 596784 5818 596840
rect 5886 596784 5942 596840
rect 5514 580294 5570 580350
rect 5638 580294 5694 580350
rect 5762 580294 5818 580350
rect 5886 580294 5942 580350
rect 5514 580170 5570 580226
rect 5638 580170 5694 580226
rect 5762 580170 5818 580226
rect 5886 580170 5942 580226
rect 5514 580046 5570 580102
rect 5638 580046 5694 580102
rect 5762 580046 5818 580102
rect 5886 580046 5942 580102
rect 5514 579922 5570 579978
rect 5638 579922 5694 579978
rect 5762 579922 5818 579978
rect 5886 579922 5942 579978
rect 5514 562294 5570 562350
rect 5638 562294 5694 562350
rect 5762 562294 5818 562350
rect 5886 562294 5942 562350
rect 5514 562170 5570 562226
rect 5638 562170 5694 562226
rect 5762 562170 5818 562226
rect 5886 562170 5942 562226
rect 5514 562046 5570 562102
rect 5638 562046 5694 562102
rect 5762 562046 5818 562102
rect 5886 562046 5942 562102
rect 5514 561922 5570 561978
rect 5638 561922 5694 561978
rect 5762 561922 5818 561978
rect 5886 561922 5942 561978
rect 5514 544294 5570 544350
rect 5638 544294 5694 544350
rect 5762 544294 5818 544350
rect 5886 544294 5942 544350
rect 5514 544170 5570 544226
rect 5638 544170 5694 544226
rect 5762 544170 5818 544226
rect 5886 544170 5942 544226
rect 5514 544046 5570 544102
rect 5638 544046 5694 544102
rect 5762 544046 5818 544102
rect 5886 544046 5942 544102
rect 5514 543922 5570 543978
rect 5638 543922 5694 543978
rect 5762 543922 5818 543978
rect 5886 543922 5942 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect 28 273482 84 273538
rect 1596 361322 1652 361378
rect 140 271862 196 271918
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect 28 267902 84 267958
rect 140 266462 196 266518
rect 5514 526294 5570 526350
rect 5638 526294 5694 526350
rect 5762 526294 5818 526350
rect 5886 526294 5942 526350
rect 5514 526170 5570 526226
rect 5638 526170 5694 526226
rect 5762 526170 5818 526226
rect 5886 526170 5942 526226
rect 5514 526046 5570 526102
rect 5638 526046 5694 526102
rect 5762 526046 5818 526102
rect 5886 526046 5942 526102
rect 5514 525922 5570 525978
rect 5638 525922 5694 525978
rect 5762 525922 5818 525978
rect 5886 525922 5942 525978
rect 5514 508294 5570 508350
rect 5638 508294 5694 508350
rect 5762 508294 5818 508350
rect 5886 508294 5942 508350
rect 5514 508170 5570 508226
rect 5638 508170 5694 508226
rect 5762 508170 5818 508226
rect 5886 508170 5942 508226
rect 5514 508046 5570 508102
rect 5638 508046 5694 508102
rect 5762 508046 5818 508102
rect 5886 508046 5942 508102
rect 5514 507922 5570 507978
rect 5638 507922 5694 507978
rect 5762 507922 5818 507978
rect 5886 507922 5942 507978
rect 5514 490294 5570 490350
rect 5638 490294 5694 490350
rect 5762 490294 5818 490350
rect 5886 490294 5942 490350
rect 5514 490170 5570 490226
rect 5638 490170 5694 490226
rect 5762 490170 5818 490226
rect 5886 490170 5942 490226
rect 5514 490046 5570 490102
rect 5638 490046 5694 490102
rect 5762 490046 5818 490102
rect 5886 490046 5942 490102
rect 5514 489922 5570 489978
rect 5638 489922 5694 489978
rect 5762 489922 5818 489978
rect 5886 489922 5942 489978
rect 2492 273662 2548 273718
rect 2940 366362 2996 366418
rect 3052 331982 3108 332038
rect 3052 281582 3108 281638
rect 5514 472294 5570 472350
rect 5638 472294 5694 472350
rect 5762 472294 5818 472350
rect 5886 472294 5942 472350
rect 5514 472170 5570 472226
rect 5638 472170 5694 472226
rect 5762 472170 5818 472226
rect 5886 472170 5942 472226
rect 5514 472046 5570 472102
rect 5638 472046 5694 472102
rect 5762 472046 5818 472102
rect 5886 472046 5942 472102
rect 5514 471922 5570 471978
rect 5638 471922 5694 471978
rect 5762 471922 5818 471978
rect 5886 471922 5942 471978
rect 5514 454294 5570 454350
rect 5638 454294 5694 454350
rect 5762 454294 5818 454350
rect 5886 454294 5942 454350
rect 5514 454170 5570 454226
rect 5638 454170 5694 454226
rect 5762 454170 5818 454226
rect 5886 454170 5942 454226
rect 5514 454046 5570 454102
rect 5638 454046 5694 454102
rect 5762 454046 5818 454102
rect 5886 454046 5942 454102
rect 5514 453922 5570 453978
rect 5638 453922 5694 453978
rect 5762 453922 5818 453978
rect 5886 453922 5942 453978
rect 4284 272042 4340 272098
rect 5514 436294 5570 436350
rect 5638 436294 5694 436350
rect 5762 436294 5818 436350
rect 5886 436294 5942 436350
rect 5514 436170 5570 436226
rect 5638 436170 5694 436226
rect 5762 436170 5818 436226
rect 5886 436170 5942 436226
rect 5514 436046 5570 436102
rect 5638 436046 5694 436102
rect 5762 436046 5818 436102
rect 5886 436046 5942 436102
rect 5514 435922 5570 435978
rect 5638 435922 5694 435978
rect 5762 435922 5818 435978
rect 5886 435922 5942 435978
rect 5514 418294 5570 418350
rect 5638 418294 5694 418350
rect 5762 418294 5818 418350
rect 5886 418294 5942 418350
rect 5514 418170 5570 418226
rect 5638 418170 5694 418226
rect 5762 418170 5818 418226
rect 5886 418170 5942 418226
rect 5514 418046 5570 418102
rect 5638 418046 5694 418102
rect 5762 418046 5818 418102
rect 5886 418046 5942 418102
rect 5514 417922 5570 417978
rect 5638 417922 5694 417978
rect 5762 417922 5818 417978
rect 5886 417922 5942 417978
rect 5514 400294 5570 400350
rect 5638 400294 5694 400350
rect 5762 400294 5818 400350
rect 5886 400294 5942 400350
rect 5514 400170 5570 400226
rect 5638 400170 5694 400226
rect 5762 400170 5818 400226
rect 5886 400170 5942 400226
rect 5514 400046 5570 400102
rect 5638 400046 5694 400102
rect 5762 400046 5818 400102
rect 5886 400046 5942 400102
rect 5514 399922 5570 399978
rect 5638 399922 5694 399978
rect 5762 399922 5818 399978
rect 5886 399922 5942 399978
rect 5514 382294 5570 382350
rect 5638 382294 5694 382350
rect 5762 382294 5818 382350
rect 5886 382294 5942 382350
rect 5514 382170 5570 382226
rect 5638 382170 5694 382226
rect 5762 382170 5818 382226
rect 5886 382170 5942 382226
rect 5514 382046 5570 382102
rect 5638 382046 5694 382102
rect 5762 382046 5818 382102
rect 5886 382046 5942 382102
rect 5514 381922 5570 381978
rect 5638 381922 5694 381978
rect 5762 381922 5818 381978
rect 5886 381922 5942 381978
rect 5514 364294 5570 364350
rect 5638 364294 5694 364350
rect 5762 364294 5818 364350
rect 5886 364294 5942 364350
rect 5514 364170 5570 364226
rect 5638 364170 5694 364226
rect 5762 364170 5818 364226
rect 5886 364170 5942 364226
rect 5514 364046 5570 364102
rect 5638 364046 5694 364102
rect 5762 364046 5818 364102
rect 5886 364046 5942 364102
rect 5514 363922 5570 363978
rect 5638 363922 5694 363978
rect 5762 363922 5818 363978
rect 5886 363922 5942 363978
rect 5514 346294 5570 346350
rect 5638 346294 5694 346350
rect 5762 346294 5818 346350
rect 5886 346294 5942 346350
rect 5514 346170 5570 346226
rect 5638 346170 5694 346226
rect 5762 346170 5818 346226
rect 5886 346170 5942 346226
rect 5514 346046 5570 346102
rect 5638 346046 5694 346102
rect 5762 346046 5818 346102
rect 5886 346046 5942 346102
rect 5514 345922 5570 345978
rect 5638 345922 5694 345978
rect 5762 345922 5818 345978
rect 5886 345922 5942 345978
rect 5068 331802 5124 331858
rect 4732 290780 4788 290818
rect 4732 290762 4788 290780
rect 9234 598116 9290 598172
rect 9358 598116 9414 598172
rect 9482 598116 9538 598172
rect 9606 598116 9662 598172
rect 9234 597992 9290 598048
rect 9358 597992 9414 598048
rect 9482 597992 9538 598048
rect 9606 597992 9662 598048
rect 9234 597868 9290 597924
rect 9358 597868 9414 597924
rect 9482 597868 9538 597924
rect 9606 597868 9662 597924
rect 9234 597744 9290 597800
rect 9358 597744 9414 597800
rect 9482 597744 9538 597800
rect 9606 597744 9662 597800
rect 9234 586294 9290 586350
rect 9358 586294 9414 586350
rect 9482 586294 9538 586350
rect 9606 586294 9662 586350
rect 9234 586170 9290 586226
rect 9358 586170 9414 586226
rect 9482 586170 9538 586226
rect 9606 586170 9662 586226
rect 9234 586046 9290 586102
rect 9358 586046 9414 586102
rect 9482 586046 9538 586102
rect 9606 586046 9662 586102
rect 9234 585922 9290 585978
rect 9358 585922 9414 585978
rect 9482 585922 9538 585978
rect 9606 585922 9662 585978
rect 9234 568294 9290 568350
rect 9358 568294 9414 568350
rect 9482 568294 9538 568350
rect 9606 568294 9662 568350
rect 9234 568170 9290 568226
rect 9358 568170 9414 568226
rect 9482 568170 9538 568226
rect 9606 568170 9662 568226
rect 9234 568046 9290 568102
rect 9358 568046 9414 568102
rect 9482 568046 9538 568102
rect 9606 568046 9662 568102
rect 9234 567922 9290 567978
rect 9358 567922 9414 567978
rect 9482 567922 9538 567978
rect 9606 567922 9662 567978
rect 9234 550294 9290 550350
rect 9358 550294 9414 550350
rect 9482 550294 9538 550350
rect 9606 550294 9662 550350
rect 9234 550170 9290 550226
rect 9358 550170 9414 550226
rect 9482 550170 9538 550226
rect 9606 550170 9662 550226
rect 9234 550046 9290 550102
rect 9358 550046 9414 550102
rect 9482 550046 9538 550102
rect 9606 550046 9662 550102
rect 9234 549922 9290 549978
rect 9358 549922 9414 549978
rect 9482 549922 9538 549978
rect 9606 549922 9662 549978
rect 9234 532294 9290 532350
rect 9358 532294 9414 532350
rect 9482 532294 9538 532350
rect 9606 532294 9662 532350
rect 9234 532170 9290 532226
rect 9358 532170 9414 532226
rect 9482 532170 9538 532226
rect 9606 532170 9662 532226
rect 9234 532046 9290 532102
rect 9358 532046 9414 532102
rect 9482 532046 9538 532102
rect 9606 532046 9662 532102
rect 9234 531922 9290 531978
rect 9358 531922 9414 531978
rect 9482 531922 9538 531978
rect 9606 531922 9662 531978
rect 9234 514294 9290 514350
rect 9358 514294 9414 514350
rect 9482 514294 9538 514350
rect 9606 514294 9662 514350
rect 9234 514170 9290 514226
rect 9358 514170 9414 514226
rect 9482 514170 9538 514226
rect 9606 514170 9662 514226
rect 9234 514046 9290 514102
rect 9358 514046 9414 514102
rect 9482 514046 9538 514102
rect 9606 514046 9662 514102
rect 9234 513922 9290 513978
rect 9358 513922 9414 513978
rect 9482 513922 9538 513978
rect 9606 513922 9662 513978
rect 9234 496294 9290 496350
rect 9358 496294 9414 496350
rect 9482 496294 9538 496350
rect 9606 496294 9662 496350
rect 9234 496170 9290 496226
rect 9358 496170 9414 496226
rect 9482 496170 9538 496226
rect 9606 496170 9662 496226
rect 9234 496046 9290 496102
rect 9358 496046 9414 496102
rect 9482 496046 9538 496102
rect 9606 496046 9662 496102
rect 9234 495922 9290 495978
rect 9358 495922 9414 495978
rect 9482 495922 9538 495978
rect 9606 495922 9662 495978
rect 9234 478294 9290 478350
rect 9358 478294 9414 478350
rect 9482 478294 9538 478350
rect 9606 478294 9662 478350
rect 9234 478170 9290 478226
rect 9358 478170 9414 478226
rect 9482 478170 9538 478226
rect 9606 478170 9662 478226
rect 9234 478046 9290 478102
rect 9358 478046 9414 478102
rect 9482 478046 9538 478102
rect 9606 478046 9662 478102
rect 9234 477922 9290 477978
rect 9358 477922 9414 477978
rect 9482 477922 9538 477978
rect 9606 477922 9662 477978
rect 9234 460294 9290 460350
rect 9358 460294 9414 460350
rect 9482 460294 9538 460350
rect 9606 460294 9662 460350
rect 9234 460170 9290 460226
rect 9358 460170 9414 460226
rect 9482 460170 9538 460226
rect 9606 460170 9662 460226
rect 9234 460046 9290 460102
rect 9358 460046 9414 460102
rect 9482 460046 9538 460102
rect 9606 460046 9662 460102
rect 9234 459922 9290 459978
rect 9358 459922 9414 459978
rect 9482 459922 9538 459978
rect 9606 459922 9662 459978
rect 9234 442294 9290 442350
rect 9358 442294 9414 442350
rect 9482 442294 9538 442350
rect 9606 442294 9662 442350
rect 9234 442170 9290 442226
rect 9358 442170 9414 442226
rect 9482 442170 9538 442226
rect 9606 442170 9662 442226
rect 9234 442046 9290 442102
rect 9358 442046 9414 442102
rect 9482 442046 9538 442102
rect 9606 442046 9662 442102
rect 9234 441922 9290 441978
rect 9358 441922 9414 441978
rect 9482 441922 9538 441978
rect 9606 441922 9662 441978
rect 9234 424294 9290 424350
rect 9358 424294 9414 424350
rect 9482 424294 9538 424350
rect 9606 424294 9662 424350
rect 9234 424170 9290 424226
rect 9358 424170 9414 424226
rect 9482 424170 9538 424226
rect 9606 424170 9662 424226
rect 9234 424046 9290 424102
rect 9358 424046 9414 424102
rect 9482 424046 9538 424102
rect 9606 424046 9662 424102
rect 9234 423922 9290 423978
rect 9358 423922 9414 423978
rect 9482 423922 9538 423978
rect 9606 423922 9662 423978
rect 9234 406294 9290 406350
rect 9358 406294 9414 406350
rect 9482 406294 9538 406350
rect 9606 406294 9662 406350
rect 9234 406170 9290 406226
rect 9358 406170 9414 406226
rect 9482 406170 9538 406226
rect 9606 406170 9662 406226
rect 9234 406046 9290 406102
rect 9358 406046 9414 406102
rect 9482 406046 9538 406102
rect 9606 406046 9662 406102
rect 9234 405922 9290 405978
rect 9358 405922 9414 405978
rect 9482 405922 9538 405978
rect 9606 405922 9662 405978
rect 9234 388294 9290 388350
rect 9358 388294 9414 388350
rect 9482 388294 9538 388350
rect 9606 388294 9662 388350
rect 9234 388170 9290 388226
rect 9358 388170 9414 388226
rect 9482 388170 9538 388226
rect 9606 388170 9662 388226
rect 9234 388046 9290 388102
rect 9358 388046 9414 388102
rect 9482 388046 9538 388102
rect 9606 388046 9662 388102
rect 9234 387922 9290 387978
rect 9358 387922 9414 387978
rect 9482 387922 9538 387978
rect 9606 387922 9662 387978
rect 9234 370294 9290 370350
rect 9358 370294 9414 370350
rect 9482 370294 9538 370350
rect 9606 370294 9662 370350
rect 9234 370170 9290 370226
rect 9358 370170 9414 370226
rect 9482 370170 9538 370226
rect 9606 370170 9662 370226
rect 9234 370046 9290 370102
rect 9358 370046 9414 370102
rect 9482 370046 9538 370102
rect 9606 370046 9662 370102
rect 9234 369922 9290 369978
rect 9358 369922 9414 369978
rect 9482 369922 9538 369978
rect 9606 369922 9662 369978
rect 9234 352294 9290 352350
rect 9358 352294 9414 352350
rect 9482 352294 9538 352350
rect 9606 352294 9662 352350
rect 9234 352170 9290 352226
rect 9358 352170 9414 352226
rect 9482 352170 9538 352226
rect 9606 352170 9662 352226
rect 9234 352046 9290 352102
rect 9358 352046 9414 352102
rect 9482 352046 9538 352102
rect 9606 352046 9662 352102
rect 9234 351922 9290 351978
rect 9358 351922 9414 351978
rect 9482 351922 9538 351978
rect 9606 351922 9662 351978
rect 5514 328294 5570 328350
rect 5638 328294 5694 328350
rect 5762 328294 5818 328350
rect 5886 328294 5942 328350
rect 5514 328170 5570 328226
rect 5638 328170 5694 328226
rect 5762 328170 5818 328226
rect 5886 328170 5942 328226
rect 5514 328046 5570 328102
rect 5638 328046 5694 328102
rect 5762 328046 5818 328102
rect 5886 328046 5942 328102
rect 5514 327922 5570 327978
rect 5638 327922 5694 327978
rect 5762 327922 5818 327978
rect 5886 327922 5942 327978
rect 5292 324962 5348 325018
rect 5514 310294 5570 310350
rect 5638 310294 5694 310350
rect 5762 310294 5818 310350
rect 5886 310294 5942 310350
rect 5514 310170 5570 310226
rect 5638 310170 5694 310226
rect 5762 310170 5818 310226
rect 5886 310170 5942 310226
rect 5514 310046 5570 310102
rect 5638 310046 5694 310102
rect 5762 310046 5818 310102
rect 5886 310046 5942 310102
rect 5514 309922 5570 309978
rect 5638 309922 5694 309978
rect 5762 309922 5818 309978
rect 5886 309922 5942 309978
rect 5292 308942 5348 308998
rect 9234 334294 9290 334350
rect 9358 334294 9414 334350
rect 9482 334294 9538 334350
rect 9606 334294 9662 334350
rect 9234 334170 9290 334226
rect 9358 334170 9414 334226
rect 9482 334170 9538 334226
rect 9606 334170 9662 334226
rect 9234 334046 9290 334102
rect 9358 334046 9414 334102
rect 9482 334046 9538 334102
rect 9606 334046 9662 334102
rect 9234 333922 9290 333978
rect 9358 333922 9414 333978
rect 9482 333922 9538 333978
rect 9606 333922 9662 333978
rect 36234 597156 36290 597212
rect 36358 597156 36414 597212
rect 36482 597156 36538 597212
rect 36606 597156 36662 597212
rect 36234 597032 36290 597088
rect 36358 597032 36414 597088
rect 36482 597032 36538 597088
rect 36606 597032 36662 597088
rect 36234 596908 36290 596964
rect 36358 596908 36414 596964
rect 36482 596908 36538 596964
rect 36606 596908 36662 596964
rect 36234 596784 36290 596840
rect 36358 596784 36414 596840
rect 36482 596784 36538 596840
rect 36606 596784 36662 596840
rect 36234 580294 36290 580350
rect 36358 580294 36414 580350
rect 36482 580294 36538 580350
rect 36606 580294 36662 580350
rect 36234 580170 36290 580226
rect 36358 580170 36414 580226
rect 36482 580170 36538 580226
rect 36606 580170 36662 580226
rect 36234 580046 36290 580102
rect 36358 580046 36414 580102
rect 36482 580046 36538 580102
rect 36606 580046 36662 580102
rect 36234 579922 36290 579978
rect 36358 579922 36414 579978
rect 36482 579922 36538 579978
rect 36606 579922 36662 579978
rect 36234 562294 36290 562350
rect 36358 562294 36414 562350
rect 36482 562294 36538 562350
rect 36606 562294 36662 562350
rect 36234 562170 36290 562226
rect 36358 562170 36414 562226
rect 36482 562170 36538 562226
rect 36606 562170 36662 562226
rect 36234 562046 36290 562102
rect 36358 562046 36414 562102
rect 36482 562046 36538 562102
rect 36606 562046 36662 562102
rect 36234 561922 36290 561978
rect 36358 561922 36414 561978
rect 36482 561922 36538 561978
rect 36606 561922 36662 561978
rect 36234 544294 36290 544350
rect 36358 544294 36414 544350
rect 36482 544294 36538 544350
rect 36606 544294 36662 544350
rect 36234 544170 36290 544226
rect 36358 544170 36414 544226
rect 36482 544170 36538 544226
rect 36606 544170 36662 544226
rect 36234 544046 36290 544102
rect 36358 544046 36414 544102
rect 36482 544046 36538 544102
rect 36606 544046 36662 544102
rect 36234 543922 36290 543978
rect 36358 543922 36414 543978
rect 36482 543922 36538 543978
rect 36606 543922 36662 543978
rect 36234 526294 36290 526350
rect 36358 526294 36414 526350
rect 36482 526294 36538 526350
rect 36606 526294 36662 526350
rect 36234 526170 36290 526226
rect 36358 526170 36414 526226
rect 36482 526170 36538 526226
rect 36606 526170 36662 526226
rect 36234 526046 36290 526102
rect 36358 526046 36414 526102
rect 36482 526046 36538 526102
rect 36606 526046 36662 526102
rect 36234 525922 36290 525978
rect 36358 525922 36414 525978
rect 36482 525922 36538 525978
rect 36606 525922 36662 525978
rect 36234 508294 36290 508350
rect 36358 508294 36414 508350
rect 36482 508294 36538 508350
rect 36606 508294 36662 508350
rect 36234 508170 36290 508226
rect 36358 508170 36414 508226
rect 36482 508170 36538 508226
rect 36606 508170 36662 508226
rect 36234 508046 36290 508102
rect 36358 508046 36414 508102
rect 36482 508046 36538 508102
rect 36606 508046 36662 508102
rect 36234 507922 36290 507978
rect 36358 507922 36414 507978
rect 36482 507922 36538 507978
rect 36606 507922 36662 507978
rect 36234 490294 36290 490350
rect 36358 490294 36414 490350
rect 36482 490294 36538 490350
rect 36606 490294 36662 490350
rect 36234 490170 36290 490226
rect 36358 490170 36414 490226
rect 36482 490170 36538 490226
rect 36606 490170 36662 490226
rect 36234 490046 36290 490102
rect 36358 490046 36414 490102
rect 36482 490046 36538 490102
rect 36606 490046 36662 490102
rect 36234 489922 36290 489978
rect 36358 489922 36414 489978
rect 36482 489922 36538 489978
rect 36606 489922 36662 489978
rect 36234 472294 36290 472350
rect 36358 472294 36414 472350
rect 36482 472294 36538 472350
rect 36606 472294 36662 472350
rect 36234 472170 36290 472226
rect 36358 472170 36414 472226
rect 36482 472170 36538 472226
rect 36606 472170 36662 472226
rect 36234 472046 36290 472102
rect 36358 472046 36414 472102
rect 36482 472046 36538 472102
rect 36606 472046 36662 472102
rect 36234 471922 36290 471978
rect 36358 471922 36414 471978
rect 36482 471922 36538 471978
rect 36606 471922 36662 471978
rect 36234 454294 36290 454350
rect 36358 454294 36414 454350
rect 36482 454294 36538 454350
rect 36606 454294 36662 454350
rect 36234 454170 36290 454226
rect 36358 454170 36414 454226
rect 36482 454170 36538 454226
rect 36606 454170 36662 454226
rect 36234 454046 36290 454102
rect 36358 454046 36414 454102
rect 36482 454046 36538 454102
rect 36606 454046 36662 454102
rect 36234 453922 36290 453978
rect 36358 453922 36414 453978
rect 36482 453922 36538 453978
rect 36606 453922 36662 453978
rect 36234 436294 36290 436350
rect 36358 436294 36414 436350
rect 36482 436294 36538 436350
rect 36606 436294 36662 436350
rect 36234 436170 36290 436226
rect 36358 436170 36414 436226
rect 36482 436170 36538 436226
rect 36606 436170 36662 436226
rect 36234 436046 36290 436102
rect 36358 436046 36414 436102
rect 36482 436046 36538 436102
rect 36606 436046 36662 436102
rect 36234 435922 36290 435978
rect 36358 435922 36414 435978
rect 36482 435922 36538 435978
rect 36606 435922 36662 435978
rect 36234 418294 36290 418350
rect 36358 418294 36414 418350
rect 36482 418294 36538 418350
rect 36606 418294 36662 418350
rect 36234 418170 36290 418226
rect 36358 418170 36414 418226
rect 36482 418170 36538 418226
rect 36606 418170 36662 418226
rect 36234 418046 36290 418102
rect 36358 418046 36414 418102
rect 36482 418046 36538 418102
rect 36606 418046 36662 418102
rect 36234 417922 36290 417978
rect 36358 417922 36414 417978
rect 36482 417922 36538 417978
rect 36606 417922 36662 417978
rect 36234 400294 36290 400350
rect 36358 400294 36414 400350
rect 36482 400294 36538 400350
rect 36606 400294 36662 400350
rect 36234 400170 36290 400226
rect 36358 400170 36414 400226
rect 36482 400170 36538 400226
rect 36606 400170 36662 400226
rect 36234 400046 36290 400102
rect 36358 400046 36414 400102
rect 36482 400046 36538 400102
rect 36606 400046 36662 400102
rect 36234 399922 36290 399978
rect 36358 399922 36414 399978
rect 36482 399922 36538 399978
rect 36606 399922 36662 399978
rect 36234 382294 36290 382350
rect 36358 382294 36414 382350
rect 36482 382294 36538 382350
rect 36606 382294 36662 382350
rect 36234 382170 36290 382226
rect 36358 382170 36414 382226
rect 36482 382170 36538 382226
rect 36606 382170 36662 382226
rect 36234 382046 36290 382102
rect 36358 382046 36414 382102
rect 36482 382046 36538 382102
rect 36606 382046 36662 382102
rect 36234 381922 36290 381978
rect 36358 381922 36414 381978
rect 36482 381922 36538 381978
rect 36606 381922 36662 381978
rect 36234 364294 36290 364350
rect 36358 364294 36414 364350
rect 36482 364294 36538 364350
rect 36606 364294 36662 364350
rect 36234 364170 36290 364226
rect 36358 364170 36414 364226
rect 36482 364170 36538 364226
rect 36606 364170 36662 364226
rect 36234 364046 36290 364102
rect 36358 364046 36414 364102
rect 36482 364046 36538 364102
rect 36606 364046 36662 364102
rect 36234 363922 36290 363978
rect 36358 363922 36414 363978
rect 36482 363922 36538 363978
rect 36606 363922 36662 363978
rect 36234 346294 36290 346350
rect 36358 346294 36414 346350
rect 36482 346294 36538 346350
rect 36606 346294 36662 346350
rect 36234 346170 36290 346226
rect 36358 346170 36414 346226
rect 36482 346170 36538 346226
rect 36606 346170 36662 346226
rect 36234 346046 36290 346102
rect 36358 346046 36414 346102
rect 36482 346046 36538 346102
rect 36606 346046 36662 346102
rect 36234 345922 36290 345978
rect 36358 345922 36414 345978
rect 36482 345922 36538 345978
rect 36606 345922 36662 345978
rect 39954 598116 40010 598172
rect 40078 598116 40134 598172
rect 40202 598116 40258 598172
rect 40326 598116 40382 598172
rect 39954 597992 40010 598048
rect 40078 597992 40134 598048
rect 40202 597992 40258 598048
rect 40326 597992 40382 598048
rect 39954 597868 40010 597924
rect 40078 597868 40134 597924
rect 40202 597868 40258 597924
rect 40326 597868 40382 597924
rect 39954 597744 40010 597800
rect 40078 597744 40134 597800
rect 40202 597744 40258 597800
rect 40326 597744 40382 597800
rect 66954 597156 67010 597212
rect 67078 597156 67134 597212
rect 67202 597156 67258 597212
rect 67326 597156 67382 597212
rect 66954 597032 67010 597088
rect 67078 597032 67134 597088
rect 67202 597032 67258 597088
rect 67326 597032 67382 597088
rect 66954 596908 67010 596964
rect 67078 596908 67134 596964
rect 67202 596908 67258 596964
rect 67326 596908 67382 596964
rect 66954 596784 67010 596840
rect 67078 596784 67134 596840
rect 67202 596784 67258 596840
rect 67326 596784 67382 596840
rect 39954 586294 40010 586350
rect 40078 586294 40134 586350
rect 40202 586294 40258 586350
rect 40326 586294 40382 586350
rect 39954 586170 40010 586226
rect 40078 586170 40134 586226
rect 40202 586170 40258 586226
rect 40326 586170 40382 586226
rect 39954 586046 40010 586102
rect 40078 586046 40134 586102
rect 40202 586046 40258 586102
rect 40326 586046 40382 586102
rect 39954 585922 40010 585978
rect 40078 585922 40134 585978
rect 40202 585922 40258 585978
rect 40326 585922 40382 585978
rect 39954 568294 40010 568350
rect 40078 568294 40134 568350
rect 40202 568294 40258 568350
rect 40326 568294 40382 568350
rect 39954 568170 40010 568226
rect 40078 568170 40134 568226
rect 40202 568170 40258 568226
rect 40326 568170 40382 568226
rect 39954 568046 40010 568102
rect 40078 568046 40134 568102
rect 40202 568046 40258 568102
rect 40326 568046 40382 568102
rect 39954 567922 40010 567978
rect 40078 567922 40134 567978
rect 40202 567922 40258 567978
rect 40326 567922 40382 567978
rect 39954 550294 40010 550350
rect 40078 550294 40134 550350
rect 40202 550294 40258 550350
rect 40326 550294 40382 550350
rect 39954 550170 40010 550226
rect 40078 550170 40134 550226
rect 40202 550170 40258 550226
rect 40326 550170 40382 550226
rect 39954 550046 40010 550102
rect 40078 550046 40134 550102
rect 40202 550046 40258 550102
rect 40326 550046 40382 550102
rect 39954 549922 40010 549978
rect 40078 549922 40134 549978
rect 40202 549922 40258 549978
rect 40326 549922 40382 549978
rect 39954 532294 40010 532350
rect 40078 532294 40134 532350
rect 40202 532294 40258 532350
rect 40326 532294 40382 532350
rect 39954 532170 40010 532226
rect 40078 532170 40134 532226
rect 40202 532170 40258 532226
rect 40326 532170 40382 532226
rect 39954 532046 40010 532102
rect 40078 532046 40134 532102
rect 40202 532046 40258 532102
rect 40326 532046 40382 532102
rect 39954 531922 40010 531978
rect 40078 531922 40134 531978
rect 40202 531922 40258 531978
rect 40326 531922 40382 531978
rect 39954 514294 40010 514350
rect 40078 514294 40134 514350
rect 40202 514294 40258 514350
rect 40326 514294 40382 514350
rect 39954 514170 40010 514226
rect 40078 514170 40134 514226
rect 40202 514170 40258 514226
rect 40326 514170 40382 514226
rect 39954 514046 40010 514102
rect 40078 514046 40134 514102
rect 40202 514046 40258 514102
rect 40326 514046 40382 514102
rect 39954 513922 40010 513978
rect 40078 513922 40134 513978
rect 40202 513922 40258 513978
rect 40326 513922 40382 513978
rect 39954 496294 40010 496350
rect 40078 496294 40134 496350
rect 40202 496294 40258 496350
rect 40326 496294 40382 496350
rect 39954 496170 40010 496226
rect 40078 496170 40134 496226
rect 40202 496170 40258 496226
rect 40326 496170 40382 496226
rect 39954 496046 40010 496102
rect 40078 496046 40134 496102
rect 40202 496046 40258 496102
rect 40326 496046 40382 496102
rect 39954 495922 40010 495978
rect 40078 495922 40134 495978
rect 40202 495922 40258 495978
rect 40326 495922 40382 495978
rect 39954 478294 40010 478350
rect 40078 478294 40134 478350
rect 40202 478294 40258 478350
rect 40326 478294 40382 478350
rect 39954 478170 40010 478226
rect 40078 478170 40134 478226
rect 40202 478170 40258 478226
rect 40326 478170 40382 478226
rect 39954 478046 40010 478102
rect 40078 478046 40134 478102
rect 40202 478046 40258 478102
rect 40326 478046 40382 478102
rect 39954 477922 40010 477978
rect 40078 477922 40134 477978
rect 40202 477922 40258 477978
rect 40326 477922 40382 477978
rect 39954 460294 40010 460350
rect 40078 460294 40134 460350
rect 40202 460294 40258 460350
rect 40326 460294 40382 460350
rect 39954 460170 40010 460226
rect 40078 460170 40134 460226
rect 40202 460170 40258 460226
rect 40326 460170 40382 460226
rect 39954 460046 40010 460102
rect 40078 460046 40134 460102
rect 40202 460046 40258 460102
rect 40326 460046 40382 460102
rect 39954 459922 40010 459978
rect 40078 459922 40134 459978
rect 40202 459922 40258 459978
rect 40326 459922 40382 459978
rect 39954 442294 40010 442350
rect 40078 442294 40134 442350
rect 40202 442294 40258 442350
rect 40326 442294 40382 442350
rect 39954 442170 40010 442226
rect 40078 442170 40134 442226
rect 40202 442170 40258 442226
rect 40326 442170 40382 442226
rect 39954 442046 40010 442102
rect 40078 442046 40134 442102
rect 40202 442046 40258 442102
rect 40326 442046 40382 442102
rect 39954 441922 40010 441978
rect 40078 441922 40134 441978
rect 40202 441922 40258 441978
rect 40326 441922 40382 441978
rect 39954 424294 40010 424350
rect 40078 424294 40134 424350
rect 40202 424294 40258 424350
rect 40326 424294 40382 424350
rect 39954 424170 40010 424226
rect 40078 424170 40134 424226
rect 40202 424170 40258 424226
rect 40326 424170 40382 424226
rect 39954 424046 40010 424102
rect 40078 424046 40134 424102
rect 40202 424046 40258 424102
rect 40326 424046 40382 424102
rect 39954 423922 40010 423978
rect 40078 423922 40134 423978
rect 40202 423922 40258 423978
rect 40326 423922 40382 423978
rect 39954 406294 40010 406350
rect 40078 406294 40134 406350
rect 40202 406294 40258 406350
rect 40326 406294 40382 406350
rect 39954 406170 40010 406226
rect 40078 406170 40134 406226
rect 40202 406170 40258 406226
rect 40326 406170 40382 406226
rect 39954 406046 40010 406102
rect 40078 406046 40134 406102
rect 40202 406046 40258 406102
rect 40326 406046 40382 406102
rect 39954 405922 40010 405978
rect 40078 405922 40134 405978
rect 40202 405922 40258 405978
rect 40326 405922 40382 405978
rect 39954 388294 40010 388350
rect 40078 388294 40134 388350
rect 40202 388294 40258 388350
rect 40326 388294 40382 388350
rect 39954 388170 40010 388226
rect 40078 388170 40134 388226
rect 40202 388170 40258 388226
rect 40326 388170 40382 388226
rect 39954 388046 40010 388102
rect 40078 388046 40134 388102
rect 40202 388046 40258 388102
rect 40326 388046 40382 388102
rect 39954 387922 40010 387978
rect 40078 387922 40134 387978
rect 40202 387922 40258 387978
rect 40326 387922 40382 387978
rect 39954 370294 40010 370350
rect 40078 370294 40134 370350
rect 40202 370294 40258 370350
rect 40326 370294 40382 370350
rect 39954 370170 40010 370226
rect 40078 370170 40134 370226
rect 40202 370170 40258 370226
rect 40326 370170 40382 370226
rect 39954 370046 40010 370102
rect 40078 370046 40134 370102
rect 40202 370046 40258 370102
rect 40326 370046 40382 370102
rect 39954 369922 40010 369978
rect 40078 369922 40134 369978
rect 40202 369922 40258 369978
rect 40326 369922 40382 369978
rect 39954 352294 40010 352350
rect 40078 352294 40134 352350
rect 40202 352294 40258 352350
rect 40326 352294 40382 352350
rect 39954 352170 40010 352226
rect 40078 352170 40134 352226
rect 40202 352170 40258 352226
rect 40326 352170 40382 352226
rect 39954 352046 40010 352102
rect 40078 352046 40134 352102
rect 40202 352046 40258 352102
rect 40326 352046 40382 352102
rect 39954 351922 40010 351978
rect 40078 351922 40134 351978
rect 40202 351922 40258 351978
rect 40326 351922 40382 351978
rect 39954 334294 40010 334350
rect 40078 334294 40134 334350
rect 40202 334294 40258 334350
rect 40326 334294 40382 334350
rect 39954 334170 40010 334226
rect 40078 334170 40134 334226
rect 40202 334170 40258 334226
rect 40326 334170 40382 334226
rect 39954 334046 40010 334102
rect 40078 334046 40134 334102
rect 40202 334046 40258 334102
rect 40326 334046 40382 334102
rect 39954 333922 40010 333978
rect 40078 333922 40134 333978
rect 40202 333922 40258 333978
rect 40326 333922 40382 333978
rect 36234 328294 36290 328350
rect 36358 328294 36414 328350
rect 36482 328294 36538 328350
rect 36606 328294 36662 328350
rect 36234 328170 36290 328226
rect 36358 328170 36414 328226
rect 36482 328170 36538 328226
rect 36606 328170 36662 328226
rect 36234 328046 36290 328102
rect 36358 328046 36414 328102
rect 36482 328046 36538 328102
rect 36606 328046 36662 328102
rect 36234 327922 36290 327978
rect 36358 327922 36414 327978
rect 36482 327922 36538 327978
rect 36606 327922 36662 327978
rect 24878 316294 24934 316350
rect 25002 316294 25058 316350
rect 24878 316170 24934 316226
rect 25002 316170 25058 316226
rect 24878 316046 24934 316102
rect 25002 316046 25058 316102
rect 24878 315922 24934 315978
rect 25002 315922 25058 315978
rect 9518 310294 9574 310350
rect 9642 310294 9698 310350
rect 9518 310170 9574 310226
rect 9642 310170 9698 310226
rect 9518 310046 9574 310102
rect 9642 310046 9698 310102
rect 9518 309922 9574 309978
rect 9642 309922 9698 309978
rect 40238 310294 40294 310350
rect 40362 310294 40418 310350
rect 40238 310170 40294 310226
rect 40362 310170 40418 310226
rect 40238 310046 40294 310102
rect 40362 310046 40418 310102
rect 40238 309922 40294 309978
rect 40362 309922 40418 309978
rect 7532 308942 7588 308998
rect 24878 298294 24934 298350
rect 25002 298294 25058 298350
rect 24878 298170 24934 298226
rect 25002 298170 25058 298226
rect 24878 298046 24934 298102
rect 25002 298046 25058 298102
rect 24878 297922 24934 297978
rect 25002 297922 25058 297978
rect 5514 292294 5570 292350
rect 5638 292294 5694 292350
rect 5762 292294 5818 292350
rect 5886 292294 5942 292350
rect 5514 292170 5570 292226
rect 5638 292170 5694 292226
rect 5762 292170 5818 292226
rect 5886 292170 5942 292226
rect 5514 292046 5570 292102
rect 5638 292046 5694 292102
rect 5762 292046 5818 292102
rect 5886 292046 5942 292102
rect 5514 291922 5570 291978
rect 5638 291922 5694 291978
rect 5762 291922 5818 291978
rect 5886 291922 5942 291978
rect 5292 281762 5348 281818
rect 5292 281402 5348 281458
rect 4956 277982 5012 278038
rect 4396 270422 4452 270478
rect 9518 292294 9574 292350
rect 9642 292294 9698 292350
rect 9518 292170 9574 292226
rect 9642 292170 9698 292226
rect 9518 292046 9574 292102
rect 9642 292046 9698 292102
rect 9518 291922 9574 291978
rect 9642 291922 9698 291978
rect 40238 292294 40294 292350
rect 40362 292294 40418 292350
rect 40238 292170 40294 292226
rect 40362 292170 40418 292226
rect 40238 292046 40294 292102
rect 40362 292046 40418 292102
rect 40238 291922 40294 291978
rect 40362 291922 40418 291978
rect 7644 290762 7700 290818
rect 7084 275462 7140 275518
rect 5514 274294 5570 274350
rect 5638 274294 5694 274350
rect 5762 274294 5818 274350
rect 5886 274294 5942 274350
rect 5514 274170 5570 274226
rect 5638 274170 5694 274226
rect 5762 274170 5818 274226
rect 5886 274170 5942 274226
rect 5514 274046 5570 274102
rect 5638 274046 5694 274102
rect 5762 274046 5818 274102
rect 5886 274046 5942 274102
rect 5514 273922 5570 273978
rect 5638 273922 5694 273978
rect 5762 273922 5818 273978
rect 5886 273922 5942 273978
rect 4172 270242 4228 270298
rect 4284 268262 4340 268318
rect 4172 266642 4228 266698
rect 4172 206522 4228 206578
rect 4956 257822 5012 257878
rect 9234 280294 9290 280350
rect 9358 280294 9414 280350
rect 9482 280294 9538 280350
rect 9606 280294 9662 280350
rect 9234 280170 9290 280226
rect 9358 280170 9414 280226
rect 9482 280170 9538 280226
rect 9606 280170 9662 280226
rect 9234 280046 9290 280102
rect 9358 280046 9414 280102
rect 9482 280046 9538 280102
rect 9606 280046 9662 280102
rect 9234 279922 9290 279978
rect 9358 279922 9414 279978
rect 9482 279922 9538 279978
rect 9606 279922 9662 279978
rect 7756 277262 7812 277318
rect 5514 256294 5570 256350
rect 5638 256294 5694 256350
rect 5762 256294 5818 256350
rect 5886 256294 5942 256350
rect 5514 256170 5570 256226
rect 5638 256170 5694 256226
rect 5762 256170 5818 256226
rect 5886 256170 5942 256226
rect 5514 256046 5570 256102
rect 5638 256046 5694 256102
rect 5762 256046 5818 256102
rect 5886 256046 5942 256102
rect 5514 255922 5570 255978
rect 5638 255922 5694 255978
rect 5762 255922 5818 255978
rect 5886 255922 5942 255978
rect 5514 238294 5570 238350
rect 5638 238294 5694 238350
rect 5762 238294 5818 238350
rect 5886 238294 5942 238350
rect 5514 238170 5570 238226
rect 5638 238170 5694 238226
rect 5762 238170 5818 238226
rect 5886 238170 5942 238226
rect 5514 238046 5570 238102
rect 5638 238046 5694 238102
rect 5762 238046 5818 238102
rect 5886 238046 5942 238102
rect 5514 237922 5570 237978
rect 5638 237922 5694 237978
rect 5762 237922 5818 237978
rect 5886 237922 5942 237978
rect 5514 220294 5570 220350
rect 5638 220294 5694 220350
rect 5762 220294 5818 220350
rect 5886 220294 5942 220350
rect 5514 220170 5570 220226
rect 5638 220170 5694 220226
rect 5762 220170 5818 220226
rect 5886 220170 5942 220226
rect 5514 220046 5570 220102
rect 5638 220046 5694 220102
rect 5762 220046 5818 220102
rect 5886 220046 5942 220102
rect 5514 219922 5570 219978
rect 5638 219922 5694 219978
rect 5762 219922 5818 219978
rect 5886 219922 5942 219978
rect 5514 202294 5570 202350
rect 5638 202294 5694 202350
rect 5762 202294 5818 202350
rect 5886 202294 5942 202350
rect 5514 202170 5570 202226
rect 5638 202170 5694 202226
rect 5762 202170 5818 202226
rect 5886 202170 5942 202226
rect 5514 202046 5570 202102
rect 5638 202046 5694 202102
rect 5762 202046 5818 202102
rect 5886 202046 5942 202102
rect 5514 201922 5570 201978
rect 5638 201922 5694 201978
rect 5762 201922 5818 201978
rect 5886 201922 5942 201978
rect 5514 184294 5570 184350
rect 5638 184294 5694 184350
rect 5762 184294 5818 184350
rect 5886 184294 5942 184350
rect 5514 184170 5570 184226
rect 5638 184170 5694 184226
rect 5762 184170 5818 184226
rect 5886 184170 5942 184226
rect 5514 184046 5570 184102
rect 5638 184046 5694 184102
rect 5762 184046 5818 184102
rect 5886 184046 5942 184102
rect 5514 183922 5570 183978
rect 5638 183922 5694 183978
rect 5762 183922 5818 183978
rect 5886 183922 5942 183978
rect 5514 166294 5570 166350
rect 5638 166294 5694 166350
rect 5762 166294 5818 166350
rect 5886 166294 5942 166350
rect 5514 166170 5570 166226
rect 5638 166170 5694 166226
rect 5762 166170 5818 166226
rect 5886 166170 5942 166226
rect 5514 166046 5570 166102
rect 5638 166046 5694 166102
rect 5762 166046 5818 166102
rect 5886 166046 5942 166102
rect 5514 165922 5570 165978
rect 5638 165922 5694 165978
rect 5762 165922 5818 165978
rect 5886 165922 5942 165978
rect 5514 148294 5570 148350
rect 5638 148294 5694 148350
rect 5762 148294 5818 148350
rect 5886 148294 5942 148350
rect 5514 148170 5570 148226
rect 5638 148170 5694 148226
rect 5762 148170 5818 148226
rect 5886 148170 5942 148226
rect 5514 148046 5570 148102
rect 5638 148046 5694 148102
rect 5762 148046 5818 148102
rect 5886 148046 5942 148102
rect 5514 147922 5570 147978
rect 5638 147922 5694 147978
rect 5762 147922 5818 147978
rect 5886 147922 5942 147978
rect 5514 130294 5570 130350
rect 5638 130294 5694 130350
rect 5762 130294 5818 130350
rect 5886 130294 5942 130350
rect 5514 130170 5570 130226
rect 5638 130170 5694 130226
rect 5762 130170 5818 130226
rect 5886 130170 5942 130226
rect 5514 130046 5570 130102
rect 5638 130046 5694 130102
rect 5762 130046 5818 130102
rect 5886 130046 5942 130102
rect 5514 129922 5570 129978
rect 5638 129922 5694 129978
rect 5762 129922 5818 129978
rect 5886 129922 5942 129978
rect 5514 112294 5570 112350
rect 5638 112294 5694 112350
rect 5762 112294 5818 112350
rect 5886 112294 5942 112350
rect 5514 112170 5570 112226
rect 5638 112170 5694 112226
rect 5762 112170 5818 112226
rect 5886 112170 5942 112226
rect 5514 112046 5570 112102
rect 5638 112046 5694 112102
rect 5762 112046 5818 112102
rect 5886 112046 5942 112102
rect 5514 111922 5570 111978
rect 5638 111922 5694 111978
rect 5762 111922 5818 111978
rect 5886 111922 5942 111978
rect 7532 266282 7588 266338
rect 7644 264662 7700 264718
rect 9234 262294 9290 262350
rect 9358 262294 9414 262350
rect 9482 262294 9538 262350
rect 9606 262294 9662 262350
rect 9234 262170 9290 262226
rect 9358 262170 9414 262226
rect 9482 262170 9538 262226
rect 9606 262170 9662 262226
rect 9234 262046 9290 262102
rect 9358 262046 9414 262102
rect 9482 262046 9538 262102
rect 9606 262046 9662 262102
rect 9234 261922 9290 261978
rect 9358 261922 9414 261978
rect 9482 261922 9538 261978
rect 9606 261922 9662 261978
rect 9234 244294 9290 244350
rect 9358 244294 9414 244350
rect 9482 244294 9538 244350
rect 9606 244294 9662 244350
rect 9234 244170 9290 244226
rect 9358 244170 9414 244226
rect 9482 244170 9538 244226
rect 9606 244170 9662 244226
rect 9234 244046 9290 244102
rect 9358 244046 9414 244102
rect 9482 244046 9538 244102
rect 9606 244046 9662 244102
rect 9234 243922 9290 243978
rect 9358 243922 9414 243978
rect 9482 243922 9538 243978
rect 9606 243922 9662 243978
rect 9234 226294 9290 226350
rect 9358 226294 9414 226350
rect 9482 226294 9538 226350
rect 9606 226294 9662 226350
rect 9234 226170 9290 226226
rect 9358 226170 9414 226226
rect 9482 226170 9538 226226
rect 9606 226170 9662 226226
rect 9234 226046 9290 226102
rect 9358 226046 9414 226102
rect 9482 226046 9538 226102
rect 9606 226046 9662 226102
rect 9234 225922 9290 225978
rect 9358 225922 9414 225978
rect 9482 225922 9538 225978
rect 9606 225922 9662 225978
rect 9234 208294 9290 208350
rect 9358 208294 9414 208350
rect 9482 208294 9538 208350
rect 9606 208294 9662 208350
rect 9234 208170 9290 208226
rect 9358 208170 9414 208226
rect 9482 208170 9538 208226
rect 9606 208170 9662 208226
rect 9234 208046 9290 208102
rect 9358 208046 9414 208102
rect 9482 208046 9538 208102
rect 9606 208046 9662 208102
rect 9234 207922 9290 207978
rect 9358 207922 9414 207978
rect 9482 207922 9538 207978
rect 9606 207922 9662 207978
rect 10892 268082 10948 268138
rect 11004 264482 11060 264538
rect 13760 256294 13816 256350
rect 13884 256294 13940 256350
rect 14008 256294 14064 256350
rect 14132 256294 14188 256350
rect 13760 256170 13816 256226
rect 13884 256170 13940 256226
rect 14008 256170 14064 256226
rect 14132 256170 14188 256226
rect 13760 256046 13816 256102
rect 13884 256046 13940 256102
rect 14008 256046 14064 256102
rect 14132 256046 14188 256102
rect 13760 255922 13816 255978
rect 13884 255922 13940 255978
rect 14008 255922 14064 255978
rect 14132 255922 14188 255978
rect 12960 244294 13016 244350
rect 13084 244294 13140 244350
rect 13208 244294 13264 244350
rect 13332 244294 13388 244350
rect 12960 244170 13016 244226
rect 13084 244170 13140 244226
rect 13208 244170 13264 244226
rect 13332 244170 13388 244226
rect 12960 244046 13016 244102
rect 13084 244046 13140 244102
rect 13208 244046 13264 244102
rect 13332 244046 13388 244102
rect 12960 243922 13016 243978
rect 13084 243922 13140 243978
rect 13208 243922 13264 243978
rect 13332 243922 13388 243978
rect 13760 238294 13816 238350
rect 13884 238294 13940 238350
rect 14008 238294 14064 238350
rect 14132 238294 14188 238350
rect 13760 238170 13816 238226
rect 13884 238170 13940 238226
rect 14008 238170 14064 238226
rect 14132 238170 14188 238226
rect 13760 238046 13816 238102
rect 13884 238046 13940 238102
rect 14008 238046 14064 238102
rect 14132 238046 14188 238102
rect 13760 237922 13816 237978
rect 13884 237922 13940 237978
rect 14008 237922 14064 237978
rect 14132 237922 14188 237978
rect 12960 226294 13016 226350
rect 13084 226294 13140 226350
rect 13208 226294 13264 226350
rect 13332 226294 13388 226350
rect 12960 226170 13016 226226
rect 13084 226170 13140 226226
rect 13208 226170 13264 226226
rect 13332 226170 13388 226226
rect 12960 226046 13016 226102
rect 13084 226046 13140 226102
rect 13208 226046 13264 226102
rect 13332 226046 13388 226102
rect 12960 225922 13016 225978
rect 13084 225922 13140 225978
rect 13208 225922 13264 225978
rect 13332 225922 13388 225978
rect 13760 220294 13816 220350
rect 13884 220294 13940 220350
rect 14008 220294 14064 220350
rect 14132 220294 14188 220350
rect 13760 220170 13816 220226
rect 13884 220170 13940 220226
rect 14008 220170 14064 220226
rect 14132 220170 14188 220226
rect 13760 220046 13816 220102
rect 13884 220046 13940 220102
rect 14008 220046 14064 220102
rect 14132 220046 14188 220102
rect 13760 219922 13816 219978
rect 13884 219922 13940 219978
rect 14008 219922 14064 219978
rect 14132 219922 14188 219978
rect 12960 208294 13016 208350
rect 13084 208294 13140 208350
rect 13208 208294 13264 208350
rect 13332 208294 13388 208350
rect 12960 208170 13016 208226
rect 13084 208170 13140 208226
rect 13208 208170 13264 208226
rect 13332 208170 13388 208226
rect 12960 208046 13016 208102
rect 13084 208046 13140 208102
rect 13208 208046 13264 208102
rect 13332 208046 13388 208102
rect 12960 207922 13016 207978
rect 13084 207922 13140 207978
rect 13208 207922 13264 207978
rect 13332 207922 13388 207978
rect 13760 202294 13816 202350
rect 13884 202294 13940 202350
rect 14008 202294 14064 202350
rect 14132 202294 14188 202350
rect 13760 202170 13816 202226
rect 13884 202170 13940 202226
rect 14008 202170 14064 202226
rect 14132 202170 14188 202226
rect 13760 202046 13816 202102
rect 13884 202046 13940 202102
rect 14008 202046 14064 202102
rect 14132 202046 14188 202102
rect 13760 201922 13816 201978
rect 13884 201922 13940 201978
rect 14008 201922 14064 201978
rect 14132 201922 14188 201978
rect 9234 190294 9290 190350
rect 9358 190294 9414 190350
rect 9482 190294 9538 190350
rect 9606 190294 9662 190350
rect 9234 190170 9290 190226
rect 9358 190170 9414 190226
rect 9482 190170 9538 190226
rect 9606 190170 9662 190226
rect 9234 190046 9290 190102
rect 9358 190046 9414 190102
rect 9482 190046 9538 190102
rect 9606 190046 9662 190102
rect 9234 189922 9290 189978
rect 9358 189922 9414 189978
rect 9482 189922 9538 189978
rect 9606 189922 9662 189978
rect 12960 190294 13016 190350
rect 13084 190294 13140 190350
rect 13208 190294 13264 190350
rect 13332 190294 13388 190350
rect 12960 190170 13016 190226
rect 13084 190170 13140 190226
rect 13208 190170 13264 190226
rect 13332 190170 13388 190226
rect 12960 190046 13016 190102
rect 13084 190046 13140 190102
rect 13208 190046 13264 190102
rect 13332 190046 13388 190102
rect 12960 189922 13016 189978
rect 13084 189922 13140 189978
rect 13208 189922 13264 189978
rect 13332 189922 13388 189978
rect 13760 184294 13816 184350
rect 13884 184294 13940 184350
rect 14008 184294 14064 184350
rect 14132 184294 14188 184350
rect 13760 184170 13816 184226
rect 13884 184170 13940 184226
rect 14008 184170 14064 184226
rect 14132 184170 14188 184226
rect 13760 184046 13816 184102
rect 13884 184046 13940 184102
rect 14008 184046 14064 184102
rect 14132 184046 14188 184102
rect 13760 183922 13816 183978
rect 13884 183922 13940 183978
rect 14008 183922 14064 183978
rect 14132 183922 14188 183978
rect 9234 172294 9290 172350
rect 9358 172294 9414 172350
rect 9482 172294 9538 172350
rect 9606 172294 9662 172350
rect 9234 172170 9290 172226
rect 9358 172170 9414 172226
rect 9482 172170 9538 172226
rect 9606 172170 9662 172226
rect 9234 172046 9290 172102
rect 9358 172046 9414 172102
rect 9482 172046 9538 172102
rect 9606 172046 9662 172102
rect 9234 171922 9290 171978
rect 9358 171922 9414 171978
rect 9482 171922 9538 171978
rect 9606 171922 9662 171978
rect 12960 172294 13016 172350
rect 13084 172294 13140 172350
rect 13208 172294 13264 172350
rect 13332 172294 13388 172350
rect 12960 172170 13016 172226
rect 13084 172170 13140 172226
rect 13208 172170 13264 172226
rect 13332 172170 13388 172226
rect 12960 172046 13016 172102
rect 13084 172046 13140 172102
rect 13208 172046 13264 172102
rect 13332 172046 13388 172102
rect 12960 171922 13016 171978
rect 13084 171922 13140 171978
rect 13208 171922 13264 171978
rect 13332 171922 13388 171978
rect 21756 185642 21812 185698
rect 20860 162782 20916 162838
rect 39954 280294 40010 280350
rect 40078 280294 40134 280350
rect 40202 280294 40258 280350
rect 40326 280294 40382 280350
rect 39954 280170 40010 280226
rect 40078 280170 40134 280226
rect 40202 280170 40258 280226
rect 40326 280170 40382 280226
rect 39954 280046 40010 280102
rect 40078 280046 40134 280102
rect 40202 280046 40258 280102
rect 40326 280046 40382 280102
rect 39954 279922 40010 279978
rect 40078 279922 40134 279978
rect 40202 279922 40258 279978
rect 40326 279922 40382 279978
rect 36234 274294 36290 274350
rect 36358 274294 36414 274350
rect 36482 274294 36538 274350
rect 36606 274294 36662 274350
rect 36234 274170 36290 274226
rect 36358 274170 36414 274226
rect 36482 274170 36538 274226
rect 36606 274170 36662 274226
rect 36234 274046 36290 274102
rect 36358 274046 36414 274102
rect 36482 274046 36538 274102
rect 36606 274046 36662 274102
rect 36234 273922 36290 273978
rect 36358 273922 36414 273978
rect 36482 273922 36538 273978
rect 36606 273922 36662 273978
rect 26796 187262 26852 187318
rect 28476 191402 28532 191458
rect 36234 256294 36290 256350
rect 36358 256294 36414 256350
rect 36482 256294 36538 256350
rect 36606 256294 36662 256350
rect 36234 256170 36290 256226
rect 36358 256170 36414 256226
rect 36482 256170 36538 256226
rect 36606 256170 36662 256226
rect 36234 256046 36290 256102
rect 36358 256046 36414 256102
rect 36482 256046 36538 256102
rect 36606 256046 36662 256102
rect 36234 255922 36290 255978
rect 36358 255922 36414 255978
rect 36482 255922 36538 255978
rect 36606 255922 36662 255978
rect 36234 238294 36290 238350
rect 36358 238294 36414 238350
rect 36482 238294 36538 238350
rect 36606 238294 36662 238350
rect 36234 238170 36290 238226
rect 36358 238170 36414 238226
rect 36482 238170 36538 238226
rect 36606 238170 36662 238226
rect 36234 238046 36290 238102
rect 36358 238046 36414 238102
rect 36482 238046 36538 238102
rect 36606 238046 36662 238102
rect 36234 237922 36290 237978
rect 36358 237922 36414 237978
rect 36482 237922 36538 237978
rect 36606 237922 36662 237978
rect 36234 220294 36290 220350
rect 36358 220294 36414 220350
rect 36482 220294 36538 220350
rect 36606 220294 36662 220350
rect 36234 220170 36290 220226
rect 36358 220170 36414 220226
rect 36482 220170 36538 220226
rect 36606 220170 36662 220226
rect 36234 220046 36290 220102
rect 36358 220046 36414 220102
rect 36482 220046 36538 220102
rect 36606 220046 36662 220102
rect 36234 219922 36290 219978
rect 36358 219922 36414 219978
rect 36482 219922 36538 219978
rect 36606 219922 36662 219978
rect 36234 202294 36290 202350
rect 36358 202294 36414 202350
rect 36482 202294 36538 202350
rect 36606 202294 36662 202350
rect 36234 202170 36290 202226
rect 36358 202170 36414 202226
rect 36482 202170 36538 202226
rect 36606 202170 36662 202226
rect 36234 202046 36290 202102
rect 36358 202046 36414 202102
rect 36482 202046 36538 202102
rect 36606 202046 36662 202102
rect 36234 201922 36290 201978
rect 36358 201922 36414 201978
rect 36482 201922 36538 201978
rect 36606 201922 36662 201978
rect 36234 184294 36290 184350
rect 36358 184294 36414 184350
rect 36482 184294 36538 184350
rect 36606 184294 36662 184350
rect 36234 184170 36290 184226
rect 36358 184170 36414 184226
rect 36482 184170 36538 184226
rect 36606 184170 36662 184226
rect 36234 184046 36290 184102
rect 36358 184046 36414 184102
rect 36482 184046 36538 184102
rect 36606 184046 36662 184102
rect 36234 183922 36290 183978
rect 36358 183922 36414 183978
rect 36482 183922 36538 183978
rect 36606 183922 36662 183978
rect 36234 166294 36290 166350
rect 36358 166294 36414 166350
rect 36482 166294 36538 166350
rect 36606 166294 36662 166350
rect 36234 166170 36290 166226
rect 36358 166170 36414 166226
rect 36482 166170 36538 166226
rect 36606 166170 36662 166226
rect 36234 166046 36290 166102
rect 36358 166046 36414 166102
rect 36482 166046 36538 166102
rect 36606 166046 36662 166102
rect 36234 165922 36290 165978
rect 36358 165922 36414 165978
rect 36482 165922 36538 165978
rect 36606 165922 36662 165978
rect 27132 162602 27188 162658
rect 9234 154294 9290 154350
rect 9358 154294 9414 154350
rect 9482 154294 9538 154350
rect 9606 154294 9662 154350
rect 9234 154170 9290 154226
rect 9358 154170 9414 154226
rect 9482 154170 9538 154226
rect 9606 154170 9662 154226
rect 9234 154046 9290 154102
rect 9358 154046 9414 154102
rect 9482 154046 9538 154102
rect 9606 154046 9662 154102
rect 9234 153922 9290 153978
rect 9358 153922 9414 153978
rect 9482 153922 9538 153978
rect 9606 153922 9662 153978
rect 39676 193022 39732 193078
rect 45276 277116 45332 277138
rect 45276 277082 45332 277116
rect 48636 276902 48692 276958
rect 48748 276542 48804 276598
rect 39954 262294 40010 262350
rect 40078 262294 40134 262350
rect 40202 262294 40258 262350
rect 40326 262294 40382 262350
rect 39954 262170 40010 262226
rect 40078 262170 40134 262226
rect 40202 262170 40258 262226
rect 40326 262170 40382 262226
rect 39954 262046 40010 262102
rect 40078 262046 40134 262102
rect 40202 262046 40258 262102
rect 40326 262046 40382 262102
rect 39954 261922 40010 261978
rect 40078 261922 40134 261978
rect 40202 261922 40258 261978
rect 40326 261922 40382 261978
rect 39954 244294 40010 244350
rect 40078 244294 40134 244350
rect 40202 244294 40258 244350
rect 40326 244294 40382 244350
rect 39954 244170 40010 244226
rect 40078 244170 40134 244226
rect 40202 244170 40258 244226
rect 40326 244170 40382 244226
rect 39954 244046 40010 244102
rect 40078 244046 40134 244102
rect 40202 244046 40258 244102
rect 40326 244046 40382 244102
rect 39954 243922 40010 243978
rect 40078 243922 40134 243978
rect 40202 243922 40258 243978
rect 40326 243922 40382 243978
rect 39954 226294 40010 226350
rect 40078 226294 40134 226350
rect 40202 226294 40258 226350
rect 40326 226294 40382 226350
rect 39954 226170 40010 226226
rect 40078 226170 40134 226226
rect 40202 226170 40258 226226
rect 40326 226170 40382 226226
rect 39954 226046 40010 226102
rect 40078 226046 40134 226102
rect 40202 226046 40258 226102
rect 40326 226046 40382 226102
rect 39954 225922 40010 225978
rect 40078 225922 40134 225978
rect 40202 225922 40258 225978
rect 40326 225922 40382 225978
rect 39954 208294 40010 208350
rect 40078 208294 40134 208350
rect 40202 208294 40258 208350
rect 40326 208294 40382 208350
rect 39954 208170 40010 208226
rect 40078 208170 40134 208226
rect 40202 208170 40258 208226
rect 40326 208170 40382 208226
rect 39954 208046 40010 208102
rect 40078 208046 40134 208102
rect 40202 208046 40258 208102
rect 40326 208046 40382 208102
rect 39954 207922 40010 207978
rect 40078 207922 40134 207978
rect 40202 207922 40258 207978
rect 40326 207922 40382 207978
rect 39954 190294 40010 190350
rect 40078 190294 40134 190350
rect 40202 190294 40258 190350
rect 40326 190294 40382 190350
rect 39954 190170 40010 190226
rect 40078 190170 40134 190226
rect 40202 190170 40258 190226
rect 40326 190170 40382 190226
rect 39954 190046 40010 190102
rect 40078 190046 40134 190102
rect 40202 190046 40258 190102
rect 40326 190046 40382 190102
rect 39954 189922 40010 189978
rect 40078 189922 40134 189978
rect 40202 189922 40258 189978
rect 40326 189922 40382 189978
rect 39954 172294 40010 172350
rect 40078 172294 40134 172350
rect 40202 172294 40258 172350
rect 40326 172294 40382 172350
rect 39954 172170 40010 172226
rect 40078 172170 40134 172226
rect 40202 172170 40258 172226
rect 40326 172170 40382 172226
rect 39954 172046 40010 172102
rect 40078 172046 40134 172102
rect 40202 172046 40258 172102
rect 40326 172046 40382 172102
rect 39954 171922 40010 171978
rect 40078 171922 40134 171978
rect 40202 171922 40258 171978
rect 40326 171922 40382 171978
rect 36234 148294 36290 148350
rect 36358 148294 36414 148350
rect 36482 148294 36538 148350
rect 36606 148294 36662 148350
rect 36234 148170 36290 148226
rect 36358 148170 36414 148226
rect 36482 148170 36538 148226
rect 36606 148170 36662 148226
rect 36234 148046 36290 148102
rect 36358 148046 36414 148102
rect 36482 148046 36538 148102
rect 36606 148046 36662 148102
rect 36234 147922 36290 147978
rect 36358 147922 36414 147978
rect 36482 147922 36538 147978
rect 36606 147922 36662 147978
rect 9234 136294 9290 136350
rect 9358 136294 9414 136350
rect 9482 136294 9538 136350
rect 9606 136294 9662 136350
rect 9234 136170 9290 136226
rect 9358 136170 9414 136226
rect 9482 136170 9538 136226
rect 9606 136170 9662 136226
rect 9234 136046 9290 136102
rect 9358 136046 9414 136102
rect 9482 136046 9538 136102
rect 9606 136046 9662 136102
rect 9234 135922 9290 135978
rect 9358 135922 9414 135978
rect 9482 135922 9538 135978
rect 9606 135922 9662 135978
rect 11930 136294 11986 136350
rect 12054 136294 12110 136350
rect 12178 136294 12234 136350
rect 12302 136294 12358 136350
rect 11930 136170 11986 136226
rect 12054 136170 12110 136226
rect 12178 136170 12234 136226
rect 12302 136170 12358 136226
rect 11930 136046 11986 136102
rect 12054 136046 12110 136102
rect 12178 136046 12234 136102
rect 12302 136046 12358 136102
rect 11930 135922 11986 135978
rect 12054 135922 12110 135978
rect 12178 135922 12234 135978
rect 12302 135922 12358 135978
rect 11130 130294 11186 130350
rect 11254 130294 11310 130350
rect 11378 130294 11434 130350
rect 11502 130294 11558 130350
rect 11130 130170 11186 130226
rect 11254 130170 11310 130226
rect 11378 130170 11434 130226
rect 11502 130170 11558 130226
rect 11130 130046 11186 130102
rect 11254 130046 11310 130102
rect 11378 130046 11434 130102
rect 11502 130046 11558 130102
rect 11130 129922 11186 129978
rect 11254 129922 11310 129978
rect 11378 129922 11434 129978
rect 11502 129922 11558 129978
rect 36234 130294 36290 130350
rect 36358 130294 36414 130350
rect 36482 130294 36538 130350
rect 36606 130294 36662 130350
rect 36234 130170 36290 130226
rect 36358 130170 36414 130226
rect 36482 130170 36538 130226
rect 36606 130170 36662 130226
rect 36234 130046 36290 130102
rect 36358 130046 36414 130102
rect 36482 130046 36538 130102
rect 36606 130046 36662 130102
rect 36234 129922 36290 129978
rect 36358 129922 36414 129978
rect 36482 129922 36538 129978
rect 36606 129922 36662 129978
rect 9234 118294 9290 118350
rect 9358 118294 9414 118350
rect 9482 118294 9538 118350
rect 9606 118294 9662 118350
rect 9234 118170 9290 118226
rect 9358 118170 9414 118226
rect 9482 118170 9538 118226
rect 9606 118170 9662 118226
rect 9234 118046 9290 118102
rect 9358 118046 9414 118102
rect 9482 118046 9538 118102
rect 9606 118046 9662 118102
rect 9234 117922 9290 117978
rect 9358 117922 9414 117978
rect 9482 117922 9538 117978
rect 9606 117922 9662 117978
rect 5514 94294 5570 94350
rect 5638 94294 5694 94350
rect 5762 94294 5818 94350
rect 5886 94294 5942 94350
rect 5514 94170 5570 94226
rect 5638 94170 5694 94226
rect 5762 94170 5818 94226
rect 5886 94170 5942 94226
rect 5514 94046 5570 94102
rect 5638 94046 5694 94102
rect 5762 94046 5818 94102
rect 5886 94046 5942 94102
rect 5514 93922 5570 93978
rect 5638 93922 5694 93978
rect 5762 93922 5818 93978
rect 5886 93922 5942 93978
rect 5514 76294 5570 76350
rect 5638 76294 5694 76350
rect 5762 76294 5818 76350
rect 5886 76294 5942 76350
rect 5514 76170 5570 76226
rect 5638 76170 5694 76226
rect 5762 76170 5818 76226
rect 5886 76170 5942 76226
rect 5514 76046 5570 76102
rect 5638 76046 5694 76102
rect 5762 76046 5818 76102
rect 5886 76046 5942 76102
rect 5514 75922 5570 75978
rect 5638 75922 5694 75978
rect 5762 75922 5818 75978
rect 5886 75922 5942 75978
rect 5514 58294 5570 58350
rect 5638 58294 5694 58350
rect 5762 58294 5818 58350
rect 5886 58294 5942 58350
rect 5514 58170 5570 58226
rect 5638 58170 5694 58226
rect 5762 58170 5818 58226
rect 5886 58170 5942 58226
rect 5514 58046 5570 58102
rect 5638 58046 5694 58102
rect 5762 58046 5818 58102
rect 5886 58046 5942 58102
rect 5514 57922 5570 57978
rect 5638 57922 5694 57978
rect 5762 57922 5818 57978
rect 5886 57922 5942 57978
rect 5514 40294 5570 40350
rect 5638 40294 5694 40350
rect 5762 40294 5818 40350
rect 5886 40294 5942 40350
rect 5514 40170 5570 40226
rect 5638 40170 5694 40226
rect 5762 40170 5818 40226
rect 5886 40170 5942 40226
rect 5514 40046 5570 40102
rect 5638 40046 5694 40102
rect 5762 40046 5818 40102
rect 5886 40046 5942 40102
rect 5514 39922 5570 39978
rect 5638 39922 5694 39978
rect 5762 39922 5818 39978
rect 5886 39922 5942 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 5514 22294 5570 22350
rect 5638 22294 5694 22350
rect 5762 22294 5818 22350
rect 5886 22294 5942 22350
rect 5514 22170 5570 22226
rect 5638 22170 5694 22226
rect 5762 22170 5818 22226
rect 5886 22170 5942 22226
rect 5514 22046 5570 22102
rect 5638 22046 5694 22102
rect 5762 22046 5818 22102
rect 5886 22046 5942 22102
rect 5514 21922 5570 21978
rect 5638 21922 5694 21978
rect 5762 21922 5818 21978
rect 5886 21922 5942 21978
rect 5514 4294 5570 4350
rect 5638 4294 5694 4350
rect 5762 4294 5818 4350
rect 5886 4294 5942 4350
rect 5514 4170 5570 4226
rect 5638 4170 5694 4226
rect 5762 4170 5818 4226
rect 5886 4170 5942 4226
rect 5514 4046 5570 4102
rect 5638 4046 5694 4102
rect 5762 4046 5818 4102
rect 5886 4046 5942 4102
rect 5514 3922 5570 3978
rect 5638 3922 5694 3978
rect 5762 3922 5818 3978
rect 5886 3922 5942 3978
rect 5514 -216 5570 -160
rect 5638 -216 5694 -160
rect 5762 -216 5818 -160
rect 5886 -216 5942 -160
rect 5514 -340 5570 -284
rect 5638 -340 5694 -284
rect 5762 -340 5818 -284
rect 5886 -340 5942 -284
rect 5514 -464 5570 -408
rect 5638 -464 5694 -408
rect 5762 -464 5818 -408
rect 5886 -464 5942 -408
rect 5514 -588 5570 -532
rect 5638 -588 5694 -532
rect 5762 -588 5818 -532
rect 5886 -588 5942 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 11930 118294 11986 118350
rect 12054 118294 12110 118350
rect 12178 118294 12234 118350
rect 12302 118294 12358 118350
rect 11930 118170 11986 118226
rect 12054 118170 12110 118226
rect 12178 118170 12234 118226
rect 12302 118170 12358 118226
rect 11930 118046 11986 118102
rect 12054 118046 12110 118102
rect 12178 118046 12234 118102
rect 12302 118046 12358 118102
rect 11930 117922 11986 117978
rect 12054 117922 12110 117978
rect 12178 117922 12234 117978
rect 12302 117922 12358 117978
rect 11130 112294 11186 112350
rect 11254 112294 11310 112350
rect 11378 112294 11434 112350
rect 11502 112294 11558 112350
rect 11130 112170 11186 112226
rect 11254 112170 11310 112226
rect 11378 112170 11434 112226
rect 11502 112170 11558 112226
rect 11130 112046 11186 112102
rect 11254 112046 11310 112102
rect 11378 112046 11434 112102
rect 11502 112046 11558 112102
rect 11130 111922 11186 111978
rect 11254 111922 11310 111978
rect 11378 111922 11434 111978
rect 11502 111922 11558 111978
rect 36234 112294 36290 112350
rect 36358 112294 36414 112350
rect 36482 112294 36538 112350
rect 36606 112294 36662 112350
rect 36234 112170 36290 112226
rect 36358 112170 36414 112226
rect 36482 112170 36538 112226
rect 36606 112170 36662 112226
rect 36234 112046 36290 112102
rect 36358 112046 36414 112102
rect 36482 112046 36538 112102
rect 36606 112046 36662 112102
rect 36234 111922 36290 111978
rect 36358 111922 36414 111978
rect 36482 111922 36538 111978
rect 36606 111922 36662 111978
rect 9234 100294 9290 100350
rect 9358 100294 9414 100350
rect 9482 100294 9538 100350
rect 9606 100294 9662 100350
rect 9234 100170 9290 100226
rect 9358 100170 9414 100226
rect 9482 100170 9538 100226
rect 9606 100170 9662 100226
rect 9234 100046 9290 100102
rect 9358 100046 9414 100102
rect 9482 100046 9538 100102
rect 9606 100046 9662 100102
rect 9234 99922 9290 99978
rect 9358 99922 9414 99978
rect 9482 99922 9538 99978
rect 9606 99922 9662 99978
rect 11930 100294 11986 100350
rect 12054 100294 12110 100350
rect 12178 100294 12234 100350
rect 12302 100294 12358 100350
rect 11930 100170 11986 100226
rect 12054 100170 12110 100226
rect 12178 100170 12234 100226
rect 12302 100170 12358 100226
rect 11930 100046 11986 100102
rect 12054 100046 12110 100102
rect 12178 100046 12234 100102
rect 12302 100046 12358 100102
rect 11930 99922 11986 99978
rect 12054 99922 12110 99978
rect 12178 99922 12234 99978
rect 12302 99922 12358 99978
rect 11130 94294 11186 94350
rect 11254 94294 11310 94350
rect 11378 94294 11434 94350
rect 11502 94294 11558 94350
rect 11130 94170 11186 94226
rect 11254 94170 11310 94226
rect 11378 94170 11434 94226
rect 11502 94170 11558 94226
rect 11130 94046 11186 94102
rect 11254 94046 11310 94102
rect 11378 94046 11434 94102
rect 11502 94046 11558 94102
rect 11130 93922 11186 93978
rect 11254 93922 11310 93978
rect 11378 93922 11434 93978
rect 11502 93922 11558 93978
rect 36234 94294 36290 94350
rect 36358 94294 36414 94350
rect 36482 94294 36538 94350
rect 36606 94294 36662 94350
rect 36234 94170 36290 94226
rect 36358 94170 36414 94226
rect 36482 94170 36538 94226
rect 36606 94170 36662 94226
rect 36234 94046 36290 94102
rect 36358 94046 36414 94102
rect 36482 94046 36538 94102
rect 36606 94046 36662 94102
rect 36234 93922 36290 93978
rect 36358 93922 36414 93978
rect 36482 93922 36538 93978
rect 36606 93922 36662 93978
rect 9234 82294 9290 82350
rect 9358 82294 9414 82350
rect 9482 82294 9538 82350
rect 9606 82294 9662 82350
rect 9234 82170 9290 82226
rect 9358 82170 9414 82226
rect 9482 82170 9538 82226
rect 9606 82170 9662 82226
rect 9234 82046 9290 82102
rect 9358 82046 9414 82102
rect 9482 82046 9538 82102
rect 9606 82046 9662 82102
rect 9234 81922 9290 81978
rect 9358 81922 9414 81978
rect 9482 81922 9538 81978
rect 9606 81922 9662 81978
rect 11930 82294 11986 82350
rect 12054 82294 12110 82350
rect 12178 82294 12234 82350
rect 12302 82294 12358 82350
rect 11930 82170 11986 82226
rect 12054 82170 12110 82226
rect 12178 82170 12234 82226
rect 12302 82170 12358 82226
rect 11930 82046 11986 82102
rect 12054 82046 12110 82102
rect 12178 82046 12234 82102
rect 12302 82046 12358 82102
rect 11930 81922 11986 81978
rect 12054 81922 12110 81978
rect 12178 81922 12234 81978
rect 12302 81922 12358 81978
rect 11130 76294 11186 76350
rect 11254 76294 11310 76350
rect 11378 76294 11434 76350
rect 11502 76294 11558 76350
rect 11130 76170 11186 76226
rect 11254 76170 11310 76226
rect 11378 76170 11434 76226
rect 11502 76170 11558 76226
rect 11130 76046 11186 76102
rect 11254 76046 11310 76102
rect 11378 76046 11434 76102
rect 11502 76046 11558 76102
rect 11130 75922 11186 75978
rect 11254 75922 11310 75978
rect 11378 75922 11434 75978
rect 11502 75922 11558 75978
rect 36234 76294 36290 76350
rect 36358 76294 36414 76350
rect 36482 76294 36538 76350
rect 36606 76294 36662 76350
rect 36234 76170 36290 76226
rect 36358 76170 36414 76226
rect 36482 76170 36538 76226
rect 36606 76170 36662 76226
rect 36234 76046 36290 76102
rect 36358 76046 36414 76102
rect 36482 76046 36538 76102
rect 36606 76046 36662 76102
rect 36234 75922 36290 75978
rect 36358 75922 36414 75978
rect 36482 75922 36538 75978
rect 36606 75922 36662 75978
rect 9234 64294 9290 64350
rect 9358 64294 9414 64350
rect 9482 64294 9538 64350
rect 9606 64294 9662 64350
rect 9234 64170 9290 64226
rect 9358 64170 9414 64226
rect 9482 64170 9538 64226
rect 9606 64170 9662 64226
rect 9234 64046 9290 64102
rect 9358 64046 9414 64102
rect 9482 64046 9538 64102
rect 9606 64046 9662 64102
rect 9234 63922 9290 63978
rect 9358 63922 9414 63978
rect 9482 63922 9538 63978
rect 9606 63922 9662 63978
rect 11930 64294 11986 64350
rect 12054 64294 12110 64350
rect 12178 64294 12234 64350
rect 12302 64294 12358 64350
rect 11930 64170 11986 64226
rect 12054 64170 12110 64226
rect 12178 64170 12234 64226
rect 12302 64170 12358 64226
rect 11930 64046 11986 64102
rect 12054 64046 12110 64102
rect 12178 64046 12234 64102
rect 12302 64046 12358 64102
rect 11930 63922 11986 63978
rect 12054 63922 12110 63978
rect 12178 63922 12234 63978
rect 12302 63922 12358 63978
rect 11130 58294 11186 58350
rect 11254 58294 11310 58350
rect 11378 58294 11434 58350
rect 11502 58294 11558 58350
rect 11130 58170 11186 58226
rect 11254 58170 11310 58226
rect 11378 58170 11434 58226
rect 11502 58170 11558 58226
rect 11130 58046 11186 58102
rect 11254 58046 11310 58102
rect 11378 58046 11434 58102
rect 11502 58046 11558 58102
rect 11130 57922 11186 57978
rect 11254 57922 11310 57978
rect 11378 57922 11434 57978
rect 11502 57922 11558 57978
rect 36234 58294 36290 58350
rect 36358 58294 36414 58350
rect 36482 58294 36538 58350
rect 36606 58294 36662 58350
rect 36234 58170 36290 58226
rect 36358 58170 36414 58226
rect 36482 58170 36538 58226
rect 36606 58170 36662 58226
rect 36234 58046 36290 58102
rect 36358 58046 36414 58102
rect 36482 58046 36538 58102
rect 36606 58046 36662 58102
rect 36234 57922 36290 57978
rect 36358 57922 36414 57978
rect 36482 57922 36538 57978
rect 36606 57922 36662 57978
rect 9234 46294 9290 46350
rect 9358 46294 9414 46350
rect 9482 46294 9538 46350
rect 9606 46294 9662 46350
rect 9234 46170 9290 46226
rect 9358 46170 9414 46226
rect 9482 46170 9538 46226
rect 9606 46170 9662 46226
rect 9234 46046 9290 46102
rect 9358 46046 9414 46102
rect 9482 46046 9538 46102
rect 9606 46046 9662 46102
rect 9234 45922 9290 45978
rect 9358 45922 9414 45978
rect 9482 45922 9538 45978
rect 9606 45922 9662 45978
rect 9234 28294 9290 28350
rect 9358 28294 9414 28350
rect 9482 28294 9538 28350
rect 9606 28294 9662 28350
rect 9234 28170 9290 28226
rect 9358 28170 9414 28226
rect 9482 28170 9538 28226
rect 9606 28170 9662 28226
rect 9234 28046 9290 28102
rect 9358 28046 9414 28102
rect 9482 28046 9538 28102
rect 9606 28046 9662 28102
rect 9234 27922 9290 27978
rect 9358 27922 9414 27978
rect 9482 27922 9538 27978
rect 9606 27922 9662 27978
rect 9234 10294 9290 10350
rect 9358 10294 9414 10350
rect 9482 10294 9538 10350
rect 9606 10294 9662 10350
rect 9234 10170 9290 10226
rect 9358 10170 9414 10226
rect 9482 10170 9538 10226
rect 9606 10170 9662 10226
rect 9234 10046 9290 10102
rect 9358 10046 9414 10102
rect 9482 10046 9538 10102
rect 9606 10046 9662 10102
rect 9234 9922 9290 9978
rect 9358 9922 9414 9978
rect 9482 9922 9538 9978
rect 9606 9922 9662 9978
rect 9234 -1176 9290 -1120
rect 9358 -1176 9414 -1120
rect 9482 -1176 9538 -1120
rect 9606 -1176 9662 -1120
rect 9234 -1300 9290 -1244
rect 9358 -1300 9414 -1244
rect 9482 -1300 9538 -1244
rect 9606 -1300 9662 -1244
rect 9234 -1424 9290 -1368
rect 9358 -1424 9414 -1368
rect 9482 -1424 9538 -1368
rect 9606 -1424 9662 -1368
rect 9234 -1548 9290 -1492
rect 9358 -1548 9414 -1492
rect 9482 -1548 9538 -1492
rect 9606 -1548 9662 -1492
rect 36234 40294 36290 40350
rect 36358 40294 36414 40350
rect 36482 40294 36538 40350
rect 36606 40294 36662 40350
rect 36234 40170 36290 40226
rect 36358 40170 36414 40226
rect 36482 40170 36538 40226
rect 36606 40170 36662 40226
rect 36234 40046 36290 40102
rect 36358 40046 36414 40102
rect 36482 40046 36538 40102
rect 36606 40046 36662 40102
rect 36234 39922 36290 39978
rect 36358 39922 36414 39978
rect 36482 39922 36538 39978
rect 36606 39922 36662 39978
rect 36234 22294 36290 22350
rect 36358 22294 36414 22350
rect 36482 22294 36538 22350
rect 36606 22294 36662 22350
rect 36234 22170 36290 22226
rect 36358 22170 36414 22226
rect 36482 22170 36538 22226
rect 36606 22170 36662 22226
rect 36234 22046 36290 22102
rect 36358 22046 36414 22102
rect 36482 22046 36538 22102
rect 36606 22046 36662 22102
rect 36234 21922 36290 21978
rect 36358 21922 36414 21978
rect 36482 21922 36538 21978
rect 36606 21922 36662 21978
rect 36234 4294 36290 4350
rect 36358 4294 36414 4350
rect 36482 4294 36538 4350
rect 36606 4294 36662 4350
rect 36234 4170 36290 4226
rect 36358 4170 36414 4226
rect 36482 4170 36538 4226
rect 36606 4170 36662 4226
rect 36234 4046 36290 4102
rect 36358 4046 36414 4102
rect 36482 4046 36538 4102
rect 36606 4046 36662 4102
rect 36234 3922 36290 3978
rect 36358 3922 36414 3978
rect 36482 3922 36538 3978
rect 36606 3922 36662 3978
rect 36234 -216 36290 -160
rect 36358 -216 36414 -160
rect 36482 -216 36538 -160
rect 36606 -216 36662 -160
rect 36234 -340 36290 -284
rect 36358 -340 36414 -284
rect 36482 -340 36538 -284
rect 36606 -340 36662 -284
rect 36234 -464 36290 -408
rect 36358 -464 36414 -408
rect 36482 -464 36538 -408
rect 36606 -464 36662 -408
rect 36234 -588 36290 -532
rect 36358 -588 36414 -532
rect 36482 -588 36538 -532
rect 36606 -588 36662 -532
rect 39954 154294 40010 154350
rect 40078 154294 40134 154350
rect 40202 154294 40258 154350
rect 40326 154294 40382 154350
rect 39954 154170 40010 154226
rect 40078 154170 40134 154226
rect 40202 154170 40258 154226
rect 40326 154170 40382 154226
rect 39954 154046 40010 154102
rect 40078 154046 40134 154102
rect 40202 154046 40258 154102
rect 40326 154046 40382 154102
rect 39954 153922 40010 153978
rect 40078 153922 40134 153978
rect 40202 153922 40258 153978
rect 40326 153922 40382 153978
rect 66954 580294 67010 580350
rect 67078 580294 67134 580350
rect 67202 580294 67258 580350
rect 67326 580294 67382 580350
rect 66954 580170 67010 580226
rect 67078 580170 67134 580226
rect 67202 580170 67258 580226
rect 67326 580170 67382 580226
rect 66954 580046 67010 580102
rect 67078 580046 67134 580102
rect 67202 580046 67258 580102
rect 67326 580046 67382 580102
rect 66954 579922 67010 579978
rect 67078 579922 67134 579978
rect 67202 579922 67258 579978
rect 67326 579922 67382 579978
rect 66954 562294 67010 562350
rect 67078 562294 67134 562350
rect 67202 562294 67258 562350
rect 67326 562294 67382 562350
rect 66954 562170 67010 562226
rect 67078 562170 67134 562226
rect 67202 562170 67258 562226
rect 67326 562170 67382 562226
rect 66954 562046 67010 562102
rect 67078 562046 67134 562102
rect 67202 562046 67258 562102
rect 67326 562046 67382 562102
rect 66954 561922 67010 561978
rect 67078 561922 67134 561978
rect 67202 561922 67258 561978
rect 67326 561922 67382 561978
rect 66954 544294 67010 544350
rect 67078 544294 67134 544350
rect 67202 544294 67258 544350
rect 67326 544294 67382 544350
rect 66954 544170 67010 544226
rect 67078 544170 67134 544226
rect 67202 544170 67258 544226
rect 67326 544170 67382 544226
rect 66954 544046 67010 544102
rect 67078 544046 67134 544102
rect 67202 544046 67258 544102
rect 67326 544046 67382 544102
rect 66954 543922 67010 543978
rect 67078 543922 67134 543978
rect 67202 543922 67258 543978
rect 67326 543922 67382 543978
rect 57036 324962 57092 325018
rect 57932 283382 57988 283438
rect 56476 283022 56532 283078
rect 56364 281942 56420 281998
rect 58156 284642 58212 284698
rect 58716 307502 58772 307558
rect 58380 286442 58436 286498
rect 59724 368702 59780 368758
rect 58716 287342 58772 287398
rect 58716 283922 58772 283978
rect 58492 283202 58548 283258
rect 58716 282302 58772 282358
rect 58268 282122 58324 282178
rect 66954 526294 67010 526350
rect 67078 526294 67134 526350
rect 67202 526294 67258 526350
rect 67326 526294 67382 526350
rect 66954 526170 67010 526226
rect 67078 526170 67134 526226
rect 67202 526170 67258 526226
rect 67326 526170 67382 526226
rect 66954 526046 67010 526102
rect 67078 526046 67134 526102
rect 67202 526046 67258 526102
rect 67326 526046 67382 526102
rect 66954 525922 67010 525978
rect 67078 525922 67134 525978
rect 67202 525922 67258 525978
rect 67326 525922 67382 525978
rect 66954 508294 67010 508350
rect 67078 508294 67134 508350
rect 67202 508294 67258 508350
rect 67326 508294 67382 508350
rect 66954 508170 67010 508226
rect 67078 508170 67134 508226
rect 67202 508170 67258 508226
rect 67326 508170 67382 508226
rect 66954 508046 67010 508102
rect 67078 508046 67134 508102
rect 67202 508046 67258 508102
rect 67326 508046 67382 508102
rect 66954 507922 67010 507978
rect 67078 507922 67134 507978
rect 67202 507922 67258 507978
rect 67326 507922 67382 507978
rect 66954 490294 67010 490350
rect 67078 490294 67134 490350
rect 67202 490294 67258 490350
rect 67326 490294 67382 490350
rect 66954 490170 67010 490226
rect 67078 490170 67134 490226
rect 67202 490170 67258 490226
rect 67326 490170 67382 490226
rect 66954 490046 67010 490102
rect 67078 490046 67134 490102
rect 67202 490046 67258 490102
rect 67326 490046 67382 490102
rect 66954 489922 67010 489978
rect 67078 489922 67134 489978
rect 67202 489922 67258 489978
rect 67326 489922 67382 489978
rect 60172 321020 60228 321058
rect 60172 321002 60228 321020
rect 58044 276362 58100 276418
rect 66954 472294 67010 472350
rect 67078 472294 67134 472350
rect 67202 472294 67258 472350
rect 67326 472294 67382 472350
rect 66954 472170 67010 472226
rect 67078 472170 67134 472226
rect 67202 472170 67258 472226
rect 67326 472170 67382 472226
rect 66954 472046 67010 472102
rect 67078 472046 67134 472102
rect 67202 472046 67258 472102
rect 67326 472046 67382 472102
rect 66954 471922 67010 471978
rect 67078 471922 67134 471978
rect 67202 471922 67258 471978
rect 67326 471922 67382 471978
rect 66954 454294 67010 454350
rect 67078 454294 67134 454350
rect 67202 454294 67258 454350
rect 67326 454294 67382 454350
rect 66954 454170 67010 454226
rect 67078 454170 67134 454226
rect 67202 454170 67258 454226
rect 67326 454170 67382 454226
rect 66954 454046 67010 454102
rect 67078 454046 67134 454102
rect 67202 454046 67258 454102
rect 67326 454046 67382 454102
rect 66954 453922 67010 453978
rect 67078 453922 67134 453978
rect 67202 453922 67258 453978
rect 67326 453922 67382 453978
rect 66954 436294 67010 436350
rect 67078 436294 67134 436350
rect 67202 436294 67258 436350
rect 67326 436294 67382 436350
rect 66954 436170 67010 436226
rect 67078 436170 67134 436226
rect 67202 436170 67258 436226
rect 67326 436170 67382 436226
rect 66954 436046 67010 436102
rect 67078 436046 67134 436102
rect 67202 436046 67258 436102
rect 67326 436046 67382 436102
rect 66954 435922 67010 435978
rect 67078 435922 67134 435978
rect 67202 435922 67258 435978
rect 67326 435922 67382 435978
rect 66954 418294 67010 418350
rect 67078 418294 67134 418350
rect 67202 418294 67258 418350
rect 67326 418294 67382 418350
rect 66954 418170 67010 418226
rect 67078 418170 67134 418226
rect 67202 418170 67258 418226
rect 67326 418170 67382 418226
rect 66954 418046 67010 418102
rect 67078 418046 67134 418102
rect 67202 418046 67258 418102
rect 67326 418046 67382 418102
rect 66954 417922 67010 417978
rect 67078 417922 67134 417978
rect 67202 417922 67258 417978
rect 67326 417922 67382 417978
rect 66954 400294 67010 400350
rect 67078 400294 67134 400350
rect 67202 400294 67258 400350
rect 67326 400294 67382 400350
rect 66954 400170 67010 400226
rect 67078 400170 67134 400226
rect 67202 400170 67258 400226
rect 67326 400170 67382 400226
rect 66954 400046 67010 400102
rect 67078 400046 67134 400102
rect 67202 400046 67258 400102
rect 67326 400046 67382 400102
rect 66954 399922 67010 399978
rect 67078 399922 67134 399978
rect 67202 399922 67258 399978
rect 67326 399922 67382 399978
rect 66954 382294 67010 382350
rect 67078 382294 67134 382350
rect 67202 382294 67258 382350
rect 67326 382294 67382 382350
rect 66954 382170 67010 382226
rect 67078 382170 67134 382226
rect 67202 382170 67258 382226
rect 67326 382170 67382 382226
rect 66954 382046 67010 382102
rect 67078 382046 67134 382102
rect 67202 382046 67258 382102
rect 67326 382046 67382 382102
rect 66954 381922 67010 381978
rect 67078 381922 67134 381978
rect 67202 381922 67258 381978
rect 67326 381922 67382 381978
rect 66954 364294 67010 364350
rect 67078 364294 67134 364350
rect 67202 364294 67258 364350
rect 67326 364294 67382 364350
rect 66954 364170 67010 364226
rect 67078 364170 67134 364226
rect 67202 364170 67258 364226
rect 67326 364170 67382 364226
rect 66954 364046 67010 364102
rect 67078 364046 67134 364102
rect 67202 364046 67258 364102
rect 67326 364046 67382 364102
rect 66954 363922 67010 363978
rect 67078 363922 67134 363978
rect 67202 363922 67258 363978
rect 67326 363922 67382 363978
rect 61292 321002 61348 321058
rect 60396 276002 60452 276058
rect 62972 307502 63028 307558
rect 62188 276542 62244 276598
rect 63532 276902 63588 276958
rect 66954 346294 67010 346350
rect 67078 346294 67134 346350
rect 67202 346294 67258 346350
rect 67326 346294 67382 346350
rect 66954 346170 67010 346226
rect 67078 346170 67134 346226
rect 67202 346170 67258 346226
rect 67326 346170 67382 346226
rect 66954 346046 67010 346102
rect 67078 346046 67134 346102
rect 67202 346046 67258 346102
rect 67326 346046 67382 346102
rect 66954 345922 67010 345978
rect 67078 345922 67134 345978
rect 67202 345922 67258 345978
rect 67326 345922 67382 345978
rect 70674 598116 70730 598172
rect 70798 598116 70854 598172
rect 70922 598116 70978 598172
rect 71046 598116 71102 598172
rect 70674 597992 70730 598048
rect 70798 597992 70854 598048
rect 70922 597992 70978 598048
rect 71046 597992 71102 598048
rect 70674 597868 70730 597924
rect 70798 597868 70854 597924
rect 70922 597868 70978 597924
rect 71046 597868 71102 597924
rect 70674 597744 70730 597800
rect 70798 597744 70854 597800
rect 70922 597744 70978 597800
rect 71046 597744 71102 597800
rect 70674 586294 70730 586350
rect 70798 586294 70854 586350
rect 70922 586294 70978 586350
rect 71046 586294 71102 586350
rect 70674 586170 70730 586226
rect 70798 586170 70854 586226
rect 70922 586170 70978 586226
rect 71046 586170 71102 586226
rect 70674 586046 70730 586102
rect 70798 586046 70854 586102
rect 70922 586046 70978 586102
rect 71046 586046 71102 586102
rect 70674 585922 70730 585978
rect 70798 585922 70854 585978
rect 70922 585922 70978 585978
rect 71046 585922 71102 585978
rect 70674 568294 70730 568350
rect 70798 568294 70854 568350
rect 70922 568294 70978 568350
rect 71046 568294 71102 568350
rect 70674 568170 70730 568226
rect 70798 568170 70854 568226
rect 70922 568170 70978 568226
rect 71046 568170 71102 568226
rect 70674 568046 70730 568102
rect 70798 568046 70854 568102
rect 70922 568046 70978 568102
rect 71046 568046 71102 568102
rect 70674 567922 70730 567978
rect 70798 567922 70854 567978
rect 70922 567922 70978 567978
rect 71046 567922 71102 567978
rect 70674 550294 70730 550350
rect 70798 550294 70854 550350
rect 70922 550294 70978 550350
rect 71046 550294 71102 550350
rect 70674 550170 70730 550226
rect 70798 550170 70854 550226
rect 70922 550170 70978 550226
rect 71046 550170 71102 550226
rect 70674 550046 70730 550102
rect 70798 550046 70854 550102
rect 70922 550046 70978 550102
rect 71046 550046 71102 550102
rect 70674 549922 70730 549978
rect 70798 549922 70854 549978
rect 70922 549922 70978 549978
rect 71046 549922 71102 549978
rect 70674 532294 70730 532350
rect 70798 532294 70854 532350
rect 70922 532294 70978 532350
rect 71046 532294 71102 532350
rect 70674 532170 70730 532226
rect 70798 532170 70854 532226
rect 70922 532170 70978 532226
rect 71046 532170 71102 532226
rect 70674 532046 70730 532102
rect 70798 532046 70854 532102
rect 70922 532046 70978 532102
rect 71046 532046 71102 532102
rect 70674 531922 70730 531978
rect 70798 531922 70854 531978
rect 70922 531922 70978 531978
rect 71046 531922 71102 531978
rect 70674 514294 70730 514350
rect 70798 514294 70854 514350
rect 70922 514294 70978 514350
rect 71046 514294 71102 514350
rect 70674 514170 70730 514226
rect 70798 514170 70854 514226
rect 70922 514170 70978 514226
rect 71046 514170 71102 514226
rect 70674 514046 70730 514102
rect 70798 514046 70854 514102
rect 70922 514046 70978 514102
rect 71046 514046 71102 514102
rect 70674 513922 70730 513978
rect 70798 513922 70854 513978
rect 70922 513922 70978 513978
rect 71046 513922 71102 513978
rect 70674 496294 70730 496350
rect 70798 496294 70854 496350
rect 70922 496294 70978 496350
rect 71046 496294 71102 496350
rect 70674 496170 70730 496226
rect 70798 496170 70854 496226
rect 70922 496170 70978 496226
rect 71046 496170 71102 496226
rect 70674 496046 70730 496102
rect 70798 496046 70854 496102
rect 70922 496046 70978 496102
rect 71046 496046 71102 496102
rect 70674 495922 70730 495978
rect 70798 495922 70854 495978
rect 70922 495922 70978 495978
rect 71046 495922 71102 495978
rect 70674 478294 70730 478350
rect 70798 478294 70854 478350
rect 70922 478294 70978 478350
rect 71046 478294 71102 478350
rect 70674 478170 70730 478226
rect 70798 478170 70854 478226
rect 70922 478170 70978 478226
rect 71046 478170 71102 478226
rect 70674 478046 70730 478102
rect 70798 478046 70854 478102
rect 70922 478046 70978 478102
rect 71046 478046 71102 478102
rect 70674 477922 70730 477978
rect 70798 477922 70854 477978
rect 70922 477922 70978 477978
rect 71046 477922 71102 477978
rect 70674 460294 70730 460350
rect 70798 460294 70854 460350
rect 70922 460294 70978 460350
rect 71046 460294 71102 460350
rect 70674 460170 70730 460226
rect 70798 460170 70854 460226
rect 70922 460170 70978 460226
rect 71046 460170 71102 460226
rect 70674 460046 70730 460102
rect 70798 460046 70854 460102
rect 70922 460046 70978 460102
rect 71046 460046 71102 460102
rect 70674 459922 70730 459978
rect 70798 459922 70854 459978
rect 70922 459922 70978 459978
rect 71046 459922 71102 459978
rect 70674 442294 70730 442350
rect 70798 442294 70854 442350
rect 70922 442294 70978 442350
rect 71046 442294 71102 442350
rect 70674 442170 70730 442226
rect 70798 442170 70854 442226
rect 70922 442170 70978 442226
rect 71046 442170 71102 442226
rect 70674 442046 70730 442102
rect 70798 442046 70854 442102
rect 70922 442046 70978 442102
rect 71046 442046 71102 442102
rect 70674 441922 70730 441978
rect 70798 441922 70854 441978
rect 70922 441922 70978 441978
rect 71046 441922 71102 441978
rect 70674 424294 70730 424350
rect 70798 424294 70854 424350
rect 70922 424294 70978 424350
rect 71046 424294 71102 424350
rect 70674 424170 70730 424226
rect 70798 424170 70854 424226
rect 70922 424170 70978 424226
rect 71046 424170 71102 424226
rect 70674 424046 70730 424102
rect 70798 424046 70854 424102
rect 70922 424046 70978 424102
rect 71046 424046 71102 424102
rect 70674 423922 70730 423978
rect 70798 423922 70854 423978
rect 70922 423922 70978 423978
rect 71046 423922 71102 423978
rect 70674 406294 70730 406350
rect 70798 406294 70854 406350
rect 70922 406294 70978 406350
rect 71046 406294 71102 406350
rect 70674 406170 70730 406226
rect 70798 406170 70854 406226
rect 70922 406170 70978 406226
rect 71046 406170 71102 406226
rect 70674 406046 70730 406102
rect 70798 406046 70854 406102
rect 70922 406046 70978 406102
rect 71046 406046 71102 406102
rect 70674 405922 70730 405978
rect 70798 405922 70854 405978
rect 70922 405922 70978 405978
rect 71046 405922 71102 405978
rect 70674 388294 70730 388350
rect 70798 388294 70854 388350
rect 70922 388294 70978 388350
rect 71046 388294 71102 388350
rect 70674 388170 70730 388226
rect 70798 388170 70854 388226
rect 70922 388170 70978 388226
rect 71046 388170 71102 388226
rect 70674 388046 70730 388102
rect 70798 388046 70854 388102
rect 70922 388046 70978 388102
rect 71046 388046 71102 388102
rect 70674 387922 70730 387978
rect 70798 387922 70854 387978
rect 70922 387922 70978 387978
rect 71046 387922 71102 387978
rect 70674 370294 70730 370350
rect 70798 370294 70854 370350
rect 70922 370294 70978 370350
rect 71046 370294 71102 370350
rect 70674 370170 70730 370226
rect 70798 370170 70854 370226
rect 70922 370170 70978 370226
rect 71046 370170 71102 370226
rect 70674 370046 70730 370102
rect 70798 370046 70854 370102
rect 70922 370046 70978 370102
rect 71046 370046 71102 370102
rect 70674 369922 70730 369978
rect 70798 369922 70854 369978
rect 70922 369922 70978 369978
rect 71046 369922 71102 369978
rect 70674 352294 70730 352350
rect 70798 352294 70854 352350
rect 70922 352294 70978 352350
rect 71046 352294 71102 352350
rect 70674 352170 70730 352226
rect 70798 352170 70854 352226
rect 70922 352170 70978 352226
rect 71046 352170 71102 352226
rect 70674 352046 70730 352102
rect 70798 352046 70854 352102
rect 70922 352046 70978 352102
rect 71046 352046 71102 352102
rect 70674 351922 70730 351978
rect 70798 351922 70854 351978
rect 70922 351922 70978 351978
rect 71046 351922 71102 351978
rect 97674 597156 97730 597212
rect 97798 597156 97854 597212
rect 97922 597156 97978 597212
rect 98046 597156 98102 597212
rect 97674 597032 97730 597088
rect 97798 597032 97854 597088
rect 97922 597032 97978 597088
rect 98046 597032 98102 597088
rect 97674 596908 97730 596964
rect 97798 596908 97854 596964
rect 97922 596908 97978 596964
rect 98046 596908 98102 596964
rect 97674 596784 97730 596840
rect 97798 596784 97854 596840
rect 97922 596784 97978 596840
rect 98046 596784 98102 596840
rect 97674 580294 97730 580350
rect 97798 580294 97854 580350
rect 97922 580294 97978 580350
rect 98046 580294 98102 580350
rect 97674 580170 97730 580226
rect 97798 580170 97854 580226
rect 97922 580170 97978 580226
rect 98046 580170 98102 580226
rect 97674 580046 97730 580102
rect 97798 580046 97854 580102
rect 97922 580046 97978 580102
rect 98046 580046 98102 580102
rect 97674 579922 97730 579978
rect 97798 579922 97854 579978
rect 97922 579922 97978 579978
rect 98046 579922 98102 579978
rect 97674 562294 97730 562350
rect 97798 562294 97854 562350
rect 97922 562294 97978 562350
rect 98046 562294 98102 562350
rect 97674 562170 97730 562226
rect 97798 562170 97854 562226
rect 97922 562170 97978 562226
rect 98046 562170 98102 562226
rect 97674 562046 97730 562102
rect 97798 562046 97854 562102
rect 97922 562046 97978 562102
rect 98046 562046 98102 562102
rect 97674 561922 97730 561978
rect 97798 561922 97854 561978
rect 97922 561922 97978 561978
rect 98046 561922 98102 561978
rect 97674 544294 97730 544350
rect 97798 544294 97854 544350
rect 97922 544294 97978 544350
rect 98046 544294 98102 544350
rect 97674 544170 97730 544226
rect 97798 544170 97854 544226
rect 97922 544170 97978 544226
rect 98046 544170 98102 544226
rect 97674 544046 97730 544102
rect 97798 544046 97854 544102
rect 97922 544046 97978 544102
rect 98046 544046 98102 544102
rect 97674 543922 97730 543978
rect 97798 543922 97854 543978
rect 97922 543922 97978 543978
rect 98046 543922 98102 543978
rect 97674 526294 97730 526350
rect 97798 526294 97854 526350
rect 97922 526294 97978 526350
rect 98046 526294 98102 526350
rect 97674 526170 97730 526226
rect 97798 526170 97854 526226
rect 97922 526170 97978 526226
rect 98046 526170 98102 526226
rect 97674 526046 97730 526102
rect 97798 526046 97854 526102
rect 97922 526046 97978 526102
rect 98046 526046 98102 526102
rect 97674 525922 97730 525978
rect 97798 525922 97854 525978
rect 97922 525922 97978 525978
rect 98046 525922 98102 525978
rect 97674 508294 97730 508350
rect 97798 508294 97854 508350
rect 97922 508294 97978 508350
rect 98046 508294 98102 508350
rect 97674 508170 97730 508226
rect 97798 508170 97854 508226
rect 97922 508170 97978 508226
rect 98046 508170 98102 508226
rect 97674 508046 97730 508102
rect 97798 508046 97854 508102
rect 97922 508046 97978 508102
rect 98046 508046 98102 508102
rect 97674 507922 97730 507978
rect 97798 507922 97854 507978
rect 97922 507922 97978 507978
rect 98046 507922 98102 507978
rect 97674 490294 97730 490350
rect 97798 490294 97854 490350
rect 97922 490294 97978 490350
rect 98046 490294 98102 490350
rect 97674 490170 97730 490226
rect 97798 490170 97854 490226
rect 97922 490170 97978 490226
rect 98046 490170 98102 490226
rect 97674 490046 97730 490102
rect 97798 490046 97854 490102
rect 97922 490046 97978 490102
rect 98046 490046 98102 490102
rect 97674 489922 97730 489978
rect 97798 489922 97854 489978
rect 97922 489922 97978 489978
rect 98046 489922 98102 489978
rect 97674 472294 97730 472350
rect 97798 472294 97854 472350
rect 97922 472294 97978 472350
rect 98046 472294 98102 472350
rect 97674 472170 97730 472226
rect 97798 472170 97854 472226
rect 97922 472170 97978 472226
rect 98046 472170 98102 472226
rect 97674 472046 97730 472102
rect 97798 472046 97854 472102
rect 97922 472046 97978 472102
rect 98046 472046 98102 472102
rect 97674 471922 97730 471978
rect 97798 471922 97854 471978
rect 97922 471922 97978 471978
rect 98046 471922 98102 471978
rect 97674 454294 97730 454350
rect 97798 454294 97854 454350
rect 97922 454294 97978 454350
rect 98046 454294 98102 454350
rect 97674 454170 97730 454226
rect 97798 454170 97854 454226
rect 97922 454170 97978 454226
rect 98046 454170 98102 454226
rect 97674 454046 97730 454102
rect 97798 454046 97854 454102
rect 97922 454046 97978 454102
rect 98046 454046 98102 454102
rect 97674 453922 97730 453978
rect 97798 453922 97854 453978
rect 97922 453922 97978 453978
rect 98046 453922 98102 453978
rect 97674 436294 97730 436350
rect 97798 436294 97854 436350
rect 97922 436294 97978 436350
rect 98046 436294 98102 436350
rect 97674 436170 97730 436226
rect 97798 436170 97854 436226
rect 97922 436170 97978 436226
rect 98046 436170 98102 436226
rect 97674 436046 97730 436102
rect 97798 436046 97854 436102
rect 97922 436046 97978 436102
rect 98046 436046 98102 436102
rect 97674 435922 97730 435978
rect 97798 435922 97854 435978
rect 97922 435922 97978 435978
rect 98046 435922 98102 435978
rect 97674 418294 97730 418350
rect 97798 418294 97854 418350
rect 97922 418294 97978 418350
rect 98046 418294 98102 418350
rect 97674 418170 97730 418226
rect 97798 418170 97854 418226
rect 97922 418170 97978 418226
rect 98046 418170 98102 418226
rect 97674 418046 97730 418102
rect 97798 418046 97854 418102
rect 97922 418046 97978 418102
rect 98046 418046 98102 418102
rect 97674 417922 97730 417978
rect 97798 417922 97854 417978
rect 97922 417922 97978 417978
rect 98046 417922 98102 417978
rect 97674 400294 97730 400350
rect 97798 400294 97854 400350
rect 97922 400294 97978 400350
rect 98046 400294 98102 400350
rect 97674 400170 97730 400226
rect 97798 400170 97854 400226
rect 97922 400170 97978 400226
rect 98046 400170 98102 400226
rect 97674 400046 97730 400102
rect 97798 400046 97854 400102
rect 97922 400046 97978 400102
rect 98046 400046 98102 400102
rect 97674 399922 97730 399978
rect 97798 399922 97854 399978
rect 97922 399922 97978 399978
rect 98046 399922 98102 399978
rect 97674 382294 97730 382350
rect 97798 382294 97854 382350
rect 97922 382294 97978 382350
rect 98046 382294 98102 382350
rect 97674 382170 97730 382226
rect 97798 382170 97854 382226
rect 97922 382170 97978 382226
rect 98046 382170 98102 382226
rect 97674 382046 97730 382102
rect 97798 382046 97854 382102
rect 97922 382046 97978 382102
rect 98046 382046 98102 382102
rect 97674 381922 97730 381978
rect 97798 381922 97854 381978
rect 97922 381922 97978 381978
rect 98046 381922 98102 381978
rect 97674 364294 97730 364350
rect 97798 364294 97854 364350
rect 97922 364294 97978 364350
rect 98046 364294 98102 364350
rect 97674 364170 97730 364226
rect 97798 364170 97854 364226
rect 97922 364170 97978 364226
rect 98046 364170 98102 364226
rect 97674 364046 97730 364102
rect 97798 364046 97854 364102
rect 97922 364046 97978 364102
rect 98046 364046 98102 364102
rect 97674 363922 97730 363978
rect 97798 363922 97854 363978
rect 97922 363922 97978 363978
rect 98046 363922 98102 363978
rect 70674 334294 70730 334350
rect 70798 334294 70854 334350
rect 70922 334294 70978 334350
rect 71046 334294 71102 334350
rect 70674 334170 70730 334226
rect 70798 334170 70854 334226
rect 70922 334170 70978 334226
rect 71046 334170 71102 334226
rect 70674 334046 70730 334102
rect 70798 334046 70854 334102
rect 70922 334046 70978 334102
rect 71046 334046 71102 334102
rect 70674 333922 70730 333978
rect 70798 333922 70854 333978
rect 70922 333922 70978 333978
rect 71046 333922 71102 333978
rect 97674 346294 97730 346350
rect 97798 346294 97854 346350
rect 97922 346294 97978 346350
rect 98046 346294 98102 346350
rect 97674 346170 97730 346226
rect 97798 346170 97854 346226
rect 97922 346170 97978 346226
rect 98046 346170 98102 346226
rect 97674 346046 97730 346102
rect 97798 346046 97854 346102
rect 97922 346046 97978 346102
rect 98046 346046 98102 346102
rect 97674 345922 97730 345978
rect 97798 345922 97854 345978
rect 97922 345922 97978 345978
rect 98046 345922 98102 345978
rect 101394 598116 101450 598172
rect 101518 598116 101574 598172
rect 101642 598116 101698 598172
rect 101766 598116 101822 598172
rect 101394 597992 101450 598048
rect 101518 597992 101574 598048
rect 101642 597992 101698 598048
rect 101766 597992 101822 598048
rect 101394 597868 101450 597924
rect 101518 597868 101574 597924
rect 101642 597868 101698 597924
rect 101766 597868 101822 597924
rect 101394 597744 101450 597800
rect 101518 597744 101574 597800
rect 101642 597744 101698 597800
rect 101766 597744 101822 597800
rect 128394 597156 128450 597212
rect 128518 597156 128574 597212
rect 128642 597156 128698 597212
rect 128766 597156 128822 597212
rect 128394 597032 128450 597088
rect 128518 597032 128574 597088
rect 128642 597032 128698 597088
rect 128766 597032 128822 597088
rect 128394 596908 128450 596964
rect 128518 596908 128574 596964
rect 128642 596908 128698 596964
rect 128766 596908 128822 596964
rect 128394 596784 128450 596840
rect 128518 596784 128574 596840
rect 128642 596784 128698 596840
rect 128766 596784 128822 596840
rect 101394 586294 101450 586350
rect 101518 586294 101574 586350
rect 101642 586294 101698 586350
rect 101766 586294 101822 586350
rect 101394 586170 101450 586226
rect 101518 586170 101574 586226
rect 101642 586170 101698 586226
rect 101766 586170 101822 586226
rect 101394 586046 101450 586102
rect 101518 586046 101574 586102
rect 101642 586046 101698 586102
rect 101766 586046 101822 586102
rect 101394 585922 101450 585978
rect 101518 585922 101574 585978
rect 101642 585922 101698 585978
rect 101766 585922 101822 585978
rect 101394 568294 101450 568350
rect 101518 568294 101574 568350
rect 101642 568294 101698 568350
rect 101766 568294 101822 568350
rect 101394 568170 101450 568226
rect 101518 568170 101574 568226
rect 101642 568170 101698 568226
rect 101766 568170 101822 568226
rect 101394 568046 101450 568102
rect 101518 568046 101574 568102
rect 101642 568046 101698 568102
rect 101766 568046 101822 568102
rect 101394 567922 101450 567978
rect 101518 567922 101574 567978
rect 101642 567922 101698 567978
rect 101766 567922 101822 567978
rect 101394 550294 101450 550350
rect 101518 550294 101574 550350
rect 101642 550294 101698 550350
rect 101766 550294 101822 550350
rect 101394 550170 101450 550226
rect 101518 550170 101574 550226
rect 101642 550170 101698 550226
rect 101766 550170 101822 550226
rect 101394 550046 101450 550102
rect 101518 550046 101574 550102
rect 101642 550046 101698 550102
rect 101766 550046 101822 550102
rect 101394 549922 101450 549978
rect 101518 549922 101574 549978
rect 101642 549922 101698 549978
rect 101766 549922 101822 549978
rect 101394 532294 101450 532350
rect 101518 532294 101574 532350
rect 101642 532294 101698 532350
rect 101766 532294 101822 532350
rect 101394 532170 101450 532226
rect 101518 532170 101574 532226
rect 101642 532170 101698 532226
rect 101766 532170 101822 532226
rect 101394 532046 101450 532102
rect 101518 532046 101574 532102
rect 101642 532046 101698 532102
rect 101766 532046 101822 532102
rect 101394 531922 101450 531978
rect 101518 531922 101574 531978
rect 101642 531922 101698 531978
rect 101766 531922 101822 531978
rect 101394 514294 101450 514350
rect 101518 514294 101574 514350
rect 101642 514294 101698 514350
rect 101766 514294 101822 514350
rect 101394 514170 101450 514226
rect 101518 514170 101574 514226
rect 101642 514170 101698 514226
rect 101766 514170 101822 514226
rect 101394 514046 101450 514102
rect 101518 514046 101574 514102
rect 101642 514046 101698 514102
rect 101766 514046 101822 514102
rect 101394 513922 101450 513978
rect 101518 513922 101574 513978
rect 101642 513922 101698 513978
rect 101766 513922 101822 513978
rect 101394 496294 101450 496350
rect 101518 496294 101574 496350
rect 101642 496294 101698 496350
rect 101766 496294 101822 496350
rect 101394 496170 101450 496226
rect 101518 496170 101574 496226
rect 101642 496170 101698 496226
rect 101766 496170 101822 496226
rect 101394 496046 101450 496102
rect 101518 496046 101574 496102
rect 101642 496046 101698 496102
rect 101766 496046 101822 496102
rect 101394 495922 101450 495978
rect 101518 495922 101574 495978
rect 101642 495922 101698 495978
rect 101766 495922 101822 495978
rect 101394 478294 101450 478350
rect 101518 478294 101574 478350
rect 101642 478294 101698 478350
rect 101766 478294 101822 478350
rect 101394 478170 101450 478226
rect 101518 478170 101574 478226
rect 101642 478170 101698 478226
rect 101766 478170 101822 478226
rect 101394 478046 101450 478102
rect 101518 478046 101574 478102
rect 101642 478046 101698 478102
rect 101766 478046 101822 478102
rect 101394 477922 101450 477978
rect 101518 477922 101574 477978
rect 101642 477922 101698 477978
rect 101766 477922 101822 477978
rect 101394 460294 101450 460350
rect 101518 460294 101574 460350
rect 101642 460294 101698 460350
rect 101766 460294 101822 460350
rect 101394 460170 101450 460226
rect 101518 460170 101574 460226
rect 101642 460170 101698 460226
rect 101766 460170 101822 460226
rect 101394 460046 101450 460102
rect 101518 460046 101574 460102
rect 101642 460046 101698 460102
rect 101766 460046 101822 460102
rect 101394 459922 101450 459978
rect 101518 459922 101574 459978
rect 101642 459922 101698 459978
rect 101766 459922 101822 459978
rect 101394 442294 101450 442350
rect 101518 442294 101574 442350
rect 101642 442294 101698 442350
rect 101766 442294 101822 442350
rect 101394 442170 101450 442226
rect 101518 442170 101574 442226
rect 101642 442170 101698 442226
rect 101766 442170 101822 442226
rect 101394 442046 101450 442102
rect 101518 442046 101574 442102
rect 101642 442046 101698 442102
rect 101766 442046 101822 442102
rect 101394 441922 101450 441978
rect 101518 441922 101574 441978
rect 101642 441922 101698 441978
rect 101766 441922 101822 441978
rect 101394 424294 101450 424350
rect 101518 424294 101574 424350
rect 101642 424294 101698 424350
rect 101766 424294 101822 424350
rect 101394 424170 101450 424226
rect 101518 424170 101574 424226
rect 101642 424170 101698 424226
rect 101766 424170 101822 424226
rect 101394 424046 101450 424102
rect 101518 424046 101574 424102
rect 101642 424046 101698 424102
rect 101766 424046 101822 424102
rect 101394 423922 101450 423978
rect 101518 423922 101574 423978
rect 101642 423922 101698 423978
rect 101766 423922 101822 423978
rect 101394 406294 101450 406350
rect 101518 406294 101574 406350
rect 101642 406294 101698 406350
rect 101766 406294 101822 406350
rect 101394 406170 101450 406226
rect 101518 406170 101574 406226
rect 101642 406170 101698 406226
rect 101766 406170 101822 406226
rect 101394 406046 101450 406102
rect 101518 406046 101574 406102
rect 101642 406046 101698 406102
rect 101766 406046 101822 406102
rect 101394 405922 101450 405978
rect 101518 405922 101574 405978
rect 101642 405922 101698 405978
rect 101766 405922 101822 405978
rect 101394 388294 101450 388350
rect 101518 388294 101574 388350
rect 101642 388294 101698 388350
rect 101766 388294 101822 388350
rect 101394 388170 101450 388226
rect 101518 388170 101574 388226
rect 101642 388170 101698 388226
rect 101766 388170 101822 388226
rect 101394 388046 101450 388102
rect 101518 388046 101574 388102
rect 101642 388046 101698 388102
rect 101766 388046 101822 388102
rect 101394 387922 101450 387978
rect 101518 387922 101574 387978
rect 101642 387922 101698 387978
rect 101766 387922 101822 387978
rect 101394 370294 101450 370350
rect 101518 370294 101574 370350
rect 101642 370294 101698 370350
rect 101766 370294 101822 370350
rect 101394 370170 101450 370226
rect 101518 370170 101574 370226
rect 101642 370170 101698 370226
rect 101766 370170 101822 370226
rect 101394 370046 101450 370102
rect 101518 370046 101574 370102
rect 101642 370046 101698 370102
rect 101766 370046 101822 370102
rect 101394 369922 101450 369978
rect 101518 369922 101574 369978
rect 101642 369922 101698 369978
rect 101766 369922 101822 369978
rect 101394 352294 101450 352350
rect 101518 352294 101574 352350
rect 101642 352294 101698 352350
rect 101766 352294 101822 352350
rect 101394 352170 101450 352226
rect 101518 352170 101574 352226
rect 101642 352170 101698 352226
rect 101766 352170 101822 352226
rect 101394 352046 101450 352102
rect 101518 352046 101574 352102
rect 101642 352046 101698 352102
rect 101766 352046 101822 352102
rect 101394 351922 101450 351978
rect 101518 351922 101574 351978
rect 101642 351922 101698 351978
rect 101766 351922 101822 351978
rect 101394 334294 101450 334350
rect 101518 334294 101574 334350
rect 101642 334294 101698 334350
rect 101766 334294 101822 334350
rect 101394 334170 101450 334226
rect 101518 334170 101574 334226
rect 101642 334170 101698 334226
rect 101766 334170 101822 334226
rect 101394 334046 101450 334102
rect 101518 334046 101574 334102
rect 101642 334046 101698 334102
rect 101766 334046 101822 334102
rect 101394 333922 101450 333978
rect 101518 333922 101574 333978
rect 101642 333922 101698 333978
rect 101766 333922 101822 333978
rect 79878 316294 79934 316350
rect 80002 316294 80058 316350
rect 79878 316170 79934 316226
rect 80002 316170 80058 316226
rect 79878 316046 79934 316102
rect 80002 316046 80058 316102
rect 79878 315922 79934 315978
rect 80002 315922 80058 315978
rect 64518 310294 64574 310350
rect 64642 310294 64698 310350
rect 64518 310170 64574 310226
rect 64642 310170 64698 310226
rect 64518 310046 64574 310102
rect 64642 310046 64698 310102
rect 64518 309922 64574 309978
rect 64642 309922 64698 309978
rect 95238 310294 95294 310350
rect 95362 310294 95418 310350
rect 95238 310170 95294 310226
rect 95362 310170 95418 310226
rect 95238 310046 95294 310102
rect 95362 310046 95418 310102
rect 95238 309922 95294 309978
rect 95362 309922 95418 309978
rect 79878 298294 79934 298350
rect 80002 298294 80058 298350
rect 79878 298170 79934 298226
rect 80002 298170 80058 298226
rect 79878 298046 79934 298102
rect 80002 298046 80058 298102
rect 79878 297922 79934 297978
rect 80002 297922 80058 297978
rect 64518 292294 64574 292350
rect 64642 292294 64698 292350
rect 64518 292170 64574 292226
rect 64642 292170 64698 292226
rect 64518 292046 64574 292102
rect 64642 292046 64698 292102
rect 64518 291922 64574 291978
rect 64642 291922 64698 291978
rect 95238 292294 95294 292350
rect 95362 292294 95418 292350
rect 95238 292170 95294 292226
rect 95362 292170 95418 292226
rect 95238 292046 95294 292102
rect 95362 292046 95418 292102
rect 95238 291922 95294 291978
rect 95362 291922 95418 291978
rect 68796 287342 68852 287398
rect 63644 277082 63700 277138
rect 63868 277262 63924 277318
rect 64204 276724 64260 276778
rect 64204 276722 64260 276724
rect 63644 276182 63700 276238
rect 63420 275462 63476 275518
rect 77532 286622 77588 286678
rect 70674 280294 70730 280350
rect 70798 280294 70854 280350
rect 70922 280294 70978 280350
rect 71046 280294 71102 280350
rect 70674 280170 70730 280226
rect 70798 280170 70854 280226
rect 70922 280170 70978 280226
rect 71046 280170 71102 280226
rect 70674 280046 70730 280102
rect 70798 280046 70854 280102
rect 70922 280046 70978 280102
rect 71046 280046 71102 280102
rect 106652 286622 106708 286678
rect 106764 326042 106820 326098
rect 101394 280294 101450 280350
rect 101518 280294 101574 280350
rect 101642 280294 101698 280350
rect 101766 280294 101822 280350
rect 101394 280170 101450 280226
rect 101518 280170 101574 280226
rect 101642 280170 101698 280226
rect 101766 280170 101822 280226
rect 101394 280046 101450 280102
rect 101518 280046 101574 280102
rect 101642 280046 101698 280102
rect 101766 280046 101822 280102
rect 70674 279922 70730 279978
rect 70798 279922 70854 279978
rect 70922 279922 70978 279978
rect 71046 279922 71102 279978
rect 70364 276724 70420 276778
rect 70364 276722 70420 276724
rect 66954 274294 67010 274350
rect 67078 274294 67134 274350
rect 67202 274294 67258 274350
rect 67326 274294 67382 274350
rect 66954 274170 67010 274226
rect 67078 274170 67134 274226
rect 67202 274170 67258 274226
rect 67326 274170 67382 274226
rect 66954 274046 67010 274102
rect 67078 274046 67134 274102
rect 67202 274046 67258 274102
rect 67326 274046 67382 274102
rect 66954 273922 67010 273978
rect 67078 273922 67134 273978
rect 67202 273922 67258 273978
rect 67326 273922 67382 273978
rect 61404 260342 61460 260398
rect 66954 256294 67010 256350
rect 67078 256294 67134 256350
rect 67202 256294 67258 256350
rect 67326 256294 67382 256350
rect 66954 256170 67010 256226
rect 67078 256170 67134 256226
rect 67202 256170 67258 256226
rect 67326 256170 67382 256226
rect 66954 256046 67010 256102
rect 67078 256046 67134 256102
rect 67202 256046 67258 256102
rect 67326 256046 67382 256102
rect 66954 255922 67010 255978
rect 67078 255922 67134 255978
rect 67202 255922 67258 255978
rect 67326 255922 67382 255978
rect 66954 238294 67010 238350
rect 67078 238294 67134 238350
rect 67202 238294 67258 238350
rect 67326 238294 67382 238350
rect 66954 238170 67010 238226
rect 67078 238170 67134 238226
rect 67202 238170 67258 238226
rect 67326 238170 67382 238226
rect 66954 238046 67010 238102
rect 67078 238046 67134 238102
rect 67202 238046 67258 238102
rect 67326 238046 67382 238102
rect 66954 237922 67010 237978
rect 67078 237922 67134 237978
rect 67202 237922 67258 237978
rect 67326 237922 67382 237978
rect 66954 220294 67010 220350
rect 67078 220294 67134 220350
rect 67202 220294 67258 220350
rect 67326 220294 67382 220350
rect 66954 220170 67010 220226
rect 67078 220170 67134 220226
rect 67202 220170 67258 220226
rect 67326 220170 67382 220226
rect 66954 220046 67010 220102
rect 67078 220046 67134 220102
rect 67202 220046 67258 220102
rect 67326 220046 67382 220102
rect 66954 219922 67010 219978
rect 67078 219922 67134 219978
rect 67202 219922 67258 219978
rect 67326 219922 67382 219978
rect 66954 202294 67010 202350
rect 67078 202294 67134 202350
rect 67202 202294 67258 202350
rect 67326 202294 67382 202350
rect 66954 202170 67010 202226
rect 67078 202170 67134 202226
rect 67202 202170 67258 202226
rect 67326 202170 67382 202226
rect 66954 202046 67010 202102
rect 67078 202046 67134 202102
rect 67202 202046 67258 202102
rect 67326 202046 67382 202102
rect 66954 201922 67010 201978
rect 67078 201922 67134 201978
rect 67202 201922 67258 201978
rect 67326 201922 67382 201978
rect 66954 184294 67010 184350
rect 67078 184294 67134 184350
rect 67202 184294 67258 184350
rect 67326 184294 67382 184350
rect 66954 184170 67010 184226
rect 67078 184170 67134 184226
rect 67202 184170 67258 184226
rect 67326 184170 67382 184226
rect 66954 184046 67010 184102
rect 67078 184046 67134 184102
rect 67202 184046 67258 184102
rect 67326 184046 67382 184102
rect 66954 183922 67010 183978
rect 67078 183922 67134 183978
rect 67202 183922 67258 183978
rect 67326 183922 67382 183978
rect 66954 166294 67010 166350
rect 67078 166294 67134 166350
rect 67202 166294 67258 166350
rect 67326 166294 67382 166350
rect 66954 166170 67010 166226
rect 67078 166170 67134 166226
rect 67202 166170 67258 166226
rect 67326 166170 67382 166226
rect 66954 166046 67010 166102
rect 67078 166046 67134 166102
rect 67202 166046 67258 166102
rect 67326 166046 67382 166102
rect 66954 165922 67010 165978
rect 67078 165922 67134 165978
rect 67202 165922 67258 165978
rect 67326 165922 67382 165978
rect 39954 136294 40010 136350
rect 40078 136294 40134 136350
rect 40202 136294 40258 136350
rect 40326 136294 40382 136350
rect 39954 136170 40010 136226
rect 40078 136170 40134 136226
rect 40202 136170 40258 136226
rect 40326 136170 40382 136226
rect 39954 136046 40010 136102
rect 40078 136046 40134 136102
rect 40202 136046 40258 136102
rect 40326 136046 40382 136102
rect 39954 135922 40010 135978
rect 40078 135922 40134 135978
rect 40202 135922 40258 135978
rect 40326 135922 40382 135978
rect 39954 118294 40010 118350
rect 40078 118294 40134 118350
rect 40202 118294 40258 118350
rect 40326 118294 40382 118350
rect 39954 118170 40010 118226
rect 40078 118170 40134 118226
rect 40202 118170 40258 118226
rect 40326 118170 40382 118226
rect 39954 118046 40010 118102
rect 40078 118046 40134 118102
rect 40202 118046 40258 118102
rect 40326 118046 40382 118102
rect 39954 117922 40010 117978
rect 40078 117922 40134 117978
rect 40202 117922 40258 117978
rect 40326 117922 40382 117978
rect 39954 100294 40010 100350
rect 40078 100294 40134 100350
rect 40202 100294 40258 100350
rect 40326 100294 40382 100350
rect 39954 100170 40010 100226
rect 40078 100170 40134 100226
rect 40202 100170 40258 100226
rect 40326 100170 40382 100226
rect 39954 100046 40010 100102
rect 40078 100046 40134 100102
rect 40202 100046 40258 100102
rect 40326 100046 40382 100102
rect 39954 99922 40010 99978
rect 40078 99922 40134 99978
rect 40202 99922 40258 99978
rect 40326 99922 40382 99978
rect 39954 82294 40010 82350
rect 40078 82294 40134 82350
rect 40202 82294 40258 82350
rect 40326 82294 40382 82350
rect 39954 82170 40010 82226
rect 40078 82170 40134 82226
rect 40202 82170 40258 82226
rect 40326 82170 40382 82226
rect 39954 82046 40010 82102
rect 40078 82046 40134 82102
rect 40202 82046 40258 82102
rect 40326 82046 40382 82102
rect 39954 81922 40010 81978
rect 40078 81922 40134 81978
rect 40202 81922 40258 81978
rect 40326 81922 40382 81978
rect 39954 64294 40010 64350
rect 40078 64294 40134 64350
rect 40202 64294 40258 64350
rect 40326 64294 40382 64350
rect 39954 64170 40010 64226
rect 40078 64170 40134 64226
rect 40202 64170 40258 64226
rect 40326 64170 40382 64226
rect 39954 64046 40010 64102
rect 40078 64046 40134 64102
rect 40202 64046 40258 64102
rect 40326 64046 40382 64102
rect 39954 63922 40010 63978
rect 40078 63922 40134 63978
rect 40202 63922 40258 63978
rect 40326 63922 40382 63978
rect 39954 46294 40010 46350
rect 40078 46294 40134 46350
rect 40202 46294 40258 46350
rect 40326 46294 40382 46350
rect 39954 46170 40010 46226
rect 40078 46170 40134 46226
rect 40202 46170 40258 46226
rect 40326 46170 40382 46226
rect 39954 46046 40010 46102
rect 40078 46046 40134 46102
rect 40202 46046 40258 46102
rect 40326 46046 40382 46102
rect 39954 45922 40010 45978
rect 40078 45922 40134 45978
rect 40202 45922 40258 45978
rect 40326 45922 40382 45978
rect 39954 28294 40010 28350
rect 40078 28294 40134 28350
rect 40202 28294 40258 28350
rect 40326 28294 40382 28350
rect 39954 28170 40010 28226
rect 40078 28170 40134 28226
rect 40202 28170 40258 28226
rect 40326 28170 40382 28226
rect 39954 28046 40010 28102
rect 40078 28046 40134 28102
rect 40202 28046 40258 28102
rect 40326 28046 40382 28102
rect 39954 27922 40010 27978
rect 40078 27922 40134 27978
rect 40202 27922 40258 27978
rect 40326 27922 40382 27978
rect 39954 10294 40010 10350
rect 40078 10294 40134 10350
rect 40202 10294 40258 10350
rect 40326 10294 40382 10350
rect 39954 10170 40010 10226
rect 40078 10170 40134 10226
rect 40202 10170 40258 10226
rect 40326 10170 40382 10226
rect 39954 10046 40010 10102
rect 40078 10046 40134 10102
rect 40202 10046 40258 10102
rect 40326 10046 40382 10102
rect 39954 9922 40010 9978
rect 40078 9922 40134 9978
rect 40202 9922 40258 9978
rect 40326 9922 40382 9978
rect 39954 -1176 40010 -1120
rect 40078 -1176 40134 -1120
rect 40202 -1176 40258 -1120
rect 40326 -1176 40382 -1120
rect 39954 -1300 40010 -1244
rect 40078 -1300 40134 -1244
rect 40202 -1300 40258 -1244
rect 40326 -1300 40382 -1244
rect 39954 -1424 40010 -1368
rect 40078 -1424 40134 -1368
rect 40202 -1424 40258 -1368
rect 40326 -1424 40382 -1368
rect 39954 -1548 40010 -1492
rect 40078 -1548 40134 -1492
rect 40202 -1548 40258 -1492
rect 40326 -1548 40382 -1492
rect 69692 276182 69748 276238
rect 70364 276002 70420 276058
rect 70364 271322 70420 271378
rect 101394 279922 101450 279978
rect 101518 279922 101574 279978
rect 101642 279922 101698 279978
rect 101766 279922 101822 279978
rect 74172 278162 74228 278218
rect 73052 276902 73108 276958
rect 70674 262294 70730 262350
rect 70798 262294 70854 262350
rect 70922 262294 70978 262350
rect 71046 262294 71102 262350
rect 70674 262170 70730 262226
rect 70798 262170 70854 262226
rect 70922 262170 70978 262226
rect 71046 262170 71102 262226
rect 70674 262046 70730 262102
rect 70798 262046 70854 262102
rect 70922 262046 70978 262102
rect 71046 262046 71102 262102
rect 70674 261922 70730 261978
rect 70798 261922 70854 261978
rect 70922 261922 70978 261978
rect 71046 261922 71102 261978
rect 70674 244294 70730 244350
rect 70798 244294 70854 244350
rect 70922 244294 70978 244350
rect 71046 244294 71102 244350
rect 70674 244170 70730 244226
rect 70798 244170 70854 244226
rect 70922 244170 70978 244226
rect 71046 244170 71102 244226
rect 70674 244046 70730 244102
rect 70798 244046 70854 244102
rect 70922 244046 70978 244102
rect 71046 244046 71102 244102
rect 70674 243922 70730 243978
rect 70798 243922 70854 243978
rect 70922 243922 70978 243978
rect 71046 243922 71102 243978
rect 70674 226294 70730 226350
rect 70798 226294 70854 226350
rect 70922 226294 70978 226350
rect 71046 226294 71102 226350
rect 70674 226170 70730 226226
rect 70798 226170 70854 226226
rect 70922 226170 70978 226226
rect 71046 226170 71102 226226
rect 70674 226046 70730 226102
rect 70798 226046 70854 226102
rect 70922 226046 70978 226102
rect 71046 226046 71102 226102
rect 70674 225922 70730 225978
rect 70798 225922 70854 225978
rect 70922 225922 70978 225978
rect 71046 225922 71102 225978
rect 70674 208294 70730 208350
rect 70798 208294 70854 208350
rect 70922 208294 70978 208350
rect 71046 208294 71102 208350
rect 70674 208170 70730 208226
rect 70798 208170 70854 208226
rect 70922 208170 70978 208226
rect 71046 208170 71102 208226
rect 70674 208046 70730 208102
rect 70798 208046 70854 208102
rect 70922 208046 70978 208102
rect 71046 208046 71102 208102
rect 70674 207922 70730 207978
rect 70798 207922 70854 207978
rect 70922 207922 70978 207978
rect 71046 207922 71102 207978
rect 70674 190294 70730 190350
rect 70798 190294 70854 190350
rect 70922 190294 70978 190350
rect 71046 190294 71102 190350
rect 70674 190170 70730 190226
rect 70798 190170 70854 190226
rect 70922 190170 70978 190226
rect 71046 190170 71102 190226
rect 70674 190046 70730 190102
rect 70798 190046 70854 190102
rect 70922 190046 70978 190102
rect 71046 190046 71102 190102
rect 70674 189922 70730 189978
rect 70798 189922 70854 189978
rect 70922 189922 70978 189978
rect 71046 189922 71102 189978
rect 70674 172294 70730 172350
rect 70798 172294 70854 172350
rect 70922 172294 70978 172350
rect 71046 172294 71102 172350
rect 70674 172170 70730 172226
rect 70798 172170 70854 172226
rect 70922 172170 70978 172226
rect 71046 172170 71102 172226
rect 70674 172046 70730 172102
rect 70798 172046 70854 172102
rect 70922 172046 70978 172102
rect 71046 172046 71102 172102
rect 70674 171922 70730 171978
rect 70798 171922 70854 171978
rect 70922 171922 70978 171978
rect 71046 171922 71102 171978
rect 72156 195722 72212 195778
rect 74732 276362 74788 276418
rect 70674 154294 70730 154350
rect 70798 154294 70854 154350
rect 70922 154294 70978 154350
rect 71046 154294 71102 154350
rect 70674 154170 70730 154226
rect 70798 154170 70854 154226
rect 70922 154170 70978 154226
rect 71046 154170 71102 154226
rect 70674 154046 70730 154102
rect 70798 154046 70854 154102
rect 70922 154046 70978 154102
rect 71046 154046 71102 154102
rect 70674 153922 70730 153978
rect 70798 153922 70854 153978
rect 70922 153922 70978 153978
rect 71046 153922 71102 153978
rect 66954 148294 67010 148350
rect 67078 148294 67134 148350
rect 67202 148294 67258 148350
rect 67326 148294 67382 148350
rect 66954 148170 67010 148226
rect 67078 148170 67134 148226
rect 67202 148170 67258 148226
rect 67326 148170 67382 148226
rect 66954 148046 67010 148102
rect 67078 148046 67134 148102
rect 67202 148046 67258 148102
rect 67326 148046 67382 148102
rect 66954 147922 67010 147978
rect 67078 147922 67134 147978
rect 67202 147922 67258 147978
rect 67326 147922 67382 147978
rect 66954 130294 67010 130350
rect 67078 130294 67134 130350
rect 67202 130294 67258 130350
rect 67326 130294 67382 130350
rect 66954 130170 67010 130226
rect 67078 130170 67134 130226
rect 67202 130170 67258 130226
rect 67326 130170 67382 130226
rect 66954 130046 67010 130102
rect 67078 130046 67134 130102
rect 67202 130046 67258 130102
rect 67326 130046 67382 130102
rect 66954 129922 67010 129978
rect 67078 129922 67134 129978
rect 67202 129922 67258 129978
rect 67326 129922 67382 129978
rect 66954 112294 67010 112350
rect 67078 112294 67134 112350
rect 67202 112294 67258 112350
rect 67326 112294 67382 112350
rect 66954 112170 67010 112226
rect 67078 112170 67134 112226
rect 67202 112170 67258 112226
rect 67326 112170 67382 112226
rect 66954 112046 67010 112102
rect 67078 112046 67134 112102
rect 67202 112046 67258 112102
rect 67326 112046 67382 112102
rect 66954 111922 67010 111978
rect 67078 111922 67134 111978
rect 67202 111922 67258 111978
rect 67326 111922 67382 111978
rect 66954 94294 67010 94350
rect 67078 94294 67134 94350
rect 67202 94294 67258 94350
rect 67326 94294 67382 94350
rect 66954 94170 67010 94226
rect 67078 94170 67134 94226
rect 67202 94170 67258 94226
rect 67326 94170 67382 94226
rect 66954 94046 67010 94102
rect 67078 94046 67134 94102
rect 67202 94046 67258 94102
rect 67326 94046 67382 94102
rect 66954 93922 67010 93978
rect 67078 93922 67134 93978
rect 67202 93922 67258 93978
rect 67326 93922 67382 93978
rect 66954 76294 67010 76350
rect 67078 76294 67134 76350
rect 67202 76294 67258 76350
rect 67326 76294 67382 76350
rect 66954 76170 67010 76226
rect 67078 76170 67134 76226
rect 67202 76170 67258 76226
rect 67326 76170 67382 76226
rect 66954 76046 67010 76102
rect 67078 76046 67134 76102
rect 67202 76046 67258 76102
rect 67326 76046 67382 76102
rect 66954 75922 67010 75978
rect 67078 75922 67134 75978
rect 67202 75922 67258 75978
rect 67326 75922 67382 75978
rect 66954 58294 67010 58350
rect 67078 58294 67134 58350
rect 67202 58294 67258 58350
rect 67326 58294 67382 58350
rect 66954 58170 67010 58226
rect 67078 58170 67134 58226
rect 67202 58170 67258 58226
rect 67326 58170 67382 58226
rect 66954 58046 67010 58102
rect 67078 58046 67134 58102
rect 67202 58046 67258 58102
rect 67326 58046 67382 58102
rect 66954 57922 67010 57978
rect 67078 57922 67134 57978
rect 67202 57922 67258 57978
rect 67326 57922 67382 57978
rect 66954 40294 67010 40350
rect 67078 40294 67134 40350
rect 67202 40294 67258 40350
rect 67326 40294 67382 40350
rect 66954 40170 67010 40226
rect 67078 40170 67134 40226
rect 67202 40170 67258 40226
rect 67326 40170 67382 40226
rect 66954 40046 67010 40102
rect 67078 40046 67134 40102
rect 67202 40046 67258 40102
rect 67326 40046 67382 40102
rect 66954 39922 67010 39978
rect 67078 39922 67134 39978
rect 67202 39922 67258 39978
rect 67326 39922 67382 39978
rect 66954 22294 67010 22350
rect 67078 22294 67134 22350
rect 67202 22294 67258 22350
rect 67326 22294 67382 22350
rect 66954 22170 67010 22226
rect 67078 22170 67134 22226
rect 67202 22170 67258 22226
rect 67326 22170 67382 22226
rect 66954 22046 67010 22102
rect 67078 22046 67134 22102
rect 67202 22046 67258 22102
rect 67326 22046 67382 22102
rect 66954 21922 67010 21978
rect 67078 21922 67134 21978
rect 67202 21922 67258 21978
rect 67326 21922 67382 21978
rect 66954 4294 67010 4350
rect 67078 4294 67134 4350
rect 67202 4294 67258 4350
rect 67326 4294 67382 4350
rect 66954 4170 67010 4226
rect 67078 4170 67134 4226
rect 67202 4170 67258 4226
rect 67326 4170 67382 4226
rect 66954 4046 67010 4102
rect 67078 4046 67134 4102
rect 67202 4046 67258 4102
rect 67326 4046 67382 4102
rect 66954 3922 67010 3978
rect 67078 3922 67134 3978
rect 67202 3922 67258 3978
rect 67326 3922 67382 3978
rect 66954 -216 67010 -160
rect 67078 -216 67134 -160
rect 67202 -216 67258 -160
rect 67326 -216 67382 -160
rect 66954 -340 67010 -284
rect 67078 -340 67134 -284
rect 67202 -340 67258 -284
rect 67326 -340 67382 -284
rect 66954 -464 67010 -408
rect 67078 -464 67134 -408
rect 67202 -464 67258 -408
rect 67326 -464 67382 -408
rect 66954 -588 67010 -532
rect 67078 -588 67134 -532
rect 67202 -588 67258 -532
rect 67326 -588 67382 -532
rect 72044 149462 72100 149518
rect 82236 198962 82292 199018
rect 81452 149282 81508 149338
rect 84812 201482 84868 201538
rect 98442 256294 98498 256350
rect 98566 256294 98622 256350
rect 98690 256294 98746 256350
rect 98814 256294 98870 256350
rect 98442 256170 98498 256226
rect 98566 256170 98622 256226
rect 98690 256170 98746 256226
rect 98814 256170 98870 256226
rect 98442 256046 98498 256102
rect 98566 256046 98622 256102
rect 98690 256046 98746 256102
rect 98814 256046 98870 256102
rect 98442 255922 98498 255978
rect 98566 255922 98622 255978
rect 98690 255922 98746 255978
rect 98814 255922 98870 255978
rect 97642 244294 97698 244350
rect 97766 244294 97822 244350
rect 97890 244294 97946 244350
rect 98014 244294 98070 244350
rect 97642 244170 97698 244226
rect 97766 244170 97822 244226
rect 97890 244170 97946 244226
rect 98014 244170 98070 244226
rect 97642 244046 97698 244102
rect 97766 244046 97822 244102
rect 97890 244046 97946 244102
rect 98014 244046 98070 244102
rect 97642 243922 97698 243978
rect 97766 243922 97822 243978
rect 97890 243922 97946 243978
rect 98014 243922 98070 243978
rect 98442 238294 98498 238350
rect 98566 238294 98622 238350
rect 98690 238294 98746 238350
rect 98814 238294 98870 238350
rect 98442 238170 98498 238226
rect 98566 238170 98622 238226
rect 98690 238170 98746 238226
rect 98814 238170 98870 238226
rect 98442 238046 98498 238102
rect 98566 238046 98622 238102
rect 98690 238046 98746 238102
rect 98814 238046 98870 238102
rect 98442 237922 98498 237978
rect 98566 237922 98622 237978
rect 98690 237922 98746 237978
rect 98814 237922 98870 237978
rect 97642 226294 97698 226350
rect 97766 226294 97822 226350
rect 97890 226294 97946 226350
rect 98014 226294 98070 226350
rect 97642 226170 97698 226226
rect 97766 226170 97822 226226
rect 97890 226170 97946 226226
rect 98014 226170 98070 226226
rect 97642 226046 97698 226102
rect 97766 226046 97822 226102
rect 97890 226046 97946 226102
rect 98014 226046 98070 226102
rect 97642 225922 97698 225978
rect 97766 225922 97822 225978
rect 97890 225922 97946 225978
rect 98014 225922 98070 225978
rect 98442 220294 98498 220350
rect 98566 220294 98622 220350
rect 98690 220294 98746 220350
rect 98814 220294 98870 220350
rect 98442 220170 98498 220226
rect 98566 220170 98622 220226
rect 98690 220170 98746 220226
rect 98814 220170 98870 220226
rect 98442 220046 98498 220102
rect 98566 220046 98622 220102
rect 98690 220046 98746 220102
rect 98814 220046 98870 220102
rect 98442 219922 98498 219978
rect 98566 219922 98622 219978
rect 98690 219922 98746 219978
rect 98814 219922 98870 219978
rect 97642 208294 97698 208350
rect 97766 208294 97822 208350
rect 97890 208294 97946 208350
rect 98014 208294 98070 208350
rect 97642 208170 97698 208226
rect 97766 208170 97822 208226
rect 97890 208170 97946 208226
rect 98014 208170 98070 208226
rect 97642 208046 97698 208102
rect 97766 208046 97822 208102
rect 97890 208046 97946 208102
rect 98014 208046 98070 208102
rect 97642 207922 97698 207978
rect 97766 207922 97822 207978
rect 97890 207922 97946 207978
rect 98014 207922 98070 207978
rect 94892 204902 94948 204958
rect 98442 202294 98498 202350
rect 98566 202294 98622 202350
rect 98690 202294 98746 202350
rect 98814 202294 98870 202350
rect 98442 202170 98498 202226
rect 98566 202170 98622 202226
rect 98690 202170 98746 202226
rect 98814 202170 98870 202226
rect 98442 202046 98498 202102
rect 98566 202046 98622 202102
rect 98690 202046 98746 202102
rect 98814 202046 98870 202102
rect 98442 201922 98498 201978
rect 98566 201922 98622 201978
rect 98690 201922 98746 201978
rect 98814 201922 98870 201978
rect 97642 190294 97698 190350
rect 97766 190294 97822 190350
rect 97890 190294 97946 190350
rect 98014 190294 98070 190350
rect 97642 190170 97698 190226
rect 97766 190170 97822 190226
rect 97890 190170 97946 190226
rect 98014 190170 98070 190226
rect 97642 190046 97698 190102
rect 97766 190046 97822 190102
rect 97890 190046 97946 190102
rect 98014 190046 98070 190102
rect 97642 189922 97698 189978
rect 97766 189922 97822 189978
rect 97890 189922 97946 189978
rect 98014 189922 98070 189978
rect 98442 184294 98498 184350
rect 98566 184294 98622 184350
rect 98690 184294 98746 184350
rect 98814 184294 98870 184350
rect 98442 184170 98498 184226
rect 98566 184170 98622 184226
rect 98690 184170 98746 184226
rect 98814 184170 98870 184226
rect 98442 184046 98498 184102
rect 98566 184046 98622 184102
rect 98690 184046 98746 184102
rect 98814 184046 98870 184102
rect 98442 183922 98498 183978
rect 98566 183922 98622 183978
rect 98690 183922 98746 183978
rect 98814 183922 98870 183978
rect 100044 178802 100100 178858
rect 106652 279602 106708 279658
rect 101394 262294 101450 262350
rect 101518 262294 101574 262350
rect 101642 262294 101698 262350
rect 101766 262294 101822 262350
rect 101394 262170 101450 262226
rect 101518 262170 101574 262226
rect 101642 262170 101698 262226
rect 101766 262170 101822 262226
rect 101394 262046 101450 262102
rect 101518 262046 101574 262102
rect 101642 262046 101698 262102
rect 101766 262046 101822 262102
rect 101394 261922 101450 261978
rect 101518 261922 101574 261978
rect 101642 261922 101698 261978
rect 101766 261922 101822 261978
rect 101394 244294 101450 244350
rect 101518 244294 101574 244350
rect 101642 244294 101698 244350
rect 101766 244294 101822 244350
rect 101394 244170 101450 244226
rect 101518 244170 101574 244226
rect 101642 244170 101698 244226
rect 101766 244170 101822 244226
rect 101394 244046 101450 244102
rect 101518 244046 101574 244102
rect 101642 244046 101698 244102
rect 101766 244046 101822 244102
rect 101394 243922 101450 243978
rect 101518 243922 101574 243978
rect 101642 243922 101698 243978
rect 101766 243922 101822 243978
rect 101394 226294 101450 226350
rect 101518 226294 101574 226350
rect 101642 226294 101698 226350
rect 101766 226294 101822 226350
rect 101394 226170 101450 226226
rect 101518 226170 101574 226226
rect 101642 226170 101698 226226
rect 101766 226170 101822 226226
rect 101394 226046 101450 226102
rect 101518 226046 101574 226102
rect 101642 226046 101698 226102
rect 101766 226046 101822 226102
rect 101394 225922 101450 225978
rect 101518 225922 101574 225978
rect 101642 225922 101698 225978
rect 101766 225922 101822 225978
rect 101394 208294 101450 208350
rect 101518 208294 101574 208350
rect 101642 208294 101698 208350
rect 101766 208294 101822 208350
rect 101394 208170 101450 208226
rect 101518 208170 101574 208226
rect 101642 208170 101698 208226
rect 101766 208170 101822 208226
rect 101394 208046 101450 208102
rect 101518 208046 101574 208102
rect 101642 208046 101698 208102
rect 101766 208046 101822 208102
rect 101394 207922 101450 207978
rect 101518 207922 101574 207978
rect 101642 207922 101698 207978
rect 101766 207922 101822 207978
rect 101394 190294 101450 190350
rect 101518 190294 101574 190350
rect 101642 190294 101698 190350
rect 101766 190294 101822 190350
rect 101394 190170 101450 190226
rect 101518 190170 101574 190226
rect 101642 190170 101698 190226
rect 101766 190170 101822 190226
rect 101394 190046 101450 190102
rect 101518 190046 101574 190102
rect 101642 190046 101698 190102
rect 101766 190046 101822 190102
rect 101394 189922 101450 189978
rect 101518 189922 101574 189978
rect 101642 189922 101698 189978
rect 101766 189922 101822 189978
rect 99932 173762 99988 173818
rect 97642 172294 97698 172350
rect 97766 172294 97822 172350
rect 97890 172294 97946 172350
rect 98014 172294 98070 172350
rect 97642 172170 97698 172226
rect 97766 172170 97822 172226
rect 97890 172170 97946 172226
rect 98014 172170 98070 172226
rect 97642 172046 97698 172102
rect 97766 172046 97822 172102
rect 97890 172046 97946 172102
rect 98014 172046 98070 172102
rect 97642 171922 97698 171978
rect 97766 171922 97822 171978
rect 97890 171922 97946 171978
rect 98014 171922 98070 171978
rect 101394 172294 101450 172350
rect 101518 172294 101574 172350
rect 101642 172294 101698 172350
rect 101766 172294 101822 172350
rect 101394 172170 101450 172226
rect 101518 172170 101574 172226
rect 101642 172170 101698 172226
rect 101766 172170 101822 172226
rect 101394 172046 101450 172102
rect 101518 172046 101574 172102
rect 101642 172046 101698 172102
rect 101766 172046 101822 172102
rect 101394 171922 101450 171978
rect 101518 171922 101574 171978
rect 101642 171922 101698 171978
rect 101766 171922 101822 171978
rect 97674 166294 97730 166350
rect 97798 166294 97854 166350
rect 97922 166294 97978 166350
rect 98046 166294 98102 166350
rect 97674 166170 97730 166226
rect 97798 166170 97854 166226
rect 97922 166170 97978 166226
rect 98046 166170 98102 166226
rect 97674 166046 97730 166102
rect 97798 166046 97854 166102
rect 97922 166046 97978 166102
rect 98046 166046 98102 166102
rect 97674 165922 97730 165978
rect 97798 165922 97854 165978
rect 97922 165922 97978 165978
rect 98046 165922 98102 165978
rect 97674 148294 97730 148350
rect 97798 148294 97854 148350
rect 97922 148294 97978 148350
rect 98046 148294 98102 148350
rect 97674 148170 97730 148226
rect 97798 148170 97854 148226
rect 97922 148170 97978 148226
rect 98046 148170 98102 148226
rect 97674 148046 97730 148102
rect 97798 148046 97854 148102
rect 97922 148046 97978 148102
rect 98046 148046 98102 148102
rect 97674 147922 97730 147978
rect 97798 147922 97854 147978
rect 97922 147922 97978 147978
rect 98046 147922 98102 147978
rect 70674 136294 70730 136350
rect 70798 136294 70854 136350
rect 70922 136294 70978 136350
rect 71046 136294 71102 136350
rect 70674 136170 70730 136226
rect 70798 136170 70854 136226
rect 70922 136170 70978 136226
rect 71046 136170 71102 136226
rect 70674 136046 70730 136102
rect 70798 136046 70854 136102
rect 70922 136046 70978 136102
rect 71046 136046 71102 136102
rect 70674 135922 70730 135978
rect 70798 135922 70854 135978
rect 70922 135922 70978 135978
rect 71046 135922 71102 135978
rect 96612 136294 96668 136350
rect 96736 136294 96792 136350
rect 96860 136294 96916 136350
rect 96984 136294 97040 136350
rect 96612 136170 96668 136226
rect 96736 136170 96792 136226
rect 96860 136170 96916 136226
rect 96984 136170 97040 136226
rect 96612 136046 96668 136102
rect 96736 136046 96792 136102
rect 96860 136046 96916 136102
rect 96984 136046 97040 136102
rect 96612 135922 96668 135978
rect 96736 135922 96792 135978
rect 96860 135922 96916 135978
rect 96984 135922 97040 135978
rect 95812 130294 95868 130350
rect 95936 130294 95992 130350
rect 96060 130294 96116 130350
rect 96184 130294 96240 130350
rect 95812 130170 95868 130226
rect 95936 130170 95992 130226
rect 96060 130170 96116 130226
rect 96184 130170 96240 130226
rect 95812 130046 95868 130102
rect 95936 130046 95992 130102
rect 96060 130046 96116 130102
rect 96184 130046 96240 130102
rect 95812 129922 95868 129978
rect 95936 129922 95992 129978
rect 96060 129922 96116 129978
rect 96184 129922 96240 129978
rect 97674 130294 97730 130350
rect 97798 130294 97854 130350
rect 97922 130294 97978 130350
rect 98046 130294 98102 130350
rect 97674 130170 97730 130226
rect 97798 130170 97854 130226
rect 97922 130170 97978 130226
rect 98046 130170 98102 130226
rect 97674 130046 97730 130102
rect 97798 130046 97854 130102
rect 97922 130046 97978 130102
rect 98046 130046 98102 130102
rect 97674 129922 97730 129978
rect 97798 129922 97854 129978
rect 97922 129922 97978 129978
rect 98046 129922 98102 129978
rect 70674 118294 70730 118350
rect 70798 118294 70854 118350
rect 70922 118294 70978 118350
rect 71046 118294 71102 118350
rect 70674 118170 70730 118226
rect 70798 118170 70854 118226
rect 70922 118170 70978 118226
rect 71046 118170 71102 118226
rect 70674 118046 70730 118102
rect 70798 118046 70854 118102
rect 70922 118046 70978 118102
rect 71046 118046 71102 118102
rect 70674 117922 70730 117978
rect 70798 117922 70854 117978
rect 70922 117922 70978 117978
rect 71046 117922 71102 117978
rect 96612 118294 96668 118350
rect 96736 118294 96792 118350
rect 96860 118294 96916 118350
rect 96984 118294 97040 118350
rect 96612 118170 96668 118226
rect 96736 118170 96792 118226
rect 96860 118170 96916 118226
rect 96984 118170 97040 118226
rect 96612 118046 96668 118102
rect 96736 118046 96792 118102
rect 96860 118046 96916 118102
rect 96984 118046 97040 118102
rect 96612 117922 96668 117978
rect 96736 117922 96792 117978
rect 96860 117922 96916 117978
rect 96984 117922 97040 117978
rect 95812 112294 95868 112350
rect 95936 112294 95992 112350
rect 96060 112294 96116 112350
rect 96184 112294 96240 112350
rect 95812 112170 95868 112226
rect 95936 112170 95992 112226
rect 96060 112170 96116 112226
rect 96184 112170 96240 112226
rect 95812 112046 95868 112102
rect 95936 112046 95992 112102
rect 96060 112046 96116 112102
rect 96184 112046 96240 112102
rect 95812 111922 95868 111978
rect 95936 111922 95992 111978
rect 96060 111922 96116 111978
rect 96184 111922 96240 111978
rect 97674 112294 97730 112350
rect 97798 112294 97854 112350
rect 97922 112294 97978 112350
rect 98046 112294 98102 112350
rect 97674 112170 97730 112226
rect 97798 112170 97854 112226
rect 97922 112170 97978 112226
rect 98046 112170 98102 112226
rect 97674 112046 97730 112102
rect 97798 112046 97854 112102
rect 97922 112046 97978 112102
rect 98046 112046 98102 112102
rect 97674 111922 97730 111978
rect 97798 111922 97854 111978
rect 97922 111922 97978 111978
rect 98046 111922 98102 111978
rect 70674 100294 70730 100350
rect 70798 100294 70854 100350
rect 70922 100294 70978 100350
rect 71046 100294 71102 100350
rect 70674 100170 70730 100226
rect 70798 100170 70854 100226
rect 70922 100170 70978 100226
rect 71046 100170 71102 100226
rect 70674 100046 70730 100102
rect 70798 100046 70854 100102
rect 70922 100046 70978 100102
rect 71046 100046 71102 100102
rect 70674 99922 70730 99978
rect 70798 99922 70854 99978
rect 70922 99922 70978 99978
rect 71046 99922 71102 99978
rect 96612 100294 96668 100350
rect 96736 100294 96792 100350
rect 96860 100294 96916 100350
rect 96984 100294 97040 100350
rect 96612 100170 96668 100226
rect 96736 100170 96792 100226
rect 96860 100170 96916 100226
rect 96984 100170 97040 100226
rect 96612 100046 96668 100102
rect 96736 100046 96792 100102
rect 96860 100046 96916 100102
rect 96984 100046 97040 100102
rect 96612 99922 96668 99978
rect 96736 99922 96792 99978
rect 96860 99922 96916 99978
rect 96984 99922 97040 99978
rect 95812 94294 95868 94350
rect 95936 94294 95992 94350
rect 96060 94294 96116 94350
rect 96184 94294 96240 94350
rect 95812 94170 95868 94226
rect 95936 94170 95992 94226
rect 96060 94170 96116 94226
rect 96184 94170 96240 94226
rect 95812 94046 95868 94102
rect 95936 94046 95992 94102
rect 96060 94046 96116 94102
rect 96184 94046 96240 94102
rect 95812 93922 95868 93978
rect 95936 93922 95992 93978
rect 96060 93922 96116 93978
rect 96184 93922 96240 93978
rect 97674 94294 97730 94350
rect 97798 94294 97854 94350
rect 97922 94294 97978 94350
rect 98046 94294 98102 94350
rect 97674 94170 97730 94226
rect 97798 94170 97854 94226
rect 97922 94170 97978 94226
rect 98046 94170 98102 94226
rect 97674 94046 97730 94102
rect 97798 94046 97854 94102
rect 97922 94046 97978 94102
rect 98046 94046 98102 94102
rect 97674 93922 97730 93978
rect 97798 93922 97854 93978
rect 97922 93922 97978 93978
rect 98046 93922 98102 93978
rect 70674 82294 70730 82350
rect 70798 82294 70854 82350
rect 70922 82294 70978 82350
rect 71046 82294 71102 82350
rect 70674 82170 70730 82226
rect 70798 82170 70854 82226
rect 70922 82170 70978 82226
rect 71046 82170 71102 82226
rect 70674 82046 70730 82102
rect 70798 82046 70854 82102
rect 70922 82046 70978 82102
rect 71046 82046 71102 82102
rect 70674 81922 70730 81978
rect 70798 81922 70854 81978
rect 70922 81922 70978 81978
rect 71046 81922 71102 81978
rect 96612 82294 96668 82350
rect 96736 82294 96792 82350
rect 96860 82294 96916 82350
rect 96984 82294 97040 82350
rect 96612 82170 96668 82226
rect 96736 82170 96792 82226
rect 96860 82170 96916 82226
rect 96984 82170 97040 82226
rect 96612 82046 96668 82102
rect 96736 82046 96792 82102
rect 96860 82046 96916 82102
rect 96984 82046 97040 82102
rect 96612 81922 96668 81978
rect 96736 81922 96792 81978
rect 96860 81922 96916 81978
rect 96984 81922 97040 81978
rect 95812 76294 95868 76350
rect 95936 76294 95992 76350
rect 96060 76294 96116 76350
rect 96184 76294 96240 76350
rect 95812 76170 95868 76226
rect 95936 76170 95992 76226
rect 96060 76170 96116 76226
rect 96184 76170 96240 76226
rect 95812 76046 95868 76102
rect 95936 76046 95992 76102
rect 96060 76046 96116 76102
rect 96184 76046 96240 76102
rect 95812 75922 95868 75978
rect 95936 75922 95992 75978
rect 96060 75922 96116 75978
rect 96184 75922 96240 75978
rect 97674 76294 97730 76350
rect 97798 76294 97854 76350
rect 97922 76294 97978 76350
rect 98046 76294 98102 76350
rect 97674 76170 97730 76226
rect 97798 76170 97854 76226
rect 97922 76170 97978 76226
rect 98046 76170 98102 76226
rect 97674 76046 97730 76102
rect 97798 76046 97854 76102
rect 97922 76046 97978 76102
rect 98046 76046 98102 76102
rect 97674 75922 97730 75978
rect 97798 75922 97854 75978
rect 97922 75922 97978 75978
rect 98046 75922 98102 75978
rect 70674 64294 70730 64350
rect 70798 64294 70854 64350
rect 70922 64294 70978 64350
rect 71046 64294 71102 64350
rect 70674 64170 70730 64226
rect 70798 64170 70854 64226
rect 70922 64170 70978 64226
rect 71046 64170 71102 64226
rect 70674 64046 70730 64102
rect 70798 64046 70854 64102
rect 70922 64046 70978 64102
rect 71046 64046 71102 64102
rect 70674 63922 70730 63978
rect 70798 63922 70854 63978
rect 70922 63922 70978 63978
rect 71046 63922 71102 63978
rect 96612 64294 96668 64350
rect 96736 64294 96792 64350
rect 96860 64294 96916 64350
rect 96984 64294 97040 64350
rect 96612 64170 96668 64226
rect 96736 64170 96792 64226
rect 96860 64170 96916 64226
rect 96984 64170 97040 64226
rect 96612 64046 96668 64102
rect 96736 64046 96792 64102
rect 96860 64046 96916 64102
rect 96984 64046 97040 64102
rect 96612 63922 96668 63978
rect 96736 63922 96792 63978
rect 96860 63922 96916 63978
rect 96984 63922 97040 63978
rect 95812 58294 95868 58350
rect 95936 58294 95992 58350
rect 96060 58294 96116 58350
rect 96184 58294 96240 58350
rect 95812 58170 95868 58226
rect 95936 58170 95992 58226
rect 96060 58170 96116 58226
rect 96184 58170 96240 58226
rect 95812 58046 95868 58102
rect 95936 58046 95992 58102
rect 96060 58046 96116 58102
rect 96184 58046 96240 58102
rect 95812 57922 95868 57978
rect 95936 57922 95992 57978
rect 96060 57922 96116 57978
rect 96184 57922 96240 57978
rect 97674 58294 97730 58350
rect 97798 58294 97854 58350
rect 97922 58294 97978 58350
rect 98046 58294 98102 58350
rect 97674 58170 97730 58226
rect 97798 58170 97854 58226
rect 97922 58170 97978 58226
rect 98046 58170 98102 58226
rect 97674 58046 97730 58102
rect 97798 58046 97854 58102
rect 97922 58046 97978 58102
rect 98046 58046 98102 58102
rect 97674 57922 97730 57978
rect 97798 57922 97854 57978
rect 97922 57922 97978 57978
rect 98046 57922 98102 57978
rect 70674 46294 70730 46350
rect 70798 46294 70854 46350
rect 70922 46294 70978 46350
rect 71046 46294 71102 46350
rect 70674 46170 70730 46226
rect 70798 46170 70854 46226
rect 70922 46170 70978 46226
rect 71046 46170 71102 46226
rect 70674 46046 70730 46102
rect 70798 46046 70854 46102
rect 70922 46046 70978 46102
rect 71046 46046 71102 46102
rect 70674 45922 70730 45978
rect 70798 45922 70854 45978
rect 70922 45922 70978 45978
rect 71046 45922 71102 45978
rect 70674 28294 70730 28350
rect 70798 28294 70854 28350
rect 70922 28294 70978 28350
rect 71046 28294 71102 28350
rect 70674 28170 70730 28226
rect 70798 28170 70854 28226
rect 70922 28170 70978 28226
rect 71046 28170 71102 28226
rect 70674 28046 70730 28102
rect 70798 28046 70854 28102
rect 70922 28046 70978 28102
rect 71046 28046 71102 28102
rect 70674 27922 70730 27978
rect 70798 27922 70854 27978
rect 70922 27922 70978 27978
rect 71046 27922 71102 27978
rect 97674 40294 97730 40350
rect 97798 40294 97854 40350
rect 97922 40294 97978 40350
rect 98046 40294 98102 40350
rect 97674 40170 97730 40226
rect 97798 40170 97854 40226
rect 97922 40170 97978 40226
rect 98046 40170 98102 40226
rect 97674 40046 97730 40102
rect 97798 40046 97854 40102
rect 97922 40046 97978 40102
rect 98046 40046 98102 40102
rect 97674 39922 97730 39978
rect 97798 39922 97854 39978
rect 97922 39922 97978 39978
rect 98046 39922 98102 39978
rect 85906 22294 85962 22350
rect 86030 22294 86086 22350
rect 85906 22170 85962 22226
rect 86030 22170 86086 22226
rect 85906 22046 85962 22102
rect 86030 22046 86086 22102
rect 85906 21922 85962 21978
rect 86030 21922 86086 21978
rect 97674 22294 97730 22350
rect 97798 22294 97854 22350
rect 97922 22294 97978 22350
rect 98046 22294 98102 22350
rect 97674 22170 97730 22226
rect 97798 22170 97854 22226
rect 97922 22170 97978 22226
rect 98046 22170 98102 22226
rect 97674 22046 97730 22102
rect 97798 22046 97854 22102
rect 97922 22046 97978 22102
rect 98046 22046 98102 22102
rect 97674 21922 97730 21978
rect 97798 21922 97854 21978
rect 97922 21922 97978 21978
rect 98046 21922 98102 21978
rect 70674 10294 70730 10350
rect 70798 10294 70854 10350
rect 70922 10294 70978 10350
rect 71046 10294 71102 10350
rect 70674 10170 70730 10226
rect 70798 10170 70854 10226
rect 70922 10170 70978 10226
rect 71046 10170 71102 10226
rect 70674 10046 70730 10102
rect 70798 10046 70854 10102
rect 70922 10046 70978 10102
rect 71046 10046 71102 10102
rect 70674 9922 70730 9978
rect 70798 9922 70854 9978
rect 70922 9922 70978 9978
rect 71046 9922 71102 9978
rect 70674 -1176 70730 -1120
rect 70798 -1176 70854 -1120
rect 70922 -1176 70978 -1120
rect 71046 -1176 71102 -1120
rect 70674 -1300 70730 -1244
rect 70798 -1300 70854 -1244
rect 70922 -1300 70978 -1244
rect 71046 -1300 71102 -1244
rect 70674 -1424 70730 -1368
rect 70798 -1424 70854 -1368
rect 70922 -1424 70978 -1368
rect 71046 -1424 71102 -1368
rect 70674 -1548 70730 -1492
rect 70798 -1548 70854 -1492
rect 70922 -1548 70978 -1492
rect 71046 -1548 71102 -1492
rect 97674 4294 97730 4350
rect 97798 4294 97854 4350
rect 97922 4294 97978 4350
rect 98046 4294 98102 4350
rect 97674 4170 97730 4226
rect 97798 4170 97854 4226
rect 97922 4170 97978 4226
rect 98046 4170 98102 4226
rect 97674 4046 97730 4102
rect 97798 4046 97854 4102
rect 97922 4046 97978 4102
rect 98046 4046 98102 4102
rect 97674 3922 97730 3978
rect 97798 3922 97854 3978
rect 97922 3922 97978 3978
rect 98046 3922 98102 3978
rect 97674 -216 97730 -160
rect 97798 -216 97854 -160
rect 97922 -216 97978 -160
rect 98046 -216 98102 -160
rect 97674 -340 97730 -284
rect 97798 -340 97854 -284
rect 97922 -340 97978 -284
rect 98046 -340 98102 -284
rect 97674 -464 97730 -408
rect 97798 -464 97854 -408
rect 97922 -464 97978 -408
rect 98046 -464 98102 -408
rect 97674 -588 97730 -532
rect 97798 -588 97854 -532
rect 97922 -588 97978 -532
rect 98046 -588 98102 -532
rect 101394 154294 101450 154350
rect 101518 154294 101574 154350
rect 101642 154294 101698 154350
rect 101766 154294 101822 154350
rect 101394 154170 101450 154226
rect 101518 154170 101574 154226
rect 101642 154170 101698 154226
rect 101766 154170 101822 154226
rect 101394 154046 101450 154102
rect 101518 154046 101574 154102
rect 101642 154046 101698 154102
rect 101766 154046 101822 154102
rect 101394 153922 101450 153978
rect 101518 153922 101574 153978
rect 101642 153922 101698 153978
rect 101766 153922 101822 153978
rect 103292 264842 103348 264898
rect 103516 271322 103572 271378
rect 103628 205802 103684 205858
rect 104972 181502 105028 181558
rect 103516 177182 103572 177238
rect 103404 162602 103460 162658
rect 109116 365102 109172 365158
rect 108332 273302 108388 273358
rect 108444 357542 108500 357598
rect 108332 266822 108388 266878
rect 108556 279422 108612 279478
rect 110012 278342 110068 278398
rect 110124 366542 110180 366598
rect 110012 268442 110068 268498
rect 101394 136294 101450 136350
rect 101518 136294 101574 136350
rect 101642 136294 101698 136350
rect 101766 136294 101822 136350
rect 101394 136170 101450 136226
rect 101518 136170 101574 136226
rect 101642 136170 101698 136226
rect 101766 136170 101822 136226
rect 101394 136046 101450 136102
rect 101518 136046 101574 136102
rect 101642 136046 101698 136102
rect 101766 136046 101822 136102
rect 101394 135922 101450 135978
rect 101518 135922 101574 135978
rect 101642 135922 101698 135978
rect 101766 135922 101822 135978
rect 101394 118294 101450 118350
rect 101518 118294 101574 118350
rect 101642 118294 101698 118350
rect 101766 118294 101822 118350
rect 101394 118170 101450 118226
rect 101518 118170 101574 118226
rect 101642 118170 101698 118226
rect 101766 118170 101822 118226
rect 101394 118046 101450 118102
rect 101518 118046 101574 118102
rect 101642 118046 101698 118102
rect 101766 118046 101822 118102
rect 101394 117922 101450 117978
rect 101518 117922 101574 117978
rect 101642 117922 101698 117978
rect 101766 117922 101822 117978
rect 101394 100294 101450 100350
rect 101518 100294 101574 100350
rect 101642 100294 101698 100350
rect 101766 100294 101822 100350
rect 101394 100170 101450 100226
rect 101518 100170 101574 100226
rect 101642 100170 101698 100226
rect 101766 100170 101822 100226
rect 101394 100046 101450 100102
rect 101518 100046 101574 100102
rect 101642 100046 101698 100102
rect 101766 100046 101822 100102
rect 101394 99922 101450 99978
rect 101518 99922 101574 99978
rect 101642 99922 101698 99978
rect 101766 99922 101822 99978
rect 101394 82294 101450 82350
rect 101518 82294 101574 82350
rect 101642 82294 101698 82350
rect 101766 82294 101822 82350
rect 101394 82170 101450 82226
rect 101518 82170 101574 82226
rect 101642 82170 101698 82226
rect 101766 82170 101822 82226
rect 101394 82046 101450 82102
rect 101518 82046 101574 82102
rect 101642 82046 101698 82102
rect 101766 82046 101822 82102
rect 101394 81922 101450 81978
rect 101518 81922 101574 81978
rect 101642 81922 101698 81978
rect 101766 81922 101822 81978
rect 101394 64294 101450 64350
rect 101518 64294 101574 64350
rect 101642 64294 101698 64350
rect 101766 64294 101822 64350
rect 101394 64170 101450 64226
rect 101518 64170 101574 64226
rect 101642 64170 101698 64226
rect 101766 64170 101822 64226
rect 101394 64046 101450 64102
rect 101518 64046 101574 64102
rect 101642 64046 101698 64102
rect 101766 64046 101822 64102
rect 101394 63922 101450 63978
rect 101518 63922 101574 63978
rect 101642 63922 101698 63978
rect 101766 63922 101822 63978
rect 101394 46294 101450 46350
rect 101518 46294 101574 46350
rect 101642 46294 101698 46350
rect 101766 46294 101822 46350
rect 101394 46170 101450 46226
rect 101518 46170 101574 46226
rect 101642 46170 101698 46226
rect 101766 46170 101822 46226
rect 101394 46046 101450 46102
rect 101518 46046 101574 46102
rect 101642 46046 101698 46102
rect 101766 46046 101822 46102
rect 101394 45922 101450 45978
rect 101518 45922 101574 45978
rect 101642 45922 101698 45978
rect 101766 45922 101822 45978
rect 110124 149462 110180 149518
rect 110236 360062 110292 360118
rect 110348 357902 110404 357958
rect 110908 278162 110964 278218
rect 111692 271682 111748 271738
rect 112364 359882 112420 359938
rect 111804 269882 111860 269938
rect 111916 274562 111972 274618
rect 111692 206522 111748 206578
rect 111916 162782 111972 162838
rect 110348 149282 110404 149338
rect 114156 331982 114212 332038
rect 113036 312542 113092 312598
rect 119196 364922 119252 364978
rect 117516 362222 117572 362278
rect 114268 310940 114324 310978
rect 114268 310922 114324 310940
rect 115948 326042 116004 326098
rect 115052 277262 115108 277318
rect 113372 262862 113428 262918
rect 112700 261602 112756 261658
rect 113760 256294 113816 256350
rect 113884 256294 113940 256350
rect 114008 256294 114064 256350
rect 114132 256294 114188 256350
rect 113760 256170 113816 256226
rect 113884 256170 113940 256226
rect 114008 256170 114064 256226
rect 114132 256170 114188 256226
rect 113760 256046 113816 256102
rect 113884 256046 113940 256102
rect 114008 256046 114064 256102
rect 114132 256046 114188 256102
rect 113760 255922 113816 255978
rect 113884 255922 113940 255978
rect 114008 255922 114064 255978
rect 114132 255922 114188 255978
rect 115052 255302 115108 255358
rect 112960 244294 113016 244350
rect 113084 244294 113140 244350
rect 113208 244294 113264 244350
rect 113332 244294 113388 244350
rect 112960 244170 113016 244226
rect 113084 244170 113140 244226
rect 113208 244170 113264 244226
rect 113332 244170 113388 244226
rect 112960 244046 113016 244102
rect 113084 244046 113140 244102
rect 113208 244046 113264 244102
rect 113332 244046 113388 244102
rect 112960 243922 113016 243978
rect 113084 243922 113140 243978
rect 113208 243922 113264 243978
rect 113332 243922 113388 243978
rect 113760 238294 113816 238350
rect 113884 238294 113940 238350
rect 114008 238294 114064 238350
rect 114132 238294 114188 238350
rect 113760 238170 113816 238226
rect 113884 238170 113940 238226
rect 114008 238170 114064 238226
rect 114132 238170 114188 238226
rect 113760 238046 113816 238102
rect 113884 238046 113940 238102
rect 114008 238046 114064 238102
rect 114132 238046 114188 238102
rect 113760 237922 113816 237978
rect 113884 237922 113940 237978
rect 114008 237922 114064 237978
rect 114132 237922 114188 237978
rect 112960 226294 113016 226350
rect 113084 226294 113140 226350
rect 113208 226294 113264 226350
rect 113332 226294 113388 226350
rect 112960 226170 113016 226226
rect 113084 226170 113140 226226
rect 113208 226170 113264 226226
rect 113332 226170 113388 226226
rect 112960 226046 113016 226102
rect 113084 226046 113140 226102
rect 113208 226046 113264 226102
rect 113332 226046 113388 226102
rect 112960 225922 113016 225978
rect 113084 225922 113140 225978
rect 113208 225922 113264 225978
rect 113332 225922 113388 225978
rect 113760 220294 113816 220350
rect 113884 220294 113940 220350
rect 114008 220294 114064 220350
rect 114132 220294 114188 220350
rect 113760 220170 113816 220226
rect 113884 220170 113940 220226
rect 114008 220170 114064 220226
rect 114132 220170 114188 220226
rect 113760 220046 113816 220102
rect 113884 220046 113940 220102
rect 114008 220046 114064 220102
rect 114132 220046 114188 220102
rect 113760 219922 113816 219978
rect 113884 219922 113940 219978
rect 114008 219922 114064 219978
rect 114132 219922 114188 219978
rect 112960 208294 113016 208350
rect 113084 208294 113140 208350
rect 113208 208294 113264 208350
rect 113332 208294 113388 208350
rect 112960 208170 113016 208226
rect 113084 208170 113140 208226
rect 113208 208170 113264 208226
rect 113332 208170 113388 208226
rect 112960 208046 113016 208102
rect 113084 208046 113140 208102
rect 113208 208046 113264 208102
rect 113332 208046 113388 208102
rect 112960 207922 113016 207978
rect 113084 207922 113140 207978
rect 113208 207922 113264 207978
rect 113332 207922 113388 207978
rect 113760 202294 113816 202350
rect 113884 202294 113940 202350
rect 114008 202294 114064 202350
rect 114132 202294 114188 202350
rect 113760 202170 113816 202226
rect 113884 202170 113940 202226
rect 114008 202170 114064 202226
rect 114132 202170 114188 202226
rect 113760 202046 113816 202102
rect 113884 202046 113940 202102
rect 114008 202046 114064 202102
rect 114132 202046 114188 202102
rect 113760 201922 113816 201978
rect 113884 201922 113940 201978
rect 114008 201922 114064 201978
rect 114132 201922 114188 201978
rect 112960 190294 113016 190350
rect 113084 190294 113140 190350
rect 113208 190294 113264 190350
rect 113332 190294 113388 190350
rect 112960 190170 113016 190226
rect 113084 190170 113140 190226
rect 113208 190170 113264 190226
rect 113332 190170 113388 190226
rect 112960 190046 113016 190102
rect 113084 190046 113140 190102
rect 113208 190046 113264 190102
rect 113332 190046 113388 190102
rect 112960 189922 113016 189978
rect 113084 189922 113140 189978
rect 113208 189922 113264 189978
rect 113332 189922 113388 189978
rect 113760 184294 113816 184350
rect 113884 184294 113940 184350
rect 114008 184294 114064 184350
rect 114132 184294 114188 184350
rect 113760 184170 113816 184226
rect 113884 184170 113940 184226
rect 114008 184170 114064 184226
rect 114132 184170 114188 184226
rect 113760 184046 113816 184102
rect 113884 184046 113940 184102
rect 114008 184046 114064 184102
rect 114132 184046 114188 184102
rect 113760 183922 113816 183978
rect 113884 183922 113940 183978
rect 114008 183922 114064 183978
rect 114132 183922 114188 183978
rect 112960 172294 113016 172350
rect 113084 172294 113140 172350
rect 113208 172294 113264 172350
rect 113332 172294 113388 172350
rect 112960 172170 113016 172226
rect 113084 172170 113140 172226
rect 113208 172170 113264 172226
rect 113332 172170 113388 172226
rect 112960 172046 113016 172102
rect 113084 172046 113140 172102
rect 113208 172046 113264 172102
rect 113332 172046 113388 172102
rect 112960 171922 113016 171978
rect 113084 171922 113140 171978
rect 113208 171922 113264 171978
rect 113332 171922 113388 171978
rect 117516 331802 117572 331858
rect 117404 312542 117460 312598
rect 118412 319022 118468 319078
rect 118636 278522 118692 278578
rect 118748 277082 118804 277138
rect 119308 283922 119364 283978
rect 119980 286442 120036 286498
rect 119868 276902 119924 276958
rect 119644 276722 119700 276778
rect 119196 276542 119252 276598
rect 118860 270062 118916 270118
rect 118636 181502 118692 181558
rect 112476 149462 112532 149518
rect 118748 149462 118804 149518
rect 128394 580294 128450 580350
rect 128518 580294 128574 580350
rect 128642 580294 128698 580350
rect 128766 580294 128822 580350
rect 128394 580170 128450 580226
rect 128518 580170 128574 580226
rect 128642 580170 128698 580226
rect 128766 580170 128822 580226
rect 128394 580046 128450 580102
rect 128518 580046 128574 580102
rect 128642 580046 128698 580102
rect 128766 580046 128822 580102
rect 128394 579922 128450 579978
rect 128518 579922 128574 579978
rect 128642 579922 128698 579978
rect 128766 579922 128822 579978
rect 128394 562294 128450 562350
rect 128518 562294 128574 562350
rect 128642 562294 128698 562350
rect 128766 562294 128822 562350
rect 128394 562170 128450 562226
rect 128518 562170 128574 562226
rect 128642 562170 128698 562226
rect 128766 562170 128822 562226
rect 128394 562046 128450 562102
rect 128518 562046 128574 562102
rect 128642 562046 128698 562102
rect 128766 562046 128822 562102
rect 128394 561922 128450 561978
rect 128518 561922 128574 561978
rect 128642 561922 128698 561978
rect 128766 561922 128822 561978
rect 128394 544294 128450 544350
rect 128518 544294 128574 544350
rect 128642 544294 128698 544350
rect 128766 544294 128822 544350
rect 128394 544170 128450 544226
rect 128518 544170 128574 544226
rect 128642 544170 128698 544226
rect 128766 544170 128822 544226
rect 128394 544046 128450 544102
rect 128518 544046 128574 544102
rect 128642 544046 128698 544102
rect 128766 544046 128822 544102
rect 128394 543922 128450 543978
rect 128518 543922 128574 543978
rect 128642 543922 128698 543978
rect 128766 543922 128822 543978
rect 128394 526294 128450 526350
rect 128518 526294 128574 526350
rect 128642 526294 128698 526350
rect 128766 526294 128822 526350
rect 128394 526170 128450 526226
rect 128518 526170 128574 526226
rect 128642 526170 128698 526226
rect 128766 526170 128822 526226
rect 128394 526046 128450 526102
rect 128518 526046 128574 526102
rect 128642 526046 128698 526102
rect 128766 526046 128822 526102
rect 128394 525922 128450 525978
rect 128518 525922 128574 525978
rect 128642 525922 128698 525978
rect 128766 525922 128822 525978
rect 128394 508294 128450 508350
rect 128518 508294 128574 508350
rect 128642 508294 128698 508350
rect 128766 508294 128822 508350
rect 128394 508170 128450 508226
rect 128518 508170 128574 508226
rect 128642 508170 128698 508226
rect 128766 508170 128822 508226
rect 128394 508046 128450 508102
rect 128518 508046 128574 508102
rect 128642 508046 128698 508102
rect 128766 508046 128822 508102
rect 128394 507922 128450 507978
rect 128518 507922 128574 507978
rect 128642 507922 128698 507978
rect 128766 507922 128822 507978
rect 128394 490294 128450 490350
rect 128518 490294 128574 490350
rect 128642 490294 128698 490350
rect 128766 490294 128822 490350
rect 128394 490170 128450 490226
rect 128518 490170 128574 490226
rect 128642 490170 128698 490226
rect 128766 490170 128822 490226
rect 128394 490046 128450 490102
rect 128518 490046 128574 490102
rect 128642 490046 128698 490102
rect 128766 490046 128822 490102
rect 128394 489922 128450 489978
rect 128518 489922 128574 489978
rect 128642 489922 128698 489978
rect 128766 489922 128822 489978
rect 128394 472294 128450 472350
rect 128518 472294 128574 472350
rect 128642 472294 128698 472350
rect 128766 472294 128822 472350
rect 128394 472170 128450 472226
rect 128518 472170 128574 472226
rect 128642 472170 128698 472226
rect 128766 472170 128822 472226
rect 128394 472046 128450 472102
rect 128518 472046 128574 472102
rect 128642 472046 128698 472102
rect 128766 472046 128822 472102
rect 128394 471922 128450 471978
rect 128518 471922 128574 471978
rect 128642 471922 128698 471978
rect 128766 471922 128822 471978
rect 128394 454294 128450 454350
rect 128518 454294 128574 454350
rect 128642 454294 128698 454350
rect 128766 454294 128822 454350
rect 128394 454170 128450 454226
rect 128518 454170 128574 454226
rect 128642 454170 128698 454226
rect 128766 454170 128822 454226
rect 128394 454046 128450 454102
rect 128518 454046 128574 454102
rect 128642 454046 128698 454102
rect 128766 454046 128822 454102
rect 128394 453922 128450 453978
rect 128518 453922 128574 453978
rect 128642 453922 128698 453978
rect 128766 453922 128822 453978
rect 128394 436294 128450 436350
rect 128518 436294 128574 436350
rect 128642 436294 128698 436350
rect 128766 436294 128822 436350
rect 128394 436170 128450 436226
rect 128518 436170 128574 436226
rect 128642 436170 128698 436226
rect 128766 436170 128822 436226
rect 128394 436046 128450 436102
rect 128518 436046 128574 436102
rect 128642 436046 128698 436102
rect 128766 436046 128822 436102
rect 128394 435922 128450 435978
rect 128518 435922 128574 435978
rect 128642 435922 128698 435978
rect 128766 435922 128822 435978
rect 128394 418294 128450 418350
rect 128518 418294 128574 418350
rect 128642 418294 128698 418350
rect 128766 418294 128822 418350
rect 128394 418170 128450 418226
rect 128518 418170 128574 418226
rect 128642 418170 128698 418226
rect 128766 418170 128822 418226
rect 128394 418046 128450 418102
rect 128518 418046 128574 418102
rect 128642 418046 128698 418102
rect 128766 418046 128822 418102
rect 128394 417922 128450 417978
rect 128518 417922 128574 417978
rect 128642 417922 128698 417978
rect 128766 417922 128822 417978
rect 128394 400294 128450 400350
rect 128518 400294 128574 400350
rect 128642 400294 128698 400350
rect 128766 400294 128822 400350
rect 128394 400170 128450 400226
rect 128518 400170 128574 400226
rect 128642 400170 128698 400226
rect 128766 400170 128822 400226
rect 128394 400046 128450 400102
rect 128518 400046 128574 400102
rect 128642 400046 128698 400102
rect 128766 400046 128822 400102
rect 128394 399922 128450 399978
rect 128518 399922 128574 399978
rect 128642 399922 128698 399978
rect 128766 399922 128822 399978
rect 128394 382294 128450 382350
rect 128518 382294 128574 382350
rect 128642 382294 128698 382350
rect 128766 382294 128822 382350
rect 128394 382170 128450 382226
rect 128518 382170 128574 382226
rect 128642 382170 128698 382226
rect 128766 382170 128822 382226
rect 128394 382046 128450 382102
rect 128518 382046 128574 382102
rect 128642 382046 128698 382102
rect 128766 382046 128822 382102
rect 128394 381922 128450 381978
rect 128518 381922 128574 381978
rect 128642 381922 128698 381978
rect 128766 381922 128822 381978
rect 128394 364294 128450 364350
rect 128518 364294 128574 364350
rect 128642 364294 128698 364350
rect 128766 364294 128822 364350
rect 128394 364170 128450 364226
rect 128518 364170 128574 364226
rect 128642 364170 128698 364226
rect 128766 364170 128822 364226
rect 128394 364046 128450 364102
rect 128518 364046 128574 364102
rect 128642 364046 128698 364102
rect 128766 364046 128822 364102
rect 128394 363922 128450 363978
rect 128518 363922 128574 363978
rect 128642 363922 128698 363978
rect 128766 363922 128822 363978
rect 132114 598116 132170 598172
rect 132238 598116 132294 598172
rect 132362 598116 132418 598172
rect 132486 598116 132542 598172
rect 132114 597992 132170 598048
rect 132238 597992 132294 598048
rect 132362 597992 132418 598048
rect 132486 597992 132542 598048
rect 132114 597868 132170 597924
rect 132238 597868 132294 597924
rect 132362 597868 132418 597924
rect 132486 597868 132542 597924
rect 132114 597744 132170 597800
rect 132238 597744 132294 597800
rect 132362 597744 132418 597800
rect 132486 597744 132542 597800
rect 132114 586294 132170 586350
rect 132238 586294 132294 586350
rect 132362 586294 132418 586350
rect 132486 586294 132542 586350
rect 132114 586170 132170 586226
rect 132238 586170 132294 586226
rect 132362 586170 132418 586226
rect 132486 586170 132542 586226
rect 132114 586046 132170 586102
rect 132238 586046 132294 586102
rect 132362 586046 132418 586102
rect 132486 586046 132542 586102
rect 132114 585922 132170 585978
rect 132238 585922 132294 585978
rect 132362 585922 132418 585978
rect 132486 585922 132542 585978
rect 132114 568294 132170 568350
rect 132238 568294 132294 568350
rect 132362 568294 132418 568350
rect 132486 568294 132542 568350
rect 132114 568170 132170 568226
rect 132238 568170 132294 568226
rect 132362 568170 132418 568226
rect 132486 568170 132542 568226
rect 132114 568046 132170 568102
rect 132238 568046 132294 568102
rect 132362 568046 132418 568102
rect 132486 568046 132542 568102
rect 132114 567922 132170 567978
rect 132238 567922 132294 567978
rect 132362 567922 132418 567978
rect 132486 567922 132542 567978
rect 132114 550294 132170 550350
rect 132238 550294 132294 550350
rect 132362 550294 132418 550350
rect 132486 550294 132542 550350
rect 132114 550170 132170 550226
rect 132238 550170 132294 550226
rect 132362 550170 132418 550226
rect 132486 550170 132542 550226
rect 132114 550046 132170 550102
rect 132238 550046 132294 550102
rect 132362 550046 132418 550102
rect 132486 550046 132542 550102
rect 132114 549922 132170 549978
rect 132238 549922 132294 549978
rect 132362 549922 132418 549978
rect 132486 549922 132542 549978
rect 132114 532294 132170 532350
rect 132238 532294 132294 532350
rect 132362 532294 132418 532350
rect 132486 532294 132542 532350
rect 132114 532170 132170 532226
rect 132238 532170 132294 532226
rect 132362 532170 132418 532226
rect 132486 532170 132542 532226
rect 132114 532046 132170 532102
rect 132238 532046 132294 532102
rect 132362 532046 132418 532102
rect 132486 532046 132542 532102
rect 132114 531922 132170 531978
rect 132238 531922 132294 531978
rect 132362 531922 132418 531978
rect 132486 531922 132542 531978
rect 132114 514294 132170 514350
rect 132238 514294 132294 514350
rect 132362 514294 132418 514350
rect 132486 514294 132542 514350
rect 132114 514170 132170 514226
rect 132238 514170 132294 514226
rect 132362 514170 132418 514226
rect 132486 514170 132542 514226
rect 132114 514046 132170 514102
rect 132238 514046 132294 514102
rect 132362 514046 132418 514102
rect 132486 514046 132542 514102
rect 132114 513922 132170 513978
rect 132238 513922 132294 513978
rect 132362 513922 132418 513978
rect 132486 513922 132542 513978
rect 132114 496294 132170 496350
rect 132238 496294 132294 496350
rect 132362 496294 132418 496350
rect 132486 496294 132542 496350
rect 132114 496170 132170 496226
rect 132238 496170 132294 496226
rect 132362 496170 132418 496226
rect 132486 496170 132542 496226
rect 132114 496046 132170 496102
rect 132238 496046 132294 496102
rect 132362 496046 132418 496102
rect 132486 496046 132542 496102
rect 132114 495922 132170 495978
rect 132238 495922 132294 495978
rect 132362 495922 132418 495978
rect 132486 495922 132542 495978
rect 132114 478294 132170 478350
rect 132238 478294 132294 478350
rect 132362 478294 132418 478350
rect 132486 478294 132542 478350
rect 132114 478170 132170 478226
rect 132238 478170 132294 478226
rect 132362 478170 132418 478226
rect 132486 478170 132542 478226
rect 132114 478046 132170 478102
rect 132238 478046 132294 478102
rect 132362 478046 132418 478102
rect 132486 478046 132542 478102
rect 132114 477922 132170 477978
rect 132238 477922 132294 477978
rect 132362 477922 132418 477978
rect 132486 477922 132542 477978
rect 132114 460294 132170 460350
rect 132238 460294 132294 460350
rect 132362 460294 132418 460350
rect 132486 460294 132542 460350
rect 132114 460170 132170 460226
rect 132238 460170 132294 460226
rect 132362 460170 132418 460226
rect 132486 460170 132542 460226
rect 132114 460046 132170 460102
rect 132238 460046 132294 460102
rect 132362 460046 132418 460102
rect 132486 460046 132542 460102
rect 132114 459922 132170 459978
rect 132238 459922 132294 459978
rect 132362 459922 132418 459978
rect 132486 459922 132542 459978
rect 132114 442294 132170 442350
rect 132238 442294 132294 442350
rect 132362 442294 132418 442350
rect 132486 442294 132542 442350
rect 132114 442170 132170 442226
rect 132238 442170 132294 442226
rect 132362 442170 132418 442226
rect 132486 442170 132542 442226
rect 132114 442046 132170 442102
rect 132238 442046 132294 442102
rect 132362 442046 132418 442102
rect 132486 442046 132542 442102
rect 132114 441922 132170 441978
rect 132238 441922 132294 441978
rect 132362 441922 132418 441978
rect 132486 441922 132542 441978
rect 132114 424294 132170 424350
rect 132238 424294 132294 424350
rect 132362 424294 132418 424350
rect 132486 424294 132542 424350
rect 132114 424170 132170 424226
rect 132238 424170 132294 424226
rect 132362 424170 132418 424226
rect 132486 424170 132542 424226
rect 132114 424046 132170 424102
rect 132238 424046 132294 424102
rect 132362 424046 132418 424102
rect 132486 424046 132542 424102
rect 132114 423922 132170 423978
rect 132238 423922 132294 423978
rect 132362 423922 132418 423978
rect 132486 423922 132542 423978
rect 132114 406294 132170 406350
rect 132238 406294 132294 406350
rect 132362 406294 132418 406350
rect 132486 406294 132542 406350
rect 132114 406170 132170 406226
rect 132238 406170 132294 406226
rect 132362 406170 132418 406226
rect 132486 406170 132542 406226
rect 132114 406046 132170 406102
rect 132238 406046 132294 406102
rect 132362 406046 132418 406102
rect 132486 406046 132542 406102
rect 132114 405922 132170 405978
rect 132238 405922 132294 405978
rect 132362 405922 132418 405978
rect 132486 405922 132542 405978
rect 132114 388294 132170 388350
rect 132238 388294 132294 388350
rect 132362 388294 132418 388350
rect 132486 388294 132542 388350
rect 132114 388170 132170 388226
rect 132238 388170 132294 388226
rect 132362 388170 132418 388226
rect 132486 388170 132542 388226
rect 132114 388046 132170 388102
rect 132238 388046 132294 388102
rect 132362 388046 132418 388102
rect 132486 388046 132542 388102
rect 132114 387922 132170 387978
rect 132238 387922 132294 387978
rect 132362 387922 132418 387978
rect 132486 387922 132542 387978
rect 132114 370294 132170 370350
rect 132238 370294 132294 370350
rect 132362 370294 132418 370350
rect 132486 370294 132542 370350
rect 132114 370170 132170 370226
rect 132238 370170 132294 370226
rect 132362 370170 132418 370226
rect 132486 370170 132542 370226
rect 132114 370046 132170 370102
rect 132238 370046 132294 370102
rect 132362 370046 132418 370102
rect 132486 370046 132542 370102
rect 132114 369922 132170 369978
rect 132238 369922 132294 369978
rect 132362 369922 132418 369978
rect 132486 369922 132542 369978
rect 159114 597156 159170 597212
rect 159238 597156 159294 597212
rect 159362 597156 159418 597212
rect 159486 597156 159542 597212
rect 159114 597032 159170 597088
rect 159238 597032 159294 597088
rect 159362 597032 159418 597088
rect 159486 597032 159542 597088
rect 159114 596908 159170 596964
rect 159238 596908 159294 596964
rect 159362 596908 159418 596964
rect 159486 596908 159542 596964
rect 159114 596784 159170 596840
rect 159238 596784 159294 596840
rect 159362 596784 159418 596840
rect 159486 596784 159542 596840
rect 159114 580294 159170 580350
rect 159238 580294 159294 580350
rect 159362 580294 159418 580350
rect 159486 580294 159542 580350
rect 159114 580170 159170 580226
rect 159238 580170 159294 580226
rect 159362 580170 159418 580226
rect 159486 580170 159542 580226
rect 159114 580046 159170 580102
rect 159238 580046 159294 580102
rect 159362 580046 159418 580102
rect 159486 580046 159542 580102
rect 159114 579922 159170 579978
rect 159238 579922 159294 579978
rect 159362 579922 159418 579978
rect 159486 579922 159542 579978
rect 159114 562294 159170 562350
rect 159238 562294 159294 562350
rect 159362 562294 159418 562350
rect 159486 562294 159542 562350
rect 159114 562170 159170 562226
rect 159238 562170 159294 562226
rect 159362 562170 159418 562226
rect 159486 562170 159542 562226
rect 159114 562046 159170 562102
rect 159238 562046 159294 562102
rect 159362 562046 159418 562102
rect 159486 562046 159542 562102
rect 159114 561922 159170 561978
rect 159238 561922 159294 561978
rect 159362 561922 159418 561978
rect 159486 561922 159542 561978
rect 159114 544294 159170 544350
rect 159238 544294 159294 544350
rect 159362 544294 159418 544350
rect 159486 544294 159542 544350
rect 159114 544170 159170 544226
rect 159238 544170 159294 544226
rect 159362 544170 159418 544226
rect 159486 544170 159542 544226
rect 159114 544046 159170 544102
rect 159238 544046 159294 544102
rect 159362 544046 159418 544102
rect 159486 544046 159542 544102
rect 159114 543922 159170 543978
rect 159238 543922 159294 543978
rect 159362 543922 159418 543978
rect 159486 543922 159542 543978
rect 159114 526294 159170 526350
rect 159238 526294 159294 526350
rect 159362 526294 159418 526350
rect 159486 526294 159542 526350
rect 159114 526170 159170 526226
rect 159238 526170 159294 526226
rect 159362 526170 159418 526226
rect 159486 526170 159542 526226
rect 159114 526046 159170 526102
rect 159238 526046 159294 526102
rect 159362 526046 159418 526102
rect 159486 526046 159542 526102
rect 159114 525922 159170 525978
rect 159238 525922 159294 525978
rect 159362 525922 159418 525978
rect 159486 525922 159542 525978
rect 159114 508294 159170 508350
rect 159238 508294 159294 508350
rect 159362 508294 159418 508350
rect 159486 508294 159542 508350
rect 159114 508170 159170 508226
rect 159238 508170 159294 508226
rect 159362 508170 159418 508226
rect 159486 508170 159542 508226
rect 159114 508046 159170 508102
rect 159238 508046 159294 508102
rect 159362 508046 159418 508102
rect 159486 508046 159542 508102
rect 159114 507922 159170 507978
rect 159238 507922 159294 507978
rect 159362 507922 159418 507978
rect 159486 507922 159542 507978
rect 159114 490294 159170 490350
rect 159238 490294 159294 490350
rect 159362 490294 159418 490350
rect 159486 490294 159542 490350
rect 159114 490170 159170 490226
rect 159238 490170 159294 490226
rect 159362 490170 159418 490226
rect 159486 490170 159542 490226
rect 159114 490046 159170 490102
rect 159238 490046 159294 490102
rect 159362 490046 159418 490102
rect 159486 490046 159542 490102
rect 159114 489922 159170 489978
rect 159238 489922 159294 489978
rect 159362 489922 159418 489978
rect 159486 489922 159542 489978
rect 159114 472294 159170 472350
rect 159238 472294 159294 472350
rect 159362 472294 159418 472350
rect 159486 472294 159542 472350
rect 159114 472170 159170 472226
rect 159238 472170 159294 472226
rect 159362 472170 159418 472226
rect 159486 472170 159542 472226
rect 159114 472046 159170 472102
rect 159238 472046 159294 472102
rect 159362 472046 159418 472102
rect 159486 472046 159542 472102
rect 159114 471922 159170 471978
rect 159238 471922 159294 471978
rect 159362 471922 159418 471978
rect 159486 471922 159542 471978
rect 159114 454294 159170 454350
rect 159238 454294 159294 454350
rect 159362 454294 159418 454350
rect 159486 454294 159542 454350
rect 159114 454170 159170 454226
rect 159238 454170 159294 454226
rect 159362 454170 159418 454226
rect 159486 454170 159542 454226
rect 159114 454046 159170 454102
rect 159238 454046 159294 454102
rect 159362 454046 159418 454102
rect 159486 454046 159542 454102
rect 159114 453922 159170 453978
rect 159238 453922 159294 453978
rect 159362 453922 159418 453978
rect 159486 453922 159542 453978
rect 159114 436294 159170 436350
rect 159238 436294 159294 436350
rect 159362 436294 159418 436350
rect 159486 436294 159542 436350
rect 159114 436170 159170 436226
rect 159238 436170 159294 436226
rect 159362 436170 159418 436226
rect 159486 436170 159542 436226
rect 159114 436046 159170 436102
rect 159238 436046 159294 436102
rect 159362 436046 159418 436102
rect 159486 436046 159542 436102
rect 159114 435922 159170 435978
rect 159238 435922 159294 435978
rect 159362 435922 159418 435978
rect 159486 435922 159542 435978
rect 159114 418294 159170 418350
rect 159238 418294 159294 418350
rect 159362 418294 159418 418350
rect 159486 418294 159542 418350
rect 159114 418170 159170 418226
rect 159238 418170 159294 418226
rect 159362 418170 159418 418226
rect 159486 418170 159542 418226
rect 159114 418046 159170 418102
rect 159238 418046 159294 418102
rect 159362 418046 159418 418102
rect 159486 418046 159542 418102
rect 159114 417922 159170 417978
rect 159238 417922 159294 417978
rect 159362 417922 159418 417978
rect 159486 417922 159542 417978
rect 159114 400294 159170 400350
rect 159238 400294 159294 400350
rect 159362 400294 159418 400350
rect 159486 400294 159542 400350
rect 159114 400170 159170 400226
rect 159238 400170 159294 400226
rect 159362 400170 159418 400226
rect 159486 400170 159542 400226
rect 159114 400046 159170 400102
rect 159238 400046 159294 400102
rect 159362 400046 159418 400102
rect 159486 400046 159542 400102
rect 159114 399922 159170 399978
rect 159238 399922 159294 399978
rect 159362 399922 159418 399978
rect 159486 399922 159542 399978
rect 159114 382294 159170 382350
rect 159238 382294 159294 382350
rect 159362 382294 159418 382350
rect 159486 382294 159542 382350
rect 159114 382170 159170 382226
rect 159238 382170 159294 382226
rect 159362 382170 159418 382226
rect 159486 382170 159542 382226
rect 159114 382046 159170 382102
rect 159238 382046 159294 382102
rect 159362 382046 159418 382102
rect 159486 382046 159542 382102
rect 159114 381922 159170 381978
rect 159238 381922 159294 381978
rect 159362 381922 159418 381978
rect 159486 381922 159542 381978
rect 156156 364742 156212 364798
rect 151340 363122 151396 363178
rect 152012 362964 152068 362998
rect 152012 362942 152068 362964
rect 157836 364562 157892 364618
rect 162834 598116 162890 598172
rect 162958 598116 163014 598172
rect 163082 598116 163138 598172
rect 163206 598116 163262 598172
rect 162834 597992 162890 598048
rect 162958 597992 163014 598048
rect 163082 597992 163138 598048
rect 163206 597992 163262 598048
rect 162834 597868 162890 597924
rect 162958 597868 163014 597924
rect 163082 597868 163138 597924
rect 163206 597868 163262 597924
rect 162834 597744 162890 597800
rect 162958 597744 163014 597800
rect 163082 597744 163138 597800
rect 163206 597744 163262 597800
rect 162834 586294 162890 586350
rect 162958 586294 163014 586350
rect 163082 586294 163138 586350
rect 163206 586294 163262 586350
rect 162834 586170 162890 586226
rect 162958 586170 163014 586226
rect 163082 586170 163138 586226
rect 163206 586170 163262 586226
rect 162834 586046 162890 586102
rect 162958 586046 163014 586102
rect 163082 586046 163138 586102
rect 163206 586046 163262 586102
rect 162834 585922 162890 585978
rect 162958 585922 163014 585978
rect 163082 585922 163138 585978
rect 163206 585922 163262 585978
rect 162834 568294 162890 568350
rect 162958 568294 163014 568350
rect 163082 568294 163138 568350
rect 163206 568294 163262 568350
rect 162834 568170 162890 568226
rect 162958 568170 163014 568226
rect 163082 568170 163138 568226
rect 163206 568170 163262 568226
rect 162834 568046 162890 568102
rect 162958 568046 163014 568102
rect 163082 568046 163138 568102
rect 163206 568046 163262 568102
rect 162834 567922 162890 567978
rect 162958 567922 163014 567978
rect 163082 567922 163138 567978
rect 163206 567922 163262 567978
rect 162834 550294 162890 550350
rect 162958 550294 163014 550350
rect 163082 550294 163138 550350
rect 163206 550294 163262 550350
rect 162834 550170 162890 550226
rect 162958 550170 163014 550226
rect 163082 550170 163138 550226
rect 163206 550170 163262 550226
rect 162834 550046 162890 550102
rect 162958 550046 163014 550102
rect 163082 550046 163138 550102
rect 163206 550046 163262 550102
rect 162834 549922 162890 549978
rect 162958 549922 163014 549978
rect 163082 549922 163138 549978
rect 163206 549922 163262 549978
rect 162834 532294 162890 532350
rect 162958 532294 163014 532350
rect 163082 532294 163138 532350
rect 163206 532294 163262 532350
rect 162834 532170 162890 532226
rect 162958 532170 163014 532226
rect 163082 532170 163138 532226
rect 163206 532170 163262 532226
rect 162834 532046 162890 532102
rect 162958 532046 163014 532102
rect 163082 532046 163138 532102
rect 163206 532046 163262 532102
rect 162834 531922 162890 531978
rect 162958 531922 163014 531978
rect 163082 531922 163138 531978
rect 163206 531922 163262 531978
rect 162834 514294 162890 514350
rect 162958 514294 163014 514350
rect 163082 514294 163138 514350
rect 163206 514294 163262 514350
rect 162834 514170 162890 514226
rect 162958 514170 163014 514226
rect 163082 514170 163138 514226
rect 163206 514170 163262 514226
rect 162834 514046 162890 514102
rect 162958 514046 163014 514102
rect 163082 514046 163138 514102
rect 163206 514046 163262 514102
rect 162834 513922 162890 513978
rect 162958 513922 163014 513978
rect 163082 513922 163138 513978
rect 163206 513922 163262 513978
rect 162834 496294 162890 496350
rect 162958 496294 163014 496350
rect 163082 496294 163138 496350
rect 163206 496294 163262 496350
rect 162834 496170 162890 496226
rect 162958 496170 163014 496226
rect 163082 496170 163138 496226
rect 163206 496170 163262 496226
rect 162834 496046 162890 496102
rect 162958 496046 163014 496102
rect 163082 496046 163138 496102
rect 163206 496046 163262 496102
rect 162834 495922 162890 495978
rect 162958 495922 163014 495978
rect 163082 495922 163138 495978
rect 163206 495922 163262 495978
rect 162834 478294 162890 478350
rect 162958 478294 163014 478350
rect 163082 478294 163138 478350
rect 163206 478294 163262 478350
rect 162834 478170 162890 478226
rect 162958 478170 163014 478226
rect 163082 478170 163138 478226
rect 163206 478170 163262 478226
rect 162834 478046 162890 478102
rect 162958 478046 163014 478102
rect 163082 478046 163138 478102
rect 163206 478046 163262 478102
rect 162834 477922 162890 477978
rect 162958 477922 163014 477978
rect 163082 477922 163138 477978
rect 163206 477922 163262 477978
rect 162834 460294 162890 460350
rect 162958 460294 163014 460350
rect 163082 460294 163138 460350
rect 163206 460294 163262 460350
rect 162834 460170 162890 460226
rect 162958 460170 163014 460226
rect 163082 460170 163138 460226
rect 163206 460170 163262 460226
rect 162834 460046 162890 460102
rect 162958 460046 163014 460102
rect 163082 460046 163138 460102
rect 163206 460046 163262 460102
rect 162834 459922 162890 459978
rect 162958 459922 163014 459978
rect 163082 459922 163138 459978
rect 163206 459922 163262 459978
rect 162834 442294 162890 442350
rect 162958 442294 163014 442350
rect 163082 442294 163138 442350
rect 163206 442294 163262 442350
rect 162834 442170 162890 442226
rect 162958 442170 163014 442226
rect 163082 442170 163138 442226
rect 163206 442170 163262 442226
rect 162834 442046 162890 442102
rect 162958 442046 163014 442102
rect 163082 442046 163138 442102
rect 163206 442046 163262 442102
rect 162834 441922 162890 441978
rect 162958 441922 163014 441978
rect 163082 441922 163138 441978
rect 163206 441922 163262 441978
rect 162834 424294 162890 424350
rect 162958 424294 163014 424350
rect 163082 424294 163138 424350
rect 163206 424294 163262 424350
rect 162834 424170 162890 424226
rect 162958 424170 163014 424226
rect 163082 424170 163138 424226
rect 163206 424170 163262 424226
rect 162834 424046 162890 424102
rect 162958 424046 163014 424102
rect 163082 424046 163138 424102
rect 163206 424046 163262 424102
rect 162834 423922 162890 423978
rect 162958 423922 163014 423978
rect 163082 423922 163138 423978
rect 163206 423922 163262 423978
rect 162834 406294 162890 406350
rect 162958 406294 163014 406350
rect 163082 406294 163138 406350
rect 163206 406294 163262 406350
rect 162834 406170 162890 406226
rect 162958 406170 163014 406226
rect 163082 406170 163138 406226
rect 163206 406170 163262 406226
rect 162834 406046 162890 406102
rect 162958 406046 163014 406102
rect 163082 406046 163138 406102
rect 163206 406046 163262 406102
rect 162834 405922 162890 405978
rect 162958 405922 163014 405978
rect 163082 405922 163138 405978
rect 163206 405922 163262 405978
rect 162834 388294 162890 388350
rect 162958 388294 163014 388350
rect 163082 388294 163138 388350
rect 163206 388294 163262 388350
rect 162834 388170 162890 388226
rect 162958 388170 163014 388226
rect 163082 388170 163138 388226
rect 163206 388170 163262 388226
rect 162834 388046 162890 388102
rect 162958 388046 163014 388102
rect 163082 388046 163138 388102
rect 163206 388046 163262 388102
rect 162834 387922 162890 387978
rect 162958 387922 163014 387978
rect 163082 387922 163138 387978
rect 163206 387922 163262 387978
rect 162834 370294 162890 370350
rect 162958 370294 163014 370350
rect 163082 370294 163138 370350
rect 163206 370294 163262 370350
rect 162834 370170 162890 370226
rect 162958 370170 163014 370226
rect 163082 370170 163138 370226
rect 163206 370170 163262 370226
rect 162834 370046 162890 370102
rect 162958 370046 163014 370102
rect 163082 370046 163138 370102
rect 163206 370046 163262 370102
rect 162834 369922 162890 369978
rect 162958 369922 163014 369978
rect 163082 369922 163138 369978
rect 163206 369922 163262 369978
rect 159114 364294 159170 364350
rect 159238 364294 159294 364350
rect 159362 364294 159418 364350
rect 159486 364294 159542 364350
rect 159114 364170 159170 364226
rect 159238 364170 159294 364226
rect 159362 364170 159418 364226
rect 159486 364170 159542 364226
rect 159114 364046 159170 364102
rect 159238 364046 159294 364102
rect 159362 364046 159418 364102
rect 159486 364046 159542 364102
rect 159114 363922 159170 363978
rect 159238 363922 159294 363978
rect 159362 363922 159418 363978
rect 159486 363922 159542 363978
rect 150668 362042 150724 362098
rect 160748 365102 160804 365158
rect 161420 361502 161476 361558
rect 189834 597156 189890 597212
rect 189958 597156 190014 597212
rect 190082 597156 190138 597212
rect 190206 597156 190262 597212
rect 189834 597032 189890 597088
rect 189958 597032 190014 597088
rect 190082 597032 190138 597088
rect 190206 597032 190262 597088
rect 189834 596908 189890 596964
rect 189958 596908 190014 596964
rect 190082 596908 190138 596964
rect 190206 596908 190262 596964
rect 189834 596784 189890 596840
rect 189958 596784 190014 596840
rect 190082 596784 190138 596840
rect 190206 596784 190262 596840
rect 189834 580294 189890 580350
rect 189958 580294 190014 580350
rect 190082 580294 190138 580350
rect 190206 580294 190262 580350
rect 189834 580170 189890 580226
rect 189958 580170 190014 580226
rect 190082 580170 190138 580226
rect 190206 580170 190262 580226
rect 189834 580046 189890 580102
rect 189958 580046 190014 580102
rect 190082 580046 190138 580102
rect 190206 580046 190262 580102
rect 189834 579922 189890 579978
rect 189958 579922 190014 579978
rect 190082 579922 190138 579978
rect 190206 579922 190262 579978
rect 189834 562294 189890 562350
rect 189958 562294 190014 562350
rect 190082 562294 190138 562350
rect 190206 562294 190262 562350
rect 189834 562170 189890 562226
rect 189958 562170 190014 562226
rect 190082 562170 190138 562226
rect 190206 562170 190262 562226
rect 189834 562046 189890 562102
rect 189958 562046 190014 562102
rect 190082 562046 190138 562102
rect 190206 562046 190262 562102
rect 189834 561922 189890 561978
rect 189958 561922 190014 561978
rect 190082 561922 190138 561978
rect 190206 561922 190262 561978
rect 189834 544294 189890 544350
rect 189958 544294 190014 544350
rect 190082 544294 190138 544350
rect 190206 544294 190262 544350
rect 189834 544170 189890 544226
rect 189958 544170 190014 544226
rect 190082 544170 190138 544226
rect 190206 544170 190262 544226
rect 189834 544046 189890 544102
rect 189958 544046 190014 544102
rect 190082 544046 190138 544102
rect 190206 544046 190262 544102
rect 189834 543922 189890 543978
rect 189958 543922 190014 543978
rect 190082 543922 190138 543978
rect 190206 543922 190262 543978
rect 189834 526294 189890 526350
rect 189958 526294 190014 526350
rect 190082 526294 190138 526350
rect 190206 526294 190262 526350
rect 189834 526170 189890 526226
rect 189958 526170 190014 526226
rect 190082 526170 190138 526226
rect 190206 526170 190262 526226
rect 189834 526046 189890 526102
rect 189958 526046 190014 526102
rect 190082 526046 190138 526102
rect 190206 526046 190262 526102
rect 189834 525922 189890 525978
rect 189958 525922 190014 525978
rect 190082 525922 190138 525978
rect 190206 525922 190262 525978
rect 189834 508294 189890 508350
rect 189958 508294 190014 508350
rect 190082 508294 190138 508350
rect 190206 508294 190262 508350
rect 189834 508170 189890 508226
rect 189958 508170 190014 508226
rect 190082 508170 190138 508226
rect 190206 508170 190262 508226
rect 189834 508046 189890 508102
rect 189958 508046 190014 508102
rect 190082 508046 190138 508102
rect 190206 508046 190262 508102
rect 189834 507922 189890 507978
rect 189958 507922 190014 507978
rect 190082 507922 190138 507978
rect 190206 507922 190262 507978
rect 189834 490294 189890 490350
rect 189958 490294 190014 490350
rect 190082 490294 190138 490350
rect 190206 490294 190262 490350
rect 189834 490170 189890 490226
rect 189958 490170 190014 490226
rect 190082 490170 190138 490226
rect 190206 490170 190262 490226
rect 189834 490046 189890 490102
rect 189958 490046 190014 490102
rect 190082 490046 190138 490102
rect 190206 490046 190262 490102
rect 189834 489922 189890 489978
rect 189958 489922 190014 489978
rect 190082 489922 190138 489978
rect 190206 489922 190262 489978
rect 189834 472294 189890 472350
rect 189958 472294 190014 472350
rect 190082 472294 190138 472350
rect 190206 472294 190262 472350
rect 189834 472170 189890 472226
rect 189958 472170 190014 472226
rect 190082 472170 190138 472226
rect 190206 472170 190262 472226
rect 189834 472046 189890 472102
rect 189958 472046 190014 472102
rect 190082 472046 190138 472102
rect 190206 472046 190262 472102
rect 189834 471922 189890 471978
rect 189958 471922 190014 471978
rect 190082 471922 190138 471978
rect 190206 471922 190262 471978
rect 189834 454294 189890 454350
rect 189958 454294 190014 454350
rect 190082 454294 190138 454350
rect 190206 454294 190262 454350
rect 189834 454170 189890 454226
rect 189958 454170 190014 454226
rect 190082 454170 190138 454226
rect 190206 454170 190262 454226
rect 189834 454046 189890 454102
rect 189958 454046 190014 454102
rect 190082 454046 190138 454102
rect 190206 454046 190262 454102
rect 189834 453922 189890 453978
rect 189958 453922 190014 453978
rect 190082 453922 190138 453978
rect 190206 453922 190262 453978
rect 189834 436294 189890 436350
rect 189958 436294 190014 436350
rect 190082 436294 190138 436350
rect 190206 436294 190262 436350
rect 189834 436170 189890 436226
rect 189958 436170 190014 436226
rect 190082 436170 190138 436226
rect 190206 436170 190262 436226
rect 189834 436046 189890 436102
rect 189958 436046 190014 436102
rect 190082 436046 190138 436102
rect 190206 436046 190262 436102
rect 189834 435922 189890 435978
rect 189958 435922 190014 435978
rect 190082 435922 190138 435978
rect 190206 435922 190262 435978
rect 189834 418294 189890 418350
rect 189958 418294 190014 418350
rect 190082 418294 190138 418350
rect 190206 418294 190262 418350
rect 189834 418170 189890 418226
rect 189958 418170 190014 418226
rect 190082 418170 190138 418226
rect 190206 418170 190262 418226
rect 189834 418046 189890 418102
rect 189958 418046 190014 418102
rect 190082 418046 190138 418102
rect 190206 418046 190262 418102
rect 189834 417922 189890 417978
rect 189958 417922 190014 417978
rect 190082 417922 190138 417978
rect 190206 417922 190262 417978
rect 189834 400294 189890 400350
rect 189958 400294 190014 400350
rect 190082 400294 190138 400350
rect 190206 400294 190262 400350
rect 189834 400170 189890 400226
rect 189958 400170 190014 400226
rect 190082 400170 190138 400226
rect 190206 400170 190262 400226
rect 189834 400046 189890 400102
rect 189958 400046 190014 400102
rect 190082 400046 190138 400102
rect 190206 400046 190262 400102
rect 189834 399922 189890 399978
rect 189958 399922 190014 399978
rect 190082 399922 190138 399978
rect 190206 399922 190262 399978
rect 189834 382294 189890 382350
rect 189958 382294 190014 382350
rect 190082 382294 190138 382350
rect 190206 382294 190262 382350
rect 189834 382170 189890 382226
rect 189958 382170 190014 382226
rect 190082 382170 190138 382226
rect 190206 382170 190262 382226
rect 189834 382046 189890 382102
rect 189958 382046 190014 382102
rect 190082 382046 190138 382102
rect 190206 382046 190262 382102
rect 189834 381922 189890 381978
rect 189958 381922 190014 381978
rect 190082 381922 190138 381978
rect 190206 381922 190262 381978
rect 171276 366722 171332 366778
rect 164668 364922 164724 364978
rect 189834 364294 189890 364350
rect 189958 364294 190014 364350
rect 190082 364294 190138 364350
rect 190206 364294 190262 364350
rect 189834 364170 189890 364226
rect 189958 364170 190014 364226
rect 190082 364170 190138 364226
rect 190206 364170 190262 364226
rect 189834 364046 189890 364102
rect 189958 364046 190014 364102
rect 190082 364046 190138 364102
rect 190206 364046 190262 364102
rect 189834 363922 189890 363978
rect 189958 363922 190014 363978
rect 190082 363922 190138 363978
rect 190206 363922 190262 363978
rect 163436 362222 163492 362278
rect 173516 360242 173572 360298
rect 182252 358982 182308 359038
rect 166124 358622 166180 358678
rect 193554 598116 193610 598172
rect 193678 598116 193734 598172
rect 193802 598116 193858 598172
rect 193926 598116 193982 598172
rect 193554 597992 193610 598048
rect 193678 597992 193734 598048
rect 193802 597992 193858 598048
rect 193926 597992 193982 598048
rect 193554 597868 193610 597924
rect 193678 597868 193734 597924
rect 193802 597868 193858 597924
rect 193926 597868 193982 597924
rect 193554 597744 193610 597800
rect 193678 597744 193734 597800
rect 193802 597744 193858 597800
rect 193926 597744 193982 597800
rect 220554 597156 220610 597212
rect 220678 597156 220734 597212
rect 220802 597156 220858 597212
rect 220926 597156 220982 597212
rect 220554 597032 220610 597088
rect 220678 597032 220734 597088
rect 220802 597032 220858 597088
rect 220926 597032 220982 597088
rect 220554 596908 220610 596964
rect 220678 596908 220734 596964
rect 220802 596908 220858 596964
rect 220926 596908 220982 596964
rect 220554 596784 220610 596840
rect 220678 596784 220734 596840
rect 220802 596784 220858 596840
rect 220926 596784 220982 596840
rect 193554 586294 193610 586350
rect 193678 586294 193734 586350
rect 193802 586294 193858 586350
rect 193926 586294 193982 586350
rect 193554 586170 193610 586226
rect 193678 586170 193734 586226
rect 193802 586170 193858 586226
rect 193926 586170 193982 586226
rect 193554 586046 193610 586102
rect 193678 586046 193734 586102
rect 193802 586046 193858 586102
rect 193926 586046 193982 586102
rect 193554 585922 193610 585978
rect 193678 585922 193734 585978
rect 193802 585922 193858 585978
rect 193926 585922 193982 585978
rect 193554 568294 193610 568350
rect 193678 568294 193734 568350
rect 193802 568294 193858 568350
rect 193926 568294 193982 568350
rect 193554 568170 193610 568226
rect 193678 568170 193734 568226
rect 193802 568170 193858 568226
rect 193926 568170 193982 568226
rect 193554 568046 193610 568102
rect 193678 568046 193734 568102
rect 193802 568046 193858 568102
rect 193926 568046 193982 568102
rect 193554 567922 193610 567978
rect 193678 567922 193734 567978
rect 193802 567922 193858 567978
rect 193926 567922 193982 567978
rect 193554 550294 193610 550350
rect 193678 550294 193734 550350
rect 193802 550294 193858 550350
rect 193926 550294 193982 550350
rect 193554 550170 193610 550226
rect 193678 550170 193734 550226
rect 193802 550170 193858 550226
rect 193926 550170 193982 550226
rect 193554 550046 193610 550102
rect 193678 550046 193734 550102
rect 193802 550046 193858 550102
rect 193926 550046 193982 550102
rect 193554 549922 193610 549978
rect 193678 549922 193734 549978
rect 193802 549922 193858 549978
rect 193926 549922 193982 549978
rect 193554 532294 193610 532350
rect 193678 532294 193734 532350
rect 193802 532294 193858 532350
rect 193926 532294 193982 532350
rect 193554 532170 193610 532226
rect 193678 532170 193734 532226
rect 193802 532170 193858 532226
rect 193926 532170 193982 532226
rect 193554 532046 193610 532102
rect 193678 532046 193734 532102
rect 193802 532046 193858 532102
rect 193926 532046 193982 532102
rect 193554 531922 193610 531978
rect 193678 531922 193734 531978
rect 193802 531922 193858 531978
rect 193926 531922 193982 531978
rect 193554 514294 193610 514350
rect 193678 514294 193734 514350
rect 193802 514294 193858 514350
rect 193926 514294 193982 514350
rect 193554 514170 193610 514226
rect 193678 514170 193734 514226
rect 193802 514170 193858 514226
rect 193926 514170 193982 514226
rect 193554 514046 193610 514102
rect 193678 514046 193734 514102
rect 193802 514046 193858 514102
rect 193926 514046 193982 514102
rect 193554 513922 193610 513978
rect 193678 513922 193734 513978
rect 193802 513922 193858 513978
rect 193926 513922 193982 513978
rect 193554 496294 193610 496350
rect 193678 496294 193734 496350
rect 193802 496294 193858 496350
rect 193926 496294 193982 496350
rect 193554 496170 193610 496226
rect 193678 496170 193734 496226
rect 193802 496170 193858 496226
rect 193926 496170 193982 496226
rect 193554 496046 193610 496102
rect 193678 496046 193734 496102
rect 193802 496046 193858 496102
rect 193926 496046 193982 496102
rect 193554 495922 193610 495978
rect 193678 495922 193734 495978
rect 193802 495922 193858 495978
rect 193926 495922 193982 495978
rect 193554 478294 193610 478350
rect 193678 478294 193734 478350
rect 193802 478294 193858 478350
rect 193926 478294 193982 478350
rect 193554 478170 193610 478226
rect 193678 478170 193734 478226
rect 193802 478170 193858 478226
rect 193926 478170 193982 478226
rect 193554 478046 193610 478102
rect 193678 478046 193734 478102
rect 193802 478046 193858 478102
rect 193926 478046 193982 478102
rect 193554 477922 193610 477978
rect 193678 477922 193734 477978
rect 193802 477922 193858 477978
rect 193926 477922 193982 477978
rect 193554 460294 193610 460350
rect 193678 460294 193734 460350
rect 193802 460294 193858 460350
rect 193926 460294 193982 460350
rect 193554 460170 193610 460226
rect 193678 460170 193734 460226
rect 193802 460170 193858 460226
rect 193926 460170 193982 460226
rect 193554 460046 193610 460102
rect 193678 460046 193734 460102
rect 193802 460046 193858 460102
rect 193926 460046 193982 460102
rect 193554 459922 193610 459978
rect 193678 459922 193734 459978
rect 193802 459922 193858 459978
rect 193926 459922 193982 459978
rect 193554 442294 193610 442350
rect 193678 442294 193734 442350
rect 193802 442294 193858 442350
rect 193926 442294 193982 442350
rect 193554 442170 193610 442226
rect 193678 442170 193734 442226
rect 193802 442170 193858 442226
rect 193926 442170 193982 442226
rect 193554 442046 193610 442102
rect 193678 442046 193734 442102
rect 193802 442046 193858 442102
rect 193926 442046 193982 442102
rect 193554 441922 193610 441978
rect 193678 441922 193734 441978
rect 193802 441922 193858 441978
rect 193926 441922 193982 441978
rect 193554 424294 193610 424350
rect 193678 424294 193734 424350
rect 193802 424294 193858 424350
rect 193926 424294 193982 424350
rect 193554 424170 193610 424226
rect 193678 424170 193734 424226
rect 193802 424170 193858 424226
rect 193926 424170 193982 424226
rect 193554 424046 193610 424102
rect 193678 424046 193734 424102
rect 193802 424046 193858 424102
rect 193926 424046 193982 424102
rect 193554 423922 193610 423978
rect 193678 423922 193734 423978
rect 193802 423922 193858 423978
rect 193926 423922 193982 423978
rect 193554 406294 193610 406350
rect 193678 406294 193734 406350
rect 193802 406294 193858 406350
rect 193926 406294 193982 406350
rect 193554 406170 193610 406226
rect 193678 406170 193734 406226
rect 193802 406170 193858 406226
rect 193926 406170 193982 406226
rect 193554 406046 193610 406102
rect 193678 406046 193734 406102
rect 193802 406046 193858 406102
rect 193926 406046 193982 406102
rect 193554 405922 193610 405978
rect 193678 405922 193734 405978
rect 193802 405922 193858 405978
rect 193926 405922 193982 405978
rect 193554 388294 193610 388350
rect 193678 388294 193734 388350
rect 193802 388294 193858 388350
rect 193926 388294 193982 388350
rect 193554 388170 193610 388226
rect 193678 388170 193734 388226
rect 193802 388170 193858 388226
rect 193926 388170 193982 388226
rect 193554 388046 193610 388102
rect 193678 388046 193734 388102
rect 193802 388046 193858 388102
rect 193926 388046 193982 388102
rect 193554 387922 193610 387978
rect 193678 387922 193734 387978
rect 193802 387922 193858 387978
rect 193926 387922 193982 387978
rect 193554 370294 193610 370350
rect 193678 370294 193734 370350
rect 193802 370294 193858 370350
rect 193926 370294 193982 370350
rect 193554 370170 193610 370226
rect 193678 370170 193734 370226
rect 193802 370170 193858 370226
rect 193926 370170 193982 370226
rect 193554 370046 193610 370102
rect 193678 370046 193734 370102
rect 193802 370046 193858 370102
rect 193926 370046 193982 370102
rect 193554 369922 193610 369978
rect 193678 369922 193734 369978
rect 193802 369922 193858 369978
rect 193926 369922 193982 369978
rect 190988 359702 191044 359758
rect 190764 359548 190820 359578
rect 190764 359522 190820 359548
rect 189532 358802 189588 358858
rect 186956 357002 187012 357058
rect 149222 352294 149278 352350
rect 149346 352294 149402 352350
rect 149222 352170 149278 352226
rect 149346 352170 149402 352226
rect 149222 352046 149278 352102
rect 149346 352046 149402 352102
rect 149222 351922 149278 351978
rect 149346 351922 149402 351978
rect 179942 352294 179998 352350
rect 180066 352294 180122 352350
rect 179942 352170 179998 352226
rect 180066 352170 180122 352226
rect 179942 352046 179998 352102
rect 180066 352046 180122 352102
rect 179942 351922 179998 351978
rect 180066 351922 180122 351978
rect 133862 346294 133918 346350
rect 133986 346294 134042 346350
rect 133862 346170 133918 346226
rect 133986 346170 134042 346226
rect 133862 346046 133918 346102
rect 133986 346046 134042 346102
rect 133862 345922 133918 345978
rect 133986 345922 134042 345978
rect 164582 346294 164638 346350
rect 164706 346294 164762 346350
rect 164582 346170 164638 346226
rect 164706 346170 164762 346226
rect 164582 346046 164638 346102
rect 164706 346046 164762 346102
rect 164582 345922 164638 345978
rect 164706 345922 164762 345978
rect 120204 278162 120260 278218
rect 120092 271502 120148 271558
rect 120092 205802 120148 205858
rect 149222 334294 149278 334350
rect 149346 334294 149402 334350
rect 149222 334170 149278 334226
rect 149346 334170 149402 334226
rect 149222 334046 149278 334102
rect 149346 334046 149402 334102
rect 149222 333922 149278 333978
rect 149346 333922 149402 333978
rect 179942 334294 179998 334350
rect 180066 334294 180122 334350
rect 179942 334170 179998 334226
rect 180066 334170 180122 334226
rect 179942 334046 179998 334102
rect 180066 334046 180122 334102
rect 179942 333922 179998 333978
rect 180066 333922 180122 333978
rect 133862 328294 133918 328350
rect 133986 328294 134042 328350
rect 133862 328170 133918 328226
rect 133986 328170 134042 328226
rect 133862 328046 133918 328102
rect 133986 328046 134042 328102
rect 133862 327922 133918 327978
rect 133986 327922 134042 327978
rect 164582 328294 164638 328350
rect 164706 328294 164762 328350
rect 164582 328170 164638 328226
rect 164706 328170 164762 328226
rect 164582 328046 164638 328102
rect 164706 328046 164762 328102
rect 164582 327922 164638 327978
rect 164706 327922 164762 327978
rect 121772 319022 121828 319078
rect 121660 310922 121716 310978
rect 121436 283382 121492 283438
rect 121548 281762 121604 281818
rect 120540 276362 120596 276418
rect 149222 316294 149278 316350
rect 149346 316294 149402 316350
rect 149222 316170 149278 316226
rect 149346 316170 149402 316226
rect 149222 316046 149278 316102
rect 149346 316046 149402 316102
rect 149222 315922 149278 315978
rect 149346 315922 149402 315978
rect 179942 316294 179998 316350
rect 180066 316294 180122 316350
rect 179942 316170 179998 316226
rect 180066 316170 180122 316226
rect 179942 316046 179998 316102
rect 180066 316046 180122 316102
rect 179942 315922 179998 315978
rect 180066 315922 180122 315978
rect 133862 310294 133918 310350
rect 133986 310294 134042 310350
rect 133862 310170 133918 310226
rect 133986 310170 134042 310226
rect 133862 310046 133918 310102
rect 133986 310046 134042 310102
rect 133862 309922 133918 309978
rect 133986 309922 134042 309978
rect 164582 310294 164638 310350
rect 164706 310294 164762 310350
rect 164582 310170 164638 310226
rect 164706 310170 164762 310226
rect 164582 310046 164638 310102
rect 164706 310046 164762 310102
rect 164582 309922 164638 309978
rect 164706 309922 164762 309978
rect 149222 298294 149278 298350
rect 149346 298294 149402 298350
rect 149222 298170 149278 298226
rect 149346 298170 149402 298226
rect 149222 298046 149278 298102
rect 149346 298046 149402 298102
rect 149222 297922 149278 297978
rect 149346 297922 149402 297978
rect 179942 298294 179998 298350
rect 180066 298294 180122 298350
rect 179942 298170 179998 298226
rect 180066 298170 180122 298226
rect 179942 298046 179998 298102
rect 180066 298046 180122 298102
rect 179942 297922 179998 297978
rect 180066 297922 180122 297978
rect 133862 292294 133918 292350
rect 133986 292294 134042 292350
rect 133862 292170 133918 292226
rect 133986 292170 134042 292226
rect 133862 292046 133918 292102
rect 133986 292046 134042 292102
rect 133862 291922 133918 291978
rect 133986 291922 134042 291978
rect 164582 292294 164638 292350
rect 164706 292294 164762 292350
rect 164582 292170 164638 292226
rect 164706 292170 164762 292226
rect 164582 292046 164638 292102
rect 164706 292046 164762 292102
rect 164582 291922 164638 291978
rect 164706 291922 164762 291978
rect 121884 284642 121940 284698
rect 141036 283202 141092 283258
rect 139692 283022 139748 283078
rect 122332 282302 122388 282358
rect 127708 281582 127764 281638
rect 133644 281402 133700 281458
rect 128394 274294 128450 274350
rect 128518 274294 128574 274350
rect 128642 274294 128698 274350
rect 128766 274294 128822 274350
rect 128394 274170 128450 274226
rect 128518 274170 128574 274226
rect 128642 274170 128698 274226
rect 128766 274170 128822 274226
rect 128394 274046 128450 274102
rect 128518 274046 128574 274102
rect 128642 274046 128698 274102
rect 128766 274046 128822 274102
rect 128394 273922 128450 273978
rect 128518 273922 128574 273978
rect 128642 273922 128698 273978
rect 128766 273922 128822 273978
rect 127596 265022 127652 265078
rect 126812 178082 126868 178138
rect 126252 162782 126308 162838
rect 128394 256294 128450 256350
rect 128518 256294 128574 256350
rect 128642 256294 128698 256350
rect 128766 256294 128822 256350
rect 128394 256170 128450 256226
rect 128518 256170 128574 256226
rect 128642 256170 128698 256226
rect 128766 256170 128822 256226
rect 128394 256046 128450 256102
rect 128518 256046 128574 256102
rect 128642 256046 128698 256102
rect 128766 256046 128822 256102
rect 128394 255922 128450 255978
rect 128518 255922 128574 255978
rect 128642 255922 128698 255978
rect 128766 255922 128822 255978
rect 128394 238294 128450 238350
rect 128518 238294 128574 238350
rect 128642 238294 128698 238350
rect 128766 238294 128822 238350
rect 128394 238170 128450 238226
rect 128518 238170 128574 238226
rect 128642 238170 128698 238226
rect 128766 238170 128822 238226
rect 128394 238046 128450 238102
rect 128518 238046 128574 238102
rect 128642 238046 128698 238102
rect 128766 238046 128822 238102
rect 128394 237922 128450 237978
rect 128518 237922 128574 237978
rect 128642 237922 128698 237978
rect 128766 237922 128822 237978
rect 128394 220294 128450 220350
rect 128518 220294 128574 220350
rect 128642 220294 128698 220350
rect 128766 220294 128822 220350
rect 128394 220170 128450 220226
rect 128518 220170 128574 220226
rect 128642 220170 128698 220226
rect 128766 220170 128822 220226
rect 128394 220046 128450 220102
rect 128518 220046 128574 220102
rect 128642 220046 128698 220102
rect 128766 220046 128822 220102
rect 128394 219922 128450 219978
rect 128518 219922 128574 219978
rect 128642 219922 128698 219978
rect 128766 219922 128822 219978
rect 128394 202294 128450 202350
rect 128518 202294 128574 202350
rect 128642 202294 128698 202350
rect 128766 202294 128822 202350
rect 128394 202170 128450 202226
rect 128518 202170 128574 202226
rect 128642 202170 128698 202226
rect 128766 202170 128822 202226
rect 128394 202046 128450 202102
rect 128518 202046 128574 202102
rect 128642 202046 128698 202102
rect 128766 202046 128822 202102
rect 128394 201922 128450 201978
rect 128518 201922 128574 201978
rect 128642 201922 128698 201978
rect 128766 201922 128822 201978
rect 128394 184294 128450 184350
rect 128518 184294 128574 184350
rect 128642 184294 128698 184350
rect 128766 184294 128822 184350
rect 128394 184170 128450 184226
rect 128518 184170 128574 184226
rect 128642 184170 128698 184226
rect 128766 184170 128822 184226
rect 128394 184046 128450 184102
rect 128518 184046 128574 184102
rect 128642 184046 128698 184102
rect 128766 184046 128822 184102
rect 128394 183922 128450 183978
rect 128518 183922 128574 183978
rect 128642 183922 128698 183978
rect 128766 183922 128822 183978
rect 146412 282122 146468 282178
rect 163660 281942 163716 281998
rect 132114 280294 132170 280350
rect 132238 280294 132294 280350
rect 132362 280294 132418 280350
rect 132486 280294 132542 280350
rect 132114 280170 132170 280226
rect 132238 280170 132294 280226
rect 132362 280170 132418 280226
rect 132486 280170 132542 280226
rect 132114 280046 132170 280102
rect 132238 280046 132294 280102
rect 132362 280046 132418 280102
rect 132486 280046 132542 280102
rect 132114 279922 132170 279978
rect 132238 279922 132294 279978
rect 132362 279922 132418 279978
rect 132486 279922 132542 279978
rect 137004 277982 137060 278038
rect 132114 262294 132170 262350
rect 132238 262294 132294 262350
rect 132362 262294 132418 262350
rect 132486 262294 132542 262350
rect 132114 262170 132170 262226
rect 132238 262170 132294 262226
rect 132362 262170 132418 262226
rect 132486 262170 132542 262226
rect 132114 262046 132170 262102
rect 132238 262046 132294 262102
rect 132362 262046 132418 262102
rect 132486 262046 132542 262102
rect 132114 261922 132170 261978
rect 132238 261922 132294 261978
rect 132362 261922 132418 261978
rect 132486 261922 132542 261978
rect 132114 244294 132170 244350
rect 132238 244294 132294 244350
rect 132362 244294 132418 244350
rect 132486 244294 132542 244350
rect 132114 244170 132170 244226
rect 132238 244170 132294 244226
rect 132362 244170 132418 244226
rect 132486 244170 132542 244226
rect 132114 244046 132170 244102
rect 132238 244046 132294 244102
rect 132362 244046 132418 244102
rect 132486 244046 132542 244102
rect 132114 243922 132170 243978
rect 132238 243922 132294 243978
rect 132362 243922 132418 243978
rect 132486 243922 132542 243978
rect 132114 226294 132170 226350
rect 132238 226294 132294 226350
rect 132362 226294 132418 226350
rect 132486 226294 132542 226350
rect 132114 226170 132170 226226
rect 132238 226170 132294 226226
rect 132362 226170 132418 226226
rect 132486 226170 132542 226226
rect 132114 226046 132170 226102
rect 132238 226046 132294 226102
rect 132362 226046 132418 226102
rect 132486 226046 132542 226102
rect 132114 225922 132170 225978
rect 132238 225922 132294 225978
rect 132362 225922 132418 225978
rect 132486 225922 132542 225978
rect 132114 208294 132170 208350
rect 132238 208294 132294 208350
rect 132362 208294 132418 208350
rect 132486 208294 132542 208350
rect 132114 208170 132170 208226
rect 132238 208170 132294 208226
rect 132362 208170 132418 208226
rect 132486 208170 132542 208226
rect 132114 208046 132170 208102
rect 132238 208046 132294 208102
rect 132362 208046 132418 208102
rect 132486 208046 132542 208102
rect 132114 207922 132170 207978
rect 132238 207922 132294 207978
rect 132362 207922 132418 207978
rect 132486 207922 132542 207978
rect 132114 190294 132170 190350
rect 132238 190294 132294 190350
rect 132362 190294 132418 190350
rect 132486 190294 132542 190350
rect 132114 190170 132170 190226
rect 132238 190170 132294 190226
rect 132362 190170 132418 190226
rect 132486 190170 132542 190226
rect 132114 190046 132170 190102
rect 132238 190046 132294 190102
rect 132362 190046 132418 190102
rect 132486 190046 132542 190102
rect 132114 189922 132170 189978
rect 132238 189922 132294 189978
rect 132362 189922 132418 189978
rect 132486 189922 132542 189978
rect 128394 166294 128450 166350
rect 128518 166294 128574 166350
rect 128642 166294 128698 166350
rect 128766 166294 128822 166350
rect 128394 166170 128450 166226
rect 128518 166170 128574 166226
rect 128642 166170 128698 166226
rect 128766 166170 128822 166226
rect 128394 166046 128450 166102
rect 128518 166046 128574 166102
rect 128642 166046 128698 166102
rect 128766 166046 128822 166102
rect 128394 165922 128450 165978
rect 128518 165922 128574 165978
rect 128642 165922 128698 165978
rect 128766 165922 128822 165978
rect 129052 176462 129108 176518
rect 132114 172294 132170 172350
rect 132238 172294 132294 172350
rect 132362 172294 132418 172350
rect 132486 172294 132542 172350
rect 132114 172170 132170 172226
rect 132238 172170 132294 172226
rect 132362 172170 132418 172226
rect 132486 172170 132542 172226
rect 132114 172046 132170 172102
rect 132238 172046 132294 172102
rect 132362 172046 132418 172102
rect 132486 172046 132542 172102
rect 132114 171922 132170 171978
rect 132238 171922 132294 171978
rect 132362 171922 132418 171978
rect 132486 171922 132542 171978
rect 128394 148294 128450 148350
rect 128518 148294 128574 148350
rect 128642 148294 128698 148350
rect 128766 148294 128822 148350
rect 128394 148170 128450 148226
rect 128518 148170 128574 148226
rect 128642 148170 128698 148226
rect 128766 148170 128822 148226
rect 128394 148046 128450 148102
rect 128518 148046 128574 148102
rect 128642 148046 128698 148102
rect 128766 148046 128822 148102
rect 128394 147922 128450 147978
rect 128518 147922 128574 147978
rect 128642 147922 128698 147978
rect 128766 147922 128822 147978
rect 111930 136294 111986 136350
rect 112054 136294 112110 136350
rect 112178 136294 112234 136350
rect 112302 136294 112358 136350
rect 111930 136170 111986 136226
rect 112054 136170 112110 136226
rect 112178 136170 112234 136226
rect 112302 136170 112358 136226
rect 111930 136046 111986 136102
rect 112054 136046 112110 136102
rect 112178 136046 112234 136102
rect 112302 136046 112358 136102
rect 111930 135922 111986 135978
rect 112054 135922 112110 135978
rect 112178 135922 112234 135978
rect 112302 135922 112358 135978
rect 111130 130294 111186 130350
rect 111254 130294 111310 130350
rect 111378 130294 111434 130350
rect 111502 130294 111558 130350
rect 111130 130170 111186 130226
rect 111254 130170 111310 130226
rect 111378 130170 111434 130226
rect 111502 130170 111558 130226
rect 111130 130046 111186 130102
rect 111254 130046 111310 130102
rect 111378 130046 111434 130102
rect 111502 130046 111558 130102
rect 111130 129922 111186 129978
rect 111254 129922 111310 129978
rect 111378 129922 111434 129978
rect 111502 129922 111558 129978
rect 128394 130294 128450 130350
rect 128518 130294 128574 130350
rect 128642 130294 128698 130350
rect 128766 130294 128822 130350
rect 128394 130170 128450 130226
rect 128518 130170 128574 130226
rect 128642 130170 128698 130226
rect 128766 130170 128822 130226
rect 128394 130046 128450 130102
rect 128518 130046 128574 130102
rect 128642 130046 128698 130102
rect 128766 130046 128822 130102
rect 128394 129922 128450 129978
rect 128518 129922 128574 129978
rect 128642 129922 128698 129978
rect 128766 129922 128822 129978
rect 111930 118294 111986 118350
rect 112054 118294 112110 118350
rect 112178 118294 112234 118350
rect 112302 118294 112358 118350
rect 111930 118170 111986 118226
rect 112054 118170 112110 118226
rect 112178 118170 112234 118226
rect 112302 118170 112358 118226
rect 111930 118046 111986 118102
rect 112054 118046 112110 118102
rect 112178 118046 112234 118102
rect 112302 118046 112358 118102
rect 111930 117922 111986 117978
rect 112054 117922 112110 117978
rect 112178 117922 112234 117978
rect 112302 117922 112358 117978
rect 111130 112294 111186 112350
rect 111254 112294 111310 112350
rect 111378 112294 111434 112350
rect 111502 112294 111558 112350
rect 111130 112170 111186 112226
rect 111254 112170 111310 112226
rect 111378 112170 111434 112226
rect 111502 112170 111558 112226
rect 111130 112046 111186 112102
rect 111254 112046 111310 112102
rect 111378 112046 111434 112102
rect 111502 112046 111558 112102
rect 111130 111922 111186 111978
rect 111254 111922 111310 111978
rect 111378 111922 111434 111978
rect 111502 111922 111558 111978
rect 128394 112294 128450 112350
rect 128518 112294 128574 112350
rect 128642 112294 128698 112350
rect 128766 112294 128822 112350
rect 128394 112170 128450 112226
rect 128518 112170 128574 112226
rect 128642 112170 128698 112226
rect 128766 112170 128822 112226
rect 128394 112046 128450 112102
rect 128518 112046 128574 112102
rect 128642 112046 128698 112102
rect 128766 112046 128822 112102
rect 128394 111922 128450 111978
rect 128518 111922 128574 111978
rect 128642 111922 128698 111978
rect 128766 111922 128822 111978
rect 111930 100294 111986 100350
rect 112054 100294 112110 100350
rect 112178 100294 112234 100350
rect 112302 100294 112358 100350
rect 111930 100170 111986 100226
rect 112054 100170 112110 100226
rect 112178 100170 112234 100226
rect 112302 100170 112358 100226
rect 111930 100046 111986 100102
rect 112054 100046 112110 100102
rect 112178 100046 112234 100102
rect 112302 100046 112358 100102
rect 111930 99922 111986 99978
rect 112054 99922 112110 99978
rect 112178 99922 112234 99978
rect 112302 99922 112358 99978
rect 111130 94294 111186 94350
rect 111254 94294 111310 94350
rect 111378 94294 111434 94350
rect 111502 94294 111558 94350
rect 111130 94170 111186 94226
rect 111254 94170 111310 94226
rect 111378 94170 111434 94226
rect 111502 94170 111558 94226
rect 111130 94046 111186 94102
rect 111254 94046 111310 94102
rect 111378 94046 111434 94102
rect 111502 94046 111558 94102
rect 111130 93922 111186 93978
rect 111254 93922 111310 93978
rect 111378 93922 111434 93978
rect 111502 93922 111558 93978
rect 128394 94294 128450 94350
rect 128518 94294 128574 94350
rect 128642 94294 128698 94350
rect 128766 94294 128822 94350
rect 128394 94170 128450 94226
rect 128518 94170 128574 94226
rect 128642 94170 128698 94226
rect 128766 94170 128822 94226
rect 128394 94046 128450 94102
rect 128518 94046 128574 94102
rect 128642 94046 128698 94102
rect 128766 94046 128822 94102
rect 128394 93922 128450 93978
rect 128518 93922 128574 93978
rect 128642 93922 128698 93978
rect 128766 93922 128822 93978
rect 111930 82294 111986 82350
rect 112054 82294 112110 82350
rect 112178 82294 112234 82350
rect 112302 82294 112358 82350
rect 111930 82170 111986 82226
rect 112054 82170 112110 82226
rect 112178 82170 112234 82226
rect 112302 82170 112358 82226
rect 111930 82046 111986 82102
rect 112054 82046 112110 82102
rect 112178 82046 112234 82102
rect 112302 82046 112358 82102
rect 111930 81922 111986 81978
rect 112054 81922 112110 81978
rect 112178 81922 112234 81978
rect 112302 81922 112358 81978
rect 111130 76294 111186 76350
rect 111254 76294 111310 76350
rect 111378 76294 111434 76350
rect 111502 76294 111558 76350
rect 111130 76170 111186 76226
rect 111254 76170 111310 76226
rect 111378 76170 111434 76226
rect 111502 76170 111558 76226
rect 111130 76046 111186 76102
rect 111254 76046 111310 76102
rect 111378 76046 111434 76102
rect 111502 76046 111558 76102
rect 111130 75922 111186 75978
rect 111254 75922 111310 75978
rect 111378 75922 111434 75978
rect 111502 75922 111558 75978
rect 128394 76294 128450 76350
rect 128518 76294 128574 76350
rect 128642 76294 128698 76350
rect 128766 76294 128822 76350
rect 128394 76170 128450 76226
rect 128518 76170 128574 76226
rect 128642 76170 128698 76226
rect 128766 76170 128822 76226
rect 128394 76046 128450 76102
rect 128518 76046 128574 76102
rect 128642 76046 128698 76102
rect 128766 76046 128822 76102
rect 128394 75922 128450 75978
rect 128518 75922 128574 75978
rect 128642 75922 128698 75978
rect 128766 75922 128822 75978
rect 111930 64294 111986 64350
rect 112054 64294 112110 64350
rect 112178 64294 112234 64350
rect 112302 64294 112358 64350
rect 111930 64170 111986 64226
rect 112054 64170 112110 64226
rect 112178 64170 112234 64226
rect 112302 64170 112358 64226
rect 111930 64046 111986 64102
rect 112054 64046 112110 64102
rect 112178 64046 112234 64102
rect 112302 64046 112358 64102
rect 111930 63922 111986 63978
rect 112054 63922 112110 63978
rect 112178 63922 112234 63978
rect 112302 63922 112358 63978
rect 111130 58294 111186 58350
rect 111254 58294 111310 58350
rect 111378 58294 111434 58350
rect 111502 58294 111558 58350
rect 111130 58170 111186 58226
rect 111254 58170 111310 58226
rect 111378 58170 111434 58226
rect 111502 58170 111558 58226
rect 111130 58046 111186 58102
rect 111254 58046 111310 58102
rect 111378 58046 111434 58102
rect 111502 58046 111558 58102
rect 111130 57922 111186 57978
rect 111254 57922 111310 57978
rect 111378 57922 111434 57978
rect 111502 57922 111558 57978
rect 128394 58294 128450 58350
rect 128518 58294 128574 58350
rect 128642 58294 128698 58350
rect 128766 58294 128822 58350
rect 128394 58170 128450 58226
rect 128518 58170 128574 58226
rect 128642 58170 128698 58226
rect 128766 58170 128822 58226
rect 128394 58046 128450 58102
rect 128518 58046 128574 58102
rect 128642 58046 128698 58102
rect 128766 58046 128822 58102
rect 128394 57922 128450 57978
rect 128518 57922 128574 57978
rect 128642 57922 128698 57978
rect 128766 57922 128822 57978
rect 128394 40294 128450 40350
rect 128518 40294 128574 40350
rect 128642 40294 128698 40350
rect 128766 40294 128822 40350
rect 128394 40170 128450 40226
rect 128518 40170 128574 40226
rect 128642 40170 128698 40226
rect 128766 40170 128822 40226
rect 128394 40046 128450 40102
rect 128518 40046 128574 40102
rect 128642 40046 128698 40102
rect 128766 40046 128822 40102
rect 128394 39922 128450 39978
rect 128518 39922 128574 39978
rect 128642 39922 128698 39978
rect 128766 39922 128822 39978
rect 101394 28294 101450 28350
rect 101518 28294 101574 28350
rect 101642 28294 101698 28350
rect 101766 28294 101822 28350
rect 101394 28170 101450 28226
rect 101518 28170 101574 28226
rect 101642 28170 101698 28226
rect 101766 28170 101822 28226
rect 101394 28046 101450 28102
rect 101518 28046 101574 28102
rect 101642 28046 101698 28102
rect 101766 28046 101822 28102
rect 101394 27922 101450 27978
rect 101518 27922 101574 27978
rect 101642 27922 101698 27978
rect 101766 27922 101822 27978
rect 101394 10294 101450 10350
rect 101518 10294 101574 10350
rect 101642 10294 101698 10350
rect 101766 10294 101822 10350
rect 101394 10170 101450 10226
rect 101518 10170 101574 10226
rect 101642 10170 101698 10226
rect 101766 10170 101822 10226
rect 101394 10046 101450 10102
rect 101518 10046 101574 10102
rect 101642 10046 101698 10102
rect 101766 10046 101822 10102
rect 101394 9922 101450 9978
rect 101518 9922 101574 9978
rect 101642 9922 101698 9978
rect 101766 9922 101822 9978
rect 101394 -1176 101450 -1120
rect 101518 -1176 101574 -1120
rect 101642 -1176 101698 -1120
rect 101766 -1176 101822 -1120
rect 101394 -1300 101450 -1244
rect 101518 -1300 101574 -1244
rect 101642 -1300 101698 -1244
rect 101766 -1300 101822 -1244
rect 101394 -1424 101450 -1368
rect 101518 -1424 101574 -1368
rect 101642 -1424 101698 -1368
rect 101766 -1424 101822 -1368
rect 101394 -1548 101450 -1492
rect 101518 -1548 101574 -1492
rect 101642 -1548 101698 -1492
rect 101766 -1548 101822 -1492
rect 128394 22294 128450 22350
rect 128518 22294 128574 22350
rect 128642 22294 128698 22350
rect 128766 22294 128822 22350
rect 128394 22170 128450 22226
rect 128518 22170 128574 22226
rect 128642 22170 128698 22226
rect 128766 22170 128822 22226
rect 128394 22046 128450 22102
rect 128518 22046 128574 22102
rect 128642 22046 128698 22102
rect 128766 22046 128822 22102
rect 128394 21922 128450 21978
rect 128518 21922 128574 21978
rect 128642 21922 128698 21978
rect 128766 21922 128822 21978
rect 128394 4294 128450 4350
rect 128518 4294 128574 4350
rect 128642 4294 128698 4350
rect 128766 4294 128822 4350
rect 128394 4170 128450 4226
rect 128518 4170 128574 4226
rect 128642 4170 128698 4226
rect 128766 4170 128822 4226
rect 128394 4046 128450 4102
rect 128518 4046 128574 4102
rect 128642 4046 128698 4102
rect 128766 4046 128822 4102
rect 128394 3922 128450 3978
rect 128518 3922 128574 3978
rect 128642 3922 128698 3978
rect 128766 3922 128822 3978
rect 128394 -216 128450 -160
rect 128518 -216 128574 -160
rect 128642 -216 128698 -160
rect 128766 -216 128822 -160
rect 128394 -340 128450 -284
rect 128518 -340 128574 -284
rect 128642 -340 128698 -284
rect 128766 -340 128822 -284
rect 128394 -464 128450 -408
rect 128518 -464 128574 -408
rect 128642 -464 128698 -408
rect 128766 -464 128822 -408
rect 128394 -588 128450 -532
rect 128518 -588 128574 -532
rect 128642 -588 128698 -532
rect 128766 -588 128822 -532
rect 132114 154294 132170 154350
rect 132238 154294 132294 154350
rect 132362 154294 132418 154350
rect 132486 154294 132542 154350
rect 132114 154170 132170 154226
rect 132238 154170 132294 154226
rect 132362 154170 132418 154226
rect 132486 154170 132542 154226
rect 132114 154046 132170 154102
rect 132238 154046 132294 154102
rect 132362 154046 132418 154102
rect 132486 154046 132542 154102
rect 132114 153922 132170 153978
rect 132238 153922 132294 153978
rect 132362 153922 132418 153978
rect 132486 153922 132542 153978
rect 155372 278522 155428 278578
rect 151116 276362 151172 276418
rect 138572 173042 138628 173098
rect 157948 276542 158004 276598
rect 162834 280294 162890 280350
rect 162958 280294 163014 280350
rect 163082 280294 163138 280350
rect 163206 280294 163262 280350
rect 162834 280170 162890 280226
rect 162958 280170 163014 280226
rect 163082 280170 163138 280226
rect 163206 280170 163262 280226
rect 162834 280046 162890 280102
rect 162958 280046 163014 280102
rect 163082 280046 163138 280102
rect 163206 280046 163262 280102
rect 162834 279922 162890 279978
rect 162958 279922 163014 279978
rect 163082 279922 163138 279978
rect 163206 279922 163262 279978
rect 159964 276722 160020 276778
rect 159114 274294 159170 274350
rect 159238 274294 159294 274350
rect 159362 274294 159418 274350
rect 159486 274294 159542 274350
rect 159114 274170 159170 274226
rect 159238 274170 159294 274226
rect 159362 274170 159418 274226
rect 159486 274170 159542 274226
rect 159114 274046 159170 274102
rect 159238 274046 159294 274102
rect 159362 274046 159418 274102
rect 159486 274046 159542 274102
rect 159114 273922 159170 273978
rect 159238 273922 159294 273978
rect 159362 273922 159418 273978
rect 159486 273922 159542 273978
rect 159114 256294 159170 256350
rect 159238 256294 159294 256350
rect 159362 256294 159418 256350
rect 159486 256294 159542 256350
rect 159114 256170 159170 256226
rect 159238 256170 159294 256226
rect 159362 256170 159418 256226
rect 159486 256170 159542 256226
rect 159114 256046 159170 256102
rect 159238 256046 159294 256102
rect 159362 256046 159418 256102
rect 159486 256046 159542 256102
rect 159114 255922 159170 255978
rect 159238 255922 159294 255978
rect 159362 255922 159418 255978
rect 159486 255922 159542 255978
rect 159114 238294 159170 238350
rect 159238 238294 159294 238350
rect 159362 238294 159418 238350
rect 159486 238294 159542 238350
rect 159114 238170 159170 238226
rect 159238 238170 159294 238226
rect 159362 238170 159418 238226
rect 159486 238170 159542 238226
rect 159114 238046 159170 238102
rect 159238 238046 159294 238102
rect 159362 238046 159418 238102
rect 159486 238046 159542 238102
rect 159114 237922 159170 237978
rect 159238 237922 159294 237978
rect 159362 237922 159418 237978
rect 159486 237922 159542 237978
rect 159114 220294 159170 220350
rect 159238 220294 159294 220350
rect 159362 220294 159418 220350
rect 159486 220294 159542 220350
rect 159114 220170 159170 220226
rect 159238 220170 159294 220226
rect 159362 220170 159418 220226
rect 159486 220170 159542 220226
rect 159114 220046 159170 220102
rect 159238 220046 159294 220102
rect 159362 220046 159418 220102
rect 159486 220046 159542 220102
rect 159114 219922 159170 219978
rect 159238 219922 159294 219978
rect 159362 219922 159418 219978
rect 159486 219922 159542 219978
rect 159114 202294 159170 202350
rect 159238 202294 159294 202350
rect 159362 202294 159418 202350
rect 159486 202294 159542 202350
rect 159114 202170 159170 202226
rect 159238 202170 159294 202226
rect 159362 202170 159418 202226
rect 159486 202170 159542 202226
rect 159114 202046 159170 202102
rect 159238 202046 159294 202102
rect 159362 202046 159418 202102
rect 159486 202046 159542 202102
rect 159114 201922 159170 201978
rect 159238 201922 159294 201978
rect 159362 201922 159418 201978
rect 159486 201922 159542 201978
rect 159114 184294 159170 184350
rect 159238 184294 159294 184350
rect 159362 184294 159418 184350
rect 159486 184294 159542 184350
rect 159114 184170 159170 184226
rect 159238 184170 159294 184226
rect 159362 184170 159418 184226
rect 159486 184170 159542 184226
rect 159114 184046 159170 184102
rect 159238 184046 159294 184102
rect 159362 184046 159418 184102
rect 159486 184046 159542 184102
rect 159114 183922 159170 183978
rect 159238 183922 159294 183978
rect 159362 183922 159418 183978
rect 159486 183922 159542 183978
rect 159114 166294 159170 166350
rect 159238 166294 159294 166350
rect 159362 166294 159418 166350
rect 159486 166294 159542 166350
rect 159114 166170 159170 166226
rect 159238 166170 159294 166226
rect 159362 166170 159418 166226
rect 159486 166170 159542 166226
rect 159114 166046 159170 166102
rect 159238 166046 159294 166102
rect 159362 166046 159418 166102
rect 159486 166046 159542 166102
rect 159114 165922 159170 165978
rect 159238 165922 159294 165978
rect 159362 165922 159418 165978
rect 159486 165922 159542 165978
rect 160524 257822 160580 257878
rect 165228 276902 165284 276958
rect 163772 266642 163828 266698
rect 162834 262294 162890 262350
rect 162958 262294 163014 262350
rect 163082 262294 163138 262350
rect 163206 262294 163262 262350
rect 162834 262170 162890 262226
rect 162958 262170 163014 262226
rect 163082 262170 163138 262226
rect 163206 262170 163262 262226
rect 162834 262046 162890 262102
rect 162958 262046 163014 262102
rect 163082 262046 163138 262102
rect 163206 262046 163262 262102
rect 162834 261922 162890 261978
rect 162958 261922 163014 261978
rect 163082 261922 163138 261978
rect 163206 261922 163262 261978
rect 162834 244294 162890 244350
rect 162958 244294 163014 244350
rect 163082 244294 163138 244350
rect 163206 244294 163262 244350
rect 162834 244170 162890 244226
rect 162958 244170 163014 244226
rect 163082 244170 163138 244226
rect 163206 244170 163262 244226
rect 162834 244046 162890 244102
rect 162958 244046 163014 244102
rect 163082 244046 163138 244102
rect 163206 244046 163262 244102
rect 162834 243922 162890 243978
rect 162958 243922 163014 243978
rect 163082 243922 163138 243978
rect 163206 243922 163262 243978
rect 162834 226294 162890 226350
rect 162958 226294 163014 226350
rect 163082 226294 163138 226350
rect 163206 226294 163262 226350
rect 162834 226170 162890 226226
rect 162958 226170 163014 226226
rect 163082 226170 163138 226226
rect 163206 226170 163262 226226
rect 162834 226046 162890 226102
rect 162958 226046 163014 226102
rect 163082 226046 163138 226102
rect 163206 226046 163262 226102
rect 162834 225922 162890 225978
rect 162958 225922 163014 225978
rect 163082 225922 163138 225978
rect 163206 225922 163262 225978
rect 160524 214082 160580 214138
rect 162834 208294 162890 208350
rect 162958 208294 163014 208350
rect 163082 208294 163138 208350
rect 163206 208294 163262 208350
rect 162834 208170 162890 208226
rect 162958 208170 163014 208226
rect 163082 208170 163138 208226
rect 163206 208170 163262 208226
rect 162834 208046 162890 208102
rect 162958 208046 163014 208102
rect 163082 208046 163138 208102
rect 163206 208046 163262 208102
rect 162834 207922 162890 207978
rect 162958 207922 163014 207978
rect 163082 207922 163138 207978
rect 163206 207922 163262 207978
rect 162834 190294 162890 190350
rect 162958 190294 163014 190350
rect 163082 190294 163138 190350
rect 163206 190294 163262 190350
rect 162834 190170 162890 190226
rect 162958 190170 163014 190226
rect 163082 190170 163138 190226
rect 163206 190170 163262 190226
rect 162834 190046 162890 190102
rect 162958 190046 163014 190102
rect 163082 190046 163138 190102
rect 163206 190046 163262 190102
rect 162834 189922 162890 189978
rect 162958 189922 163014 189978
rect 163082 189922 163138 189978
rect 163206 189922 163262 189978
rect 162834 172294 162890 172350
rect 162958 172294 163014 172350
rect 163082 172294 163138 172350
rect 163206 172294 163262 172350
rect 162834 172170 162890 172226
rect 162958 172170 163014 172226
rect 163082 172170 163138 172226
rect 163206 172170 163262 172226
rect 162834 172046 162890 172102
rect 162958 172046 163014 172102
rect 163082 172046 163138 172102
rect 163206 172046 163262 172102
rect 162834 171922 162890 171978
rect 162958 171922 163014 171978
rect 163082 171922 163138 171978
rect 163206 171922 163262 171978
rect 159114 148294 159170 148350
rect 159238 148294 159294 148350
rect 159362 148294 159418 148350
rect 159486 148294 159542 148350
rect 159114 148170 159170 148226
rect 159238 148170 159294 148226
rect 159362 148170 159418 148226
rect 159486 148170 159542 148226
rect 159114 148046 159170 148102
rect 159238 148046 159294 148102
rect 159362 148046 159418 148102
rect 159486 148046 159542 148102
rect 159114 147922 159170 147978
rect 159238 147922 159294 147978
rect 159362 147922 159418 147978
rect 159486 147922 159542 147978
rect 132114 136294 132170 136350
rect 132238 136294 132294 136350
rect 132362 136294 132418 136350
rect 132486 136294 132542 136350
rect 132114 136170 132170 136226
rect 132238 136170 132294 136226
rect 132362 136170 132418 136226
rect 132486 136170 132542 136226
rect 132114 136046 132170 136102
rect 132238 136046 132294 136102
rect 132362 136046 132418 136102
rect 132486 136046 132542 136102
rect 132114 135922 132170 135978
rect 132238 135922 132294 135978
rect 132362 135922 132418 135978
rect 132486 135922 132542 135978
rect 132114 118294 132170 118350
rect 132238 118294 132294 118350
rect 132362 118294 132418 118350
rect 132486 118294 132542 118350
rect 132114 118170 132170 118226
rect 132238 118170 132294 118226
rect 132362 118170 132418 118226
rect 132486 118170 132542 118226
rect 132114 118046 132170 118102
rect 132238 118046 132294 118102
rect 132362 118046 132418 118102
rect 132486 118046 132542 118102
rect 132114 117922 132170 117978
rect 132238 117922 132294 117978
rect 132362 117922 132418 117978
rect 132486 117922 132542 117978
rect 132114 100294 132170 100350
rect 132238 100294 132294 100350
rect 132362 100294 132418 100350
rect 132486 100294 132542 100350
rect 132114 100170 132170 100226
rect 132238 100170 132294 100226
rect 132362 100170 132418 100226
rect 132486 100170 132542 100226
rect 132114 100046 132170 100102
rect 132238 100046 132294 100102
rect 132362 100046 132418 100102
rect 132486 100046 132542 100102
rect 132114 99922 132170 99978
rect 132238 99922 132294 99978
rect 132362 99922 132418 99978
rect 132486 99922 132542 99978
rect 132114 82294 132170 82350
rect 132238 82294 132294 82350
rect 132362 82294 132418 82350
rect 132486 82294 132542 82350
rect 132114 82170 132170 82226
rect 132238 82170 132294 82226
rect 132362 82170 132418 82226
rect 132486 82170 132542 82226
rect 132114 82046 132170 82102
rect 132238 82046 132294 82102
rect 132362 82046 132418 82102
rect 132486 82046 132542 82102
rect 132114 81922 132170 81978
rect 132238 81922 132294 81978
rect 132362 81922 132418 81978
rect 132486 81922 132542 81978
rect 132114 64294 132170 64350
rect 132238 64294 132294 64350
rect 132362 64294 132418 64350
rect 132486 64294 132542 64350
rect 132114 64170 132170 64226
rect 132238 64170 132294 64226
rect 132362 64170 132418 64226
rect 132486 64170 132542 64226
rect 132114 64046 132170 64102
rect 132238 64046 132294 64102
rect 132362 64046 132418 64102
rect 132486 64046 132542 64102
rect 132114 63922 132170 63978
rect 132238 63922 132294 63978
rect 132362 63922 132418 63978
rect 132486 63922 132542 63978
rect 132114 46294 132170 46350
rect 132238 46294 132294 46350
rect 132362 46294 132418 46350
rect 132486 46294 132542 46350
rect 132114 46170 132170 46226
rect 132238 46170 132294 46226
rect 132362 46170 132418 46226
rect 132486 46170 132542 46226
rect 132114 46046 132170 46102
rect 132238 46046 132294 46102
rect 132362 46046 132418 46102
rect 132486 46046 132542 46102
rect 132114 45922 132170 45978
rect 132238 45922 132294 45978
rect 132362 45922 132418 45978
rect 132486 45922 132542 45978
rect 159114 130294 159170 130350
rect 159238 130294 159294 130350
rect 159362 130294 159418 130350
rect 159486 130294 159542 130350
rect 159114 130170 159170 130226
rect 159238 130170 159294 130226
rect 159362 130170 159418 130226
rect 159486 130170 159542 130226
rect 159114 130046 159170 130102
rect 159238 130046 159294 130102
rect 159362 130046 159418 130102
rect 159486 130046 159542 130102
rect 159114 129922 159170 129978
rect 159238 129922 159294 129978
rect 159362 129922 159418 129978
rect 159486 129922 159542 129978
rect 159114 112294 159170 112350
rect 159238 112294 159294 112350
rect 159362 112294 159418 112350
rect 159486 112294 159542 112350
rect 159114 112170 159170 112226
rect 159238 112170 159294 112226
rect 159362 112170 159418 112226
rect 159486 112170 159542 112226
rect 159114 112046 159170 112102
rect 159238 112046 159294 112102
rect 159362 112046 159418 112102
rect 159486 112046 159542 112102
rect 159114 111922 159170 111978
rect 159238 111922 159294 111978
rect 159362 111922 159418 111978
rect 159486 111922 159542 111978
rect 159114 94294 159170 94350
rect 159238 94294 159294 94350
rect 159362 94294 159418 94350
rect 159486 94294 159542 94350
rect 159114 94170 159170 94226
rect 159238 94170 159294 94226
rect 159362 94170 159418 94226
rect 159486 94170 159542 94226
rect 159114 94046 159170 94102
rect 159238 94046 159294 94102
rect 159362 94046 159418 94102
rect 159486 94046 159542 94102
rect 159114 93922 159170 93978
rect 159238 93922 159294 93978
rect 159362 93922 159418 93978
rect 159486 93922 159542 93978
rect 159114 76294 159170 76350
rect 159238 76294 159294 76350
rect 159362 76294 159418 76350
rect 159486 76294 159542 76350
rect 159114 76170 159170 76226
rect 159238 76170 159294 76226
rect 159362 76170 159418 76226
rect 159486 76170 159542 76226
rect 159114 76046 159170 76102
rect 159238 76046 159294 76102
rect 159362 76046 159418 76102
rect 159486 76046 159542 76102
rect 159114 75922 159170 75978
rect 159238 75922 159294 75978
rect 159362 75922 159418 75978
rect 159486 75922 159542 75978
rect 159114 58294 159170 58350
rect 159238 58294 159294 58350
rect 159362 58294 159418 58350
rect 159486 58294 159542 58350
rect 159114 58170 159170 58226
rect 159238 58170 159294 58226
rect 159362 58170 159418 58226
rect 159486 58170 159542 58226
rect 159114 58046 159170 58102
rect 159238 58046 159294 58102
rect 159362 58046 159418 58102
rect 159486 58046 159542 58102
rect 159114 57922 159170 57978
rect 159238 57922 159294 57978
rect 159362 57922 159418 57978
rect 159486 57922 159542 57978
rect 159114 40294 159170 40350
rect 159238 40294 159294 40350
rect 159362 40294 159418 40350
rect 159486 40294 159542 40350
rect 159114 40170 159170 40226
rect 159238 40170 159294 40226
rect 159362 40170 159418 40226
rect 159486 40170 159542 40226
rect 159114 40046 159170 40102
rect 159238 40046 159294 40102
rect 159362 40046 159418 40102
rect 159486 40046 159542 40102
rect 159114 39922 159170 39978
rect 159238 39922 159294 39978
rect 159362 39922 159418 39978
rect 159486 39922 159542 39978
rect 132114 28294 132170 28350
rect 132238 28294 132294 28350
rect 132362 28294 132418 28350
rect 132486 28294 132542 28350
rect 132114 28170 132170 28226
rect 132238 28170 132294 28226
rect 132362 28170 132418 28226
rect 132486 28170 132542 28226
rect 132114 28046 132170 28102
rect 132238 28046 132294 28102
rect 132362 28046 132418 28102
rect 132486 28046 132542 28102
rect 132114 27922 132170 27978
rect 132238 27922 132294 27978
rect 132362 27922 132418 27978
rect 132486 27922 132542 27978
rect 150558 28294 150614 28350
rect 150682 28294 150738 28350
rect 150558 28170 150614 28226
rect 150682 28170 150738 28226
rect 150558 28046 150614 28102
rect 150682 28046 150738 28102
rect 150558 27922 150614 27978
rect 150682 27922 150738 27978
rect 159114 22294 159170 22350
rect 159238 22294 159294 22350
rect 159362 22294 159418 22350
rect 159486 22294 159542 22350
rect 159114 22170 159170 22226
rect 159238 22170 159294 22226
rect 159362 22170 159418 22226
rect 159486 22170 159542 22226
rect 159114 22046 159170 22102
rect 159238 22046 159294 22102
rect 159362 22046 159418 22102
rect 159486 22046 159542 22102
rect 159114 21922 159170 21978
rect 159238 21922 159294 21978
rect 159362 21922 159418 21978
rect 159486 21922 159542 21978
rect 132114 10294 132170 10350
rect 132238 10294 132294 10350
rect 132362 10294 132418 10350
rect 132486 10294 132542 10350
rect 132114 10170 132170 10226
rect 132238 10170 132294 10226
rect 132362 10170 132418 10226
rect 132486 10170 132542 10226
rect 132114 10046 132170 10102
rect 132238 10046 132294 10102
rect 132362 10046 132418 10102
rect 132486 10046 132542 10102
rect 132114 9922 132170 9978
rect 132238 9922 132294 9978
rect 132362 9922 132418 9978
rect 132486 9922 132542 9978
rect 150558 10294 150614 10350
rect 150682 10294 150738 10350
rect 150558 10170 150614 10226
rect 150682 10170 150738 10226
rect 150558 10046 150614 10102
rect 150682 10046 150738 10102
rect 150558 9922 150614 9978
rect 150682 9922 150738 9978
rect 132114 -1176 132170 -1120
rect 132238 -1176 132294 -1120
rect 132362 -1176 132418 -1120
rect 132486 -1176 132542 -1120
rect 132114 -1300 132170 -1244
rect 132238 -1300 132294 -1244
rect 132362 -1300 132418 -1244
rect 132486 -1300 132542 -1244
rect 132114 -1424 132170 -1368
rect 132238 -1424 132294 -1368
rect 132362 -1424 132418 -1368
rect 132486 -1424 132542 -1368
rect 132114 -1548 132170 -1492
rect 132238 -1548 132294 -1492
rect 132362 -1548 132418 -1492
rect 132486 -1548 132542 -1492
rect 159114 4294 159170 4350
rect 159238 4294 159294 4350
rect 159362 4294 159418 4350
rect 159486 4294 159542 4350
rect 159114 4170 159170 4226
rect 159238 4170 159294 4226
rect 159362 4170 159418 4226
rect 159486 4170 159542 4226
rect 159114 4046 159170 4102
rect 159238 4046 159294 4102
rect 159362 4046 159418 4102
rect 159486 4046 159542 4102
rect 159114 3922 159170 3978
rect 159238 3922 159294 3978
rect 159362 3922 159418 3978
rect 159486 3922 159542 3978
rect 159114 -216 159170 -160
rect 159238 -216 159294 -160
rect 159362 -216 159418 -160
rect 159486 -216 159542 -160
rect 159114 -340 159170 -284
rect 159238 -340 159294 -284
rect 159362 -340 159418 -284
rect 159486 -340 159542 -284
rect 159114 -464 159170 -408
rect 159238 -464 159294 -408
rect 159362 -464 159418 -408
rect 159486 -464 159542 -408
rect 159114 -588 159170 -532
rect 159238 -588 159294 -532
rect 159362 -588 159418 -532
rect 159486 -588 159542 -532
rect 165900 277116 165956 277138
rect 165900 277082 165956 277116
rect 168140 266462 168196 266518
rect 169260 268262 169316 268318
rect 169708 264662 169764 264718
rect 168028 255302 168084 255358
rect 168028 214082 168084 214138
rect 174636 278342 174692 278398
rect 175308 277262 175364 277318
rect 173852 276362 173908 276418
rect 175980 273482 176036 273538
rect 173852 261602 173908 261658
rect 177324 271502 177380 271558
rect 176540 269882 176596 269938
rect 178108 267902 178164 267958
rect 176428 218222 176484 218278
rect 173852 212462 173908 212518
rect 177212 209942 177268 209998
rect 180012 268082 180068 268138
rect 179900 266282 179956 266338
rect 179788 264842 179844 264898
rect 178892 209942 178948 209998
rect 184716 271862 184772 271918
rect 184828 270422 184884 270478
rect 183148 270242 183204 270298
rect 181468 264482 181524 264538
rect 183932 262862 183988 262918
rect 186172 260342 186228 260398
rect 183932 222542 183988 222598
rect 184716 222542 184772 222598
rect 183036 219122 183092 219178
rect 186284 201482 186340 201538
rect 187404 278162 187460 278218
rect 189532 276722 189588 276778
rect 186732 273662 186788 273718
rect 188076 272042 188132 272098
rect 188748 271682 188804 271738
rect 186396 191402 186452 191458
rect 187292 260342 187348 260398
rect 187404 225062 187460 225118
rect 187292 172682 187348 172738
rect 189532 276542 189588 276598
rect 189420 268442 189476 268498
rect 189084 168722 189140 168778
rect 189834 274294 189890 274350
rect 189958 274294 190014 274350
rect 190082 274294 190138 274350
rect 190206 274294 190262 274350
rect 189834 274170 189890 274226
rect 189958 274170 190014 274226
rect 190082 274170 190138 274226
rect 190206 274170 190262 274226
rect 189834 274046 189890 274102
rect 189958 274046 190014 274102
rect 190082 274046 190138 274102
rect 190206 274046 190262 274102
rect 189834 273922 189890 273978
rect 189958 273922 190014 273978
rect 190082 273922 190138 273978
rect 190206 273922 190262 273978
rect 190428 266822 190484 266878
rect 189834 256294 189890 256350
rect 189958 256294 190014 256350
rect 190082 256294 190138 256350
rect 190206 256294 190262 256350
rect 189834 256170 189890 256226
rect 189958 256170 190014 256226
rect 190082 256170 190138 256226
rect 190206 256170 190262 256226
rect 189834 256046 189890 256102
rect 189958 256046 190014 256102
rect 190082 256046 190138 256102
rect 190206 256046 190262 256102
rect 189834 255922 189890 255978
rect 189958 255922 190014 255978
rect 190082 255922 190138 255978
rect 190206 255922 190262 255978
rect 189834 238294 189890 238350
rect 189958 238294 190014 238350
rect 190082 238294 190138 238350
rect 190206 238294 190262 238350
rect 189834 238170 189890 238226
rect 189958 238170 190014 238226
rect 190082 238170 190138 238226
rect 190206 238170 190262 238226
rect 189834 238046 189890 238102
rect 189958 238046 190014 238102
rect 190082 238046 190138 238102
rect 190206 238046 190262 238102
rect 189834 237922 189890 237978
rect 189958 237922 190014 237978
rect 190082 237922 190138 237978
rect 190206 237922 190262 237978
rect 189834 220294 189890 220350
rect 189958 220294 190014 220350
rect 190082 220294 190138 220350
rect 190206 220294 190262 220350
rect 189834 220170 189890 220226
rect 189958 220170 190014 220226
rect 190082 220170 190138 220226
rect 190206 220170 190262 220226
rect 189834 220046 189890 220102
rect 189958 220046 190014 220102
rect 190082 220046 190138 220102
rect 190206 220046 190262 220102
rect 189834 219922 189890 219978
rect 189958 219922 190014 219978
rect 190082 219922 190138 219978
rect 190206 219922 190262 219978
rect 189834 202294 189890 202350
rect 189958 202294 190014 202350
rect 190082 202294 190138 202350
rect 190206 202294 190262 202350
rect 189834 202170 189890 202226
rect 189958 202170 190014 202226
rect 190082 202170 190138 202226
rect 190206 202170 190262 202226
rect 189834 202046 189890 202102
rect 189958 202046 190014 202102
rect 190082 202046 190138 202102
rect 190206 202046 190262 202102
rect 189834 201922 189890 201978
rect 189958 201922 190014 201978
rect 190082 201922 190138 201978
rect 190206 201922 190262 201978
rect 189834 184294 189890 184350
rect 189958 184294 190014 184350
rect 190082 184294 190138 184350
rect 190206 184294 190262 184350
rect 189834 184170 189890 184226
rect 189958 184170 190014 184226
rect 190082 184170 190138 184226
rect 190206 184170 190262 184226
rect 189834 184046 189890 184102
rect 189958 184046 190014 184102
rect 190082 184046 190138 184102
rect 190206 184046 190262 184102
rect 189834 183922 189890 183978
rect 189958 183922 190014 183978
rect 190082 183922 190138 183978
rect 190206 183922 190262 183978
rect 189834 166294 189890 166350
rect 189958 166294 190014 166350
rect 190082 166294 190138 166350
rect 190206 166294 190262 166350
rect 189834 166170 189890 166226
rect 189958 166170 190014 166226
rect 190082 166170 190138 166226
rect 190206 166170 190262 166226
rect 189834 166046 189890 166102
rect 189958 166046 190014 166102
rect 190082 166046 190138 166102
rect 190206 166046 190262 166102
rect 189834 165922 189890 165978
rect 189958 165922 190014 165978
rect 190082 165922 190138 165978
rect 190206 165922 190262 165978
rect 162834 154294 162890 154350
rect 162958 154294 163014 154350
rect 163082 154294 163138 154350
rect 163206 154294 163262 154350
rect 162834 154170 162890 154226
rect 162958 154170 163014 154226
rect 163082 154170 163138 154226
rect 163206 154170 163262 154226
rect 162834 154046 162890 154102
rect 162958 154046 163014 154102
rect 163082 154046 163138 154102
rect 163206 154046 163262 154102
rect 162834 153922 162890 153978
rect 162958 153922 163014 153978
rect 163082 153922 163138 153978
rect 163206 153922 163262 153978
rect 162834 136294 162890 136350
rect 162958 136294 163014 136350
rect 163082 136294 163138 136350
rect 163206 136294 163262 136350
rect 162834 136170 162890 136226
rect 162958 136170 163014 136226
rect 163082 136170 163138 136226
rect 163206 136170 163262 136226
rect 162834 136046 162890 136102
rect 162958 136046 163014 136102
rect 163082 136046 163138 136102
rect 163206 136046 163262 136102
rect 162834 135922 162890 135978
rect 162958 135922 163014 135978
rect 163082 135922 163138 135978
rect 163206 135922 163262 135978
rect 162834 118294 162890 118350
rect 162958 118294 163014 118350
rect 163082 118294 163138 118350
rect 163206 118294 163262 118350
rect 162834 118170 162890 118226
rect 162958 118170 163014 118226
rect 163082 118170 163138 118226
rect 163206 118170 163262 118226
rect 162834 118046 162890 118102
rect 162958 118046 163014 118102
rect 163082 118046 163138 118102
rect 163206 118046 163262 118102
rect 162834 117922 162890 117978
rect 162958 117922 163014 117978
rect 163082 117922 163138 117978
rect 163206 117922 163262 117978
rect 162834 100294 162890 100350
rect 162958 100294 163014 100350
rect 163082 100294 163138 100350
rect 163206 100294 163262 100350
rect 162834 100170 162890 100226
rect 162958 100170 163014 100226
rect 163082 100170 163138 100226
rect 163206 100170 163262 100226
rect 162834 100046 162890 100102
rect 162958 100046 163014 100102
rect 163082 100046 163138 100102
rect 163206 100046 163262 100102
rect 162834 99922 162890 99978
rect 162958 99922 163014 99978
rect 163082 99922 163138 99978
rect 163206 99922 163262 99978
rect 162834 82294 162890 82350
rect 162958 82294 163014 82350
rect 163082 82294 163138 82350
rect 163206 82294 163262 82350
rect 162834 82170 162890 82226
rect 162958 82170 163014 82226
rect 163082 82170 163138 82226
rect 163206 82170 163262 82226
rect 162834 82046 162890 82102
rect 162958 82046 163014 82102
rect 163082 82046 163138 82102
rect 163206 82046 163262 82102
rect 162834 81922 162890 81978
rect 162958 81922 163014 81978
rect 163082 81922 163138 81978
rect 163206 81922 163262 81978
rect 162834 64294 162890 64350
rect 162958 64294 163014 64350
rect 163082 64294 163138 64350
rect 163206 64294 163262 64350
rect 162834 64170 162890 64226
rect 162958 64170 163014 64226
rect 163082 64170 163138 64226
rect 163206 64170 163262 64226
rect 162834 64046 162890 64102
rect 162958 64046 163014 64102
rect 163082 64046 163138 64102
rect 163206 64046 163262 64102
rect 162834 63922 162890 63978
rect 162958 63922 163014 63978
rect 163082 63922 163138 63978
rect 163206 63922 163262 63978
rect 162834 46294 162890 46350
rect 162958 46294 163014 46350
rect 163082 46294 163138 46350
rect 163206 46294 163262 46350
rect 162834 46170 162890 46226
rect 162958 46170 163014 46226
rect 163082 46170 163138 46226
rect 163206 46170 163262 46226
rect 162834 46046 162890 46102
rect 162958 46046 163014 46102
rect 163082 46046 163138 46102
rect 163206 46046 163262 46102
rect 162834 45922 162890 45978
rect 162958 45922 163014 45978
rect 163082 45922 163138 45978
rect 163206 45922 163262 45978
rect 162834 28294 162890 28350
rect 162958 28294 163014 28350
rect 163082 28294 163138 28350
rect 163206 28294 163262 28350
rect 162834 28170 162890 28226
rect 162958 28170 163014 28226
rect 163082 28170 163138 28226
rect 163206 28170 163262 28226
rect 162834 28046 162890 28102
rect 162958 28046 163014 28102
rect 163082 28046 163138 28102
rect 163206 28046 163262 28102
rect 162834 27922 162890 27978
rect 162958 27922 163014 27978
rect 163082 27922 163138 27978
rect 163206 27922 163262 27978
rect 162834 10294 162890 10350
rect 162958 10294 163014 10350
rect 163082 10294 163138 10350
rect 163206 10294 163262 10350
rect 162834 10170 162890 10226
rect 162958 10170 163014 10226
rect 163082 10170 163138 10226
rect 163206 10170 163262 10226
rect 162834 10046 162890 10102
rect 162958 10046 163014 10102
rect 163082 10046 163138 10102
rect 163206 10046 163262 10102
rect 162834 9922 162890 9978
rect 162958 9922 163014 9978
rect 163082 9922 163138 9978
rect 163206 9922 163262 9978
rect 162834 -1176 162890 -1120
rect 162958 -1176 163014 -1120
rect 163082 -1176 163138 -1120
rect 163206 -1176 163262 -1120
rect 162834 -1300 162890 -1244
rect 162958 -1300 163014 -1244
rect 163082 -1300 163138 -1244
rect 163206 -1300 163262 -1244
rect 162834 -1424 162890 -1368
rect 162958 -1424 163014 -1368
rect 163082 -1424 163138 -1368
rect 163206 -1424 163262 -1368
rect 162834 -1548 162890 -1492
rect 162958 -1548 163014 -1492
rect 163082 -1548 163138 -1492
rect 163206 -1548 163262 -1492
rect 192332 225062 192388 225118
rect 192332 223442 192388 223498
rect 193004 357362 193060 357418
rect 193116 282122 193172 282178
rect 193554 280294 193610 280350
rect 193678 280294 193734 280350
rect 193802 280294 193858 280350
rect 193926 280294 193982 280350
rect 193554 280170 193610 280226
rect 193678 280170 193734 280226
rect 193802 280170 193858 280226
rect 193926 280170 193982 280226
rect 193554 280046 193610 280102
rect 193678 280046 193734 280102
rect 193802 280046 193858 280102
rect 193926 280046 193982 280102
rect 193554 279922 193610 279978
rect 193678 279922 193734 279978
rect 193802 279922 193858 279978
rect 193926 279922 193982 279978
rect 193554 262294 193610 262350
rect 193678 262294 193734 262350
rect 193802 262294 193858 262350
rect 193926 262294 193982 262350
rect 193554 262170 193610 262226
rect 193678 262170 193734 262226
rect 193802 262170 193858 262226
rect 193926 262170 193982 262226
rect 193554 262046 193610 262102
rect 193678 262046 193734 262102
rect 193802 262046 193858 262102
rect 193926 262046 193982 262102
rect 193554 261922 193610 261978
rect 193678 261922 193734 261978
rect 193802 261922 193858 261978
rect 193926 261922 193982 261978
rect 193554 244294 193610 244350
rect 193678 244294 193734 244350
rect 193802 244294 193858 244350
rect 193926 244294 193982 244350
rect 193554 244170 193610 244226
rect 193678 244170 193734 244226
rect 193802 244170 193858 244226
rect 193926 244170 193982 244226
rect 193554 244046 193610 244102
rect 193678 244046 193734 244102
rect 193802 244046 193858 244102
rect 193926 244046 193982 244102
rect 193554 243922 193610 243978
rect 193678 243922 193734 243978
rect 193802 243922 193858 243978
rect 193926 243922 193982 243978
rect 193554 226294 193610 226350
rect 193678 226294 193734 226350
rect 193802 226294 193858 226350
rect 193926 226294 193982 226350
rect 193554 226170 193610 226226
rect 193678 226170 193734 226226
rect 193802 226170 193858 226226
rect 193926 226170 193982 226226
rect 193554 226046 193610 226102
rect 193678 226046 193734 226102
rect 193802 226046 193858 226102
rect 193926 226046 193982 226102
rect 193554 225922 193610 225978
rect 193678 225922 193734 225978
rect 193802 225922 193858 225978
rect 193926 225922 193982 225978
rect 193554 208294 193610 208350
rect 193678 208294 193734 208350
rect 193802 208294 193858 208350
rect 193926 208294 193982 208350
rect 193554 208170 193610 208226
rect 193678 208170 193734 208226
rect 193802 208170 193858 208226
rect 193926 208170 193982 208226
rect 193554 208046 193610 208102
rect 193678 208046 193734 208102
rect 193802 208046 193858 208102
rect 193926 208046 193982 208102
rect 193554 207922 193610 207978
rect 193678 207922 193734 207978
rect 193802 207922 193858 207978
rect 193926 207922 193982 207978
rect 193554 190294 193610 190350
rect 193678 190294 193734 190350
rect 193802 190294 193858 190350
rect 193926 190294 193982 190350
rect 193554 190170 193610 190226
rect 193678 190170 193734 190226
rect 193802 190170 193858 190226
rect 193926 190170 193982 190226
rect 193554 190046 193610 190102
rect 193678 190046 193734 190102
rect 193802 190046 193858 190102
rect 193926 190046 193982 190102
rect 193554 189922 193610 189978
rect 193678 189922 193734 189978
rect 193802 189922 193858 189978
rect 193926 189922 193982 189978
rect 193554 172294 193610 172350
rect 193678 172294 193734 172350
rect 193802 172294 193858 172350
rect 193926 172294 193982 172350
rect 193554 172170 193610 172226
rect 193678 172170 193734 172226
rect 193802 172170 193858 172226
rect 193926 172170 193982 172226
rect 193554 172046 193610 172102
rect 193678 172046 193734 172102
rect 193802 172046 193858 172102
rect 193926 172046 193982 172102
rect 193554 171922 193610 171978
rect 193678 171922 193734 171978
rect 193802 171922 193858 171978
rect 193926 171922 193982 171978
rect 193554 154294 193610 154350
rect 193678 154294 193734 154350
rect 193802 154294 193858 154350
rect 193926 154294 193982 154350
rect 193554 154170 193610 154226
rect 193678 154170 193734 154226
rect 193802 154170 193858 154226
rect 193926 154170 193982 154226
rect 193554 154046 193610 154102
rect 193678 154046 193734 154102
rect 193802 154046 193858 154102
rect 193926 154046 193982 154102
rect 193554 153922 193610 153978
rect 193678 153922 193734 153978
rect 193802 153922 193858 153978
rect 193926 153922 193982 153978
rect 189834 148294 189890 148350
rect 189958 148294 190014 148350
rect 190082 148294 190138 148350
rect 190206 148294 190262 148350
rect 189834 148170 189890 148226
rect 189958 148170 190014 148226
rect 190082 148170 190138 148226
rect 190206 148170 190262 148226
rect 189834 148046 189890 148102
rect 189958 148046 190014 148102
rect 190082 148046 190138 148102
rect 190206 148046 190262 148102
rect 189834 147922 189890 147978
rect 189958 147922 190014 147978
rect 190082 147922 190138 147978
rect 190206 147922 190262 147978
rect 189834 130294 189890 130350
rect 189958 130294 190014 130350
rect 190082 130294 190138 130350
rect 190206 130294 190262 130350
rect 189834 130170 189890 130226
rect 189958 130170 190014 130226
rect 190082 130170 190138 130226
rect 190206 130170 190262 130226
rect 189834 130046 189890 130102
rect 189958 130046 190014 130102
rect 190082 130046 190138 130102
rect 190206 130046 190262 130102
rect 189834 129922 189890 129978
rect 189958 129922 190014 129978
rect 190082 129922 190138 129978
rect 190206 129922 190262 129978
rect 189834 112294 189890 112350
rect 189958 112294 190014 112350
rect 190082 112294 190138 112350
rect 190206 112294 190262 112350
rect 189834 112170 189890 112226
rect 189958 112170 190014 112226
rect 190082 112170 190138 112226
rect 190206 112170 190262 112226
rect 189834 112046 189890 112102
rect 189958 112046 190014 112102
rect 190082 112046 190138 112102
rect 190206 112046 190262 112102
rect 189834 111922 189890 111978
rect 189958 111922 190014 111978
rect 190082 111922 190138 111978
rect 190206 111922 190262 111978
rect 189834 94294 189890 94350
rect 189958 94294 190014 94350
rect 190082 94294 190138 94350
rect 190206 94294 190262 94350
rect 189834 94170 189890 94226
rect 189958 94170 190014 94226
rect 190082 94170 190138 94226
rect 190206 94170 190262 94226
rect 189834 94046 189890 94102
rect 189958 94046 190014 94102
rect 190082 94046 190138 94102
rect 190206 94046 190262 94102
rect 189834 93922 189890 93978
rect 189958 93922 190014 93978
rect 190082 93922 190138 93978
rect 190206 93922 190262 93978
rect 189834 76294 189890 76350
rect 189958 76294 190014 76350
rect 190082 76294 190138 76350
rect 190206 76294 190262 76350
rect 189834 76170 189890 76226
rect 189958 76170 190014 76226
rect 190082 76170 190138 76226
rect 190206 76170 190262 76226
rect 189834 76046 189890 76102
rect 189958 76046 190014 76102
rect 190082 76046 190138 76102
rect 190206 76046 190262 76102
rect 189834 75922 189890 75978
rect 189958 75922 190014 75978
rect 190082 75922 190138 75978
rect 190206 75922 190262 75978
rect 189834 58294 189890 58350
rect 189958 58294 190014 58350
rect 190082 58294 190138 58350
rect 190206 58294 190262 58350
rect 189834 58170 189890 58226
rect 189958 58170 190014 58226
rect 190082 58170 190138 58226
rect 190206 58170 190262 58226
rect 189834 58046 189890 58102
rect 189958 58046 190014 58102
rect 190082 58046 190138 58102
rect 190206 58046 190262 58102
rect 189834 57922 189890 57978
rect 189958 57922 190014 57978
rect 190082 57922 190138 57978
rect 190206 57922 190262 57978
rect 189834 40294 189890 40350
rect 189958 40294 190014 40350
rect 190082 40294 190138 40350
rect 190206 40294 190262 40350
rect 189834 40170 189890 40226
rect 189958 40170 190014 40226
rect 190082 40170 190138 40226
rect 190206 40170 190262 40226
rect 189834 40046 189890 40102
rect 189958 40046 190014 40102
rect 190082 40046 190138 40102
rect 190206 40046 190262 40102
rect 189834 39922 189890 39978
rect 189958 39922 190014 39978
rect 190082 39922 190138 39978
rect 190206 39922 190262 39978
rect 189834 22294 189890 22350
rect 189958 22294 190014 22350
rect 190082 22294 190138 22350
rect 190206 22294 190262 22350
rect 189834 22170 189890 22226
rect 189958 22170 190014 22226
rect 190082 22170 190138 22226
rect 190206 22170 190262 22226
rect 189834 22046 189890 22102
rect 189958 22046 190014 22102
rect 190082 22046 190138 22102
rect 190206 22046 190262 22102
rect 189834 21922 189890 21978
rect 189958 21922 190014 21978
rect 190082 21922 190138 21978
rect 190206 21922 190262 21978
rect 189834 4294 189890 4350
rect 189958 4294 190014 4350
rect 190082 4294 190138 4350
rect 190206 4294 190262 4350
rect 189834 4170 189890 4226
rect 189958 4170 190014 4226
rect 190082 4170 190138 4226
rect 190206 4170 190262 4226
rect 189834 4046 189890 4102
rect 189958 4046 190014 4102
rect 190082 4046 190138 4102
rect 190206 4046 190262 4102
rect 189834 3922 189890 3978
rect 189958 3922 190014 3978
rect 190082 3922 190138 3978
rect 190206 3922 190262 3978
rect 189834 -216 189890 -160
rect 189958 -216 190014 -160
rect 190082 -216 190138 -160
rect 190206 -216 190262 -160
rect 189834 -340 189890 -284
rect 189958 -340 190014 -284
rect 190082 -340 190138 -284
rect 190206 -340 190262 -284
rect 189834 -464 189890 -408
rect 189958 -464 190014 -408
rect 190082 -464 190138 -408
rect 190206 -464 190262 -408
rect 189834 -588 189890 -532
rect 189958 -588 190014 -532
rect 190082 -588 190138 -532
rect 190206 -588 190262 -532
rect 194348 296702 194404 296758
rect 194796 360242 194852 360298
rect 194684 282122 194740 282178
rect 194572 270116 194628 270118
rect 194572 270062 194628 270116
rect 195916 359702 195972 359758
rect 195302 346294 195358 346350
rect 195426 346294 195482 346350
rect 195302 346170 195358 346226
rect 195426 346170 195482 346226
rect 195302 346046 195358 346102
rect 195426 346046 195482 346102
rect 195302 345922 195358 345978
rect 195426 345922 195482 345978
rect 195302 328294 195358 328350
rect 195426 328294 195482 328350
rect 195302 328170 195358 328226
rect 195426 328170 195482 328226
rect 195302 328046 195358 328102
rect 195426 328046 195482 328102
rect 195302 327922 195358 327978
rect 195426 327922 195482 327978
rect 195302 310294 195358 310350
rect 195426 310294 195482 310350
rect 195302 310170 195358 310226
rect 195426 310170 195482 310226
rect 195302 310046 195358 310102
rect 195426 310046 195482 310102
rect 195302 309922 195358 309978
rect 195426 309922 195482 309978
rect 195302 292294 195358 292350
rect 195426 292294 195482 292350
rect 195302 292170 195358 292226
rect 195426 292170 195482 292226
rect 195302 292046 195358 292102
rect 195426 292046 195482 292102
rect 195302 291922 195358 291978
rect 195426 291922 195482 291978
rect 195804 296342 195860 296398
rect 196476 359522 196532 359578
rect 196476 357542 196532 357598
rect 197372 336302 197428 336358
rect 197036 273302 197092 273358
rect 197484 330182 197540 330238
rect 197596 317762 197652 317818
rect 199276 359522 199332 359578
rect 199388 357902 199444 357958
rect 199276 357182 199332 357238
rect 199276 336302 199332 336358
rect 199276 330204 199332 330238
rect 199276 330182 199332 330204
rect 199276 317772 199332 317818
rect 199276 317762 199332 317772
rect 198156 305702 198212 305758
rect 197820 287522 197876 287578
rect 199276 296716 199332 296758
rect 199276 296702 199332 296716
rect 199276 287532 199332 287578
rect 199276 287522 199332 287532
rect 197820 265022 197876 265078
rect 198442 256294 198498 256350
rect 198566 256294 198622 256350
rect 198690 256294 198746 256350
rect 198814 256294 198870 256350
rect 198442 256170 198498 256226
rect 198566 256170 198622 256226
rect 198690 256170 198746 256226
rect 198814 256170 198870 256226
rect 198442 256046 198498 256102
rect 198566 256046 198622 256102
rect 198690 256046 198746 256102
rect 198814 256046 198870 256102
rect 198442 255922 198498 255978
rect 198566 255922 198622 255978
rect 198690 255922 198746 255978
rect 198814 255922 198870 255978
rect 197642 244294 197698 244350
rect 197766 244294 197822 244350
rect 197890 244294 197946 244350
rect 198014 244294 198070 244350
rect 197642 244170 197698 244226
rect 197766 244170 197822 244226
rect 197890 244170 197946 244226
rect 198014 244170 198070 244226
rect 197642 244046 197698 244102
rect 197766 244046 197822 244102
rect 197890 244046 197946 244102
rect 198014 244046 198070 244102
rect 197642 243922 197698 243978
rect 197766 243922 197822 243978
rect 197890 243922 197946 243978
rect 198014 243922 198070 243978
rect 198442 238294 198498 238350
rect 198566 238294 198622 238350
rect 198690 238294 198746 238350
rect 198814 238294 198870 238350
rect 198442 238170 198498 238226
rect 198566 238170 198622 238226
rect 198690 238170 198746 238226
rect 198814 238170 198870 238226
rect 198442 238046 198498 238102
rect 198566 238046 198622 238102
rect 198690 238046 198746 238102
rect 198814 238046 198870 238102
rect 198442 237922 198498 237978
rect 198566 237922 198622 237978
rect 198690 237922 198746 237978
rect 198814 237922 198870 237978
rect 197642 226294 197698 226350
rect 197766 226294 197822 226350
rect 197890 226294 197946 226350
rect 198014 226294 198070 226350
rect 197642 226170 197698 226226
rect 197766 226170 197822 226226
rect 197890 226170 197946 226226
rect 198014 226170 198070 226226
rect 197642 226046 197698 226102
rect 197766 226046 197822 226102
rect 197890 226046 197946 226102
rect 198014 226046 198070 226102
rect 197642 225922 197698 225978
rect 197766 225922 197822 225978
rect 197890 225922 197946 225978
rect 198014 225922 198070 225978
rect 198442 220294 198498 220350
rect 198566 220294 198622 220350
rect 198690 220294 198746 220350
rect 198814 220294 198870 220350
rect 198442 220170 198498 220226
rect 198566 220170 198622 220226
rect 198690 220170 198746 220226
rect 198814 220170 198870 220226
rect 198442 220046 198498 220102
rect 198566 220046 198622 220102
rect 198690 220046 198746 220102
rect 198814 220046 198870 220102
rect 198442 219922 198498 219978
rect 198566 219922 198622 219978
rect 198690 219922 198746 219978
rect 198814 219922 198870 219978
rect 197642 208294 197698 208350
rect 197766 208294 197822 208350
rect 197890 208294 197946 208350
rect 198014 208294 198070 208350
rect 197642 208170 197698 208226
rect 197766 208170 197822 208226
rect 197890 208170 197946 208226
rect 198014 208170 198070 208226
rect 197642 208046 197698 208102
rect 197766 208046 197822 208102
rect 197890 208046 197946 208102
rect 198014 208046 198070 208102
rect 197642 207922 197698 207978
rect 197766 207922 197822 207978
rect 197890 207922 197946 207978
rect 198014 207922 198070 207978
rect 198442 202294 198498 202350
rect 198566 202294 198622 202350
rect 198690 202294 198746 202350
rect 198814 202294 198870 202350
rect 198442 202170 198498 202226
rect 198566 202170 198622 202226
rect 198690 202170 198746 202226
rect 198814 202170 198870 202226
rect 198442 202046 198498 202102
rect 198566 202046 198622 202102
rect 198690 202046 198746 202102
rect 198814 202046 198870 202102
rect 198442 201922 198498 201978
rect 198566 201922 198622 201978
rect 198690 201922 198746 201978
rect 198814 201922 198870 201978
rect 197642 190294 197698 190350
rect 197766 190294 197822 190350
rect 197890 190294 197946 190350
rect 198014 190294 198070 190350
rect 197642 190170 197698 190226
rect 197766 190170 197822 190226
rect 197890 190170 197946 190226
rect 198014 190170 198070 190226
rect 197642 190046 197698 190102
rect 197766 190046 197822 190102
rect 197890 190046 197946 190102
rect 198014 190046 198070 190102
rect 197642 189922 197698 189978
rect 197766 189922 197822 189978
rect 197890 189922 197946 189978
rect 198014 189922 198070 189978
rect 198442 184294 198498 184350
rect 198566 184294 198622 184350
rect 198690 184294 198746 184350
rect 198814 184294 198870 184350
rect 198442 184170 198498 184226
rect 198566 184170 198622 184226
rect 198690 184170 198746 184226
rect 198814 184170 198870 184226
rect 198442 184046 198498 184102
rect 198566 184046 198622 184102
rect 198690 184046 198746 184102
rect 198814 184046 198870 184102
rect 198442 183922 198498 183978
rect 198566 183922 198622 183978
rect 198690 183922 198746 183978
rect 198814 183922 198870 183978
rect 197642 172294 197698 172350
rect 197766 172294 197822 172350
rect 197890 172294 197946 172350
rect 198014 172294 198070 172350
rect 197642 172170 197698 172226
rect 197766 172170 197822 172226
rect 197890 172170 197946 172226
rect 198014 172170 198070 172226
rect 197642 172046 197698 172102
rect 197766 172046 197822 172102
rect 197890 172046 197946 172102
rect 198014 172046 198070 172102
rect 197642 171922 197698 171978
rect 197766 171922 197822 171978
rect 197890 171922 197946 171978
rect 198014 171922 198070 171978
rect 220554 580294 220610 580350
rect 220678 580294 220734 580350
rect 220802 580294 220858 580350
rect 220926 580294 220982 580350
rect 220554 580170 220610 580226
rect 220678 580170 220734 580226
rect 220802 580170 220858 580226
rect 220926 580170 220982 580226
rect 220554 580046 220610 580102
rect 220678 580046 220734 580102
rect 220802 580046 220858 580102
rect 220926 580046 220982 580102
rect 220554 579922 220610 579978
rect 220678 579922 220734 579978
rect 220802 579922 220858 579978
rect 220926 579922 220982 579978
rect 220554 562294 220610 562350
rect 220678 562294 220734 562350
rect 220802 562294 220858 562350
rect 220926 562294 220982 562350
rect 220554 562170 220610 562226
rect 220678 562170 220734 562226
rect 220802 562170 220858 562226
rect 220926 562170 220982 562226
rect 220554 562046 220610 562102
rect 220678 562046 220734 562102
rect 220802 562046 220858 562102
rect 220926 562046 220982 562102
rect 220554 561922 220610 561978
rect 220678 561922 220734 561978
rect 220802 561922 220858 561978
rect 220926 561922 220982 561978
rect 220554 544294 220610 544350
rect 220678 544294 220734 544350
rect 220802 544294 220858 544350
rect 220926 544294 220982 544350
rect 220554 544170 220610 544226
rect 220678 544170 220734 544226
rect 220802 544170 220858 544226
rect 220926 544170 220982 544226
rect 220554 544046 220610 544102
rect 220678 544046 220734 544102
rect 220802 544046 220858 544102
rect 220926 544046 220982 544102
rect 220554 543922 220610 543978
rect 220678 543922 220734 543978
rect 220802 543922 220858 543978
rect 220926 543922 220982 543978
rect 220554 526294 220610 526350
rect 220678 526294 220734 526350
rect 220802 526294 220858 526350
rect 220926 526294 220982 526350
rect 220554 526170 220610 526226
rect 220678 526170 220734 526226
rect 220802 526170 220858 526226
rect 220926 526170 220982 526226
rect 220554 526046 220610 526102
rect 220678 526046 220734 526102
rect 220802 526046 220858 526102
rect 220926 526046 220982 526102
rect 220554 525922 220610 525978
rect 220678 525922 220734 525978
rect 220802 525922 220858 525978
rect 220926 525922 220982 525978
rect 220554 508294 220610 508350
rect 220678 508294 220734 508350
rect 220802 508294 220858 508350
rect 220926 508294 220982 508350
rect 220554 508170 220610 508226
rect 220678 508170 220734 508226
rect 220802 508170 220858 508226
rect 220926 508170 220982 508226
rect 220554 508046 220610 508102
rect 220678 508046 220734 508102
rect 220802 508046 220858 508102
rect 220926 508046 220982 508102
rect 220554 507922 220610 507978
rect 220678 507922 220734 507978
rect 220802 507922 220858 507978
rect 220926 507922 220982 507978
rect 220554 490294 220610 490350
rect 220678 490294 220734 490350
rect 220802 490294 220858 490350
rect 220926 490294 220982 490350
rect 220554 490170 220610 490226
rect 220678 490170 220734 490226
rect 220802 490170 220858 490226
rect 220926 490170 220982 490226
rect 220554 490046 220610 490102
rect 220678 490046 220734 490102
rect 220802 490046 220858 490102
rect 220926 490046 220982 490102
rect 220554 489922 220610 489978
rect 220678 489922 220734 489978
rect 220802 489922 220858 489978
rect 220926 489922 220982 489978
rect 220554 472294 220610 472350
rect 220678 472294 220734 472350
rect 220802 472294 220858 472350
rect 220926 472294 220982 472350
rect 220554 472170 220610 472226
rect 220678 472170 220734 472226
rect 220802 472170 220858 472226
rect 220926 472170 220982 472226
rect 220554 472046 220610 472102
rect 220678 472046 220734 472102
rect 220802 472046 220858 472102
rect 220926 472046 220982 472102
rect 220554 471922 220610 471978
rect 220678 471922 220734 471978
rect 220802 471922 220858 471978
rect 220926 471922 220982 471978
rect 220554 454294 220610 454350
rect 220678 454294 220734 454350
rect 220802 454294 220858 454350
rect 220926 454294 220982 454350
rect 220554 454170 220610 454226
rect 220678 454170 220734 454226
rect 220802 454170 220858 454226
rect 220926 454170 220982 454226
rect 220554 454046 220610 454102
rect 220678 454046 220734 454102
rect 220802 454046 220858 454102
rect 220926 454046 220982 454102
rect 220554 453922 220610 453978
rect 220678 453922 220734 453978
rect 220802 453922 220858 453978
rect 220926 453922 220982 453978
rect 220554 436294 220610 436350
rect 220678 436294 220734 436350
rect 220802 436294 220858 436350
rect 220926 436294 220982 436350
rect 220554 436170 220610 436226
rect 220678 436170 220734 436226
rect 220802 436170 220858 436226
rect 220926 436170 220982 436226
rect 220554 436046 220610 436102
rect 220678 436046 220734 436102
rect 220802 436046 220858 436102
rect 220926 436046 220982 436102
rect 220554 435922 220610 435978
rect 220678 435922 220734 435978
rect 220802 435922 220858 435978
rect 220926 435922 220982 435978
rect 220554 418294 220610 418350
rect 220678 418294 220734 418350
rect 220802 418294 220858 418350
rect 220926 418294 220982 418350
rect 220554 418170 220610 418226
rect 220678 418170 220734 418226
rect 220802 418170 220858 418226
rect 220926 418170 220982 418226
rect 220554 418046 220610 418102
rect 220678 418046 220734 418102
rect 220802 418046 220858 418102
rect 220926 418046 220982 418102
rect 220554 417922 220610 417978
rect 220678 417922 220734 417978
rect 220802 417922 220858 417978
rect 220926 417922 220982 417978
rect 220554 400294 220610 400350
rect 220678 400294 220734 400350
rect 220802 400294 220858 400350
rect 220926 400294 220982 400350
rect 220554 400170 220610 400226
rect 220678 400170 220734 400226
rect 220802 400170 220858 400226
rect 220926 400170 220982 400226
rect 220554 400046 220610 400102
rect 220678 400046 220734 400102
rect 220802 400046 220858 400102
rect 220926 400046 220982 400102
rect 220554 399922 220610 399978
rect 220678 399922 220734 399978
rect 220802 399922 220858 399978
rect 220926 399922 220982 399978
rect 202412 366722 202468 366778
rect 202076 366542 202132 366598
rect 201852 366362 201908 366418
rect 201964 361322 202020 361378
rect 199836 305702 199892 305758
rect 202188 359522 202244 359578
rect 201852 296342 201908 296398
rect 201740 279602 201796 279658
rect 201516 168756 201572 168778
rect 201516 168722 201572 168756
rect 202076 279422 202132 279478
rect 202188 274562 202244 274618
rect 202412 205082 202468 205138
rect 220554 382294 220610 382350
rect 220678 382294 220734 382350
rect 220802 382294 220858 382350
rect 220926 382294 220982 382350
rect 220554 382170 220610 382226
rect 220678 382170 220734 382226
rect 220802 382170 220858 382226
rect 220926 382170 220982 382226
rect 220554 382046 220610 382102
rect 220678 382046 220734 382102
rect 220802 382046 220858 382102
rect 220926 382046 220982 382102
rect 220554 381922 220610 381978
rect 220678 381922 220734 381978
rect 220802 381922 220858 381978
rect 220926 381922 220982 381978
rect 204092 364742 204148 364798
rect 203420 187262 203476 187318
rect 203420 181502 203476 181558
rect 193554 136294 193610 136350
rect 193678 136294 193734 136350
rect 193802 136294 193858 136350
rect 193926 136294 193982 136350
rect 193554 136170 193610 136226
rect 193678 136170 193734 136226
rect 193802 136170 193858 136226
rect 193926 136170 193982 136226
rect 193554 136046 193610 136102
rect 193678 136046 193734 136102
rect 193802 136046 193858 136102
rect 193926 136046 193982 136102
rect 193554 135922 193610 135978
rect 193678 135922 193734 135978
rect 193802 135922 193858 135978
rect 193926 135922 193982 135978
rect 196612 136294 196668 136350
rect 196736 136294 196792 136350
rect 196860 136294 196916 136350
rect 196984 136294 197040 136350
rect 196612 136170 196668 136226
rect 196736 136170 196792 136226
rect 196860 136170 196916 136226
rect 196984 136170 197040 136226
rect 196612 136046 196668 136102
rect 196736 136046 196792 136102
rect 196860 136046 196916 136102
rect 196984 136046 197040 136102
rect 196612 135922 196668 135978
rect 196736 135922 196792 135978
rect 196860 135922 196916 135978
rect 196984 135922 197040 135978
rect 195812 130294 195868 130350
rect 195936 130294 195992 130350
rect 196060 130294 196116 130350
rect 196184 130294 196240 130350
rect 195812 130170 195868 130226
rect 195936 130170 195992 130226
rect 196060 130170 196116 130226
rect 196184 130170 196240 130226
rect 195812 130046 195868 130102
rect 195936 130046 195992 130102
rect 196060 130046 196116 130102
rect 196184 130046 196240 130102
rect 195812 129922 195868 129978
rect 195936 129922 195992 129978
rect 196060 129922 196116 129978
rect 196184 129922 196240 129978
rect 193554 118294 193610 118350
rect 193678 118294 193734 118350
rect 193802 118294 193858 118350
rect 193926 118294 193982 118350
rect 193554 118170 193610 118226
rect 193678 118170 193734 118226
rect 193802 118170 193858 118226
rect 193926 118170 193982 118226
rect 193554 118046 193610 118102
rect 193678 118046 193734 118102
rect 193802 118046 193858 118102
rect 193926 118046 193982 118102
rect 193554 117922 193610 117978
rect 193678 117922 193734 117978
rect 193802 117922 193858 117978
rect 193926 117922 193982 117978
rect 196612 118294 196668 118350
rect 196736 118294 196792 118350
rect 196860 118294 196916 118350
rect 196984 118294 197040 118350
rect 196612 118170 196668 118226
rect 196736 118170 196792 118226
rect 196860 118170 196916 118226
rect 196984 118170 197040 118226
rect 196612 118046 196668 118102
rect 196736 118046 196792 118102
rect 196860 118046 196916 118102
rect 196984 118046 197040 118102
rect 196612 117922 196668 117978
rect 196736 117922 196792 117978
rect 196860 117922 196916 117978
rect 196984 117922 197040 117978
rect 195812 112294 195868 112350
rect 195936 112294 195992 112350
rect 196060 112294 196116 112350
rect 196184 112294 196240 112350
rect 195812 112170 195868 112226
rect 195936 112170 195992 112226
rect 196060 112170 196116 112226
rect 196184 112170 196240 112226
rect 195812 112046 195868 112102
rect 195936 112046 195992 112102
rect 196060 112046 196116 112102
rect 196184 112046 196240 112102
rect 195812 111922 195868 111978
rect 195936 111922 195992 111978
rect 196060 111922 196116 111978
rect 196184 111922 196240 111978
rect 193554 100294 193610 100350
rect 193678 100294 193734 100350
rect 193802 100294 193858 100350
rect 193926 100294 193982 100350
rect 193554 100170 193610 100226
rect 193678 100170 193734 100226
rect 193802 100170 193858 100226
rect 193926 100170 193982 100226
rect 193554 100046 193610 100102
rect 193678 100046 193734 100102
rect 193802 100046 193858 100102
rect 193926 100046 193982 100102
rect 193554 99922 193610 99978
rect 193678 99922 193734 99978
rect 193802 99922 193858 99978
rect 193926 99922 193982 99978
rect 196612 100294 196668 100350
rect 196736 100294 196792 100350
rect 196860 100294 196916 100350
rect 196984 100294 197040 100350
rect 196612 100170 196668 100226
rect 196736 100170 196792 100226
rect 196860 100170 196916 100226
rect 196984 100170 197040 100226
rect 196612 100046 196668 100102
rect 196736 100046 196792 100102
rect 196860 100046 196916 100102
rect 196984 100046 197040 100102
rect 196612 99922 196668 99978
rect 196736 99922 196792 99978
rect 196860 99922 196916 99978
rect 196984 99922 197040 99978
rect 195812 94294 195868 94350
rect 195936 94294 195992 94350
rect 196060 94294 196116 94350
rect 196184 94294 196240 94350
rect 195812 94170 195868 94226
rect 195936 94170 195992 94226
rect 196060 94170 196116 94226
rect 196184 94170 196240 94226
rect 195812 94046 195868 94102
rect 195936 94046 195992 94102
rect 196060 94046 196116 94102
rect 196184 94046 196240 94102
rect 195812 93922 195868 93978
rect 195936 93922 195992 93978
rect 196060 93922 196116 93978
rect 196184 93922 196240 93978
rect 205884 364562 205940 364618
rect 205100 358982 205156 359038
rect 204988 357362 205044 357418
rect 204876 306602 204932 306658
rect 205772 358622 205828 358678
rect 204988 223442 205044 223498
rect 204988 222542 205044 222598
rect 204876 204902 204932 204958
rect 204988 201482 205044 201538
rect 204988 191402 205044 191458
rect 204988 185642 205044 185698
rect 204988 178082 205044 178138
rect 204988 172682 205044 172738
rect 205212 193022 205268 193078
rect 206108 363122 206164 363178
rect 207452 362042 207508 362098
rect 206668 219122 206724 219178
rect 206668 218222 206724 218278
rect 206668 214982 206724 215038
rect 206668 212462 206724 212518
rect 206668 209942 206724 209998
rect 206668 198962 206724 199018
rect 206892 195722 206948 195778
rect 206668 176462 206724 176518
rect 206892 173042 206948 173098
rect 206780 162782 206836 162838
rect 193554 82294 193610 82350
rect 193678 82294 193734 82350
rect 193802 82294 193858 82350
rect 193926 82294 193982 82350
rect 193554 82170 193610 82226
rect 193678 82170 193734 82226
rect 193802 82170 193858 82226
rect 193926 82170 193982 82226
rect 193554 82046 193610 82102
rect 193678 82046 193734 82102
rect 193802 82046 193858 82102
rect 193926 82046 193982 82102
rect 193554 81922 193610 81978
rect 193678 81922 193734 81978
rect 193802 81922 193858 81978
rect 193926 81922 193982 81978
rect 196612 82294 196668 82350
rect 196736 82294 196792 82350
rect 196860 82294 196916 82350
rect 196984 82294 197040 82350
rect 196612 82170 196668 82226
rect 196736 82170 196792 82226
rect 196860 82170 196916 82226
rect 196984 82170 197040 82226
rect 196612 82046 196668 82102
rect 196736 82046 196792 82102
rect 196860 82046 196916 82102
rect 196984 82046 197040 82102
rect 196612 81922 196668 81978
rect 196736 81922 196792 81978
rect 196860 81922 196916 81978
rect 196984 81922 197040 81978
rect 195812 76294 195868 76350
rect 195936 76294 195992 76350
rect 196060 76294 196116 76350
rect 196184 76294 196240 76350
rect 195812 76170 195868 76226
rect 195936 76170 195992 76226
rect 196060 76170 196116 76226
rect 196184 76170 196240 76226
rect 195812 76046 195868 76102
rect 195936 76046 195992 76102
rect 196060 76046 196116 76102
rect 196184 76046 196240 76102
rect 195812 75922 195868 75978
rect 195936 75922 195992 75978
rect 196060 75922 196116 75978
rect 196184 75922 196240 75978
rect 193554 64294 193610 64350
rect 193678 64294 193734 64350
rect 193802 64294 193858 64350
rect 193926 64294 193982 64350
rect 193554 64170 193610 64226
rect 193678 64170 193734 64226
rect 193802 64170 193858 64226
rect 193926 64170 193982 64226
rect 193554 64046 193610 64102
rect 193678 64046 193734 64102
rect 193802 64046 193858 64102
rect 193926 64046 193982 64102
rect 193554 63922 193610 63978
rect 193678 63922 193734 63978
rect 193802 63922 193858 63978
rect 193926 63922 193982 63978
rect 196612 64294 196668 64350
rect 196736 64294 196792 64350
rect 196860 64294 196916 64350
rect 196984 64294 197040 64350
rect 196612 64170 196668 64226
rect 196736 64170 196792 64226
rect 196860 64170 196916 64226
rect 196984 64170 197040 64226
rect 196612 64046 196668 64102
rect 196736 64046 196792 64102
rect 196860 64046 196916 64102
rect 196984 64046 197040 64102
rect 196612 63922 196668 63978
rect 196736 63922 196792 63978
rect 196860 63922 196916 63978
rect 196984 63922 197040 63978
rect 195812 58294 195868 58350
rect 195936 58294 195992 58350
rect 196060 58294 196116 58350
rect 196184 58294 196240 58350
rect 195812 58170 195868 58226
rect 195936 58170 195992 58226
rect 196060 58170 196116 58226
rect 196184 58170 196240 58226
rect 195812 58046 195868 58102
rect 195936 58046 195992 58102
rect 196060 58046 196116 58102
rect 196184 58046 196240 58102
rect 195812 57922 195868 57978
rect 195936 57922 195992 57978
rect 196060 57922 196116 57978
rect 196184 57922 196240 57978
rect 209132 361502 209188 361558
rect 208348 357182 208404 357238
rect 208460 357002 208516 357058
rect 209580 277082 209636 277138
rect 209580 276542 209636 276598
rect 210700 276362 210756 276418
rect 210700 257822 210756 257878
rect 210700 236042 210756 236098
rect 212044 358802 212100 358858
rect 212268 362942 212324 362998
rect 212156 306602 212212 306658
rect 213388 277082 213444 277138
rect 212044 276722 212100 276778
rect 211932 276542 211988 276598
rect 220554 364294 220610 364350
rect 220678 364294 220734 364350
rect 220802 364294 220858 364350
rect 220926 364294 220982 364350
rect 220554 364170 220610 364226
rect 220678 364170 220734 364226
rect 220802 364170 220858 364226
rect 220926 364170 220982 364226
rect 220554 364046 220610 364102
rect 220678 364046 220734 364102
rect 220802 364046 220858 364102
rect 220926 364046 220982 364102
rect 220554 363922 220610 363978
rect 220678 363922 220734 363978
rect 220802 363922 220858 363978
rect 220926 363922 220982 363978
rect 220554 346294 220610 346350
rect 220678 346294 220734 346350
rect 220802 346294 220858 346350
rect 220926 346294 220982 346350
rect 220554 346170 220610 346226
rect 220678 346170 220734 346226
rect 220802 346170 220858 346226
rect 220926 346170 220982 346226
rect 220554 346046 220610 346102
rect 220678 346046 220734 346102
rect 220802 346046 220858 346102
rect 220926 346046 220982 346102
rect 220554 345922 220610 345978
rect 220678 345922 220734 345978
rect 220802 345922 220858 345978
rect 220926 345922 220982 345978
rect 220554 328294 220610 328350
rect 220678 328294 220734 328350
rect 220802 328294 220858 328350
rect 220926 328294 220982 328350
rect 220554 328170 220610 328226
rect 220678 328170 220734 328226
rect 220802 328170 220858 328226
rect 220926 328170 220982 328226
rect 220554 328046 220610 328102
rect 220678 328046 220734 328102
rect 220802 328046 220858 328102
rect 220926 328046 220982 328102
rect 220554 327922 220610 327978
rect 220678 327922 220734 327978
rect 220802 327922 220858 327978
rect 220926 327922 220982 327978
rect 224274 598116 224330 598172
rect 224398 598116 224454 598172
rect 224522 598116 224578 598172
rect 224646 598116 224702 598172
rect 224274 597992 224330 598048
rect 224398 597992 224454 598048
rect 224522 597992 224578 598048
rect 224646 597992 224702 598048
rect 224274 597868 224330 597924
rect 224398 597868 224454 597924
rect 224522 597868 224578 597924
rect 224646 597868 224702 597924
rect 224274 597744 224330 597800
rect 224398 597744 224454 597800
rect 224522 597744 224578 597800
rect 224646 597744 224702 597800
rect 224274 586294 224330 586350
rect 224398 586294 224454 586350
rect 224522 586294 224578 586350
rect 224646 586294 224702 586350
rect 224274 586170 224330 586226
rect 224398 586170 224454 586226
rect 224522 586170 224578 586226
rect 224646 586170 224702 586226
rect 224274 586046 224330 586102
rect 224398 586046 224454 586102
rect 224522 586046 224578 586102
rect 224646 586046 224702 586102
rect 224274 585922 224330 585978
rect 224398 585922 224454 585978
rect 224522 585922 224578 585978
rect 224646 585922 224702 585978
rect 224274 568294 224330 568350
rect 224398 568294 224454 568350
rect 224522 568294 224578 568350
rect 224646 568294 224702 568350
rect 224274 568170 224330 568226
rect 224398 568170 224454 568226
rect 224522 568170 224578 568226
rect 224646 568170 224702 568226
rect 224274 568046 224330 568102
rect 224398 568046 224454 568102
rect 224522 568046 224578 568102
rect 224646 568046 224702 568102
rect 224274 567922 224330 567978
rect 224398 567922 224454 567978
rect 224522 567922 224578 567978
rect 224646 567922 224702 567978
rect 224274 550294 224330 550350
rect 224398 550294 224454 550350
rect 224522 550294 224578 550350
rect 224646 550294 224702 550350
rect 224274 550170 224330 550226
rect 224398 550170 224454 550226
rect 224522 550170 224578 550226
rect 224646 550170 224702 550226
rect 224274 550046 224330 550102
rect 224398 550046 224454 550102
rect 224522 550046 224578 550102
rect 224646 550046 224702 550102
rect 224274 549922 224330 549978
rect 224398 549922 224454 549978
rect 224522 549922 224578 549978
rect 224646 549922 224702 549978
rect 224274 532294 224330 532350
rect 224398 532294 224454 532350
rect 224522 532294 224578 532350
rect 224646 532294 224702 532350
rect 224274 532170 224330 532226
rect 224398 532170 224454 532226
rect 224522 532170 224578 532226
rect 224646 532170 224702 532226
rect 224274 532046 224330 532102
rect 224398 532046 224454 532102
rect 224522 532046 224578 532102
rect 224646 532046 224702 532102
rect 224274 531922 224330 531978
rect 224398 531922 224454 531978
rect 224522 531922 224578 531978
rect 224646 531922 224702 531978
rect 224274 514294 224330 514350
rect 224398 514294 224454 514350
rect 224522 514294 224578 514350
rect 224646 514294 224702 514350
rect 224274 514170 224330 514226
rect 224398 514170 224454 514226
rect 224522 514170 224578 514226
rect 224646 514170 224702 514226
rect 224274 514046 224330 514102
rect 224398 514046 224454 514102
rect 224522 514046 224578 514102
rect 224646 514046 224702 514102
rect 224274 513922 224330 513978
rect 224398 513922 224454 513978
rect 224522 513922 224578 513978
rect 224646 513922 224702 513978
rect 224274 496294 224330 496350
rect 224398 496294 224454 496350
rect 224522 496294 224578 496350
rect 224646 496294 224702 496350
rect 224274 496170 224330 496226
rect 224398 496170 224454 496226
rect 224522 496170 224578 496226
rect 224646 496170 224702 496226
rect 224274 496046 224330 496102
rect 224398 496046 224454 496102
rect 224522 496046 224578 496102
rect 224646 496046 224702 496102
rect 224274 495922 224330 495978
rect 224398 495922 224454 495978
rect 224522 495922 224578 495978
rect 224646 495922 224702 495978
rect 224274 478294 224330 478350
rect 224398 478294 224454 478350
rect 224522 478294 224578 478350
rect 224646 478294 224702 478350
rect 224274 478170 224330 478226
rect 224398 478170 224454 478226
rect 224522 478170 224578 478226
rect 224646 478170 224702 478226
rect 224274 478046 224330 478102
rect 224398 478046 224454 478102
rect 224522 478046 224578 478102
rect 224646 478046 224702 478102
rect 224274 477922 224330 477978
rect 224398 477922 224454 477978
rect 224522 477922 224578 477978
rect 224646 477922 224702 477978
rect 224274 460294 224330 460350
rect 224398 460294 224454 460350
rect 224522 460294 224578 460350
rect 224646 460294 224702 460350
rect 224274 460170 224330 460226
rect 224398 460170 224454 460226
rect 224522 460170 224578 460226
rect 224646 460170 224702 460226
rect 224274 460046 224330 460102
rect 224398 460046 224454 460102
rect 224522 460046 224578 460102
rect 224646 460046 224702 460102
rect 224274 459922 224330 459978
rect 224398 459922 224454 459978
rect 224522 459922 224578 459978
rect 224646 459922 224702 459978
rect 224274 442294 224330 442350
rect 224398 442294 224454 442350
rect 224522 442294 224578 442350
rect 224646 442294 224702 442350
rect 224274 442170 224330 442226
rect 224398 442170 224454 442226
rect 224522 442170 224578 442226
rect 224646 442170 224702 442226
rect 224274 442046 224330 442102
rect 224398 442046 224454 442102
rect 224522 442046 224578 442102
rect 224646 442046 224702 442102
rect 224274 441922 224330 441978
rect 224398 441922 224454 441978
rect 224522 441922 224578 441978
rect 224646 441922 224702 441978
rect 224274 424294 224330 424350
rect 224398 424294 224454 424350
rect 224522 424294 224578 424350
rect 224646 424294 224702 424350
rect 224274 424170 224330 424226
rect 224398 424170 224454 424226
rect 224522 424170 224578 424226
rect 224646 424170 224702 424226
rect 224274 424046 224330 424102
rect 224398 424046 224454 424102
rect 224522 424046 224578 424102
rect 224646 424046 224702 424102
rect 224274 423922 224330 423978
rect 224398 423922 224454 423978
rect 224522 423922 224578 423978
rect 224646 423922 224702 423978
rect 224274 406294 224330 406350
rect 224398 406294 224454 406350
rect 224522 406294 224578 406350
rect 224646 406294 224702 406350
rect 224274 406170 224330 406226
rect 224398 406170 224454 406226
rect 224522 406170 224578 406226
rect 224646 406170 224702 406226
rect 224274 406046 224330 406102
rect 224398 406046 224454 406102
rect 224522 406046 224578 406102
rect 224646 406046 224702 406102
rect 224274 405922 224330 405978
rect 224398 405922 224454 405978
rect 224522 405922 224578 405978
rect 224646 405922 224702 405978
rect 224274 388294 224330 388350
rect 224398 388294 224454 388350
rect 224522 388294 224578 388350
rect 224646 388294 224702 388350
rect 224274 388170 224330 388226
rect 224398 388170 224454 388226
rect 224522 388170 224578 388226
rect 224646 388170 224702 388226
rect 224274 388046 224330 388102
rect 224398 388046 224454 388102
rect 224522 388046 224578 388102
rect 224646 388046 224702 388102
rect 224274 387922 224330 387978
rect 224398 387922 224454 387978
rect 224522 387922 224578 387978
rect 224646 387922 224702 387978
rect 224274 370294 224330 370350
rect 224398 370294 224454 370350
rect 224522 370294 224578 370350
rect 224646 370294 224702 370350
rect 224274 370170 224330 370226
rect 224398 370170 224454 370226
rect 224522 370170 224578 370226
rect 224646 370170 224702 370226
rect 224274 370046 224330 370102
rect 224398 370046 224454 370102
rect 224522 370046 224578 370102
rect 224646 370046 224702 370102
rect 224274 369922 224330 369978
rect 224398 369922 224454 369978
rect 224522 369922 224578 369978
rect 224646 369922 224702 369978
rect 224274 352294 224330 352350
rect 224398 352294 224454 352350
rect 224522 352294 224578 352350
rect 224646 352294 224702 352350
rect 224274 352170 224330 352226
rect 224398 352170 224454 352226
rect 224522 352170 224578 352226
rect 224646 352170 224702 352226
rect 224274 352046 224330 352102
rect 224398 352046 224454 352102
rect 224522 352046 224578 352102
rect 224646 352046 224702 352102
rect 224274 351922 224330 351978
rect 224398 351922 224454 351978
rect 224522 351922 224578 351978
rect 224646 351922 224702 351978
rect 224274 334294 224330 334350
rect 224398 334294 224454 334350
rect 224522 334294 224578 334350
rect 224646 334294 224702 334350
rect 224274 334170 224330 334226
rect 224398 334170 224454 334226
rect 224522 334170 224578 334226
rect 224646 334170 224702 334226
rect 224274 334046 224330 334102
rect 224398 334046 224454 334102
rect 224522 334046 224578 334102
rect 224646 334046 224702 334102
rect 224274 333922 224330 333978
rect 224398 333922 224454 333978
rect 224522 333922 224578 333978
rect 224646 333922 224702 333978
rect 251274 597156 251330 597212
rect 251398 597156 251454 597212
rect 251522 597156 251578 597212
rect 251646 597156 251702 597212
rect 251274 597032 251330 597088
rect 251398 597032 251454 597088
rect 251522 597032 251578 597088
rect 251646 597032 251702 597088
rect 251274 596908 251330 596964
rect 251398 596908 251454 596964
rect 251522 596908 251578 596964
rect 251646 596908 251702 596964
rect 251274 596784 251330 596840
rect 251398 596784 251454 596840
rect 251522 596784 251578 596840
rect 251646 596784 251702 596840
rect 251274 580294 251330 580350
rect 251398 580294 251454 580350
rect 251522 580294 251578 580350
rect 251646 580294 251702 580350
rect 251274 580170 251330 580226
rect 251398 580170 251454 580226
rect 251522 580170 251578 580226
rect 251646 580170 251702 580226
rect 251274 580046 251330 580102
rect 251398 580046 251454 580102
rect 251522 580046 251578 580102
rect 251646 580046 251702 580102
rect 251274 579922 251330 579978
rect 251398 579922 251454 579978
rect 251522 579922 251578 579978
rect 251646 579922 251702 579978
rect 251274 562294 251330 562350
rect 251398 562294 251454 562350
rect 251522 562294 251578 562350
rect 251646 562294 251702 562350
rect 251274 562170 251330 562226
rect 251398 562170 251454 562226
rect 251522 562170 251578 562226
rect 251646 562170 251702 562226
rect 251274 562046 251330 562102
rect 251398 562046 251454 562102
rect 251522 562046 251578 562102
rect 251646 562046 251702 562102
rect 251274 561922 251330 561978
rect 251398 561922 251454 561978
rect 251522 561922 251578 561978
rect 251646 561922 251702 561978
rect 251274 544294 251330 544350
rect 251398 544294 251454 544350
rect 251522 544294 251578 544350
rect 251646 544294 251702 544350
rect 251274 544170 251330 544226
rect 251398 544170 251454 544226
rect 251522 544170 251578 544226
rect 251646 544170 251702 544226
rect 251274 544046 251330 544102
rect 251398 544046 251454 544102
rect 251522 544046 251578 544102
rect 251646 544046 251702 544102
rect 251274 543922 251330 543978
rect 251398 543922 251454 543978
rect 251522 543922 251578 543978
rect 251646 543922 251702 543978
rect 251274 526294 251330 526350
rect 251398 526294 251454 526350
rect 251522 526294 251578 526350
rect 251646 526294 251702 526350
rect 251274 526170 251330 526226
rect 251398 526170 251454 526226
rect 251522 526170 251578 526226
rect 251646 526170 251702 526226
rect 251274 526046 251330 526102
rect 251398 526046 251454 526102
rect 251522 526046 251578 526102
rect 251646 526046 251702 526102
rect 251274 525922 251330 525978
rect 251398 525922 251454 525978
rect 251522 525922 251578 525978
rect 251646 525922 251702 525978
rect 251274 508294 251330 508350
rect 251398 508294 251454 508350
rect 251522 508294 251578 508350
rect 251646 508294 251702 508350
rect 251274 508170 251330 508226
rect 251398 508170 251454 508226
rect 251522 508170 251578 508226
rect 251646 508170 251702 508226
rect 251274 508046 251330 508102
rect 251398 508046 251454 508102
rect 251522 508046 251578 508102
rect 251646 508046 251702 508102
rect 251274 507922 251330 507978
rect 251398 507922 251454 507978
rect 251522 507922 251578 507978
rect 251646 507922 251702 507978
rect 251274 490294 251330 490350
rect 251398 490294 251454 490350
rect 251522 490294 251578 490350
rect 251646 490294 251702 490350
rect 251274 490170 251330 490226
rect 251398 490170 251454 490226
rect 251522 490170 251578 490226
rect 251646 490170 251702 490226
rect 251274 490046 251330 490102
rect 251398 490046 251454 490102
rect 251522 490046 251578 490102
rect 251646 490046 251702 490102
rect 251274 489922 251330 489978
rect 251398 489922 251454 489978
rect 251522 489922 251578 489978
rect 251646 489922 251702 489978
rect 251274 472294 251330 472350
rect 251398 472294 251454 472350
rect 251522 472294 251578 472350
rect 251646 472294 251702 472350
rect 251274 472170 251330 472226
rect 251398 472170 251454 472226
rect 251522 472170 251578 472226
rect 251646 472170 251702 472226
rect 251274 472046 251330 472102
rect 251398 472046 251454 472102
rect 251522 472046 251578 472102
rect 251646 472046 251702 472102
rect 251274 471922 251330 471978
rect 251398 471922 251454 471978
rect 251522 471922 251578 471978
rect 251646 471922 251702 471978
rect 251274 454294 251330 454350
rect 251398 454294 251454 454350
rect 251522 454294 251578 454350
rect 251646 454294 251702 454350
rect 251274 454170 251330 454226
rect 251398 454170 251454 454226
rect 251522 454170 251578 454226
rect 251646 454170 251702 454226
rect 251274 454046 251330 454102
rect 251398 454046 251454 454102
rect 251522 454046 251578 454102
rect 251646 454046 251702 454102
rect 251274 453922 251330 453978
rect 251398 453922 251454 453978
rect 251522 453922 251578 453978
rect 251646 453922 251702 453978
rect 251274 436294 251330 436350
rect 251398 436294 251454 436350
rect 251522 436294 251578 436350
rect 251646 436294 251702 436350
rect 251274 436170 251330 436226
rect 251398 436170 251454 436226
rect 251522 436170 251578 436226
rect 251646 436170 251702 436226
rect 251274 436046 251330 436102
rect 251398 436046 251454 436102
rect 251522 436046 251578 436102
rect 251646 436046 251702 436102
rect 251274 435922 251330 435978
rect 251398 435922 251454 435978
rect 251522 435922 251578 435978
rect 251646 435922 251702 435978
rect 251274 418294 251330 418350
rect 251398 418294 251454 418350
rect 251522 418294 251578 418350
rect 251646 418294 251702 418350
rect 251274 418170 251330 418226
rect 251398 418170 251454 418226
rect 251522 418170 251578 418226
rect 251646 418170 251702 418226
rect 251274 418046 251330 418102
rect 251398 418046 251454 418102
rect 251522 418046 251578 418102
rect 251646 418046 251702 418102
rect 251274 417922 251330 417978
rect 251398 417922 251454 417978
rect 251522 417922 251578 417978
rect 251646 417922 251702 417978
rect 251274 400294 251330 400350
rect 251398 400294 251454 400350
rect 251522 400294 251578 400350
rect 251646 400294 251702 400350
rect 251274 400170 251330 400226
rect 251398 400170 251454 400226
rect 251522 400170 251578 400226
rect 251646 400170 251702 400226
rect 251274 400046 251330 400102
rect 251398 400046 251454 400102
rect 251522 400046 251578 400102
rect 251646 400046 251702 400102
rect 251274 399922 251330 399978
rect 251398 399922 251454 399978
rect 251522 399922 251578 399978
rect 251646 399922 251702 399978
rect 251274 382294 251330 382350
rect 251398 382294 251454 382350
rect 251522 382294 251578 382350
rect 251646 382294 251702 382350
rect 251274 382170 251330 382226
rect 251398 382170 251454 382226
rect 251522 382170 251578 382226
rect 251646 382170 251702 382226
rect 251274 382046 251330 382102
rect 251398 382046 251454 382102
rect 251522 382046 251578 382102
rect 251646 382046 251702 382102
rect 251274 381922 251330 381978
rect 251398 381922 251454 381978
rect 251522 381922 251578 381978
rect 251646 381922 251702 381978
rect 251274 364294 251330 364350
rect 251398 364294 251454 364350
rect 251522 364294 251578 364350
rect 251646 364294 251702 364350
rect 251274 364170 251330 364226
rect 251398 364170 251454 364226
rect 251522 364170 251578 364226
rect 251646 364170 251702 364226
rect 251274 364046 251330 364102
rect 251398 364046 251454 364102
rect 251522 364046 251578 364102
rect 251646 364046 251702 364102
rect 251274 363922 251330 363978
rect 251398 363922 251454 363978
rect 251522 363922 251578 363978
rect 251646 363922 251702 363978
rect 251274 346294 251330 346350
rect 251398 346294 251454 346350
rect 251522 346294 251578 346350
rect 251646 346294 251702 346350
rect 251274 346170 251330 346226
rect 251398 346170 251454 346226
rect 251522 346170 251578 346226
rect 251646 346170 251702 346226
rect 251274 346046 251330 346102
rect 251398 346046 251454 346102
rect 251522 346046 251578 346102
rect 251646 346046 251702 346102
rect 251274 345922 251330 345978
rect 251398 345922 251454 345978
rect 251522 345922 251578 345978
rect 251646 345922 251702 345978
rect 251274 328294 251330 328350
rect 251398 328294 251454 328350
rect 251522 328294 251578 328350
rect 251646 328294 251702 328350
rect 251274 328170 251330 328226
rect 251398 328170 251454 328226
rect 251522 328170 251578 328226
rect 251646 328170 251702 328226
rect 251274 328046 251330 328102
rect 251398 328046 251454 328102
rect 251522 328046 251578 328102
rect 251646 328046 251702 328102
rect 251274 327922 251330 327978
rect 251398 327922 251454 327978
rect 251522 327922 251578 327978
rect 251646 327922 251702 327978
rect 254994 598116 255050 598172
rect 255118 598116 255174 598172
rect 255242 598116 255298 598172
rect 255366 598116 255422 598172
rect 254994 597992 255050 598048
rect 255118 597992 255174 598048
rect 255242 597992 255298 598048
rect 255366 597992 255422 598048
rect 254994 597868 255050 597924
rect 255118 597868 255174 597924
rect 255242 597868 255298 597924
rect 255366 597868 255422 597924
rect 254994 597744 255050 597800
rect 255118 597744 255174 597800
rect 255242 597744 255298 597800
rect 255366 597744 255422 597800
rect 254994 586294 255050 586350
rect 255118 586294 255174 586350
rect 255242 586294 255298 586350
rect 255366 586294 255422 586350
rect 254994 586170 255050 586226
rect 255118 586170 255174 586226
rect 255242 586170 255298 586226
rect 255366 586170 255422 586226
rect 254994 586046 255050 586102
rect 255118 586046 255174 586102
rect 255242 586046 255298 586102
rect 255366 586046 255422 586102
rect 254994 585922 255050 585978
rect 255118 585922 255174 585978
rect 255242 585922 255298 585978
rect 255366 585922 255422 585978
rect 254994 568294 255050 568350
rect 255118 568294 255174 568350
rect 255242 568294 255298 568350
rect 255366 568294 255422 568350
rect 254994 568170 255050 568226
rect 255118 568170 255174 568226
rect 255242 568170 255298 568226
rect 255366 568170 255422 568226
rect 254994 568046 255050 568102
rect 255118 568046 255174 568102
rect 255242 568046 255298 568102
rect 255366 568046 255422 568102
rect 254994 567922 255050 567978
rect 255118 567922 255174 567978
rect 255242 567922 255298 567978
rect 255366 567922 255422 567978
rect 254994 550294 255050 550350
rect 255118 550294 255174 550350
rect 255242 550294 255298 550350
rect 255366 550294 255422 550350
rect 254994 550170 255050 550226
rect 255118 550170 255174 550226
rect 255242 550170 255298 550226
rect 255366 550170 255422 550226
rect 254994 550046 255050 550102
rect 255118 550046 255174 550102
rect 255242 550046 255298 550102
rect 255366 550046 255422 550102
rect 254994 549922 255050 549978
rect 255118 549922 255174 549978
rect 255242 549922 255298 549978
rect 255366 549922 255422 549978
rect 254994 532294 255050 532350
rect 255118 532294 255174 532350
rect 255242 532294 255298 532350
rect 255366 532294 255422 532350
rect 254994 532170 255050 532226
rect 255118 532170 255174 532226
rect 255242 532170 255298 532226
rect 255366 532170 255422 532226
rect 254994 532046 255050 532102
rect 255118 532046 255174 532102
rect 255242 532046 255298 532102
rect 255366 532046 255422 532102
rect 254994 531922 255050 531978
rect 255118 531922 255174 531978
rect 255242 531922 255298 531978
rect 255366 531922 255422 531978
rect 254994 514294 255050 514350
rect 255118 514294 255174 514350
rect 255242 514294 255298 514350
rect 255366 514294 255422 514350
rect 254994 514170 255050 514226
rect 255118 514170 255174 514226
rect 255242 514170 255298 514226
rect 255366 514170 255422 514226
rect 254994 514046 255050 514102
rect 255118 514046 255174 514102
rect 255242 514046 255298 514102
rect 255366 514046 255422 514102
rect 254994 513922 255050 513978
rect 255118 513922 255174 513978
rect 255242 513922 255298 513978
rect 255366 513922 255422 513978
rect 254994 496294 255050 496350
rect 255118 496294 255174 496350
rect 255242 496294 255298 496350
rect 255366 496294 255422 496350
rect 254994 496170 255050 496226
rect 255118 496170 255174 496226
rect 255242 496170 255298 496226
rect 255366 496170 255422 496226
rect 254994 496046 255050 496102
rect 255118 496046 255174 496102
rect 255242 496046 255298 496102
rect 255366 496046 255422 496102
rect 254994 495922 255050 495978
rect 255118 495922 255174 495978
rect 255242 495922 255298 495978
rect 255366 495922 255422 495978
rect 254994 478294 255050 478350
rect 255118 478294 255174 478350
rect 255242 478294 255298 478350
rect 255366 478294 255422 478350
rect 254994 478170 255050 478226
rect 255118 478170 255174 478226
rect 255242 478170 255298 478226
rect 255366 478170 255422 478226
rect 254994 478046 255050 478102
rect 255118 478046 255174 478102
rect 255242 478046 255298 478102
rect 255366 478046 255422 478102
rect 254994 477922 255050 477978
rect 255118 477922 255174 477978
rect 255242 477922 255298 477978
rect 255366 477922 255422 477978
rect 254994 460294 255050 460350
rect 255118 460294 255174 460350
rect 255242 460294 255298 460350
rect 255366 460294 255422 460350
rect 254994 460170 255050 460226
rect 255118 460170 255174 460226
rect 255242 460170 255298 460226
rect 255366 460170 255422 460226
rect 254994 460046 255050 460102
rect 255118 460046 255174 460102
rect 255242 460046 255298 460102
rect 255366 460046 255422 460102
rect 254994 459922 255050 459978
rect 255118 459922 255174 459978
rect 255242 459922 255298 459978
rect 255366 459922 255422 459978
rect 254994 442294 255050 442350
rect 255118 442294 255174 442350
rect 255242 442294 255298 442350
rect 255366 442294 255422 442350
rect 254994 442170 255050 442226
rect 255118 442170 255174 442226
rect 255242 442170 255298 442226
rect 255366 442170 255422 442226
rect 254994 442046 255050 442102
rect 255118 442046 255174 442102
rect 255242 442046 255298 442102
rect 255366 442046 255422 442102
rect 254994 441922 255050 441978
rect 255118 441922 255174 441978
rect 255242 441922 255298 441978
rect 255366 441922 255422 441978
rect 254994 424294 255050 424350
rect 255118 424294 255174 424350
rect 255242 424294 255298 424350
rect 255366 424294 255422 424350
rect 254994 424170 255050 424226
rect 255118 424170 255174 424226
rect 255242 424170 255298 424226
rect 255366 424170 255422 424226
rect 254994 424046 255050 424102
rect 255118 424046 255174 424102
rect 255242 424046 255298 424102
rect 255366 424046 255422 424102
rect 254994 423922 255050 423978
rect 255118 423922 255174 423978
rect 255242 423922 255298 423978
rect 255366 423922 255422 423978
rect 254994 406294 255050 406350
rect 255118 406294 255174 406350
rect 255242 406294 255298 406350
rect 255366 406294 255422 406350
rect 254994 406170 255050 406226
rect 255118 406170 255174 406226
rect 255242 406170 255298 406226
rect 255366 406170 255422 406226
rect 254994 406046 255050 406102
rect 255118 406046 255174 406102
rect 255242 406046 255298 406102
rect 255366 406046 255422 406102
rect 254994 405922 255050 405978
rect 255118 405922 255174 405978
rect 255242 405922 255298 405978
rect 255366 405922 255422 405978
rect 254994 388294 255050 388350
rect 255118 388294 255174 388350
rect 255242 388294 255298 388350
rect 255366 388294 255422 388350
rect 254994 388170 255050 388226
rect 255118 388170 255174 388226
rect 255242 388170 255298 388226
rect 255366 388170 255422 388226
rect 254994 388046 255050 388102
rect 255118 388046 255174 388102
rect 255242 388046 255298 388102
rect 255366 388046 255422 388102
rect 254994 387922 255050 387978
rect 255118 387922 255174 387978
rect 255242 387922 255298 387978
rect 255366 387922 255422 387978
rect 254994 370294 255050 370350
rect 255118 370294 255174 370350
rect 255242 370294 255298 370350
rect 255366 370294 255422 370350
rect 254994 370170 255050 370226
rect 255118 370170 255174 370226
rect 255242 370170 255298 370226
rect 255366 370170 255422 370226
rect 254994 370046 255050 370102
rect 255118 370046 255174 370102
rect 255242 370046 255298 370102
rect 255366 370046 255422 370102
rect 254994 369922 255050 369978
rect 255118 369922 255174 369978
rect 255242 369922 255298 369978
rect 255366 369922 255422 369978
rect 254994 352294 255050 352350
rect 255118 352294 255174 352350
rect 255242 352294 255298 352350
rect 255366 352294 255422 352350
rect 254994 352170 255050 352226
rect 255118 352170 255174 352226
rect 255242 352170 255298 352226
rect 255366 352170 255422 352226
rect 254994 352046 255050 352102
rect 255118 352046 255174 352102
rect 255242 352046 255298 352102
rect 255366 352046 255422 352102
rect 254994 351922 255050 351978
rect 255118 351922 255174 351978
rect 255242 351922 255298 351978
rect 255366 351922 255422 351978
rect 254994 334294 255050 334350
rect 255118 334294 255174 334350
rect 255242 334294 255298 334350
rect 255366 334294 255422 334350
rect 254994 334170 255050 334226
rect 255118 334170 255174 334226
rect 255242 334170 255298 334226
rect 255366 334170 255422 334226
rect 254994 334046 255050 334102
rect 255118 334046 255174 334102
rect 255242 334046 255298 334102
rect 255366 334046 255422 334102
rect 254994 333922 255050 333978
rect 255118 333922 255174 333978
rect 255242 333922 255298 333978
rect 255366 333922 255422 333978
rect 281994 597156 282050 597212
rect 282118 597156 282174 597212
rect 282242 597156 282298 597212
rect 282366 597156 282422 597212
rect 281994 597032 282050 597088
rect 282118 597032 282174 597088
rect 282242 597032 282298 597088
rect 282366 597032 282422 597088
rect 281994 596908 282050 596964
rect 282118 596908 282174 596964
rect 282242 596908 282298 596964
rect 282366 596908 282422 596964
rect 281994 596784 282050 596840
rect 282118 596784 282174 596840
rect 282242 596784 282298 596840
rect 282366 596784 282422 596840
rect 281994 580294 282050 580350
rect 282118 580294 282174 580350
rect 282242 580294 282298 580350
rect 282366 580294 282422 580350
rect 281994 580170 282050 580226
rect 282118 580170 282174 580226
rect 282242 580170 282298 580226
rect 282366 580170 282422 580226
rect 281994 580046 282050 580102
rect 282118 580046 282174 580102
rect 282242 580046 282298 580102
rect 282366 580046 282422 580102
rect 281994 579922 282050 579978
rect 282118 579922 282174 579978
rect 282242 579922 282298 579978
rect 282366 579922 282422 579978
rect 281994 562294 282050 562350
rect 282118 562294 282174 562350
rect 282242 562294 282298 562350
rect 282366 562294 282422 562350
rect 281994 562170 282050 562226
rect 282118 562170 282174 562226
rect 282242 562170 282298 562226
rect 282366 562170 282422 562226
rect 281994 562046 282050 562102
rect 282118 562046 282174 562102
rect 282242 562046 282298 562102
rect 282366 562046 282422 562102
rect 281994 561922 282050 561978
rect 282118 561922 282174 561978
rect 282242 561922 282298 561978
rect 282366 561922 282422 561978
rect 281994 544294 282050 544350
rect 282118 544294 282174 544350
rect 282242 544294 282298 544350
rect 282366 544294 282422 544350
rect 281994 544170 282050 544226
rect 282118 544170 282174 544226
rect 282242 544170 282298 544226
rect 282366 544170 282422 544226
rect 281994 544046 282050 544102
rect 282118 544046 282174 544102
rect 282242 544046 282298 544102
rect 282366 544046 282422 544102
rect 281994 543922 282050 543978
rect 282118 543922 282174 543978
rect 282242 543922 282298 543978
rect 282366 543922 282422 543978
rect 281994 526294 282050 526350
rect 282118 526294 282174 526350
rect 282242 526294 282298 526350
rect 282366 526294 282422 526350
rect 281994 526170 282050 526226
rect 282118 526170 282174 526226
rect 282242 526170 282298 526226
rect 282366 526170 282422 526226
rect 281994 526046 282050 526102
rect 282118 526046 282174 526102
rect 282242 526046 282298 526102
rect 282366 526046 282422 526102
rect 281994 525922 282050 525978
rect 282118 525922 282174 525978
rect 282242 525922 282298 525978
rect 282366 525922 282422 525978
rect 281994 508294 282050 508350
rect 282118 508294 282174 508350
rect 282242 508294 282298 508350
rect 282366 508294 282422 508350
rect 281994 508170 282050 508226
rect 282118 508170 282174 508226
rect 282242 508170 282298 508226
rect 282366 508170 282422 508226
rect 281994 508046 282050 508102
rect 282118 508046 282174 508102
rect 282242 508046 282298 508102
rect 282366 508046 282422 508102
rect 281994 507922 282050 507978
rect 282118 507922 282174 507978
rect 282242 507922 282298 507978
rect 282366 507922 282422 507978
rect 281994 490294 282050 490350
rect 282118 490294 282174 490350
rect 282242 490294 282298 490350
rect 282366 490294 282422 490350
rect 281994 490170 282050 490226
rect 282118 490170 282174 490226
rect 282242 490170 282298 490226
rect 282366 490170 282422 490226
rect 281994 490046 282050 490102
rect 282118 490046 282174 490102
rect 282242 490046 282298 490102
rect 282366 490046 282422 490102
rect 281994 489922 282050 489978
rect 282118 489922 282174 489978
rect 282242 489922 282298 489978
rect 282366 489922 282422 489978
rect 281994 472294 282050 472350
rect 282118 472294 282174 472350
rect 282242 472294 282298 472350
rect 282366 472294 282422 472350
rect 281994 472170 282050 472226
rect 282118 472170 282174 472226
rect 282242 472170 282298 472226
rect 282366 472170 282422 472226
rect 281994 472046 282050 472102
rect 282118 472046 282174 472102
rect 282242 472046 282298 472102
rect 282366 472046 282422 472102
rect 281994 471922 282050 471978
rect 282118 471922 282174 471978
rect 282242 471922 282298 471978
rect 282366 471922 282422 471978
rect 281994 454294 282050 454350
rect 282118 454294 282174 454350
rect 282242 454294 282298 454350
rect 282366 454294 282422 454350
rect 281994 454170 282050 454226
rect 282118 454170 282174 454226
rect 282242 454170 282298 454226
rect 282366 454170 282422 454226
rect 281994 454046 282050 454102
rect 282118 454046 282174 454102
rect 282242 454046 282298 454102
rect 282366 454046 282422 454102
rect 281994 453922 282050 453978
rect 282118 453922 282174 453978
rect 282242 453922 282298 453978
rect 282366 453922 282422 453978
rect 281994 436294 282050 436350
rect 282118 436294 282174 436350
rect 282242 436294 282298 436350
rect 282366 436294 282422 436350
rect 281994 436170 282050 436226
rect 282118 436170 282174 436226
rect 282242 436170 282298 436226
rect 282366 436170 282422 436226
rect 281994 436046 282050 436102
rect 282118 436046 282174 436102
rect 282242 436046 282298 436102
rect 282366 436046 282422 436102
rect 281994 435922 282050 435978
rect 282118 435922 282174 435978
rect 282242 435922 282298 435978
rect 282366 435922 282422 435978
rect 281994 418294 282050 418350
rect 282118 418294 282174 418350
rect 282242 418294 282298 418350
rect 282366 418294 282422 418350
rect 281994 418170 282050 418226
rect 282118 418170 282174 418226
rect 282242 418170 282298 418226
rect 282366 418170 282422 418226
rect 281994 418046 282050 418102
rect 282118 418046 282174 418102
rect 282242 418046 282298 418102
rect 282366 418046 282422 418102
rect 281994 417922 282050 417978
rect 282118 417922 282174 417978
rect 282242 417922 282298 417978
rect 282366 417922 282422 417978
rect 281994 400294 282050 400350
rect 282118 400294 282174 400350
rect 282242 400294 282298 400350
rect 282366 400294 282422 400350
rect 281994 400170 282050 400226
rect 282118 400170 282174 400226
rect 282242 400170 282298 400226
rect 282366 400170 282422 400226
rect 281994 400046 282050 400102
rect 282118 400046 282174 400102
rect 282242 400046 282298 400102
rect 282366 400046 282422 400102
rect 281994 399922 282050 399978
rect 282118 399922 282174 399978
rect 282242 399922 282298 399978
rect 282366 399922 282422 399978
rect 281994 382294 282050 382350
rect 282118 382294 282174 382350
rect 282242 382294 282298 382350
rect 282366 382294 282422 382350
rect 281994 382170 282050 382226
rect 282118 382170 282174 382226
rect 282242 382170 282298 382226
rect 282366 382170 282422 382226
rect 281994 382046 282050 382102
rect 282118 382046 282174 382102
rect 282242 382046 282298 382102
rect 282366 382046 282422 382102
rect 281994 381922 282050 381978
rect 282118 381922 282174 381978
rect 282242 381922 282298 381978
rect 282366 381922 282422 381978
rect 281994 364294 282050 364350
rect 282118 364294 282174 364350
rect 282242 364294 282298 364350
rect 282366 364294 282422 364350
rect 281994 364170 282050 364226
rect 282118 364170 282174 364226
rect 282242 364170 282298 364226
rect 282366 364170 282422 364226
rect 281994 364046 282050 364102
rect 282118 364046 282174 364102
rect 282242 364046 282298 364102
rect 282366 364046 282422 364102
rect 281994 363922 282050 363978
rect 282118 363922 282174 363978
rect 282242 363922 282298 363978
rect 282366 363922 282422 363978
rect 281994 346294 282050 346350
rect 282118 346294 282174 346350
rect 282242 346294 282298 346350
rect 282366 346294 282422 346350
rect 281994 346170 282050 346226
rect 282118 346170 282174 346226
rect 282242 346170 282298 346226
rect 282366 346170 282422 346226
rect 281994 346046 282050 346102
rect 282118 346046 282174 346102
rect 282242 346046 282298 346102
rect 282366 346046 282422 346102
rect 281994 345922 282050 345978
rect 282118 345922 282174 345978
rect 282242 345922 282298 345978
rect 282366 345922 282422 345978
rect 281994 328294 282050 328350
rect 282118 328294 282174 328350
rect 282242 328294 282298 328350
rect 282366 328294 282422 328350
rect 281994 328170 282050 328226
rect 282118 328170 282174 328226
rect 282242 328170 282298 328226
rect 282366 328170 282422 328226
rect 281994 328046 282050 328102
rect 282118 328046 282174 328102
rect 282242 328046 282298 328102
rect 282366 328046 282422 328102
rect 281994 327922 282050 327978
rect 282118 327922 282174 327978
rect 282242 327922 282298 327978
rect 282366 327922 282422 327978
rect 285714 598116 285770 598172
rect 285838 598116 285894 598172
rect 285962 598116 286018 598172
rect 286086 598116 286142 598172
rect 285714 597992 285770 598048
rect 285838 597992 285894 598048
rect 285962 597992 286018 598048
rect 286086 597992 286142 598048
rect 285714 597868 285770 597924
rect 285838 597868 285894 597924
rect 285962 597868 286018 597924
rect 286086 597868 286142 597924
rect 285714 597744 285770 597800
rect 285838 597744 285894 597800
rect 285962 597744 286018 597800
rect 286086 597744 286142 597800
rect 285714 586294 285770 586350
rect 285838 586294 285894 586350
rect 285962 586294 286018 586350
rect 286086 586294 286142 586350
rect 285714 586170 285770 586226
rect 285838 586170 285894 586226
rect 285962 586170 286018 586226
rect 286086 586170 286142 586226
rect 285714 586046 285770 586102
rect 285838 586046 285894 586102
rect 285962 586046 286018 586102
rect 286086 586046 286142 586102
rect 285714 585922 285770 585978
rect 285838 585922 285894 585978
rect 285962 585922 286018 585978
rect 286086 585922 286142 585978
rect 285714 568294 285770 568350
rect 285838 568294 285894 568350
rect 285962 568294 286018 568350
rect 286086 568294 286142 568350
rect 285714 568170 285770 568226
rect 285838 568170 285894 568226
rect 285962 568170 286018 568226
rect 286086 568170 286142 568226
rect 285714 568046 285770 568102
rect 285838 568046 285894 568102
rect 285962 568046 286018 568102
rect 286086 568046 286142 568102
rect 285714 567922 285770 567978
rect 285838 567922 285894 567978
rect 285962 567922 286018 567978
rect 286086 567922 286142 567978
rect 285714 550294 285770 550350
rect 285838 550294 285894 550350
rect 285962 550294 286018 550350
rect 286086 550294 286142 550350
rect 285714 550170 285770 550226
rect 285838 550170 285894 550226
rect 285962 550170 286018 550226
rect 286086 550170 286142 550226
rect 285714 550046 285770 550102
rect 285838 550046 285894 550102
rect 285962 550046 286018 550102
rect 286086 550046 286142 550102
rect 285714 549922 285770 549978
rect 285838 549922 285894 549978
rect 285962 549922 286018 549978
rect 286086 549922 286142 549978
rect 285714 532294 285770 532350
rect 285838 532294 285894 532350
rect 285962 532294 286018 532350
rect 286086 532294 286142 532350
rect 285714 532170 285770 532226
rect 285838 532170 285894 532226
rect 285962 532170 286018 532226
rect 286086 532170 286142 532226
rect 285714 532046 285770 532102
rect 285838 532046 285894 532102
rect 285962 532046 286018 532102
rect 286086 532046 286142 532102
rect 285714 531922 285770 531978
rect 285838 531922 285894 531978
rect 285962 531922 286018 531978
rect 286086 531922 286142 531978
rect 285714 514294 285770 514350
rect 285838 514294 285894 514350
rect 285962 514294 286018 514350
rect 286086 514294 286142 514350
rect 285714 514170 285770 514226
rect 285838 514170 285894 514226
rect 285962 514170 286018 514226
rect 286086 514170 286142 514226
rect 285714 514046 285770 514102
rect 285838 514046 285894 514102
rect 285962 514046 286018 514102
rect 286086 514046 286142 514102
rect 285714 513922 285770 513978
rect 285838 513922 285894 513978
rect 285962 513922 286018 513978
rect 286086 513922 286142 513978
rect 285714 496294 285770 496350
rect 285838 496294 285894 496350
rect 285962 496294 286018 496350
rect 286086 496294 286142 496350
rect 285714 496170 285770 496226
rect 285838 496170 285894 496226
rect 285962 496170 286018 496226
rect 286086 496170 286142 496226
rect 285714 496046 285770 496102
rect 285838 496046 285894 496102
rect 285962 496046 286018 496102
rect 286086 496046 286142 496102
rect 285714 495922 285770 495978
rect 285838 495922 285894 495978
rect 285962 495922 286018 495978
rect 286086 495922 286142 495978
rect 285714 478294 285770 478350
rect 285838 478294 285894 478350
rect 285962 478294 286018 478350
rect 286086 478294 286142 478350
rect 285714 478170 285770 478226
rect 285838 478170 285894 478226
rect 285962 478170 286018 478226
rect 286086 478170 286142 478226
rect 285714 478046 285770 478102
rect 285838 478046 285894 478102
rect 285962 478046 286018 478102
rect 286086 478046 286142 478102
rect 285714 477922 285770 477978
rect 285838 477922 285894 477978
rect 285962 477922 286018 477978
rect 286086 477922 286142 477978
rect 285714 460294 285770 460350
rect 285838 460294 285894 460350
rect 285962 460294 286018 460350
rect 286086 460294 286142 460350
rect 285714 460170 285770 460226
rect 285838 460170 285894 460226
rect 285962 460170 286018 460226
rect 286086 460170 286142 460226
rect 285714 460046 285770 460102
rect 285838 460046 285894 460102
rect 285962 460046 286018 460102
rect 286086 460046 286142 460102
rect 285714 459922 285770 459978
rect 285838 459922 285894 459978
rect 285962 459922 286018 459978
rect 286086 459922 286142 459978
rect 285714 442294 285770 442350
rect 285838 442294 285894 442350
rect 285962 442294 286018 442350
rect 286086 442294 286142 442350
rect 285714 442170 285770 442226
rect 285838 442170 285894 442226
rect 285962 442170 286018 442226
rect 286086 442170 286142 442226
rect 285714 442046 285770 442102
rect 285838 442046 285894 442102
rect 285962 442046 286018 442102
rect 286086 442046 286142 442102
rect 285714 441922 285770 441978
rect 285838 441922 285894 441978
rect 285962 441922 286018 441978
rect 286086 441922 286142 441978
rect 285714 424294 285770 424350
rect 285838 424294 285894 424350
rect 285962 424294 286018 424350
rect 286086 424294 286142 424350
rect 285714 424170 285770 424226
rect 285838 424170 285894 424226
rect 285962 424170 286018 424226
rect 286086 424170 286142 424226
rect 285714 424046 285770 424102
rect 285838 424046 285894 424102
rect 285962 424046 286018 424102
rect 286086 424046 286142 424102
rect 285714 423922 285770 423978
rect 285838 423922 285894 423978
rect 285962 423922 286018 423978
rect 286086 423922 286142 423978
rect 285714 406294 285770 406350
rect 285838 406294 285894 406350
rect 285962 406294 286018 406350
rect 286086 406294 286142 406350
rect 285714 406170 285770 406226
rect 285838 406170 285894 406226
rect 285962 406170 286018 406226
rect 286086 406170 286142 406226
rect 285714 406046 285770 406102
rect 285838 406046 285894 406102
rect 285962 406046 286018 406102
rect 286086 406046 286142 406102
rect 285714 405922 285770 405978
rect 285838 405922 285894 405978
rect 285962 405922 286018 405978
rect 286086 405922 286142 405978
rect 285714 388294 285770 388350
rect 285838 388294 285894 388350
rect 285962 388294 286018 388350
rect 286086 388294 286142 388350
rect 285714 388170 285770 388226
rect 285838 388170 285894 388226
rect 285962 388170 286018 388226
rect 286086 388170 286142 388226
rect 285714 388046 285770 388102
rect 285838 388046 285894 388102
rect 285962 388046 286018 388102
rect 286086 388046 286142 388102
rect 285714 387922 285770 387978
rect 285838 387922 285894 387978
rect 285962 387922 286018 387978
rect 286086 387922 286142 387978
rect 285714 370294 285770 370350
rect 285838 370294 285894 370350
rect 285962 370294 286018 370350
rect 286086 370294 286142 370350
rect 285714 370170 285770 370226
rect 285838 370170 285894 370226
rect 285962 370170 286018 370226
rect 286086 370170 286142 370226
rect 285714 370046 285770 370102
rect 285838 370046 285894 370102
rect 285962 370046 286018 370102
rect 286086 370046 286142 370102
rect 285714 369922 285770 369978
rect 285838 369922 285894 369978
rect 285962 369922 286018 369978
rect 286086 369922 286142 369978
rect 285714 352294 285770 352350
rect 285838 352294 285894 352350
rect 285962 352294 286018 352350
rect 286086 352294 286142 352350
rect 285714 352170 285770 352226
rect 285838 352170 285894 352226
rect 285962 352170 286018 352226
rect 286086 352170 286142 352226
rect 285714 352046 285770 352102
rect 285838 352046 285894 352102
rect 285962 352046 286018 352102
rect 286086 352046 286142 352102
rect 285714 351922 285770 351978
rect 285838 351922 285894 351978
rect 285962 351922 286018 351978
rect 286086 351922 286142 351978
rect 285714 334294 285770 334350
rect 285838 334294 285894 334350
rect 285962 334294 286018 334350
rect 286086 334294 286142 334350
rect 285714 334170 285770 334226
rect 285838 334170 285894 334226
rect 285962 334170 286018 334226
rect 286086 334170 286142 334226
rect 285714 334046 285770 334102
rect 285838 334046 285894 334102
rect 285962 334046 286018 334102
rect 286086 334046 286142 334102
rect 285714 333922 285770 333978
rect 285838 333922 285894 333978
rect 285962 333922 286018 333978
rect 286086 333922 286142 333978
rect 312714 597156 312770 597212
rect 312838 597156 312894 597212
rect 312962 597156 313018 597212
rect 313086 597156 313142 597212
rect 312714 597032 312770 597088
rect 312838 597032 312894 597088
rect 312962 597032 313018 597088
rect 313086 597032 313142 597088
rect 312714 596908 312770 596964
rect 312838 596908 312894 596964
rect 312962 596908 313018 596964
rect 313086 596908 313142 596964
rect 312714 596784 312770 596840
rect 312838 596784 312894 596840
rect 312962 596784 313018 596840
rect 313086 596784 313142 596840
rect 312714 580294 312770 580350
rect 312838 580294 312894 580350
rect 312962 580294 313018 580350
rect 313086 580294 313142 580350
rect 312714 580170 312770 580226
rect 312838 580170 312894 580226
rect 312962 580170 313018 580226
rect 313086 580170 313142 580226
rect 312714 580046 312770 580102
rect 312838 580046 312894 580102
rect 312962 580046 313018 580102
rect 313086 580046 313142 580102
rect 312714 579922 312770 579978
rect 312838 579922 312894 579978
rect 312962 579922 313018 579978
rect 313086 579922 313142 579978
rect 312714 562294 312770 562350
rect 312838 562294 312894 562350
rect 312962 562294 313018 562350
rect 313086 562294 313142 562350
rect 312714 562170 312770 562226
rect 312838 562170 312894 562226
rect 312962 562170 313018 562226
rect 313086 562170 313142 562226
rect 312714 562046 312770 562102
rect 312838 562046 312894 562102
rect 312962 562046 313018 562102
rect 313086 562046 313142 562102
rect 312714 561922 312770 561978
rect 312838 561922 312894 561978
rect 312962 561922 313018 561978
rect 313086 561922 313142 561978
rect 312714 544294 312770 544350
rect 312838 544294 312894 544350
rect 312962 544294 313018 544350
rect 313086 544294 313142 544350
rect 312714 544170 312770 544226
rect 312838 544170 312894 544226
rect 312962 544170 313018 544226
rect 313086 544170 313142 544226
rect 312714 544046 312770 544102
rect 312838 544046 312894 544102
rect 312962 544046 313018 544102
rect 313086 544046 313142 544102
rect 312714 543922 312770 543978
rect 312838 543922 312894 543978
rect 312962 543922 313018 543978
rect 313086 543922 313142 543978
rect 312714 526294 312770 526350
rect 312838 526294 312894 526350
rect 312962 526294 313018 526350
rect 313086 526294 313142 526350
rect 312714 526170 312770 526226
rect 312838 526170 312894 526226
rect 312962 526170 313018 526226
rect 313086 526170 313142 526226
rect 312714 526046 312770 526102
rect 312838 526046 312894 526102
rect 312962 526046 313018 526102
rect 313086 526046 313142 526102
rect 312714 525922 312770 525978
rect 312838 525922 312894 525978
rect 312962 525922 313018 525978
rect 313086 525922 313142 525978
rect 312714 508294 312770 508350
rect 312838 508294 312894 508350
rect 312962 508294 313018 508350
rect 313086 508294 313142 508350
rect 312714 508170 312770 508226
rect 312838 508170 312894 508226
rect 312962 508170 313018 508226
rect 313086 508170 313142 508226
rect 312714 508046 312770 508102
rect 312838 508046 312894 508102
rect 312962 508046 313018 508102
rect 313086 508046 313142 508102
rect 312714 507922 312770 507978
rect 312838 507922 312894 507978
rect 312962 507922 313018 507978
rect 313086 507922 313142 507978
rect 312714 490294 312770 490350
rect 312838 490294 312894 490350
rect 312962 490294 313018 490350
rect 313086 490294 313142 490350
rect 312714 490170 312770 490226
rect 312838 490170 312894 490226
rect 312962 490170 313018 490226
rect 313086 490170 313142 490226
rect 312714 490046 312770 490102
rect 312838 490046 312894 490102
rect 312962 490046 313018 490102
rect 313086 490046 313142 490102
rect 312714 489922 312770 489978
rect 312838 489922 312894 489978
rect 312962 489922 313018 489978
rect 313086 489922 313142 489978
rect 312714 472294 312770 472350
rect 312838 472294 312894 472350
rect 312962 472294 313018 472350
rect 313086 472294 313142 472350
rect 312714 472170 312770 472226
rect 312838 472170 312894 472226
rect 312962 472170 313018 472226
rect 313086 472170 313142 472226
rect 312714 472046 312770 472102
rect 312838 472046 312894 472102
rect 312962 472046 313018 472102
rect 313086 472046 313142 472102
rect 312714 471922 312770 471978
rect 312838 471922 312894 471978
rect 312962 471922 313018 471978
rect 313086 471922 313142 471978
rect 312714 454294 312770 454350
rect 312838 454294 312894 454350
rect 312962 454294 313018 454350
rect 313086 454294 313142 454350
rect 312714 454170 312770 454226
rect 312838 454170 312894 454226
rect 312962 454170 313018 454226
rect 313086 454170 313142 454226
rect 312714 454046 312770 454102
rect 312838 454046 312894 454102
rect 312962 454046 313018 454102
rect 313086 454046 313142 454102
rect 312714 453922 312770 453978
rect 312838 453922 312894 453978
rect 312962 453922 313018 453978
rect 313086 453922 313142 453978
rect 312714 436294 312770 436350
rect 312838 436294 312894 436350
rect 312962 436294 313018 436350
rect 313086 436294 313142 436350
rect 312714 436170 312770 436226
rect 312838 436170 312894 436226
rect 312962 436170 313018 436226
rect 313086 436170 313142 436226
rect 312714 436046 312770 436102
rect 312838 436046 312894 436102
rect 312962 436046 313018 436102
rect 313086 436046 313142 436102
rect 312714 435922 312770 435978
rect 312838 435922 312894 435978
rect 312962 435922 313018 435978
rect 313086 435922 313142 435978
rect 312714 418294 312770 418350
rect 312838 418294 312894 418350
rect 312962 418294 313018 418350
rect 313086 418294 313142 418350
rect 312714 418170 312770 418226
rect 312838 418170 312894 418226
rect 312962 418170 313018 418226
rect 313086 418170 313142 418226
rect 312714 418046 312770 418102
rect 312838 418046 312894 418102
rect 312962 418046 313018 418102
rect 313086 418046 313142 418102
rect 312714 417922 312770 417978
rect 312838 417922 312894 417978
rect 312962 417922 313018 417978
rect 313086 417922 313142 417978
rect 312714 400294 312770 400350
rect 312838 400294 312894 400350
rect 312962 400294 313018 400350
rect 313086 400294 313142 400350
rect 312714 400170 312770 400226
rect 312838 400170 312894 400226
rect 312962 400170 313018 400226
rect 313086 400170 313142 400226
rect 312714 400046 312770 400102
rect 312838 400046 312894 400102
rect 312962 400046 313018 400102
rect 313086 400046 313142 400102
rect 312714 399922 312770 399978
rect 312838 399922 312894 399978
rect 312962 399922 313018 399978
rect 313086 399922 313142 399978
rect 312714 382294 312770 382350
rect 312838 382294 312894 382350
rect 312962 382294 313018 382350
rect 313086 382294 313142 382350
rect 312714 382170 312770 382226
rect 312838 382170 312894 382226
rect 312962 382170 313018 382226
rect 313086 382170 313142 382226
rect 312714 382046 312770 382102
rect 312838 382046 312894 382102
rect 312962 382046 313018 382102
rect 313086 382046 313142 382102
rect 312714 381922 312770 381978
rect 312838 381922 312894 381978
rect 312962 381922 313018 381978
rect 313086 381922 313142 381978
rect 312714 364294 312770 364350
rect 312838 364294 312894 364350
rect 312962 364294 313018 364350
rect 313086 364294 313142 364350
rect 312714 364170 312770 364226
rect 312838 364170 312894 364226
rect 312962 364170 313018 364226
rect 313086 364170 313142 364226
rect 312714 364046 312770 364102
rect 312838 364046 312894 364102
rect 312962 364046 313018 364102
rect 313086 364046 313142 364102
rect 312714 363922 312770 363978
rect 312838 363922 312894 363978
rect 312962 363922 313018 363978
rect 313086 363922 313142 363978
rect 312714 346294 312770 346350
rect 312838 346294 312894 346350
rect 312962 346294 313018 346350
rect 313086 346294 313142 346350
rect 312714 346170 312770 346226
rect 312838 346170 312894 346226
rect 312962 346170 313018 346226
rect 313086 346170 313142 346226
rect 312714 346046 312770 346102
rect 312838 346046 312894 346102
rect 312962 346046 313018 346102
rect 313086 346046 313142 346102
rect 312714 345922 312770 345978
rect 312838 345922 312894 345978
rect 312962 345922 313018 345978
rect 313086 345922 313142 345978
rect 312714 328294 312770 328350
rect 312838 328294 312894 328350
rect 312962 328294 313018 328350
rect 313086 328294 313142 328350
rect 312714 328170 312770 328226
rect 312838 328170 312894 328226
rect 312962 328170 313018 328226
rect 313086 328170 313142 328226
rect 312714 328046 312770 328102
rect 312838 328046 312894 328102
rect 312962 328046 313018 328102
rect 313086 328046 313142 328102
rect 312714 327922 312770 327978
rect 312838 327922 312894 327978
rect 312962 327922 313018 327978
rect 313086 327922 313142 327978
rect 316434 598116 316490 598172
rect 316558 598116 316614 598172
rect 316682 598116 316738 598172
rect 316806 598116 316862 598172
rect 316434 597992 316490 598048
rect 316558 597992 316614 598048
rect 316682 597992 316738 598048
rect 316806 597992 316862 598048
rect 316434 597868 316490 597924
rect 316558 597868 316614 597924
rect 316682 597868 316738 597924
rect 316806 597868 316862 597924
rect 316434 597744 316490 597800
rect 316558 597744 316614 597800
rect 316682 597744 316738 597800
rect 316806 597744 316862 597800
rect 316434 586294 316490 586350
rect 316558 586294 316614 586350
rect 316682 586294 316738 586350
rect 316806 586294 316862 586350
rect 316434 586170 316490 586226
rect 316558 586170 316614 586226
rect 316682 586170 316738 586226
rect 316806 586170 316862 586226
rect 316434 586046 316490 586102
rect 316558 586046 316614 586102
rect 316682 586046 316738 586102
rect 316806 586046 316862 586102
rect 316434 585922 316490 585978
rect 316558 585922 316614 585978
rect 316682 585922 316738 585978
rect 316806 585922 316862 585978
rect 316434 568294 316490 568350
rect 316558 568294 316614 568350
rect 316682 568294 316738 568350
rect 316806 568294 316862 568350
rect 316434 568170 316490 568226
rect 316558 568170 316614 568226
rect 316682 568170 316738 568226
rect 316806 568170 316862 568226
rect 316434 568046 316490 568102
rect 316558 568046 316614 568102
rect 316682 568046 316738 568102
rect 316806 568046 316862 568102
rect 316434 567922 316490 567978
rect 316558 567922 316614 567978
rect 316682 567922 316738 567978
rect 316806 567922 316862 567978
rect 316434 550294 316490 550350
rect 316558 550294 316614 550350
rect 316682 550294 316738 550350
rect 316806 550294 316862 550350
rect 316434 550170 316490 550226
rect 316558 550170 316614 550226
rect 316682 550170 316738 550226
rect 316806 550170 316862 550226
rect 316434 550046 316490 550102
rect 316558 550046 316614 550102
rect 316682 550046 316738 550102
rect 316806 550046 316862 550102
rect 316434 549922 316490 549978
rect 316558 549922 316614 549978
rect 316682 549922 316738 549978
rect 316806 549922 316862 549978
rect 316434 532294 316490 532350
rect 316558 532294 316614 532350
rect 316682 532294 316738 532350
rect 316806 532294 316862 532350
rect 316434 532170 316490 532226
rect 316558 532170 316614 532226
rect 316682 532170 316738 532226
rect 316806 532170 316862 532226
rect 316434 532046 316490 532102
rect 316558 532046 316614 532102
rect 316682 532046 316738 532102
rect 316806 532046 316862 532102
rect 316434 531922 316490 531978
rect 316558 531922 316614 531978
rect 316682 531922 316738 531978
rect 316806 531922 316862 531978
rect 316434 514294 316490 514350
rect 316558 514294 316614 514350
rect 316682 514294 316738 514350
rect 316806 514294 316862 514350
rect 316434 514170 316490 514226
rect 316558 514170 316614 514226
rect 316682 514170 316738 514226
rect 316806 514170 316862 514226
rect 316434 514046 316490 514102
rect 316558 514046 316614 514102
rect 316682 514046 316738 514102
rect 316806 514046 316862 514102
rect 316434 513922 316490 513978
rect 316558 513922 316614 513978
rect 316682 513922 316738 513978
rect 316806 513922 316862 513978
rect 316434 496294 316490 496350
rect 316558 496294 316614 496350
rect 316682 496294 316738 496350
rect 316806 496294 316862 496350
rect 316434 496170 316490 496226
rect 316558 496170 316614 496226
rect 316682 496170 316738 496226
rect 316806 496170 316862 496226
rect 316434 496046 316490 496102
rect 316558 496046 316614 496102
rect 316682 496046 316738 496102
rect 316806 496046 316862 496102
rect 316434 495922 316490 495978
rect 316558 495922 316614 495978
rect 316682 495922 316738 495978
rect 316806 495922 316862 495978
rect 316434 478294 316490 478350
rect 316558 478294 316614 478350
rect 316682 478294 316738 478350
rect 316806 478294 316862 478350
rect 316434 478170 316490 478226
rect 316558 478170 316614 478226
rect 316682 478170 316738 478226
rect 316806 478170 316862 478226
rect 316434 478046 316490 478102
rect 316558 478046 316614 478102
rect 316682 478046 316738 478102
rect 316806 478046 316862 478102
rect 316434 477922 316490 477978
rect 316558 477922 316614 477978
rect 316682 477922 316738 477978
rect 316806 477922 316862 477978
rect 316434 460294 316490 460350
rect 316558 460294 316614 460350
rect 316682 460294 316738 460350
rect 316806 460294 316862 460350
rect 316434 460170 316490 460226
rect 316558 460170 316614 460226
rect 316682 460170 316738 460226
rect 316806 460170 316862 460226
rect 316434 460046 316490 460102
rect 316558 460046 316614 460102
rect 316682 460046 316738 460102
rect 316806 460046 316862 460102
rect 316434 459922 316490 459978
rect 316558 459922 316614 459978
rect 316682 459922 316738 459978
rect 316806 459922 316862 459978
rect 316434 442294 316490 442350
rect 316558 442294 316614 442350
rect 316682 442294 316738 442350
rect 316806 442294 316862 442350
rect 316434 442170 316490 442226
rect 316558 442170 316614 442226
rect 316682 442170 316738 442226
rect 316806 442170 316862 442226
rect 316434 442046 316490 442102
rect 316558 442046 316614 442102
rect 316682 442046 316738 442102
rect 316806 442046 316862 442102
rect 316434 441922 316490 441978
rect 316558 441922 316614 441978
rect 316682 441922 316738 441978
rect 316806 441922 316862 441978
rect 316434 424294 316490 424350
rect 316558 424294 316614 424350
rect 316682 424294 316738 424350
rect 316806 424294 316862 424350
rect 316434 424170 316490 424226
rect 316558 424170 316614 424226
rect 316682 424170 316738 424226
rect 316806 424170 316862 424226
rect 316434 424046 316490 424102
rect 316558 424046 316614 424102
rect 316682 424046 316738 424102
rect 316806 424046 316862 424102
rect 316434 423922 316490 423978
rect 316558 423922 316614 423978
rect 316682 423922 316738 423978
rect 316806 423922 316862 423978
rect 316434 406294 316490 406350
rect 316558 406294 316614 406350
rect 316682 406294 316738 406350
rect 316806 406294 316862 406350
rect 316434 406170 316490 406226
rect 316558 406170 316614 406226
rect 316682 406170 316738 406226
rect 316806 406170 316862 406226
rect 316434 406046 316490 406102
rect 316558 406046 316614 406102
rect 316682 406046 316738 406102
rect 316806 406046 316862 406102
rect 316434 405922 316490 405978
rect 316558 405922 316614 405978
rect 316682 405922 316738 405978
rect 316806 405922 316862 405978
rect 316434 388294 316490 388350
rect 316558 388294 316614 388350
rect 316682 388294 316738 388350
rect 316806 388294 316862 388350
rect 316434 388170 316490 388226
rect 316558 388170 316614 388226
rect 316682 388170 316738 388226
rect 316806 388170 316862 388226
rect 316434 388046 316490 388102
rect 316558 388046 316614 388102
rect 316682 388046 316738 388102
rect 316806 388046 316862 388102
rect 316434 387922 316490 387978
rect 316558 387922 316614 387978
rect 316682 387922 316738 387978
rect 316806 387922 316862 387978
rect 316434 370294 316490 370350
rect 316558 370294 316614 370350
rect 316682 370294 316738 370350
rect 316806 370294 316862 370350
rect 316434 370170 316490 370226
rect 316558 370170 316614 370226
rect 316682 370170 316738 370226
rect 316806 370170 316862 370226
rect 316434 370046 316490 370102
rect 316558 370046 316614 370102
rect 316682 370046 316738 370102
rect 316806 370046 316862 370102
rect 316434 369922 316490 369978
rect 316558 369922 316614 369978
rect 316682 369922 316738 369978
rect 316806 369922 316862 369978
rect 316434 352294 316490 352350
rect 316558 352294 316614 352350
rect 316682 352294 316738 352350
rect 316806 352294 316862 352350
rect 316434 352170 316490 352226
rect 316558 352170 316614 352226
rect 316682 352170 316738 352226
rect 316806 352170 316862 352226
rect 316434 352046 316490 352102
rect 316558 352046 316614 352102
rect 316682 352046 316738 352102
rect 316806 352046 316862 352102
rect 316434 351922 316490 351978
rect 316558 351922 316614 351978
rect 316682 351922 316738 351978
rect 316806 351922 316862 351978
rect 316434 334294 316490 334350
rect 316558 334294 316614 334350
rect 316682 334294 316738 334350
rect 316806 334294 316862 334350
rect 316434 334170 316490 334226
rect 316558 334170 316614 334226
rect 316682 334170 316738 334226
rect 316806 334170 316862 334226
rect 316434 334046 316490 334102
rect 316558 334046 316614 334102
rect 316682 334046 316738 334102
rect 316806 334046 316862 334102
rect 316434 333922 316490 333978
rect 316558 333922 316614 333978
rect 316682 333922 316738 333978
rect 316806 333922 316862 333978
rect 343434 597156 343490 597212
rect 343558 597156 343614 597212
rect 343682 597156 343738 597212
rect 343806 597156 343862 597212
rect 343434 597032 343490 597088
rect 343558 597032 343614 597088
rect 343682 597032 343738 597088
rect 343806 597032 343862 597088
rect 343434 596908 343490 596964
rect 343558 596908 343614 596964
rect 343682 596908 343738 596964
rect 343806 596908 343862 596964
rect 343434 596784 343490 596840
rect 343558 596784 343614 596840
rect 343682 596784 343738 596840
rect 343806 596784 343862 596840
rect 343434 580294 343490 580350
rect 343558 580294 343614 580350
rect 343682 580294 343738 580350
rect 343806 580294 343862 580350
rect 343434 580170 343490 580226
rect 343558 580170 343614 580226
rect 343682 580170 343738 580226
rect 343806 580170 343862 580226
rect 343434 580046 343490 580102
rect 343558 580046 343614 580102
rect 343682 580046 343738 580102
rect 343806 580046 343862 580102
rect 343434 579922 343490 579978
rect 343558 579922 343614 579978
rect 343682 579922 343738 579978
rect 343806 579922 343862 579978
rect 343434 562294 343490 562350
rect 343558 562294 343614 562350
rect 343682 562294 343738 562350
rect 343806 562294 343862 562350
rect 343434 562170 343490 562226
rect 343558 562170 343614 562226
rect 343682 562170 343738 562226
rect 343806 562170 343862 562226
rect 343434 562046 343490 562102
rect 343558 562046 343614 562102
rect 343682 562046 343738 562102
rect 343806 562046 343862 562102
rect 343434 561922 343490 561978
rect 343558 561922 343614 561978
rect 343682 561922 343738 561978
rect 343806 561922 343862 561978
rect 343434 544294 343490 544350
rect 343558 544294 343614 544350
rect 343682 544294 343738 544350
rect 343806 544294 343862 544350
rect 343434 544170 343490 544226
rect 343558 544170 343614 544226
rect 343682 544170 343738 544226
rect 343806 544170 343862 544226
rect 343434 544046 343490 544102
rect 343558 544046 343614 544102
rect 343682 544046 343738 544102
rect 343806 544046 343862 544102
rect 343434 543922 343490 543978
rect 343558 543922 343614 543978
rect 343682 543922 343738 543978
rect 343806 543922 343862 543978
rect 343434 526294 343490 526350
rect 343558 526294 343614 526350
rect 343682 526294 343738 526350
rect 343806 526294 343862 526350
rect 343434 526170 343490 526226
rect 343558 526170 343614 526226
rect 343682 526170 343738 526226
rect 343806 526170 343862 526226
rect 343434 526046 343490 526102
rect 343558 526046 343614 526102
rect 343682 526046 343738 526102
rect 343806 526046 343862 526102
rect 343434 525922 343490 525978
rect 343558 525922 343614 525978
rect 343682 525922 343738 525978
rect 343806 525922 343862 525978
rect 343434 508294 343490 508350
rect 343558 508294 343614 508350
rect 343682 508294 343738 508350
rect 343806 508294 343862 508350
rect 343434 508170 343490 508226
rect 343558 508170 343614 508226
rect 343682 508170 343738 508226
rect 343806 508170 343862 508226
rect 343434 508046 343490 508102
rect 343558 508046 343614 508102
rect 343682 508046 343738 508102
rect 343806 508046 343862 508102
rect 343434 507922 343490 507978
rect 343558 507922 343614 507978
rect 343682 507922 343738 507978
rect 343806 507922 343862 507978
rect 343434 490294 343490 490350
rect 343558 490294 343614 490350
rect 343682 490294 343738 490350
rect 343806 490294 343862 490350
rect 343434 490170 343490 490226
rect 343558 490170 343614 490226
rect 343682 490170 343738 490226
rect 343806 490170 343862 490226
rect 343434 490046 343490 490102
rect 343558 490046 343614 490102
rect 343682 490046 343738 490102
rect 343806 490046 343862 490102
rect 343434 489922 343490 489978
rect 343558 489922 343614 489978
rect 343682 489922 343738 489978
rect 343806 489922 343862 489978
rect 343434 472294 343490 472350
rect 343558 472294 343614 472350
rect 343682 472294 343738 472350
rect 343806 472294 343862 472350
rect 343434 472170 343490 472226
rect 343558 472170 343614 472226
rect 343682 472170 343738 472226
rect 343806 472170 343862 472226
rect 343434 472046 343490 472102
rect 343558 472046 343614 472102
rect 343682 472046 343738 472102
rect 343806 472046 343862 472102
rect 343434 471922 343490 471978
rect 343558 471922 343614 471978
rect 343682 471922 343738 471978
rect 343806 471922 343862 471978
rect 343434 454294 343490 454350
rect 343558 454294 343614 454350
rect 343682 454294 343738 454350
rect 343806 454294 343862 454350
rect 343434 454170 343490 454226
rect 343558 454170 343614 454226
rect 343682 454170 343738 454226
rect 343806 454170 343862 454226
rect 343434 454046 343490 454102
rect 343558 454046 343614 454102
rect 343682 454046 343738 454102
rect 343806 454046 343862 454102
rect 343434 453922 343490 453978
rect 343558 453922 343614 453978
rect 343682 453922 343738 453978
rect 343806 453922 343862 453978
rect 343434 436294 343490 436350
rect 343558 436294 343614 436350
rect 343682 436294 343738 436350
rect 343806 436294 343862 436350
rect 343434 436170 343490 436226
rect 343558 436170 343614 436226
rect 343682 436170 343738 436226
rect 343806 436170 343862 436226
rect 343434 436046 343490 436102
rect 343558 436046 343614 436102
rect 343682 436046 343738 436102
rect 343806 436046 343862 436102
rect 343434 435922 343490 435978
rect 343558 435922 343614 435978
rect 343682 435922 343738 435978
rect 343806 435922 343862 435978
rect 343434 418294 343490 418350
rect 343558 418294 343614 418350
rect 343682 418294 343738 418350
rect 343806 418294 343862 418350
rect 343434 418170 343490 418226
rect 343558 418170 343614 418226
rect 343682 418170 343738 418226
rect 343806 418170 343862 418226
rect 343434 418046 343490 418102
rect 343558 418046 343614 418102
rect 343682 418046 343738 418102
rect 343806 418046 343862 418102
rect 343434 417922 343490 417978
rect 343558 417922 343614 417978
rect 343682 417922 343738 417978
rect 343806 417922 343862 417978
rect 343434 400294 343490 400350
rect 343558 400294 343614 400350
rect 343682 400294 343738 400350
rect 343806 400294 343862 400350
rect 343434 400170 343490 400226
rect 343558 400170 343614 400226
rect 343682 400170 343738 400226
rect 343806 400170 343862 400226
rect 343434 400046 343490 400102
rect 343558 400046 343614 400102
rect 343682 400046 343738 400102
rect 343806 400046 343862 400102
rect 343434 399922 343490 399978
rect 343558 399922 343614 399978
rect 343682 399922 343738 399978
rect 343806 399922 343862 399978
rect 343434 382294 343490 382350
rect 343558 382294 343614 382350
rect 343682 382294 343738 382350
rect 343806 382294 343862 382350
rect 343434 382170 343490 382226
rect 343558 382170 343614 382226
rect 343682 382170 343738 382226
rect 343806 382170 343862 382226
rect 343434 382046 343490 382102
rect 343558 382046 343614 382102
rect 343682 382046 343738 382102
rect 343806 382046 343862 382102
rect 343434 381922 343490 381978
rect 343558 381922 343614 381978
rect 343682 381922 343738 381978
rect 343806 381922 343862 381978
rect 343434 364294 343490 364350
rect 343558 364294 343614 364350
rect 343682 364294 343738 364350
rect 343806 364294 343862 364350
rect 343434 364170 343490 364226
rect 343558 364170 343614 364226
rect 343682 364170 343738 364226
rect 343806 364170 343862 364226
rect 343434 364046 343490 364102
rect 343558 364046 343614 364102
rect 343682 364046 343738 364102
rect 343806 364046 343862 364102
rect 343434 363922 343490 363978
rect 343558 363922 343614 363978
rect 343682 363922 343738 363978
rect 343806 363922 343862 363978
rect 343434 346294 343490 346350
rect 343558 346294 343614 346350
rect 343682 346294 343738 346350
rect 343806 346294 343862 346350
rect 343434 346170 343490 346226
rect 343558 346170 343614 346226
rect 343682 346170 343738 346226
rect 343806 346170 343862 346226
rect 343434 346046 343490 346102
rect 343558 346046 343614 346102
rect 343682 346046 343738 346102
rect 343806 346046 343862 346102
rect 343434 345922 343490 345978
rect 343558 345922 343614 345978
rect 343682 345922 343738 345978
rect 343806 345922 343862 345978
rect 343434 328294 343490 328350
rect 343558 328294 343614 328350
rect 343682 328294 343738 328350
rect 343806 328294 343862 328350
rect 343434 328170 343490 328226
rect 343558 328170 343614 328226
rect 343682 328170 343738 328226
rect 343806 328170 343862 328226
rect 343434 328046 343490 328102
rect 343558 328046 343614 328102
rect 343682 328046 343738 328102
rect 343806 328046 343862 328102
rect 343434 327922 343490 327978
rect 343558 327922 343614 327978
rect 343682 327922 343738 327978
rect 343806 327922 343862 327978
rect 347154 598116 347210 598172
rect 347278 598116 347334 598172
rect 347402 598116 347458 598172
rect 347526 598116 347582 598172
rect 347154 597992 347210 598048
rect 347278 597992 347334 598048
rect 347402 597992 347458 598048
rect 347526 597992 347582 598048
rect 347154 597868 347210 597924
rect 347278 597868 347334 597924
rect 347402 597868 347458 597924
rect 347526 597868 347582 597924
rect 347154 597744 347210 597800
rect 347278 597744 347334 597800
rect 347402 597744 347458 597800
rect 347526 597744 347582 597800
rect 347154 586294 347210 586350
rect 347278 586294 347334 586350
rect 347402 586294 347458 586350
rect 347526 586294 347582 586350
rect 347154 586170 347210 586226
rect 347278 586170 347334 586226
rect 347402 586170 347458 586226
rect 347526 586170 347582 586226
rect 347154 586046 347210 586102
rect 347278 586046 347334 586102
rect 347402 586046 347458 586102
rect 347526 586046 347582 586102
rect 347154 585922 347210 585978
rect 347278 585922 347334 585978
rect 347402 585922 347458 585978
rect 347526 585922 347582 585978
rect 347154 568294 347210 568350
rect 347278 568294 347334 568350
rect 347402 568294 347458 568350
rect 347526 568294 347582 568350
rect 347154 568170 347210 568226
rect 347278 568170 347334 568226
rect 347402 568170 347458 568226
rect 347526 568170 347582 568226
rect 347154 568046 347210 568102
rect 347278 568046 347334 568102
rect 347402 568046 347458 568102
rect 347526 568046 347582 568102
rect 347154 567922 347210 567978
rect 347278 567922 347334 567978
rect 347402 567922 347458 567978
rect 347526 567922 347582 567978
rect 347154 550294 347210 550350
rect 347278 550294 347334 550350
rect 347402 550294 347458 550350
rect 347526 550294 347582 550350
rect 347154 550170 347210 550226
rect 347278 550170 347334 550226
rect 347402 550170 347458 550226
rect 347526 550170 347582 550226
rect 347154 550046 347210 550102
rect 347278 550046 347334 550102
rect 347402 550046 347458 550102
rect 347526 550046 347582 550102
rect 347154 549922 347210 549978
rect 347278 549922 347334 549978
rect 347402 549922 347458 549978
rect 347526 549922 347582 549978
rect 347154 532294 347210 532350
rect 347278 532294 347334 532350
rect 347402 532294 347458 532350
rect 347526 532294 347582 532350
rect 347154 532170 347210 532226
rect 347278 532170 347334 532226
rect 347402 532170 347458 532226
rect 347526 532170 347582 532226
rect 347154 532046 347210 532102
rect 347278 532046 347334 532102
rect 347402 532046 347458 532102
rect 347526 532046 347582 532102
rect 347154 531922 347210 531978
rect 347278 531922 347334 531978
rect 347402 531922 347458 531978
rect 347526 531922 347582 531978
rect 347154 514294 347210 514350
rect 347278 514294 347334 514350
rect 347402 514294 347458 514350
rect 347526 514294 347582 514350
rect 347154 514170 347210 514226
rect 347278 514170 347334 514226
rect 347402 514170 347458 514226
rect 347526 514170 347582 514226
rect 347154 514046 347210 514102
rect 347278 514046 347334 514102
rect 347402 514046 347458 514102
rect 347526 514046 347582 514102
rect 347154 513922 347210 513978
rect 347278 513922 347334 513978
rect 347402 513922 347458 513978
rect 347526 513922 347582 513978
rect 347154 496294 347210 496350
rect 347278 496294 347334 496350
rect 347402 496294 347458 496350
rect 347526 496294 347582 496350
rect 347154 496170 347210 496226
rect 347278 496170 347334 496226
rect 347402 496170 347458 496226
rect 347526 496170 347582 496226
rect 347154 496046 347210 496102
rect 347278 496046 347334 496102
rect 347402 496046 347458 496102
rect 347526 496046 347582 496102
rect 347154 495922 347210 495978
rect 347278 495922 347334 495978
rect 347402 495922 347458 495978
rect 347526 495922 347582 495978
rect 347154 478294 347210 478350
rect 347278 478294 347334 478350
rect 347402 478294 347458 478350
rect 347526 478294 347582 478350
rect 347154 478170 347210 478226
rect 347278 478170 347334 478226
rect 347402 478170 347458 478226
rect 347526 478170 347582 478226
rect 347154 478046 347210 478102
rect 347278 478046 347334 478102
rect 347402 478046 347458 478102
rect 347526 478046 347582 478102
rect 347154 477922 347210 477978
rect 347278 477922 347334 477978
rect 347402 477922 347458 477978
rect 347526 477922 347582 477978
rect 347154 460294 347210 460350
rect 347278 460294 347334 460350
rect 347402 460294 347458 460350
rect 347526 460294 347582 460350
rect 347154 460170 347210 460226
rect 347278 460170 347334 460226
rect 347402 460170 347458 460226
rect 347526 460170 347582 460226
rect 347154 460046 347210 460102
rect 347278 460046 347334 460102
rect 347402 460046 347458 460102
rect 347526 460046 347582 460102
rect 347154 459922 347210 459978
rect 347278 459922 347334 459978
rect 347402 459922 347458 459978
rect 347526 459922 347582 459978
rect 347154 442294 347210 442350
rect 347278 442294 347334 442350
rect 347402 442294 347458 442350
rect 347526 442294 347582 442350
rect 347154 442170 347210 442226
rect 347278 442170 347334 442226
rect 347402 442170 347458 442226
rect 347526 442170 347582 442226
rect 347154 442046 347210 442102
rect 347278 442046 347334 442102
rect 347402 442046 347458 442102
rect 347526 442046 347582 442102
rect 347154 441922 347210 441978
rect 347278 441922 347334 441978
rect 347402 441922 347458 441978
rect 347526 441922 347582 441978
rect 347154 424294 347210 424350
rect 347278 424294 347334 424350
rect 347402 424294 347458 424350
rect 347526 424294 347582 424350
rect 347154 424170 347210 424226
rect 347278 424170 347334 424226
rect 347402 424170 347458 424226
rect 347526 424170 347582 424226
rect 347154 424046 347210 424102
rect 347278 424046 347334 424102
rect 347402 424046 347458 424102
rect 347526 424046 347582 424102
rect 347154 423922 347210 423978
rect 347278 423922 347334 423978
rect 347402 423922 347458 423978
rect 347526 423922 347582 423978
rect 347154 406294 347210 406350
rect 347278 406294 347334 406350
rect 347402 406294 347458 406350
rect 347526 406294 347582 406350
rect 347154 406170 347210 406226
rect 347278 406170 347334 406226
rect 347402 406170 347458 406226
rect 347526 406170 347582 406226
rect 347154 406046 347210 406102
rect 347278 406046 347334 406102
rect 347402 406046 347458 406102
rect 347526 406046 347582 406102
rect 347154 405922 347210 405978
rect 347278 405922 347334 405978
rect 347402 405922 347458 405978
rect 347526 405922 347582 405978
rect 347154 388294 347210 388350
rect 347278 388294 347334 388350
rect 347402 388294 347458 388350
rect 347526 388294 347582 388350
rect 347154 388170 347210 388226
rect 347278 388170 347334 388226
rect 347402 388170 347458 388226
rect 347526 388170 347582 388226
rect 347154 388046 347210 388102
rect 347278 388046 347334 388102
rect 347402 388046 347458 388102
rect 347526 388046 347582 388102
rect 347154 387922 347210 387978
rect 347278 387922 347334 387978
rect 347402 387922 347458 387978
rect 347526 387922 347582 387978
rect 347154 370294 347210 370350
rect 347278 370294 347334 370350
rect 347402 370294 347458 370350
rect 347526 370294 347582 370350
rect 347154 370170 347210 370226
rect 347278 370170 347334 370226
rect 347402 370170 347458 370226
rect 347526 370170 347582 370226
rect 347154 370046 347210 370102
rect 347278 370046 347334 370102
rect 347402 370046 347458 370102
rect 347526 370046 347582 370102
rect 347154 369922 347210 369978
rect 347278 369922 347334 369978
rect 347402 369922 347458 369978
rect 347526 369922 347582 369978
rect 347154 352294 347210 352350
rect 347278 352294 347334 352350
rect 347402 352294 347458 352350
rect 347526 352294 347582 352350
rect 347154 352170 347210 352226
rect 347278 352170 347334 352226
rect 347402 352170 347458 352226
rect 347526 352170 347582 352226
rect 347154 352046 347210 352102
rect 347278 352046 347334 352102
rect 347402 352046 347458 352102
rect 347526 352046 347582 352102
rect 347154 351922 347210 351978
rect 347278 351922 347334 351978
rect 347402 351922 347458 351978
rect 347526 351922 347582 351978
rect 347154 334294 347210 334350
rect 347278 334294 347334 334350
rect 347402 334294 347458 334350
rect 347526 334294 347582 334350
rect 347154 334170 347210 334226
rect 347278 334170 347334 334226
rect 347402 334170 347458 334226
rect 347526 334170 347582 334226
rect 347154 334046 347210 334102
rect 347278 334046 347334 334102
rect 347402 334046 347458 334102
rect 347526 334046 347582 334102
rect 347154 333922 347210 333978
rect 347278 333922 347334 333978
rect 347402 333922 347458 333978
rect 347526 333922 347582 333978
rect 374154 597156 374210 597212
rect 374278 597156 374334 597212
rect 374402 597156 374458 597212
rect 374526 597156 374582 597212
rect 374154 597032 374210 597088
rect 374278 597032 374334 597088
rect 374402 597032 374458 597088
rect 374526 597032 374582 597088
rect 374154 596908 374210 596964
rect 374278 596908 374334 596964
rect 374402 596908 374458 596964
rect 374526 596908 374582 596964
rect 374154 596784 374210 596840
rect 374278 596784 374334 596840
rect 374402 596784 374458 596840
rect 374526 596784 374582 596840
rect 374154 580294 374210 580350
rect 374278 580294 374334 580350
rect 374402 580294 374458 580350
rect 374526 580294 374582 580350
rect 374154 580170 374210 580226
rect 374278 580170 374334 580226
rect 374402 580170 374458 580226
rect 374526 580170 374582 580226
rect 374154 580046 374210 580102
rect 374278 580046 374334 580102
rect 374402 580046 374458 580102
rect 374526 580046 374582 580102
rect 374154 579922 374210 579978
rect 374278 579922 374334 579978
rect 374402 579922 374458 579978
rect 374526 579922 374582 579978
rect 374154 562294 374210 562350
rect 374278 562294 374334 562350
rect 374402 562294 374458 562350
rect 374526 562294 374582 562350
rect 374154 562170 374210 562226
rect 374278 562170 374334 562226
rect 374402 562170 374458 562226
rect 374526 562170 374582 562226
rect 374154 562046 374210 562102
rect 374278 562046 374334 562102
rect 374402 562046 374458 562102
rect 374526 562046 374582 562102
rect 374154 561922 374210 561978
rect 374278 561922 374334 561978
rect 374402 561922 374458 561978
rect 374526 561922 374582 561978
rect 374154 544294 374210 544350
rect 374278 544294 374334 544350
rect 374402 544294 374458 544350
rect 374526 544294 374582 544350
rect 374154 544170 374210 544226
rect 374278 544170 374334 544226
rect 374402 544170 374458 544226
rect 374526 544170 374582 544226
rect 374154 544046 374210 544102
rect 374278 544046 374334 544102
rect 374402 544046 374458 544102
rect 374526 544046 374582 544102
rect 374154 543922 374210 543978
rect 374278 543922 374334 543978
rect 374402 543922 374458 543978
rect 374526 543922 374582 543978
rect 374154 526294 374210 526350
rect 374278 526294 374334 526350
rect 374402 526294 374458 526350
rect 374526 526294 374582 526350
rect 374154 526170 374210 526226
rect 374278 526170 374334 526226
rect 374402 526170 374458 526226
rect 374526 526170 374582 526226
rect 374154 526046 374210 526102
rect 374278 526046 374334 526102
rect 374402 526046 374458 526102
rect 374526 526046 374582 526102
rect 374154 525922 374210 525978
rect 374278 525922 374334 525978
rect 374402 525922 374458 525978
rect 374526 525922 374582 525978
rect 374154 508294 374210 508350
rect 374278 508294 374334 508350
rect 374402 508294 374458 508350
rect 374526 508294 374582 508350
rect 374154 508170 374210 508226
rect 374278 508170 374334 508226
rect 374402 508170 374458 508226
rect 374526 508170 374582 508226
rect 374154 508046 374210 508102
rect 374278 508046 374334 508102
rect 374402 508046 374458 508102
rect 374526 508046 374582 508102
rect 374154 507922 374210 507978
rect 374278 507922 374334 507978
rect 374402 507922 374458 507978
rect 374526 507922 374582 507978
rect 374154 490294 374210 490350
rect 374278 490294 374334 490350
rect 374402 490294 374458 490350
rect 374526 490294 374582 490350
rect 374154 490170 374210 490226
rect 374278 490170 374334 490226
rect 374402 490170 374458 490226
rect 374526 490170 374582 490226
rect 374154 490046 374210 490102
rect 374278 490046 374334 490102
rect 374402 490046 374458 490102
rect 374526 490046 374582 490102
rect 374154 489922 374210 489978
rect 374278 489922 374334 489978
rect 374402 489922 374458 489978
rect 374526 489922 374582 489978
rect 374154 472294 374210 472350
rect 374278 472294 374334 472350
rect 374402 472294 374458 472350
rect 374526 472294 374582 472350
rect 374154 472170 374210 472226
rect 374278 472170 374334 472226
rect 374402 472170 374458 472226
rect 374526 472170 374582 472226
rect 374154 472046 374210 472102
rect 374278 472046 374334 472102
rect 374402 472046 374458 472102
rect 374526 472046 374582 472102
rect 374154 471922 374210 471978
rect 374278 471922 374334 471978
rect 374402 471922 374458 471978
rect 374526 471922 374582 471978
rect 374154 454294 374210 454350
rect 374278 454294 374334 454350
rect 374402 454294 374458 454350
rect 374526 454294 374582 454350
rect 374154 454170 374210 454226
rect 374278 454170 374334 454226
rect 374402 454170 374458 454226
rect 374526 454170 374582 454226
rect 374154 454046 374210 454102
rect 374278 454046 374334 454102
rect 374402 454046 374458 454102
rect 374526 454046 374582 454102
rect 374154 453922 374210 453978
rect 374278 453922 374334 453978
rect 374402 453922 374458 453978
rect 374526 453922 374582 453978
rect 374154 436294 374210 436350
rect 374278 436294 374334 436350
rect 374402 436294 374458 436350
rect 374526 436294 374582 436350
rect 374154 436170 374210 436226
rect 374278 436170 374334 436226
rect 374402 436170 374458 436226
rect 374526 436170 374582 436226
rect 374154 436046 374210 436102
rect 374278 436046 374334 436102
rect 374402 436046 374458 436102
rect 374526 436046 374582 436102
rect 374154 435922 374210 435978
rect 374278 435922 374334 435978
rect 374402 435922 374458 435978
rect 374526 435922 374582 435978
rect 374154 418294 374210 418350
rect 374278 418294 374334 418350
rect 374402 418294 374458 418350
rect 374526 418294 374582 418350
rect 374154 418170 374210 418226
rect 374278 418170 374334 418226
rect 374402 418170 374458 418226
rect 374526 418170 374582 418226
rect 374154 418046 374210 418102
rect 374278 418046 374334 418102
rect 374402 418046 374458 418102
rect 374526 418046 374582 418102
rect 374154 417922 374210 417978
rect 374278 417922 374334 417978
rect 374402 417922 374458 417978
rect 374526 417922 374582 417978
rect 374154 400294 374210 400350
rect 374278 400294 374334 400350
rect 374402 400294 374458 400350
rect 374526 400294 374582 400350
rect 374154 400170 374210 400226
rect 374278 400170 374334 400226
rect 374402 400170 374458 400226
rect 374526 400170 374582 400226
rect 374154 400046 374210 400102
rect 374278 400046 374334 400102
rect 374402 400046 374458 400102
rect 374526 400046 374582 400102
rect 374154 399922 374210 399978
rect 374278 399922 374334 399978
rect 374402 399922 374458 399978
rect 374526 399922 374582 399978
rect 374154 382294 374210 382350
rect 374278 382294 374334 382350
rect 374402 382294 374458 382350
rect 374526 382294 374582 382350
rect 374154 382170 374210 382226
rect 374278 382170 374334 382226
rect 374402 382170 374458 382226
rect 374526 382170 374582 382226
rect 374154 382046 374210 382102
rect 374278 382046 374334 382102
rect 374402 382046 374458 382102
rect 374526 382046 374582 382102
rect 374154 381922 374210 381978
rect 374278 381922 374334 381978
rect 374402 381922 374458 381978
rect 374526 381922 374582 381978
rect 374154 364294 374210 364350
rect 374278 364294 374334 364350
rect 374402 364294 374458 364350
rect 374526 364294 374582 364350
rect 374154 364170 374210 364226
rect 374278 364170 374334 364226
rect 374402 364170 374458 364226
rect 374526 364170 374582 364226
rect 374154 364046 374210 364102
rect 374278 364046 374334 364102
rect 374402 364046 374458 364102
rect 374526 364046 374582 364102
rect 374154 363922 374210 363978
rect 374278 363922 374334 363978
rect 374402 363922 374458 363978
rect 374526 363922 374582 363978
rect 374154 346294 374210 346350
rect 374278 346294 374334 346350
rect 374402 346294 374458 346350
rect 374526 346294 374582 346350
rect 374154 346170 374210 346226
rect 374278 346170 374334 346226
rect 374402 346170 374458 346226
rect 374526 346170 374582 346226
rect 374154 346046 374210 346102
rect 374278 346046 374334 346102
rect 374402 346046 374458 346102
rect 374526 346046 374582 346102
rect 374154 345922 374210 345978
rect 374278 345922 374334 345978
rect 374402 345922 374458 345978
rect 374526 345922 374582 345978
rect 374154 328294 374210 328350
rect 374278 328294 374334 328350
rect 374402 328294 374458 328350
rect 374526 328294 374582 328350
rect 374154 328170 374210 328226
rect 374278 328170 374334 328226
rect 374402 328170 374458 328226
rect 374526 328170 374582 328226
rect 374154 328046 374210 328102
rect 374278 328046 374334 328102
rect 374402 328046 374458 328102
rect 374526 328046 374582 328102
rect 374154 327922 374210 327978
rect 374278 327922 374334 327978
rect 374402 327922 374458 327978
rect 374526 327922 374582 327978
rect 229878 316294 229934 316350
rect 230002 316294 230058 316350
rect 229878 316170 229934 316226
rect 230002 316170 230058 316226
rect 229878 316046 229934 316102
rect 230002 316046 230058 316102
rect 229878 315922 229934 315978
rect 230002 315922 230058 315978
rect 260598 316294 260654 316350
rect 260722 316294 260778 316350
rect 260598 316170 260654 316226
rect 260722 316170 260778 316226
rect 260598 316046 260654 316102
rect 260722 316046 260778 316102
rect 260598 315922 260654 315978
rect 260722 315922 260778 315978
rect 291318 316294 291374 316350
rect 291442 316294 291498 316350
rect 291318 316170 291374 316226
rect 291442 316170 291498 316226
rect 291318 316046 291374 316102
rect 291442 316046 291498 316102
rect 291318 315922 291374 315978
rect 291442 315922 291498 315978
rect 322038 316294 322094 316350
rect 322162 316294 322218 316350
rect 322038 316170 322094 316226
rect 322162 316170 322218 316226
rect 322038 316046 322094 316102
rect 322162 316046 322218 316102
rect 322038 315922 322094 315978
rect 322162 315922 322218 315978
rect 352758 316294 352814 316350
rect 352882 316294 352938 316350
rect 352758 316170 352814 316226
rect 352882 316170 352938 316226
rect 352758 316046 352814 316102
rect 352882 316046 352938 316102
rect 352758 315922 352814 315978
rect 352882 315922 352938 315978
rect 214518 310294 214574 310350
rect 214642 310294 214698 310350
rect 214518 310170 214574 310226
rect 214642 310170 214698 310226
rect 214518 310046 214574 310102
rect 214642 310046 214698 310102
rect 214518 309922 214574 309978
rect 214642 309922 214698 309978
rect 245238 310294 245294 310350
rect 245362 310294 245418 310350
rect 245238 310170 245294 310226
rect 245362 310170 245418 310226
rect 245238 310046 245294 310102
rect 245362 310046 245418 310102
rect 245238 309922 245294 309978
rect 245362 309922 245418 309978
rect 275958 310294 276014 310350
rect 276082 310294 276138 310350
rect 275958 310170 276014 310226
rect 276082 310170 276138 310226
rect 275958 310046 276014 310102
rect 276082 310046 276138 310102
rect 275958 309922 276014 309978
rect 276082 309922 276138 309978
rect 306678 310294 306734 310350
rect 306802 310294 306858 310350
rect 306678 310170 306734 310226
rect 306802 310170 306858 310226
rect 306678 310046 306734 310102
rect 306802 310046 306858 310102
rect 306678 309922 306734 309978
rect 306802 309922 306858 309978
rect 337398 310294 337454 310350
rect 337522 310294 337578 310350
rect 337398 310170 337454 310226
rect 337522 310170 337578 310226
rect 337398 310046 337454 310102
rect 337522 310046 337578 310102
rect 337398 309922 337454 309978
rect 337522 309922 337578 309978
rect 368118 310294 368174 310350
rect 368242 310294 368298 310350
rect 368118 310170 368174 310226
rect 368242 310170 368298 310226
rect 368118 310046 368174 310102
rect 368242 310046 368298 310102
rect 368118 309922 368174 309978
rect 368242 309922 368298 309978
rect 229878 298294 229934 298350
rect 230002 298294 230058 298350
rect 229878 298170 229934 298226
rect 230002 298170 230058 298226
rect 229878 298046 229934 298102
rect 230002 298046 230058 298102
rect 229878 297922 229934 297978
rect 230002 297922 230058 297978
rect 260598 298294 260654 298350
rect 260722 298294 260778 298350
rect 260598 298170 260654 298226
rect 260722 298170 260778 298226
rect 260598 298046 260654 298102
rect 260722 298046 260778 298102
rect 260598 297922 260654 297978
rect 260722 297922 260778 297978
rect 291318 298294 291374 298350
rect 291442 298294 291498 298350
rect 291318 298170 291374 298226
rect 291442 298170 291498 298226
rect 291318 298046 291374 298102
rect 291442 298046 291498 298102
rect 291318 297922 291374 297978
rect 291442 297922 291498 297978
rect 322038 298294 322094 298350
rect 322162 298294 322218 298350
rect 322038 298170 322094 298226
rect 322162 298170 322218 298226
rect 322038 298046 322094 298102
rect 322162 298046 322218 298102
rect 322038 297922 322094 297978
rect 322162 297922 322218 297978
rect 352758 298294 352814 298350
rect 352882 298294 352938 298350
rect 352758 298170 352814 298226
rect 352882 298170 352938 298226
rect 352758 298046 352814 298102
rect 352882 298046 352938 298102
rect 352758 297922 352814 297978
rect 352882 297922 352938 297978
rect 214518 292294 214574 292350
rect 214642 292294 214698 292350
rect 214518 292170 214574 292226
rect 214642 292170 214698 292226
rect 214518 292046 214574 292102
rect 214642 292046 214698 292102
rect 214518 291922 214574 291978
rect 214642 291922 214698 291978
rect 245238 292294 245294 292350
rect 245362 292294 245418 292350
rect 245238 292170 245294 292226
rect 245362 292170 245418 292226
rect 245238 292046 245294 292102
rect 245362 292046 245418 292102
rect 245238 291922 245294 291978
rect 245362 291922 245418 291978
rect 275958 292294 276014 292350
rect 276082 292294 276138 292350
rect 275958 292170 276014 292226
rect 276082 292170 276138 292226
rect 275958 292046 276014 292102
rect 276082 292046 276138 292102
rect 275958 291922 276014 291978
rect 276082 291922 276138 291978
rect 306678 292294 306734 292350
rect 306802 292294 306858 292350
rect 306678 292170 306734 292226
rect 306802 292170 306858 292226
rect 306678 292046 306734 292102
rect 306802 292046 306858 292102
rect 306678 291922 306734 291978
rect 306802 291922 306858 291978
rect 337398 292294 337454 292350
rect 337522 292294 337578 292350
rect 337398 292170 337454 292226
rect 337522 292170 337578 292226
rect 337398 292046 337454 292102
rect 337522 292046 337578 292102
rect 337398 291922 337454 291978
rect 337522 291922 337578 291978
rect 368118 292294 368174 292350
rect 368242 292294 368298 292350
rect 368118 292170 368174 292226
rect 368242 292170 368298 292226
rect 368118 292046 368174 292102
rect 368242 292046 368298 292102
rect 368118 291922 368174 291978
rect 368242 291922 368298 291978
rect 229878 280294 229934 280350
rect 230002 280294 230058 280350
rect 229878 280170 229934 280226
rect 230002 280170 230058 280226
rect 229878 280046 229934 280102
rect 230002 280046 230058 280102
rect 229878 279922 229934 279978
rect 230002 279922 230058 279978
rect 260598 280294 260654 280350
rect 260722 280294 260778 280350
rect 260598 280170 260654 280226
rect 260722 280170 260778 280226
rect 260598 280046 260654 280102
rect 260722 280046 260778 280102
rect 260598 279922 260654 279978
rect 260722 279922 260778 279978
rect 291318 280294 291374 280350
rect 291442 280294 291498 280350
rect 291318 280170 291374 280226
rect 291442 280170 291498 280226
rect 291318 280046 291374 280102
rect 291442 280046 291498 280102
rect 291318 279922 291374 279978
rect 291442 279922 291498 279978
rect 322038 280294 322094 280350
rect 322162 280294 322218 280350
rect 322038 280170 322094 280226
rect 322162 280170 322218 280226
rect 322038 280046 322094 280102
rect 322162 280046 322218 280102
rect 322038 279922 322094 279978
rect 322162 279922 322218 279978
rect 352758 280294 352814 280350
rect 352882 280294 352938 280350
rect 352758 280170 352814 280226
rect 352882 280170 352938 280226
rect 352758 280046 352814 280102
rect 352882 280046 352938 280102
rect 352758 279922 352814 279978
rect 352882 279922 352938 279978
rect 213500 276362 213556 276418
rect 214518 274294 214574 274350
rect 214642 274294 214698 274350
rect 214518 274170 214574 274226
rect 214642 274170 214698 274226
rect 214518 274046 214574 274102
rect 214642 274046 214698 274102
rect 214518 273922 214574 273978
rect 214642 273922 214698 273978
rect 245238 274294 245294 274350
rect 245362 274294 245418 274350
rect 245238 274170 245294 274226
rect 245362 274170 245418 274226
rect 245238 274046 245294 274102
rect 245362 274046 245418 274102
rect 245238 273922 245294 273978
rect 245362 273922 245418 273978
rect 275958 274294 276014 274350
rect 276082 274294 276138 274350
rect 275958 274170 276014 274226
rect 276082 274170 276138 274226
rect 275958 274046 276014 274102
rect 276082 274046 276138 274102
rect 275958 273922 276014 273978
rect 276082 273922 276138 273978
rect 306678 274294 306734 274350
rect 306802 274294 306858 274350
rect 306678 274170 306734 274226
rect 306802 274170 306858 274226
rect 306678 274046 306734 274102
rect 306802 274046 306858 274102
rect 306678 273922 306734 273978
rect 306802 273922 306858 273978
rect 337398 274294 337454 274350
rect 337522 274294 337578 274350
rect 337398 274170 337454 274226
rect 337522 274170 337578 274226
rect 337398 274046 337454 274102
rect 337522 274046 337578 274102
rect 337398 273922 337454 273978
rect 337522 273922 337578 273978
rect 368118 274294 368174 274350
rect 368242 274294 368298 274350
rect 368118 274170 368174 274226
rect 368242 274170 368298 274226
rect 368118 274046 368174 274102
rect 368242 274046 368298 274102
rect 368118 273922 368174 273978
rect 368242 273922 368298 273978
rect 229878 262294 229934 262350
rect 230002 262294 230058 262350
rect 229878 262170 229934 262226
rect 230002 262170 230058 262226
rect 229878 262046 229934 262102
rect 230002 262046 230058 262102
rect 229878 261922 229934 261978
rect 230002 261922 230058 261978
rect 260598 262294 260654 262350
rect 260722 262294 260778 262350
rect 260598 262170 260654 262226
rect 260722 262170 260778 262226
rect 260598 262046 260654 262102
rect 260722 262046 260778 262102
rect 260598 261922 260654 261978
rect 260722 261922 260778 261978
rect 291318 262294 291374 262350
rect 291442 262294 291498 262350
rect 291318 262170 291374 262226
rect 291442 262170 291498 262226
rect 291318 262046 291374 262102
rect 291442 262046 291498 262102
rect 291318 261922 291374 261978
rect 291442 261922 291498 261978
rect 322038 262294 322094 262350
rect 322162 262294 322218 262350
rect 322038 262170 322094 262226
rect 322162 262170 322218 262226
rect 322038 262046 322094 262102
rect 322162 262046 322218 262102
rect 322038 261922 322094 261978
rect 322162 261922 322218 261978
rect 352758 262294 352814 262350
rect 352882 262294 352938 262350
rect 352758 262170 352814 262226
rect 352882 262170 352938 262226
rect 352758 262046 352814 262102
rect 352882 262046 352938 262102
rect 352758 261922 352814 261978
rect 352882 261922 352938 261978
rect 211820 257822 211876 257878
rect 214518 256294 214574 256350
rect 214642 256294 214698 256350
rect 214518 256170 214574 256226
rect 214642 256170 214698 256226
rect 214518 256046 214574 256102
rect 214642 256046 214698 256102
rect 214518 255922 214574 255978
rect 214642 255922 214698 255978
rect 245238 256294 245294 256350
rect 245362 256294 245418 256350
rect 245238 256170 245294 256226
rect 245362 256170 245418 256226
rect 245238 256046 245294 256102
rect 245362 256046 245418 256102
rect 245238 255922 245294 255978
rect 245362 255922 245418 255978
rect 275958 256294 276014 256350
rect 276082 256294 276138 256350
rect 275958 256170 276014 256226
rect 276082 256170 276138 256226
rect 275958 256046 276014 256102
rect 276082 256046 276138 256102
rect 275958 255922 276014 255978
rect 276082 255922 276138 255978
rect 306678 256294 306734 256350
rect 306802 256294 306858 256350
rect 306678 256170 306734 256226
rect 306802 256170 306858 256226
rect 306678 256046 306734 256102
rect 306802 256046 306858 256102
rect 306678 255922 306734 255978
rect 306802 255922 306858 255978
rect 337398 256294 337454 256350
rect 337522 256294 337578 256350
rect 337398 256170 337454 256226
rect 337522 256170 337578 256226
rect 337398 256046 337454 256102
rect 337522 256046 337578 256102
rect 337398 255922 337454 255978
rect 337522 255922 337578 255978
rect 368118 256294 368174 256350
rect 368242 256294 368298 256350
rect 368118 256170 368174 256226
rect 368242 256170 368298 256226
rect 368118 256046 368174 256102
rect 368242 256046 368298 256102
rect 368118 255922 368174 255978
rect 368242 255922 368298 255978
rect 229878 244294 229934 244350
rect 230002 244294 230058 244350
rect 229878 244170 229934 244226
rect 230002 244170 230058 244226
rect 229878 244046 229934 244102
rect 230002 244046 230058 244102
rect 229878 243922 229934 243978
rect 230002 243922 230058 243978
rect 260598 244294 260654 244350
rect 260722 244294 260778 244350
rect 260598 244170 260654 244226
rect 260722 244170 260778 244226
rect 260598 244046 260654 244102
rect 260722 244046 260778 244102
rect 260598 243922 260654 243978
rect 260722 243922 260778 243978
rect 291318 244294 291374 244350
rect 291442 244294 291498 244350
rect 291318 244170 291374 244226
rect 291442 244170 291498 244226
rect 291318 244046 291374 244102
rect 291442 244046 291498 244102
rect 291318 243922 291374 243978
rect 291442 243922 291498 243978
rect 322038 244294 322094 244350
rect 322162 244294 322218 244350
rect 322038 244170 322094 244226
rect 322162 244170 322218 244226
rect 322038 244046 322094 244102
rect 322162 244046 322218 244102
rect 322038 243922 322094 243978
rect 322162 243922 322218 243978
rect 352758 244294 352814 244350
rect 352882 244294 352938 244350
rect 352758 244170 352814 244226
rect 352882 244170 352938 244226
rect 352758 244046 352814 244102
rect 352882 244046 352938 244102
rect 352758 243922 352814 243978
rect 352882 243922 352938 243978
rect 214518 238294 214574 238350
rect 214642 238294 214698 238350
rect 214518 238170 214574 238226
rect 214642 238170 214698 238226
rect 214518 238046 214574 238102
rect 214642 238046 214698 238102
rect 214518 237922 214574 237978
rect 214642 237922 214698 237978
rect 245238 238294 245294 238350
rect 245362 238294 245418 238350
rect 245238 238170 245294 238226
rect 245362 238170 245418 238226
rect 245238 238046 245294 238102
rect 245362 238046 245418 238102
rect 245238 237922 245294 237978
rect 245362 237922 245418 237978
rect 275958 238294 276014 238350
rect 276082 238294 276138 238350
rect 275958 238170 276014 238226
rect 276082 238170 276138 238226
rect 275958 238046 276014 238102
rect 276082 238046 276138 238102
rect 275958 237922 276014 237978
rect 276082 237922 276138 237978
rect 306678 238294 306734 238350
rect 306802 238294 306858 238350
rect 306678 238170 306734 238226
rect 306802 238170 306858 238226
rect 306678 238046 306734 238102
rect 306802 238046 306858 238102
rect 306678 237922 306734 237978
rect 306802 237922 306858 237978
rect 337398 238294 337454 238350
rect 337522 238294 337578 238350
rect 337398 238170 337454 238226
rect 337522 238170 337578 238226
rect 337398 238046 337454 238102
rect 337522 238046 337578 238102
rect 337398 237922 337454 237978
rect 337522 237922 337578 237978
rect 368118 238294 368174 238350
rect 368242 238294 368298 238350
rect 368118 238170 368174 238226
rect 368242 238170 368298 238226
rect 368118 238046 368174 238102
rect 368242 238046 368298 238102
rect 368118 237922 368174 237978
rect 368242 237922 368298 237978
rect 211708 236042 211764 236098
rect 229878 226294 229934 226350
rect 230002 226294 230058 226350
rect 229878 226170 229934 226226
rect 230002 226170 230058 226226
rect 229878 226046 229934 226102
rect 230002 226046 230058 226102
rect 229878 225922 229934 225978
rect 230002 225922 230058 225978
rect 260598 226294 260654 226350
rect 260722 226294 260778 226350
rect 260598 226170 260654 226226
rect 260722 226170 260778 226226
rect 260598 226046 260654 226102
rect 260722 226046 260778 226102
rect 260598 225922 260654 225978
rect 260722 225922 260778 225978
rect 291318 226294 291374 226350
rect 291442 226294 291498 226350
rect 291318 226170 291374 226226
rect 291442 226170 291498 226226
rect 291318 226046 291374 226102
rect 291442 226046 291498 226102
rect 291318 225922 291374 225978
rect 291442 225922 291498 225978
rect 322038 226294 322094 226350
rect 322162 226294 322218 226350
rect 322038 226170 322094 226226
rect 322162 226170 322218 226226
rect 322038 226046 322094 226102
rect 322162 226046 322218 226102
rect 322038 225922 322094 225978
rect 322162 225922 322218 225978
rect 352758 226294 352814 226350
rect 352882 226294 352938 226350
rect 352758 226170 352814 226226
rect 352882 226170 352938 226226
rect 352758 226046 352814 226102
rect 352882 226046 352938 226102
rect 352758 225922 352814 225978
rect 352882 225922 352938 225978
rect 214518 220294 214574 220350
rect 214642 220294 214698 220350
rect 214518 220170 214574 220226
rect 214642 220170 214698 220226
rect 214518 220046 214574 220102
rect 214642 220046 214698 220102
rect 214518 219922 214574 219978
rect 214642 219922 214698 219978
rect 245238 220294 245294 220350
rect 245362 220294 245418 220350
rect 245238 220170 245294 220226
rect 245362 220170 245418 220226
rect 245238 220046 245294 220102
rect 245362 220046 245418 220102
rect 245238 219922 245294 219978
rect 245362 219922 245418 219978
rect 275958 220294 276014 220350
rect 276082 220294 276138 220350
rect 275958 220170 276014 220226
rect 276082 220170 276138 220226
rect 275958 220046 276014 220102
rect 276082 220046 276138 220102
rect 275958 219922 276014 219978
rect 276082 219922 276138 219978
rect 306678 220294 306734 220350
rect 306802 220294 306858 220350
rect 306678 220170 306734 220226
rect 306802 220170 306858 220226
rect 306678 220046 306734 220102
rect 306802 220046 306858 220102
rect 306678 219922 306734 219978
rect 306802 219922 306858 219978
rect 337398 220294 337454 220350
rect 337522 220294 337578 220350
rect 337398 220170 337454 220226
rect 337522 220170 337578 220226
rect 337398 220046 337454 220102
rect 337522 220046 337578 220102
rect 337398 219922 337454 219978
rect 337522 219922 337578 219978
rect 368118 220294 368174 220350
rect 368242 220294 368298 220350
rect 368118 220170 368174 220226
rect 368242 220170 368298 220226
rect 368118 220046 368174 220102
rect 368242 220046 368298 220102
rect 368118 219922 368174 219978
rect 368242 219922 368298 219978
rect 369404 216602 369460 216658
rect 229878 208294 229934 208350
rect 230002 208294 230058 208350
rect 229878 208170 229934 208226
rect 230002 208170 230058 208226
rect 229878 208046 229934 208102
rect 230002 208046 230058 208102
rect 229878 207922 229934 207978
rect 230002 207922 230058 207978
rect 260598 208294 260654 208350
rect 260722 208294 260778 208350
rect 260598 208170 260654 208226
rect 260722 208170 260778 208226
rect 260598 208046 260654 208102
rect 260722 208046 260778 208102
rect 260598 207922 260654 207978
rect 260722 207922 260778 207978
rect 291318 208294 291374 208350
rect 291442 208294 291498 208350
rect 291318 208170 291374 208226
rect 291442 208170 291498 208226
rect 291318 208046 291374 208102
rect 291442 208046 291498 208102
rect 291318 207922 291374 207978
rect 291442 207922 291498 207978
rect 322038 208294 322094 208350
rect 322162 208294 322218 208350
rect 322038 208170 322094 208226
rect 322162 208170 322218 208226
rect 322038 208046 322094 208102
rect 322162 208046 322218 208102
rect 322038 207922 322094 207978
rect 322162 207922 322218 207978
rect 352758 208294 352814 208350
rect 352882 208294 352938 208350
rect 352758 208170 352814 208226
rect 352882 208170 352938 208226
rect 352758 208046 352814 208102
rect 352882 208046 352938 208102
rect 352758 207922 352814 207978
rect 352882 207922 352938 207978
rect 214518 202294 214574 202350
rect 214642 202294 214698 202350
rect 214518 202170 214574 202226
rect 214642 202170 214698 202226
rect 214518 202046 214574 202102
rect 214642 202046 214698 202102
rect 214518 201922 214574 201978
rect 214642 201922 214698 201978
rect 245238 202294 245294 202350
rect 245362 202294 245418 202350
rect 245238 202170 245294 202226
rect 245362 202170 245418 202226
rect 245238 202046 245294 202102
rect 245362 202046 245418 202102
rect 245238 201922 245294 201978
rect 245362 201922 245418 201978
rect 275958 202294 276014 202350
rect 276082 202294 276138 202350
rect 275958 202170 276014 202226
rect 276082 202170 276138 202226
rect 275958 202046 276014 202102
rect 276082 202046 276138 202102
rect 275958 201922 276014 201978
rect 276082 201922 276138 201978
rect 306678 202294 306734 202350
rect 306802 202294 306858 202350
rect 306678 202170 306734 202226
rect 306802 202170 306858 202226
rect 306678 202046 306734 202102
rect 306802 202046 306858 202102
rect 306678 201922 306734 201978
rect 306802 201922 306858 201978
rect 337398 202294 337454 202350
rect 337522 202294 337578 202350
rect 337398 202170 337454 202226
rect 337522 202170 337578 202226
rect 337398 202046 337454 202102
rect 337522 202046 337578 202102
rect 337398 201922 337454 201978
rect 337522 201922 337578 201978
rect 368118 202294 368174 202350
rect 368242 202294 368298 202350
rect 368118 202170 368174 202226
rect 368242 202170 368298 202226
rect 368118 202046 368174 202102
rect 368242 202046 368298 202102
rect 368118 201922 368174 201978
rect 368242 201922 368298 201978
rect 369516 193922 369572 193978
rect 229878 190294 229934 190350
rect 230002 190294 230058 190350
rect 229878 190170 229934 190226
rect 230002 190170 230058 190226
rect 229878 190046 229934 190102
rect 230002 190046 230058 190102
rect 229878 189922 229934 189978
rect 230002 189922 230058 189978
rect 260598 190294 260654 190350
rect 260722 190294 260778 190350
rect 260598 190170 260654 190226
rect 260722 190170 260778 190226
rect 260598 190046 260654 190102
rect 260722 190046 260778 190102
rect 260598 189922 260654 189978
rect 260722 189922 260778 189978
rect 291318 190294 291374 190350
rect 291442 190294 291498 190350
rect 291318 190170 291374 190226
rect 291442 190170 291498 190226
rect 291318 190046 291374 190102
rect 291442 190046 291498 190102
rect 291318 189922 291374 189978
rect 291442 189922 291498 189978
rect 322038 190294 322094 190350
rect 322162 190294 322218 190350
rect 322038 190170 322094 190226
rect 322162 190170 322218 190226
rect 322038 190046 322094 190102
rect 322162 190046 322218 190102
rect 322038 189922 322094 189978
rect 322162 189922 322218 189978
rect 352758 190294 352814 190350
rect 352882 190294 352938 190350
rect 352758 190170 352814 190226
rect 352882 190170 352938 190226
rect 352758 190046 352814 190102
rect 352882 190046 352938 190102
rect 352758 189922 352814 189978
rect 352882 189922 352938 189978
rect 373772 310922 373828 310978
rect 377874 598116 377930 598172
rect 377998 598116 378054 598172
rect 378122 598116 378178 598172
rect 378246 598116 378302 598172
rect 377874 597992 377930 598048
rect 377998 597992 378054 598048
rect 378122 597992 378178 598048
rect 378246 597992 378302 598048
rect 377874 597868 377930 597924
rect 377998 597868 378054 597924
rect 378122 597868 378178 597924
rect 378246 597868 378302 597924
rect 377874 597744 377930 597800
rect 377998 597744 378054 597800
rect 378122 597744 378178 597800
rect 378246 597744 378302 597800
rect 377874 586294 377930 586350
rect 377998 586294 378054 586350
rect 378122 586294 378178 586350
rect 378246 586294 378302 586350
rect 377874 586170 377930 586226
rect 377998 586170 378054 586226
rect 378122 586170 378178 586226
rect 378246 586170 378302 586226
rect 377874 586046 377930 586102
rect 377998 586046 378054 586102
rect 378122 586046 378178 586102
rect 378246 586046 378302 586102
rect 377874 585922 377930 585978
rect 377998 585922 378054 585978
rect 378122 585922 378178 585978
rect 378246 585922 378302 585978
rect 377874 568294 377930 568350
rect 377998 568294 378054 568350
rect 378122 568294 378178 568350
rect 378246 568294 378302 568350
rect 377874 568170 377930 568226
rect 377998 568170 378054 568226
rect 378122 568170 378178 568226
rect 378246 568170 378302 568226
rect 377874 568046 377930 568102
rect 377998 568046 378054 568102
rect 378122 568046 378178 568102
rect 378246 568046 378302 568102
rect 377874 567922 377930 567978
rect 377998 567922 378054 567978
rect 378122 567922 378178 567978
rect 378246 567922 378302 567978
rect 377874 550294 377930 550350
rect 377998 550294 378054 550350
rect 378122 550294 378178 550350
rect 378246 550294 378302 550350
rect 377874 550170 377930 550226
rect 377998 550170 378054 550226
rect 378122 550170 378178 550226
rect 378246 550170 378302 550226
rect 377874 550046 377930 550102
rect 377998 550046 378054 550102
rect 378122 550046 378178 550102
rect 378246 550046 378302 550102
rect 377874 549922 377930 549978
rect 377998 549922 378054 549978
rect 378122 549922 378178 549978
rect 378246 549922 378302 549978
rect 377874 532294 377930 532350
rect 377998 532294 378054 532350
rect 378122 532294 378178 532350
rect 378246 532294 378302 532350
rect 377874 532170 377930 532226
rect 377998 532170 378054 532226
rect 378122 532170 378178 532226
rect 378246 532170 378302 532226
rect 377874 532046 377930 532102
rect 377998 532046 378054 532102
rect 378122 532046 378178 532102
rect 378246 532046 378302 532102
rect 377874 531922 377930 531978
rect 377998 531922 378054 531978
rect 378122 531922 378178 531978
rect 378246 531922 378302 531978
rect 377874 514294 377930 514350
rect 377998 514294 378054 514350
rect 378122 514294 378178 514350
rect 378246 514294 378302 514350
rect 377874 514170 377930 514226
rect 377998 514170 378054 514226
rect 378122 514170 378178 514226
rect 378246 514170 378302 514226
rect 377874 514046 377930 514102
rect 377998 514046 378054 514102
rect 378122 514046 378178 514102
rect 378246 514046 378302 514102
rect 377874 513922 377930 513978
rect 377998 513922 378054 513978
rect 378122 513922 378178 513978
rect 378246 513922 378302 513978
rect 377874 496294 377930 496350
rect 377998 496294 378054 496350
rect 378122 496294 378178 496350
rect 378246 496294 378302 496350
rect 377874 496170 377930 496226
rect 377998 496170 378054 496226
rect 378122 496170 378178 496226
rect 378246 496170 378302 496226
rect 377874 496046 377930 496102
rect 377998 496046 378054 496102
rect 378122 496046 378178 496102
rect 378246 496046 378302 496102
rect 377874 495922 377930 495978
rect 377998 495922 378054 495978
rect 378122 495922 378178 495978
rect 378246 495922 378302 495978
rect 377874 478294 377930 478350
rect 377998 478294 378054 478350
rect 378122 478294 378178 478350
rect 378246 478294 378302 478350
rect 377874 478170 377930 478226
rect 377998 478170 378054 478226
rect 378122 478170 378178 478226
rect 378246 478170 378302 478226
rect 377874 478046 377930 478102
rect 377998 478046 378054 478102
rect 378122 478046 378178 478102
rect 378246 478046 378302 478102
rect 377874 477922 377930 477978
rect 377998 477922 378054 477978
rect 378122 477922 378178 477978
rect 378246 477922 378302 477978
rect 377874 460294 377930 460350
rect 377998 460294 378054 460350
rect 378122 460294 378178 460350
rect 378246 460294 378302 460350
rect 377874 460170 377930 460226
rect 377998 460170 378054 460226
rect 378122 460170 378178 460226
rect 378246 460170 378302 460226
rect 377874 460046 377930 460102
rect 377998 460046 378054 460102
rect 378122 460046 378178 460102
rect 378246 460046 378302 460102
rect 377874 459922 377930 459978
rect 377998 459922 378054 459978
rect 378122 459922 378178 459978
rect 378246 459922 378302 459978
rect 377874 442294 377930 442350
rect 377998 442294 378054 442350
rect 378122 442294 378178 442350
rect 378246 442294 378302 442350
rect 377874 442170 377930 442226
rect 377998 442170 378054 442226
rect 378122 442170 378178 442226
rect 378246 442170 378302 442226
rect 377874 442046 377930 442102
rect 377998 442046 378054 442102
rect 378122 442046 378178 442102
rect 378246 442046 378302 442102
rect 377874 441922 377930 441978
rect 377998 441922 378054 441978
rect 378122 441922 378178 441978
rect 378246 441922 378302 441978
rect 377874 424294 377930 424350
rect 377998 424294 378054 424350
rect 378122 424294 378178 424350
rect 378246 424294 378302 424350
rect 377874 424170 377930 424226
rect 377998 424170 378054 424226
rect 378122 424170 378178 424226
rect 378246 424170 378302 424226
rect 377874 424046 377930 424102
rect 377998 424046 378054 424102
rect 378122 424046 378178 424102
rect 378246 424046 378302 424102
rect 377874 423922 377930 423978
rect 377998 423922 378054 423978
rect 378122 423922 378178 423978
rect 378246 423922 378302 423978
rect 377874 406294 377930 406350
rect 377998 406294 378054 406350
rect 378122 406294 378178 406350
rect 378246 406294 378302 406350
rect 377874 406170 377930 406226
rect 377998 406170 378054 406226
rect 378122 406170 378178 406226
rect 378246 406170 378302 406226
rect 377874 406046 377930 406102
rect 377998 406046 378054 406102
rect 378122 406046 378178 406102
rect 378246 406046 378302 406102
rect 377874 405922 377930 405978
rect 377998 405922 378054 405978
rect 378122 405922 378178 405978
rect 378246 405922 378302 405978
rect 377874 388294 377930 388350
rect 377998 388294 378054 388350
rect 378122 388294 378178 388350
rect 378246 388294 378302 388350
rect 377874 388170 377930 388226
rect 377998 388170 378054 388226
rect 378122 388170 378178 388226
rect 378246 388170 378302 388226
rect 377874 388046 377930 388102
rect 377998 388046 378054 388102
rect 378122 388046 378178 388102
rect 378246 388046 378302 388102
rect 377874 387922 377930 387978
rect 377998 387922 378054 387978
rect 378122 387922 378178 387978
rect 378246 387922 378302 387978
rect 404874 597156 404930 597212
rect 404998 597156 405054 597212
rect 405122 597156 405178 597212
rect 405246 597156 405302 597212
rect 404874 597032 404930 597088
rect 404998 597032 405054 597088
rect 405122 597032 405178 597088
rect 405246 597032 405302 597088
rect 404874 596908 404930 596964
rect 404998 596908 405054 596964
rect 405122 596908 405178 596964
rect 405246 596908 405302 596964
rect 404874 596784 404930 596840
rect 404998 596784 405054 596840
rect 405122 596784 405178 596840
rect 405246 596784 405302 596840
rect 404874 580294 404930 580350
rect 404998 580294 405054 580350
rect 405122 580294 405178 580350
rect 405246 580294 405302 580350
rect 404874 580170 404930 580226
rect 404998 580170 405054 580226
rect 405122 580170 405178 580226
rect 405246 580170 405302 580226
rect 404874 580046 404930 580102
rect 404998 580046 405054 580102
rect 405122 580046 405178 580102
rect 405246 580046 405302 580102
rect 404874 579922 404930 579978
rect 404998 579922 405054 579978
rect 405122 579922 405178 579978
rect 405246 579922 405302 579978
rect 404874 562294 404930 562350
rect 404998 562294 405054 562350
rect 405122 562294 405178 562350
rect 405246 562294 405302 562350
rect 404874 562170 404930 562226
rect 404998 562170 405054 562226
rect 405122 562170 405178 562226
rect 405246 562170 405302 562226
rect 404874 562046 404930 562102
rect 404998 562046 405054 562102
rect 405122 562046 405178 562102
rect 405246 562046 405302 562102
rect 404874 561922 404930 561978
rect 404998 561922 405054 561978
rect 405122 561922 405178 561978
rect 405246 561922 405302 561978
rect 404874 544294 404930 544350
rect 404998 544294 405054 544350
rect 405122 544294 405178 544350
rect 405246 544294 405302 544350
rect 404874 544170 404930 544226
rect 404998 544170 405054 544226
rect 405122 544170 405178 544226
rect 405246 544170 405302 544226
rect 404874 544046 404930 544102
rect 404998 544046 405054 544102
rect 405122 544046 405178 544102
rect 405246 544046 405302 544102
rect 404874 543922 404930 543978
rect 404998 543922 405054 543978
rect 405122 543922 405178 543978
rect 405246 543922 405302 543978
rect 404874 526294 404930 526350
rect 404998 526294 405054 526350
rect 405122 526294 405178 526350
rect 405246 526294 405302 526350
rect 404874 526170 404930 526226
rect 404998 526170 405054 526226
rect 405122 526170 405178 526226
rect 405246 526170 405302 526226
rect 404874 526046 404930 526102
rect 404998 526046 405054 526102
rect 405122 526046 405178 526102
rect 405246 526046 405302 526102
rect 404874 525922 404930 525978
rect 404998 525922 405054 525978
rect 405122 525922 405178 525978
rect 405246 525922 405302 525978
rect 404874 508294 404930 508350
rect 404998 508294 405054 508350
rect 405122 508294 405178 508350
rect 405246 508294 405302 508350
rect 404874 508170 404930 508226
rect 404998 508170 405054 508226
rect 405122 508170 405178 508226
rect 405246 508170 405302 508226
rect 404874 508046 404930 508102
rect 404998 508046 405054 508102
rect 405122 508046 405178 508102
rect 405246 508046 405302 508102
rect 404874 507922 404930 507978
rect 404998 507922 405054 507978
rect 405122 507922 405178 507978
rect 405246 507922 405302 507978
rect 404874 490294 404930 490350
rect 404998 490294 405054 490350
rect 405122 490294 405178 490350
rect 405246 490294 405302 490350
rect 404874 490170 404930 490226
rect 404998 490170 405054 490226
rect 405122 490170 405178 490226
rect 405246 490170 405302 490226
rect 404874 490046 404930 490102
rect 404998 490046 405054 490102
rect 405122 490046 405178 490102
rect 405246 490046 405302 490102
rect 404874 489922 404930 489978
rect 404998 489922 405054 489978
rect 405122 489922 405178 489978
rect 405246 489922 405302 489978
rect 404874 472294 404930 472350
rect 404998 472294 405054 472350
rect 405122 472294 405178 472350
rect 405246 472294 405302 472350
rect 404874 472170 404930 472226
rect 404998 472170 405054 472226
rect 405122 472170 405178 472226
rect 405246 472170 405302 472226
rect 404874 472046 404930 472102
rect 404998 472046 405054 472102
rect 405122 472046 405178 472102
rect 405246 472046 405302 472102
rect 404874 471922 404930 471978
rect 404998 471922 405054 471978
rect 405122 471922 405178 471978
rect 405246 471922 405302 471978
rect 404874 454294 404930 454350
rect 404998 454294 405054 454350
rect 405122 454294 405178 454350
rect 405246 454294 405302 454350
rect 404874 454170 404930 454226
rect 404998 454170 405054 454226
rect 405122 454170 405178 454226
rect 405246 454170 405302 454226
rect 404874 454046 404930 454102
rect 404998 454046 405054 454102
rect 405122 454046 405178 454102
rect 405246 454046 405302 454102
rect 404874 453922 404930 453978
rect 404998 453922 405054 453978
rect 405122 453922 405178 453978
rect 405246 453922 405302 453978
rect 404874 436294 404930 436350
rect 404998 436294 405054 436350
rect 405122 436294 405178 436350
rect 405246 436294 405302 436350
rect 404874 436170 404930 436226
rect 404998 436170 405054 436226
rect 405122 436170 405178 436226
rect 405246 436170 405302 436226
rect 404874 436046 404930 436102
rect 404998 436046 405054 436102
rect 405122 436046 405178 436102
rect 405246 436046 405302 436102
rect 404874 435922 404930 435978
rect 404998 435922 405054 435978
rect 405122 435922 405178 435978
rect 405246 435922 405302 435978
rect 404874 418294 404930 418350
rect 404998 418294 405054 418350
rect 405122 418294 405178 418350
rect 405246 418294 405302 418350
rect 404874 418170 404930 418226
rect 404998 418170 405054 418226
rect 405122 418170 405178 418226
rect 405246 418170 405302 418226
rect 404874 418046 404930 418102
rect 404998 418046 405054 418102
rect 405122 418046 405178 418102
rect 405246 418046 405302 418102
rect 404874 417922 404930 417978
rect 404998 417922 405054 417978
rect 405122 417922 405178 417978
rect 405246 417922 405302 417978
rect 404874 400294 404930 400350
rect 404998 400294 405054 400350
rect 405122 400294 405178 400350
rect 405246 400294 405302 400350
rect 404874 400170 404930 400226
rect 404998 400170 405054 400226
rect 405122 400170 405178 400226
rect 405246 400170 405302 400226
rect 404874 400046 404930 400102
rect 404998 400046 405054 400102
rect 405122 400046 405178 400102
rect 405246 400046 405302 400102
rect 404874 399922 404930 399978
rect 404998 399922 405054 399978
rect 405122 399922 405178 399978
rect 405246 399922 405302 399978
rect 404874 382294 404930 382350
rect 404998 382294 405054 382350
rect 405122 382294 405178 382350
rect 405246 382294 405302 382350
rect 404874 382170 404930 382226
rect 404998 382170 405054 382226
rect 405122 382170 405178 382226
rect 405246 382170 405302 382226
rect 404874 382046 404930 382102
rect 404998 382046 405054 382102
rect 405122 382046 405178 382102
rect 405246 382046 405302 382102
rect 404874 381922 404930 381978
rect 404998 381922 405054 381978
rect 405122 381922 405178 381978
rect 405246 381922 405302 381978
rect 377874 370294 377930 370350
rect 377998 370294 378054 370350
rect 378122 370294 378178 370350
rect 378246 370294 378302 370350
rect 377874 370170 377930 370226
rect 377998 370170 378054 370226
rect 378122 370170 378178 370226
rect 378246 370170 378302 370226
rect 377874 370046 377930 370102
rect 377998 370046 378054 370102
rect 378122 370046 378178 370102
rect 378246 370046 378302 370102
rect 377874 369922 377930 369978
rect 377998 369922 378054 369978
rect 378122 369922 378178 369978
rect 378246 369922 378302 369978
rect 377874 352294 377930 352350
rect 377998 352294 378054 352350
rect 378122 352294 378178 352350
rect 378246 352294 378302 352350
rect 377874 352170 377930 352226
rect 377998 352170 378054 352226
rect 378122 352170 378178 352226
rect 378246 352170 378302 352226
rect 377874 352046 377930 352102
rect 377998 352046 378054 352102
rect 378122 352046 378178 352102
rect 378246 352046 378302 352102
rect 377874 351922 377930 351978
rect 377998 351922 378054 351978
rect 378122 351922 378178 351978
rect 378246 351922 378302 351978
rect 377874 334294 377930 334350
rect 377998 334294 378054 334350
rect 378122 334294 378178 334350
rect 378246 334294 378302 334350
rect 377874 334170 377930 334226
rect 377998 334170 378054 334226
rect 378122 334170 378178 334226
rect 378246 334170 378302 334226
rect 377874 334046 377930 334102
rect 377998 334046 378054 334102
rect 378122 334046 378178 334102
rect 378246 334046 378302 334102
rect 377874 333922 377930 333978
rect 377998 333922 378054 333978
rect 378122 333922 378178 333978
rect 378246 333922 378302 333978
rect 374154 310294 374210 310350
rect 374278 310294 374334 310350
rect 374402 310294 374458 310350
rect 374526 310294 374582 310350
rect 374154 310170 374210 310226
rect 374278 310170 374334 310226
rect 374402 310170 374458 310226
rect 374526 310170 374582 310226
rect 374154 310046 374210 310102
rect 374278 310046 374334 310102
rect 374402 310046 374458 310102
rect 374526 310046 374582 310102
rect 374154 309922 374210 309978
rect 374278 309922 374334 309978
rect 374402 309922 374458 309978
rect 374526 309922 374582 309978
rect 370860 270602 370916 270658
rect 214518 184294 214574 184350
rect 214642 184294 214698 184350
rect 214518 184170 214574 184226
rect 214642 184170 214698 184226
rect 214518 184046 214574 184102
rect 214642 184046 214698 184102
rect 214518 183922 214574 183978
rect 214642 183922 214698 183978
rect 245238 184294 245294 184350
rect 245362 184294 245418 184350
rect 245238 184170 245294 184226
rect 245362 184170 245418 184226
rect 245238 184046 245294 184102
rect 245362 184046 245418 184102
rect 245238 183922 245294 183978
rect 245362 183922 245418 183978
rect 275958 184294 276014 184350
rect 276082 184294 276138 184350
rect 275958 184170 276014 184226
rect 276082 184170 276138 184226
rect 275958 184046 276014 184102
rect 276082 184046 276138 184102
rect 275958 183922 276014 183978
rect 276082 183922 276138 183978
rect 306678 184294 306734 184350
rect 306802 184294 306858 184350
rect 306678 184170 306734 184226
rect 306802 184170 306858 184226
rect 306678 184046 306734 184102
rect 306802 184046 306858 184102
rect 306678 183922 306734 183978
rect 306802 183922 306858 183978
rect 337398 184294 337454 184350
rect 337522 184294 337578 184350
rect 337398 184170 337454 184226
rect 337522 184170 337578 184226
rect 337398 184046 337454 184102
rect 337522 184046 337578 184102
rect 337398 183922 337454 183978
rect 337522 183922 337578 183978
rect 368118 184294 368174 184350
rect 368242 184294 368298 184350
rect 368118 184170 368174 184226
rect 368242 184170 368298 184226
rect 368118 184046 368174 184102
rect 368242 184046 368298 184102
rect 368118 183922 368174 183978
rect 368242 183922 368298 183978
rect 229878 172294 229934 172350
rect 230002 172294 230058 172350
rect 229878 172170 229934 172226
rect 230002 172170 230058 172226
rect 229878 172046 229934 172102
rect 230002 172046 230058 172102
rect 229878 171922 229934 171978
rect 230002 171922 230058 171978
rect 260598 172294 260654 172350
rect 260722 172294 260778 172350
rect 260598 172170 260654 172226
rect 260722 172170 260778 172226
rect 260598 172046 260654 172102
rect 260722 172046 260778 172102
rect 260598 171922 260654 171978
rect 260722 171922 260778 171978
rect 291318 172294 291374 172350
rect 291442 172294 291498 172350
rect 291318 172170 291374 172226
rect 291442 172170 291498 172226
rect 291318 172046 291374 172102
rect 291442 172046 291498 172102
rect 291318 171922 291374 171978
rect 291442 171922 291498 171978
rect 322038 172294 322094 172350
rect 322162 172294 322218 172350
rect 322038 172170 322094 172226
rect 322162 172170 322218 172226
rect 322038 172046 322094 172102
rect 322162 172046 322218 172102
rect 322038 171922 322094 171978
rect 322162 171922 322218 171978
rect 352758 172294 352814 172350
rect 352882 172294 352938 172350
rect 352758 172170 352814 172226
rect 352882 172170 352938 172226
rect 352758 172046 352814 172102
rect 352882 172046 352938 172102
rect 352758 171922 352814 171978
rect 352882 171922 352938 171978
rect 214518 166294 214574 166350
rect 214642 166294 214698 166350
rect 214518 166170 214574 166226
rect 214642 166170 214698 166226
rect 214518 166046 214574 166102
rect 214642 166046 214698 166102
rect 214518 165922 214574 165978
rect 214642 165922 214698 165978
rect 245238 166294 245294 166350
rect 245362 166294 245418 166350
rect 245238 166170 245294 166226
rect 245362 166170 245418 166226
rect 245238 166046 245294 166102
rect 245362 166046 245418 166102
rect 245238 165922 245294 165978
rect 245362 165922 245418 165978
rect 275958 166294 276014 166350
rect 276082 166294 276138 166350
rect 275958 166170 276014 166226
rect 276082 166170 276138 166226
rect 275958 166046 276014 166102
rect 276082 166046 276138 166102
rect 275958 165922 276014 165978
rect 276082 165922 276138 165978
rect 306678 166294 306734 166350
rect 306802 166294 306858 166350
rect 306678 166170 306734 166226
rect 306802 166170 306858 166226
rect 306678 166046 306734 166102
rect 306802 166046 306858 166102
rect 306678 165922 306734 165978
rect 306802 165922 306858 165978
rect 337398 166294 337454 166350
rect 337522 166294 337578 166350
rect 337398 166170 337454 166226
rect 337522 166170 337578 166226
rect 337398 166046 337454 166102
rect 337522 166046 337578 166102
rect 337398 165922 337454 165978
rect 337522 165922 337578 165978
rect 368118 166294 368174 166350
rect 368242 166294 368298 166350
rect 368118 166170 368174 166226
rect 368242 166170 368298 166226
rect 368118 166046 368174 166102
rect 368242 166046 368298 166102
rect 368118 165922 368174 165978
rect 368242 165922 368298 165978
rect 229878 154294 229934 154350
rect 230002 154294 230058 154350
rect 229878 154170 229934 154226
rect 230002 154170 230058 154226
rect 229878 154046 229934 154102
rect 230002 154046 230058 154102
rect 229878 153922 229934 153978
rect 230002 153922 230058 153978
rect 260598 154294 260654 154350
rect 260722 154294 260778 154350
rect 260598 154170 260654 154226
rect 260722 154170 260778 154226
rect 260598 154046 260654 154102
rect 260722 154046 260778 154102
rect 260598 153922 260654 153978
rect 260722 153922 260778 153978
rect 291318 154294 291374 154350
rect 291442 154294 291498 154350
rect 291318 154170 291374 154226
rect 291442 154170 291498 154226
rect 291318 154046 291374 154102
rect 291442 154046 291498 154102
rect 291318 153922 291374 153978
rect 291442 153922 291498 153978
rect 322038 154294 322094 154350
rect 322162 154294 322218 154350
rect 322038 154170 322094 154226
rect 322162 154170 322218 154226
rect 322038 154046 322094 154102
rect 322162 154046 322218 154102
rect 322038 153922 322094 153978
rect 322162 153922 322218 153978
rect 352758 154294 352814 154350
rect 352882 154294 352938 154350
rect 352758 154170 352814 154226
rect 352882 154170 352938 154226
rect 352758 154046 352814 154102
rect 352882 154046 352938 154102
rect 352758 153922 352814 153978
rect 352882 153922 352938 153978
rect 214518 148294 214574 148350
rect 214642 148294 214698 148350
rect 214518 148170 214574 148226
rect 214642 148170 214698 148226
rect 214518 148046 214574 148102
rect 214642 148046 214698 148102
rect 214518 147922 214574 147978
rect 214642 147922 214698 147978
rect 245238 148294 245294 148350
rect 245362 148294 245418 148350
rect 245238 148170 245294 148226
rect 245362 148170 245418 148226
rect 245238 148046 245294 148102
rect 245362 148046 245418 148102
rect 245238 147922 245294 147978
rect 245362 147922 245418 147978
rect 275958 148294 276014 148350
rect 276082 148294 276138 148350
rect 275958 148170 276014 148226
rect 276082 148170 276138 148226
rect 275958 148046 276014 148102
rect 276082 148046 276138 148102
rect 275958 147922 276014 147978
rect 276082 147922 276138 147978
rect 306678 148294 306734 148350
rect 306802 148294 306858 148350
rect 306678 148170 306734 148226
rect 306802 148170 306858 148226
rect 306678 148046 306734 148102
rect 306802 148046 306858 148102
rect 306678 147922 306734 147978
rect 306802 147922 306858 147978
rect 337398 148294 337454 148350
rect 337522 148294 337578 148350
rect 337398 148170 337454 148226
rect 337522 148170 337578 148226
rect 337398 148046 337454 148102
rect 337522 148046 337578 148102
rect 337398 147922 337454 147978
rect 337522 147922 337578 147978
rect 368118 148294 368174 148350
rect 368242 148294 368298 148350
rect 368118 148170 368174 148226
rect 368242 148170 368298 148226
rect 368118 148046 368174 148102
rect 368242 148046 368298 148102
rect 368118 147922 368174 147978
rect 368242 147922 368298 147978
rect 229878 136294 229934 136350
rect 230002 136294 230058 136350
rect 229878 136170 229934 136226
rect 230002 136170 230058 136226
rect 229878 136046 229934 136102
rect 230002 136046 230058 136102
rect 229878 135922 229934 135978
rect 230002 135922 230058 135978
rect 260598 136294 260654 136350
rect 260722 136294 260778 136350
rect 260598 136170 260654 136226
rect 260722 136170 260778 136226
rect 260598 136046 260654 136102
rect 260722 136046 260778 136102
rect 260598 135922 260654 135978
rect 260722 135922 260778 135978
rect 291318 136294 291374 136350
rect 291442 136294 291498 136350
rect 291318 136170 291374 136226
rect 291442 136170 291498 136226
rect 291318 136046 291374 136102
rect 291442 136046 291498 136102
rect 291318 135922 291374 135978
rect 291442 135922 291498 135978
rect 322038 136294 322094 136350
rect 322162 136294 322218 136350
rect 322038 136170 322094 136226
rect 322162 136170 322218 136226
rect 322038 136046 322094 136102
rect 322162 136046 322218 136102
rect 322038 135922 322094 135978
rect 322162 135922 322218 135978
rect 352758 136294 352814 136350
rect 352882 136294 352938 136350
rect 352758 136170 352814 136226
rect 352882 136170 352938 136226
rect 352758 136046 352814 136102
rect 352882 136046 352938 136102
rect 352758 135922 352814 135978
rect 352882 135922 352938 135978
rect 214518 130294 214574 130350
rect 214642 130294 214698 130350
rect 214518 130170 214574 130226
rect 214642 130170 214698 130226
rect 214518 130046 214574 130102
rect 214642 130046 214698 130102
rect 214518 129922 214574 129978
rect 214642 129922 214698 129978
rect 245238 130294 245294 130350
rect 245362 130294 245418 130350
rect 245238 130170 245294 130226
rect 245362 130170 245418 130226
rect 245238 130046 245294 130102
rect 245362 130046 245418 130102
rect 245238 129922 245294 129978
rect 245362 129922 245418 129978
rect 275958 130294 276014 130350
rect 276082 130294 276138 130350
rect 275958 130170 276014 130226
rect 276082 130170 276138 130226
rect 275958 130046 276014 130102
rect 276082 130046 276138 130102
rect 275958 129922 276014 129978
rect 276082 129922 276138 129978
rect 306678 130294 306734 130350
rect 306802 130294 306858 130350
rect 306678 130170 306734 130226
rect 306802 130170 306858 130226
rect 306678 130046 306734 130102
rect 306802 130046 306858 130102
rect 306678 129922 306734 129978
rect 306802 129922 306858 129978
rect 337398 130294 337454 130350
rect 337522 130294 337578 130350
rect 337398 130170 337454 130226
rect 337522 130170 337578 130226
rect 337398 130046 337454 130102
rect 337522 130046 337578 130102
rect 337398 129922 337454 129978
rect 337522 129922 337578 129978
rect 368118 130294 368174 130350
rect 368242 130294 368298 130350
rect 368118 130170 368174 130226
rect 368242 130170 368298 130226
rect 368118 130046 368174 130102
rect 368242 130046 368298 130102
rect 368118 129922 368174 129978
rect 368242 129922 368298 129978
rect 229878 118294 229934 118350
rect 230002 118294 230058 118350
rect 229878 118170 229934 118226
rect 230002 118170 230058 118226
rect 229878 118046 229934 118102
rect 230002 118046 230058 118102
rect 229878 117922 229934 117978
rect 230002 117922 230058 117978
rect 260598 118294 260654 118350
rect 260722 118294 260778 118350
rect 260598 118170 260654 118226
rect 260722 118170 260778 118226
rect 260598 118046 260654 118102
rect 260722 118046 260778 118102
rect 260598 117922 260654 117978
rect 260722 117922 260778 117978
rect 291318 118294 291374 118350
rect 291442 118294 291498 118350
rect 291318 118170 291374 118226
rect 291442 118170 291498 118226
rect 291318 118046 291374 118102
rect 291442 118046 291498 118102
rect 291318 117922 291374 117978
rect 291442 117922 291498 117978
rect 322038 118294 322094 118350
rect 322162 118294 322218 118350
rect 322038 118170 322094 118226
rect 322162 118170 322218 118226
rect 322038 118046 322094 118102
rect 322162 118046 322218 118102
rect 322038 117922 322094 117978
rect 322162 117922 322218 117978
rect 352758 118294 352814 118350
rect 352882 118294 352938 118350
rect 352758 118170 352814 118226
rect 352882 118170 352938 118226
rect 352758 118046 352814 118102
rect 352882 118046 352938 118102
rect 352758 117922 352814 117978
rect 352882 117922 352938 117978
rect 214518 112294 214574 112350
rect 214642 112294 214698 112350
rect 214518 112170 214574 112226
rect 214642 112170 214698 112226
rect 214518 112046 214574 112102
rect 214642 112046 214698 112102
rect 214518 111922 214574 111978
rect 214642 111922 214698 111978
rect 245238 112294 245294 112350
rect 245362 112294 245418 112350
rect 245238 112170 245294 112226
rect 245362 112170 245418 112226
rect 245238 112046 245294 112102
rect 245362 112046 245418 112102
rect 245238 111922 245294 111978
rect 245362 111922 245418 111978
rect 275958 112294 276014 112350
rect 276082 112294 276138 112350
rect 275958 112170 276014 112226
rect 276082 112170 276138 112226
rect 275958 112046 276014 112102
rect 276082 112046 276138 112102
rect 275958 111922 276014 111978
rect 276082 111922 276138 111978
rect 306678 112294 306734 112350
rect 306802 112294 306858 112350
rect 306678 112170 306734 112226
rect 306802 112170 306858 112226
rect 306678 112046 306734 112102
rect 306802 112046 306858 112102
rect 306678 111922 306734 111978
rect 306802 111922 306858 111978
rect 337398 112294 337454 112350
rect 337522 112294 337578 112350
rect 337398 112170 337454 112226
rect 337522 112170 337578 112226
rect 337398 112046 337454 112102
rect 337522 112046 337578 112102
rect 337398 111922 337454 111978
rect 337522 111922 337578 111978
rect 368118 112294 368174 112350
rect 368242 112294 368298 112350
rect 368118 112170 368174 112226
rect 368242 112170 368298 112226
rect 368118 112046 368174 112102
rect 368242 112046 368298 112102
rect 368118 111922 368174 111978
rect 368242 111922 368298 111978
rect 229878 100294 229934 100350
rect 230002 100294 230058 100350
rect 229878 100170 229934 100226
rect 230002 100170 230058 100226
rect 229878 100046 229934 100102
rect 230002 100046 230058 100102
rect 229878 99922 229934 99978
rect 230002 99922 230058 99978
rect 260598 100294 260654 100350
rect 260722 100294 260778 100350
rect 260598 100170 260654 100226
rect 260722 100170 260778 100226
rect 260598 100046 260654 100102
rect 260722 100046 260778 100102
rect 260598 99922 260654 99978
rect 260722 99922 260778 99978
rect 291318 100294 291374 100350
rect 291442 100294 291498 100350
rect 291318 100170 291374 100226
rect 291442 100170 291498 100226
rect 291318 100046 291374 100102
rect 291442 100046 291498 100102
rect 291318 99922 291374 99978
rect 291442 99922 291498 99978
rect 322038 100294 322094 100350
rect 322162 100294 322218 100350
rect 322038 100170 322094 100226
rect 322162 100170 322218 100226
rect 322038 100046 322094 100102
rect 322162 100046 322218 100102
rect 322038 99922 322094 99978
rect 322162 99922 322218 99978
rect 352758 100294 352814 100350
rect 352882 100294 352938 100350
rect 352758 100170 352814 100226
rect 352882 100170 352938 100226
rect 352758 100046 352814 100102
rect 352882 100046 352938 100102
rect 352758 99922 352814 99978
rect 352882 99922 352938 99978
rect 214518 94294 214574 94350
rect 214642 94294 214698 94350
rect 214518 94170 214574 94226
rect 214642 94170 214698 94226
rect 214518 94046 214574 94102
rect 214642 94046 214698 94102
rect 214518 93922 214574 93978
rect 214642 93922 214698 93978
rect 245238 94294 245294 94350
rect 245362 94294 245418 94350
rect 245238 94170 245294 94226
rect 245362 94170 245418 94226
rect 245238 94046 245294 94102
rect 245362 94046 245418 94102
rect 245238 93922 245294 93978
rect 245362 93922 245418 93978
rect 275958 94294 276014 94350
rect 276082 94294 276138 94350
rect 275958 94170 276014 94226
rect 276082 94170 276138 94226
rect 275958 94046 276014 94102
rect 276082 94046 276138 94102
rect 275958 93922 276014 93978
rect 276082 93922 276138 93978
rect 306678 94294 306734 94350
rect 306802 94294 306858 94350
rect 306678 94170 306734 94226
rect 306802 94170 306858 94226
rect 306678 94046 306734 94102
rect 306802 94046 306858 94102
rect 306678 93922 306734 93978
rect 306802 93922 306858 93978
rect 337398 94294 337454 94350
rect 337522 94294 337578 94350
rect 337398 94170 337454 94226
rect 337522 94170 337578 94226
rect 337398 94046 337454 94102
rect 337522 94046 337578 94102
rect 337398 93922 337454 93978
rect 337522 93922 337578 93978
rect 368118 94294 368174 94350
rect 368242 94294 368298 94350
rect 368118 94170 368174 94226
rect 368242 94170 368298 94226
rect 368118 94046 368174 94102
rect 368242 94046 368298 94102
rect 368118 93922 368174 93978
rect 368242 93922 368298 93978
rect 229878 82294 229934 82350
rect 230002 82294 230058 82350
rect 229878 82170 229934 82226
rect 230002 82170 230058 82226
rect 229878 82046 229934 82102
rect 230002 82046 230058 82102
rect 229878 81922 229934 81978
rect 230002 81922 230058 81978
rect 260598 82294 260654 82350
rect 260722 82294 260778 82350
rect 260598 82170 260654 82226
rect 260722 82170 260778 82226
rect 260598 82046 260654 82102
rect 260722 82046 260778 82102
rect 260598 81922 260654 81978
rect 260722 81922 260778 81978
rect 291318 82294 291374 82350
rect 291442 82294 291498 82350
rect 291318 82170 291374 82226
rect 291442 82170 291498 82226
rect 291318 82046 291374 82102
rect 291442 82046 291498 82102
rect 291318 81922 291374 81978
rect 291442 81922 291498 81978
rect 322038 82294 322094 82350
rect 322162 82294 322218 82350
rect 322038 82170 322094 82226
rect 322162 82170 322218 82226
rect 322038 82046 322094 82102
rect 322162 82046 322218 82102
rect 322038 81922 322094 81978
rect 322162 81922 322218 81978
rect 352758 82294 352814 82350
rect 352882 82294 352938 82350
rect 352758 82170 352814 82226
rect 352882 82170 352938 82226
rect 352758 82046 352814 82102
rect 352882 82046 352938 82102
rect 352758 81922 352814 81978
rect 352882 81922 352938 81978
rect 214518 76294 214574 76350
rect 214642 76294 214698 76350
rect 214518 76170 214574 76226
rect 214642 76170 214698 76226
rect 214518 76046 214574 76102
rect 214642 76046 214698 76102
rect 214518 75922 214574 75978
rect 214642 75922 214698 75978
rect 245238 76294 245294 76350
rect 245362 76294 245418 76350
rect 245238 76170 245294 76226
rect 245362 76170 245418 76226
rect 245238 76046 245294 76102
rect 245362 76046 245418 76102
rect 245238 75922 245294 75978
rect 245362 75922 245418 75978
rect 275958 76294 276014 76350
rect 276082 76294 276138 76350
rect 275958 76170 276014 76226
rect 276082 76170 276138 76226
rect 275958 76046 276014 76102
rect 276082 76046 276138 76102
rect 275958 75922 276014 75978
rect 276082 75922 276138 75978
rect 306678 76294 306734 76350
rect 306802 76294 306858 76350
rect 306678 76170 306734 76226
rect 306802 76170 306858 76226
rect 306678 76046 306734 76102
rect 306802 76046 306858 76102
rect 306678 75922 306734 75978
rect 306802 75922 306858 75978
rect 337398 76294 337454 76350
rect 337522 76294 337578 76350
rect 337398 76170 337454 76226
rect 337522 76170 337578 76226
rect 337398 76046 337454 76102
rect 337522 76046 337578 76102
rect 337398 75922 337454 75978
rect 337522 75922 337578 75978
rect 368118 76294 368174 76350
rect 368242 76294 368298 76350
rect 368118 76170 368174 76226
rect 368242 76170 368298 76226
rect 368118 76046 368174 76102
rect 368242 76046 368298 76102
rect 368118 75922 368174 75978
rect 368242 75922 368298 75978
rect 370972 209042 371028 209098
rect 229878 64294 229934 64350
rect 230002 64294 230058 64350
rect 229878 64170 229934 64226
rect 230002 64170 230058 64226
rect 229878 64046 229934 64102
rect 230002 64046 230058 64102
rect 229878 63922 229934 63978
rect 230002 63922 230058 63978
rect 260598 64294 260654 64350
rect 260722 64294 260778 64350
rect 260598 64170 260654 64226
rect 260722 64170 260778 64226
rect 260598 64046 260654 64102
rect 260722 64046 260778 64102
rect 260598 63922 260654 63978
rect 260722 63922 260778 63978
rect 291318 64294 291374 64350
rect 291442 64294 291498 64350
rect 291318 64170 291374 64226
rect 291442 64170 291498 64226
rect 291318 64046 291374 64102
rect 291442 64046 291498 64102
rect 291318 63922 291374 63978
rect 291442 63922 291498 63978
rect 322038 64294 322094 64350
rect 322162 64294 322218 64350
rect 322038 64170 322094 64226
rect 322162 64170 322218 64226
rect 322038 64046 322094 64102
rect 322162 64046 322218 64102
rect 322038 63922 322094 63978
rect 322162 63922 322218 63978
rect 352758 64294 352814 64350
rect 352882 64294 352938 64350
rect 352758 64170 352814 64226
rect 352882 64170 352938 64226
rect 352758 64046 352814 64102
rect 352882 64046 352938 64102
rect 352758 63922 352814 63978
rect 352882 63922 352938 63978
rect 214518 58294 214574 58350
rect 214642 58294 214698 58350
rect 214518 58170 214574 58226
rect 214642 58170 214698 58226
rect 214518 58046 214574 58102
rect 214642 58046 214698 58102
rect 214518 57922 214574 57978
rect 214642 57922 214698 57978
rect 245238 58294 245294 58350
rect 245362 58294 245418 58350
rect 245238 58170 245294 58226
rect 245362 58170 245418 58226
rect 245238 58046 245294 58102
rect 245362 58046 245418 58102
rect 245238 57922 245294 57978
rect 245362 57922 245418 57978
rect 275958 58294 276014 58350
rect 276082 58294 276138 58350
rect 275958 58170 276014 58226
rect 276082 58170 276138 58226
rect 275958 58046 276014 58102
rect 276082 58046 276138 58102
rect 275958 57922 276014 57978
rect 276082 57922 276138 57978
rect 306678 58294 306734 58350
rect 306802 58294 306858 58350
rect 306678 58170 306734 58226
rect 306802 58170 306858 58226
rect 306678 58046 306734 58102
rect 306802 58046 306858 58102
rect 306678 57922 306734 57978
rect 306802 57922 306858 57978
rect 337398 58294 337454 58350
rect 337522 58294 337578 58350
rect 337398 58170 337454 58226
rect 337522 58170 337578 58226
rect 337398 58046 337454 58102
rect 337522 58046 337578 58102
rect 337398 57922 337454 57978
rect 337522 57922 337578 57978
rect 368118 58294 368174 58350
rect 368242 58294 368298 58350
rect 368118 58170 368174 58226
rect 368242 58170 368298 58226
rect 368118 58046 368174 58102
rect 368242 58046 368298 58102
rect 368118 57922 368174 57978
rect 368242 57922 368298 57978
rect 209916 56942 209972 56998
rect 370412 56942 370468 56998
rect 193554 46294 193610 46350
rect 193678 46294 193734 46350
rect 193802 46294 193858 46350
rect 193926 46294 193982 46350
rect 193554 46170 193610 46226
rect 193678 46170 193734 46226
rect 193802 46170 193858 46226
rect 193926 46170 193982 46226
rect 193554 46046 193610 46102
rect 193678 46046 193734 46102
rect 193802 46046 193858 46102
rect 193926 46046 193982 46102
rect 193554 45922 193610 45978
rect 193678 45922 193734 45978
rect 193802 45922 193858 45978
rect 193926 45922 193982 45978
rect 193554 28294 193610 28350
rect 193678 28294 193734 28350
rect 193802 28294 193858 28350
rect 193926 28294 193982 28350
rect 193554 28170 193610 28226
rect 193678 28170 193734 28226
rect 193802 28170 193858 28226
rect 193926 28170 193982 28226
rect 193554 28046 193610 28102
rect 193678 28046 193734 28102
rect 193802 28046 193858 28102
rect 193926 28046 193982 28102
rect 193554 27922 193610 27978
rect 193678 27922 193734 27978
rect 193802 27922 193858 27978
rect 193926 27922 193982 27978
rect 220554 40294 220610 40350
rect 220678 40294 220734 40350
rect 220802 40294 220858 40350
rect 220926 40294 220982 40350
rect 220554 40170 220610 40226
rect 220678 40170 220734 40226
rect 220802 40170 220858 40226
rect 220926 40170 220982 40226
rect 220554 40046 220610 40102
rect 220678 40046 220734 40102
rect 220802 40046 220858 40102
rect 220926 40046 220982 40102
rect 220554 39922 220610 39978
rect 220678 39922 220734 39978
rect 220802 39922 220858 39978
rect 220926 39922 220982 39978
rect 215210 22294 215266 22350
rect 215334 22294 215390 22350
rect 215210 22170 215266 22226
rect 215334 22170 215390 22226
rect 215210 22046 215266 22102
rect 215334 22046 215390 22102
rect 215210 21922 215266 21978
rect 215334 21922 215390 21978
rect 220554 22294 220610 22350
rect 220678 22294 220734 22350
rect 220802 22294 220858 22350
rect 220926 22294 220982 22350
rect 220554 22170 220610 22226
rect 220678 22170 220734 22226
rect 220802 22170 220858 22226
rect 220926 22170 220982 22226
rect 220554 22046 220610 22102
rect 220678 22046 220734 22102
rect 220802 22046 220858 22102
rect 220926 22046 220982 22102
rect 220554 21922 220610 21978
rect 220678 21922 220734 21978
rect 220802 21922 220858 21978
rect 220926 21922 220982 21978
rect 193554 10294 193610 10350
rect 193678 10294 193734 10350
rect 193802 10294 193858 10350
rect 193926 10294 193982 10350
rect 193554 10170 193610 10226
rect 193678 10170 193734 10226
rect 193802 10170 193858 10226
rect 193926 10170 193982 10226
rect 193554 10046 193610 10102
rect 193678 10046 193734 10102
rect 193802 10046 193858 10102
rect 193926 10046 193982 10102
rect 193554 9922 193610 9978
rect 193678 9922 193734 9978
rect 193802 9922 193858 9978
rect 193926 9922 193982 9978
rect 193554 -1176 193610 -1120
rect 193678 -1176 193734 -1120
rect 193802 -1176 193858 -1120
rect 193926 -1176 193982 -1120
rect 193554 -1300 193610 -1244
rect 193678 -1300 193734 -1244
rect 193802 -1300 193858 -1244
rect 193926 -1300 193982 -1244
rect 193554 -1424 193610 -1368
rect 193678 -1424 193734 -1368
rect 193802 -1424 193858 -1368
rect 193926 -1424 193982 -1368
rect 193554 -1548 193610 -1492
rect 193678 -1548 193734 -1492
rect 193802 -1548 193858 -1492
rect 193926 -1548 193982 -1492
rect 220554 4294 220610 4350
rect 220678 4294 220734 4350
rect 220802 4294 220858 4350
rect 220926 4294 220982 4350
rect 220554 4170 220610 4226
rect 220678 4170 220734 4226
rect 220802 4170 220858 4226
rect 220926 4170 220982 4226
rect 220554 4046 220610 4102
rect 220678 4046 220734 4102
rect 220802 4046 220858 4102
rect 220926 4046 220982 4102
rect 220554 3922 220610 3978
rect 220678 3922 220734 3978
rect 220802 3922 220858 3978
rect 220926 3922 220982 3978
rect 220554 -216 220610 -160
rect 220678 -216 220734 -160
rect 220802 -216 220858 -160
rect 220926 -216 220982 -160
rect 220554 -340 220610 -284
rect 220678 -340 220734 -284
rect 220802 -340 220858 -284
rect 220926 -340 220982 -284
rect 220554 -464 220610 -408
rect 220678 -464 220734 -408
rect 220802 -464 220858 -408
rect 220926 -464 220982 -408
rect 220554 -588 220610 -532
rect 220678 -588 220734 -532
rect 220802 -588 220858 -532
rect 220926 -588 220982 -532
rect 224274 46294 224330 46350
rect 224398 46294 224454 46350
rect 224522 46294 224578 46350
rect 224646 46294 224702 46350
rect 224274 46170 224330 46226
rect 224398 46170 224454 46226
rect 224522 46170 224578 46226
rect 224646 46170 224702 46226
rect 224274 46046 224330 46102
rect 224398 46046 224454 46102
rect 224522 46046 224578 46102
rect 224646 46046 224702 46102
rect 224274 45922 224330 45978
rect 224398 45922 224454 45978
rect 224522 45922 224578 45978
rect 224646 45922 224702 45978
rect 224274 28294 224330 28350
rect 224398 28294 224454 28350
rect 224522 28294 224578 28350
rect 224646 28294 224702 28350
rect 224274 28170 224330 28226
rect 224398 28170 224454 28226
rect 224522 28170 224578 28226
rect 224646 28170 224702 28226
rect 224274 28046 224330 28102
rect 224398 28046 224454 28102
rect 224522 28046 224578 28102
rect 224646 28046 224702 28102
rect 224274 27922 224330 27978
rect 224398 27922 224454 27978
rect 224522 27922 224578 27978
rect 224646 27922 224702 27978
rect 224274 10294 224330 10350
rect 224398 10294 224454 10350
rect 224522 10294 224578 10350
rect 224646 10294 224702 10350
rect 224274 10170 224330 10226
rect 224398 10170 224454 10226
rect 224522 10170 224578 10226
rect 224646 10170 224702 10226
rect 224274 10046 224330 10102
rect 224398 10046 224454 10102
rect 224522 10046 224578 10102
rect 224646 10046 224702 10102
rect 224274 9922 224330 9978
rect 224398 9922 224454 9978
rect 224522 9922 224578 9978
rect 224646 9922 224702 9978
rect 224274 -1176 224330 -1120
rect 224398 -1176 224454 -1120
rect 224522 -1176 224578 -1120
rect 224646 -1176 224702 -1120
rect 224274 -1300 224330 -1244
rect 224398 -1300 224454 -1244
rect 224522 -1300 224578 -1244
rect 224646 -1300 224702 -1244
rect 224274 -1424 224330 -1368
rect 224398 -1424 224454 -1368
rect 224522 -1424 224578 -1368
rect 224646 -1424 224702 -1368
rect 224274 -1548 224330 -1492
rect 224398 -1548 224454 -1492
rect 224522 -1548 224578 -1492
rect 224646 -1548 224702 -1492
rect 251274 40294 251330 40350
rect 251398 40294 251454 40350
rect 251522 40294 251578 40350
rect 251646 40294 251702 40350
rect 251274 40170 251330 40226
rect 251398 40170 251454 40226
rect 251522 40170 251578 40226
rect 251646 40170 251702 40226
rect 251274 40046 251330 40102
rect 251398 40046 251454 40102
rect 251522 40046 251578 40102
rect 251646 40046 251702 40102
rect 251274 39922 251330 39978
rect 251398 39922 251454 39978
rect 251522 39922 251578 39978
rect 251646 39922 251702 39978
rect 251274 22294 251330 22350
rect 251398 22294 251454 22350
rect 251522 22294 251578 22350
rect 251646 22294 251702 22350
rect 251274 22170 251330 22226
rect 251398 22170 251454 22226
rect 251522 22170 251578 22226
rect 251646 22170 251702 22226
rect 251274 22046 251330 22102
rect 251398 22046 251454 22102
rect 251522 22046 251578 22102
rect 251646 22046 251702 22102
rect 251274 21922 251330 21978
rect 251398 21922 251454 21978
rect 251522 21922 251578 21978
rect 251646 21922 251702 21978
rect 251274 4294 251330 4350
rect 251398 4294 251454 4350
rect 251522 4294 251578 4350
rect 251646 4294 251702 4350
rect 251274 4170 251330 4226
rect 251398 4170 251454 4226
rect 251522 4170 251578 4226
rect 251646 4170 251702 4226
rect 251274 4046 251330 4102
rect 251398 4046 251454 4102
rect 251522 4046 251578 4102
rect 251646 4046 251702 4102
rect 251274 3922 251330 3978
rect 251398 3922 251454 3978
rect 251522 3922 251578 3978
rect 251646 3922 251702 3978
rect 251274 -216 251330 -160
rect 251398 -216 251454 -160
rect 251522 -216 251578 -160
rect 251646 -216 251702 -160
rect 251274 -340 251330 -284
rect 251398 -340 251454 -284
rect 251522 -340 251578 -284
rect 251646 -340 251702 -284
rect 251274 -464 251330 -408
rect 251398 -464 251454 -408
rect 251522 -464 251578 -408
rect 251646 -464 251702 -408
rect 251274 -588 251330 -532
rect 251398 -588 251454 -532
rect 251522 -588 251578 -532
rect 251646 -588 251702 -532
rect 254994 46294 255050 46350
rect 255118 46294 255174 46350
rect 255242 46294 255298 46350
rect 255366 46294 255422 46350
rect 254994 46170 255050 46226
rect 255118 46170 255174 46226
rect 255242 46170 255298 46226
rect 255366 46170 255422 46226
rect 254994 46046 255050 46102
rect 255118 46046 255174 46102
rect 255242 46046 255298 46102
rect 255366 46046 255422 46102
rect 254994 45922 255050 45978
rect 255118 45922 255174 45978
rect 255242 45922 255298 45978
rect 255366 45922 255422 45978
rect 281994 40294 282050 40350
rect 282118 40294 282174 40350
rect 282242 40294 282298 40350
rect 282366 40294 282422 40350
rect 281994 40170 282050 40226
rect 282118 40170 282174 40226
rect 282242 40170 282298 40226
rect 282366 40170 282422 40226
rect 281994 40046 282050 40102
rect 282118 40046 282174 40102
rect 282242 40046 282298 40102
rect 282366 40046 282422 40102
rect 281994 39922 282050 39978
rect 282118 39922 282174 39978
rect 282242 39922 282298 39978
rect 282366 39922 282422 39978
rect 254994 28294 255050 28350
rect 255118 28294 255174 28350
rect 255242 28294 255298 28350
rect 255366 28294 255422 28350
rect 254994 28170 255050 28226
rect 255118 28170 255174 28226
rect 255242 28170 255298 28226
rect 255366 28170 255422 28226
rect 254994 28046 255050 28102
rect 255118 28046 255174 28102
rect 255242 28046 255298 28102
rect 255366 28046 255422 28102
rect 254994 27922 255050 27978
rect 255118 27922 255174 27978
rect 255242 27922 255298 27978
rect 255366 27922 255422 27978
rect 279862 28294 279918 28350
rect 279986 28294 280042 28350
rect 279862 28170 279918 28226
rect 279986 28170 280042 28226
rect 279862 28046 279918 28102
rect 279986 28046 280042 28102
rect 279862 27922 279918 27978
rect 279986 27922 280042 27978
rect 281994 22294 282050 22350
rect 282118 22294 282174 22350
rect 282242 22294 282298 22350
rect 282366 22294 282422 22350
rect 281994 22170 282050 22226
rect 282118 22170 282174 22226
rect 282242 22170 282298 22226
rect 282366 22170 282422 22226
rect 281994 22046 282050 22102
rect 282118 22046 282174 22102
rect 282242 22046 282298 22102
rect 282366 22046 282422 22102
rect 281994 21922 282050 21978
rect 282118 21922 282174 21978
rect 282242 21922 282298 21978
rect 282366 21922 282422 21978
rect 254994 10294 255050 10350
rect 255118 10294 255174 10350
rect 255242 10294 255298 10350
rect 255366 10294 255422 10350
rect 254994 10170 255050 10226
rect 255118 10170 255174 10226
rect 255242 10170 255298 10226
rect 255366 10170 255422 10226
rect 254994 10046 255050 10102
rect 255118 10046 255174 10102
rect 255242 10046 255298 10102
rect 255366 10046 255422 10102
rect 254994 9922 255050 9978
rect 255118 9922 255174 9978
rect 255242 9922 255298 9978
rect 255366 9922 255422 9978
rect 279862 10294 279918 10350
rect 279986 10294 280042 10350
rect 279862 10170 279918 10226
rect 279986 10170 280042 10226
rect 279862 10046 279918 10102
rect 279986 10046 280042 10102
rect 279862 9922 279918 9978
rect 279986 9922 280042 9978
rect 254994 -1176 255050 -1120
rect 255118 -1176 255174 -1120
rect 255242 -1176 255298 -1120
rect 255366 -1176 255422 -1120
rect 254994 -1300 255050 -1244
rect 255118 -1300 255174 -1244
rect 255242 -1300 255298 -1244
rect 255366 -1300 255422 -1244
rect 254994 -1424 255050 -1368
rect 255118 -1424 255174 -1368
rect 255242 -1424 255298 -1368
rect 255366 -1424 255422 -1368
rect 254994 -1548 255050 -1492
rect 255118 -1548 255174 -1492
rect 255242 -1548 255298 -1492
rect 255366 -1548 255422 -1492
rect 281994 4294 282050 4350
rect 282118 4294 282174 4350
rect 282242 4294 282298 4350
rect 282366 4294 282422 4350
rect 281994 4170 282050 4226
rect 282118 4170 282174 4226
rect 282242 4170 282298 4226
rect 282366 4170 282422 4226
rect 281994 4046 282050 4102
rect 282118 4046 282174 4102
rect 282242 4046 282298 4102
rect 282366 4046 282422 4102
rect 281994 3922 282050 3978
rect 282118 3922 282174 3978
rect 282242 3922 282298 3978
rect 282366 3922 282422 3978
rect 281994 -216 282050 -160
rect 282118 -216 282174 -160
rect 282242 -216 282298 -160
rect 282366 -216 282422 -160
rect 281994 -340 282050 -284
rect 282118 -340 282174 -284
rect 282242 -340 282298 -284
rect 282366 -340 282422 -284
rect 281994 -464 282050 -408
rect 282118 -464 282174 -408
rect 282242 -464 282298 -408
rect 282366 -464 282422 -408
rect 281994 -588 282050 -532
rect 282118 -588 282174 -532
rect 282242 -588 282298 -532
rect 282366 -588 282422 -532
rect 285714 46294 285770 46350
rect 285838 46294 285894 46350
rect 285962 46294 286018 46350
rect 286086 46294 286142 46350
rect 285714 46170 285770 46226
rect 285838 46170 285894 46226
rect 285962 46170 286018 46226
rect 286086 46170 286142 46226
rect 285714 46046 285770 46102
rect 285838 46046 285894 46102
rect 285962 46046 286018 46102
rect 286086 46046 286142 46102
rect 285714 45922 285770 45978
rect 285838 45922 285894 45978
rect 285962 45922 286018 45978
rect 286086 45922 286142 45978
rect 285714 28294 285770 28350
rect 285838 28294 285894 28350
rect 285962 28294 286018 28350
rect 286086 28294 286142 28350
rect 285714 28170 285770 28226
rect 285838 28170 285894 28226
rect 285962 28170 286018 28226
rect 286086 28170 286142 28226
rect 285714 28046 285770 28102
rect 285838 28046 285894 28102
rect 285962 28046 286018 28102
rect 286086 28046 286142 28102
rect 285714 27922 285770 27978
rect 285838 27922 285894 27978
rect 285962 27922 286018 27978
rect 286086 27922 286142 27978
rect 285714 10294 285770 10350
rect 285838 10294 285894 10350
rect 285962 10294 286018 10350
rect 286086 10294 286142 10350
rect 285714 10170 285770 10226
rect 285838 10170 285894 10226
rect 285962 10170 286018 10226
rect 286086 10170 286142 10226
rect 285714 10046 285770 10102
rect 285838 10046 285894 10102
rect 285962 10046 286018 10102
rect 286086 10046 286142 10102
rect 285714 9922 285770 9978
rect 285838 9922 285894 9978
rect 285962 9922 286018 9978
rect 286086 9922 286142 9978
rect 285714 -1176 285770 -1120
rect 285838 -1176 285894 -1120
rect 285962 -1176 286018 -1120
rect 286086 -1176 286142 -1120
rect 285714 -1300 285770 -1244
rect 285838 -1300 285894 -1244
rect 285962 -1300 286018 -1244
rect 286086 -1300 286142 -1244
rect 285714 -1424 285770 -1368
rect 285838 -1424 285894 -1368
rect 285962 -1424 286018 -1368
rect 286086 -1424 286142 -1368
rect 285714 -1548 285770 -1492
rect 285838 -1548 285894 -1492
rect 285962 -1548 286018 -1492
rect 286086 -1548 286142 -1492
rect 312714 40294 312770 40350
rect 312838 40294 312894 40350
rect 312962 40294 313018 40350
rect 313086 40294 313142 40350
rect 312714 40170 312770 40226
rect 312838 40170 312894 40226
rect 312962 40170 313018 40226
rect 313086 40170 313142 40226
rect 312714 40046 312770 40102
rect 312838 40046 312894 40102
rect 312962 40046 313018 40102
rect 313086 40046 313142 40102
rect 312714 39922 312770 39978
rect 312838 39922 312894 39978
rect 312962 39922 313018 39978
rect 313086 39922 313142 39978
rect 312714 22294 312770 22350
rect 312838 22294 312894 22350
rect 312962 22294 313018 22350
rect 313086 22294 313142 22350
rect 312714 22170 312770 22226
rect 312838 22170 312894 22226
rect 312962 22170 313018 22226
rect 313086 22170 313142 22226
rect 312714 22046 312770 22102
rect 312838 22046 312894 22102
rect 312962 22046 313018 22102
rect 313086 22046 313142 22102
rect 312714 21922 312770 21978
rect 312838 21922 312894 21978
rect 312962 21922 313018 21978
rect 313086 21922 313142 21978
rect 312714 4294 312770 4350
rect 312838 4294 312894 4350
rect 312962 4294 313018 4350
rect 313086 4294 313142 4350
rect 312714 4170 312770 4226
rect 312838 4170 312894 4226
rect 312962 4170 313018 4226
rect 313086 4170 313142 4226
rect 312714 4046 312770 4102
rect 312838 4046 312894 4102
rect 312962 4046 313018 4102
rect 313086 4046 313142 4102
rect 312714 3922 312770 3978
rect 312838 3922 312894 3978
rect 312962 3922 313018 3978
rect 313086 3922 313142 3978
rect 312714 -216 312770 -160
rect 312838 -216 312894 -160
rect 312962 -216 313018 -160
rect 313086 -216 313142 -160
rect 312714 -340 312770 -284
rect 312838 -340 312894 -284
rect 312962 -340 313018 -284
rect 313086 -340 313142 -284
rect 312714 -464 312770 -408
rect 312838 -464 312894 -408
rect 312962 -464 313018 -408
rect 313086 -464 313142 -408
rect 312714 -588 312770 -532
rect 312838 -588 312894 -532
rect 312962 -588 313018 -532
rect 313086 -588 313142 -532
rect 316434 46294 316490 46350
rect 316558 46294 316614 46350
rect 316682 46294 316738 46350
rect 316806 46294 316862 46350
rect 316434 46170 316490 46226
rect 316558 46170 316614 46226
rect 316682 46170 316738 46226
rect 316806 46170 316862 46226
rect 316434 46046 316490 46102
rect 316558 46046 316614 46102
rect 316682 46046 316738 46102
rect 316806 46046 316862 46102
rect 316434 45922 316490 45978
rect 316558 45922 316614 45978
rect 316682 45922 316738 45978
rect 316806 45922 316862 45978
rect 316434 28294 316490 28350
rect 316558 28294 316614 28350
rect 316682 28294 316738 28350
rect 316806 28294 316862 28350
rect 316434 28170 316490 28226
rect 316558 28170 316614 28226
rect 316682 28170 316738 28226
rect 316806 28170 316862 28226
rect 316434 28046 316490 28102
rect 316558 28046 316614 28102
rect 316682 28046 316738 28102
rect 316806 28046 316862 28102
rect 316434 27922 316490 27978
rect 316558 27922 316614 27978
rect 316682 27922 316738 27978
rect 316806 27922 316862 27978
rect 316434 10294 316490 10350
rect 316558 10294 316614 10350
rect 316682 10294 316738 10350
rect 316806 10294 316862 10350
rect 316434 10170 316490 10226
rect 316558 10170 316614 10226
rect 316682 10170 316738 10226
rect 316806 10170 316862 10226
rect 316434 10046 316490 10102
rect 316558 10046 316614 10102
rect 316682 10046 316738 10102
rect 316806 10046 316862 10102
rect 316434 9922 316490 9978
rect 316558 9922 316614 9978
rect 316682 9922 316738 9978
rect 316806 9922 316862 9978
rect 316434 -1176 316490 -1120
rect 316558 -1176 316614 -1120
rect 316682 -1176 316738 -1120
rect 316806 -1176 316862 -1120
rect 316434 -1300 316490 -1244
rect 316558 -1300 316614 -1244
rect 316682 -1300 316738 -1244
rect 316806 -1300 316862 -1244
rect 316434 -1424 316490 -1368
rect 316558 -1424 316614 -1368
rect 316682 -1424 316738 -1368
rect 316806 -1424 316862 -1368
rect 316434 -1548 316490 -1492
rect 316558 -1548 316614 -1492
rect 316682 -1548 316738 -1492
rect 316806 -1548 316862 -1492
rect 343434 40294 343490 40350
rect 343558 40294 343614 40350
rect 343682 40294 343738 40350
rect 343806 40294 343862 40350
rect 343434 40170 343490 40226
rect 343558 40170 343614 40226
rect 343682 40170 343738 40226
rect 343806 40170 343862 40226
rect 343434 40046 343490 40102
rect 343558 40046 343614 40102
rect 343682 40046 343738 40102
rect 343806 40046 343862 40102
rect 343434 39922 343490 39978
rect 343558 39922 343614 39978
rect 343682 39922 343738 39978
rect 343806 39922 343862 39978
rect 372428 210842 372484 210898
rect 374154 292294 374210 292350
rect 374278 292294 374334 292350
rect 374402 292294 374458 292350
rect 374526 292294 374582 292350
rect 374154 292170 374210 292226
rect 374278 292170 374334 292226
rect 374402 292170 374458 292226
rect 374526 292170 374582 292226
rect 374154 292046 374210 292102
rect 374278 292046 374334 292102
rect 374402 292046 374458 292102
rect 374526 292046 374582 292102
rect 374154 291922 374210 291978
rect 374278 291922 374334 291978
rect 374402 291922 374458 291978
rect 374526 291922 374582 291978
rect 374154 274294 374210 274350
rect 374278 274294 374334 274350
rect 374402 274294 374458 274350
rect 374526 274294 374582 274350
rect 374154 274170 374210 274226
rect 374278 274170 374334 274226
rect 374402 274170 374458 274226
rect 374526 274170 374582 274226
rect 374154 274046 374210 274102
rect 374278 274046 374334 274102
rect 374402 274046 374458 274102
rect 374526 274046 374582 274102
rect 374154 273922 374210 273978
rect 374278 273922 374334 273978
rect 374402 273922 374458 273978
rect 374526 273922 374582 273978
rect 374154 256294 374210 256350
rect 374278 256294 374334 256350
rect 374402 256294 374458 256350
rect 374526 256294 374582 256350
rect 374154 256170 374210 256226
rect 374278 256170 374334 256226
rect 374402 256170 374458 256226
rect 374526 256170 374582 256226
rect 374154 256046 374210 256102
rect 374278 256046 374334 256102
rect 374402 256046 374458 256102
rect 374526 256046 374582 256102
rect 374154 255922 374210 255978
rect 374278 255922 374334 255978
rect 374402 255922 374458 255978
rect 374526 255922 374582 255978
rect 372876 217502 372932 217558
rect 372764 209222 372820 209278
rect 374154 238294 374210 238350
rect 374278 238294 374334 238350
rect 374402 238294 374458 238350
rect 374526 238294 374582 238350
rect 374154 238170 374210 238226
rect 374278 238170 374334 238226
rect 374402 238170 374458 238226
rect 374526 238170 374582 238226
rect 374154 238046 374210 238102
rect 374278 238046 374334 238102
rect 374402 238046 374458 238102
rect 374526 238046 374582 238102
rect 374154 237922 374210 237978
rect 374278 237922 374334 237978
rect 374402 237922 374458 237978
rect 374526 237922 374582 237978
rect 374154 220294 374210 220350
rect 374278 220294 374334 220350
rect 374402 220294 374458 220350
rect 374526 220294 374582 220350
rect 374154 220170 374210 220226
rect 374278 220170 374334 220226
rect 374402 220170 374458 220226
rect 374526 220170 374582 220226
rect 374154 220046 374210 220102
rect 374278 220046 374334 220102
rect 374402 220046 374458 220102
rect 374526 220046 374582 220102
rect 374154 219922 374210 219978
rect 374278 219922 374334 219978
rect 374402 219922 374458 219978
rect 374526 219922 374582 219978
rect 373884 218428 373940 218458
rect 373884 218402 373940 218428
rect 373660 214262 373716 214318
rect 373772 216602 373828 216658
rect 373436 187802 373492 187858
rect 373884 213362 373940 213418
rect 373884 211922 373940 211978
rect 374154 202294 374210 202350
rect 374278 202294 374334 202350
rect 374402 202294 374458 202350
rect 374526 202294 374582 202350
rect 374154 202170 374210 202226
rect 374278 202170 374334 202226
rect 374402 202170 374458 202226
rect 374526 202170 374582 202226
rect 374154 202046 374210 202102
rect 374278 202046 374334 202102
rect 374402 202046 374458 202102
rect 374526 202046 374582 202102
rect 374154 201922 374210 201978
rect 374278 201922 374334 201978
rect 374402 201922 374458 201978
rect 374526 201922 374582 201978
rect 373884 184922 373940 184978
rect 374154 184294 374210 184350
rect 374278 184294 374334 184350
rect 374402 184294 374458 184350
rect 374526 184294 374582 184350
rect 374154 184170 374210 184226
rect 374278 184170 374334 184226
rect 374402 184170 374458 184226
rect 374526 184170 374582 184226
rect 374154 184046 374210 184102
rect 374278 184046 374334 184102
rect 374402 184046 374458 184102
rect 374526 184046 374582 184102
rect 374154 183922 374210 183978
rect 374278 183922 374334 183978
rect 374402 183922 374458 183978
rect 374526 183922 374582 183978
rect 375452 268802 375508 268858
rect 375004 213182 375060 213238
rect 375228 187982 375284 188038
rect 374154 166294 374210 166350
rect 374278 166294 374334 166350
rect 374402 166294 374458 166350
rect 374526 166294 374582 166350
rect 374154 166170 374210 166226
rect 374278 166170 374334 166226
rect 374402 166170 374458 166226
rect 374526 166170 374582 166226
rect 374154 166046 374210 166102
rect 374278 166046 374334 166102
rect 374402 166046 374458 166102
rect 374526 166046 374582 166102
rect 374154 165922 374210 165978
rect 374278 165922 374334 165978
rect 374402 165922 374458 165978
rect 374526 165922 374582 165978
rect 374154 148294 374210 148350
rect 374278 148294 374334 148350
rect 374402 148294 374458 148350
rect 374526 148294 374582 148350
rect 374154 148170 374210 148226
rect 374278 148170 374334 148226
rect 374402 148170 374458 148226
rect 374526 148170 374582 148226
rect 374154 148046 374210 148102
rect 374278 148046 374334 148102
rect 374402 148046 374458 148102
rect 374526 148046 374582 148102
rect 374154 147922 374210 147978
rect 374278 147922 374334 147978
rect 374402 147922 374458 147978
rect 374526 147922 374582 147978
rect 375340 133442 375396 133498
rect 374154 130294 374210 130350
rect 374278 130294 374334 130350
rect 374402 130294 374458 130350
rect 374526 130294 374582 130350
rect 374154 130170 374210 130226
rect 374278 130170 374334 130226
rect 374402 130170 374458 130226
rect 374526 130170 374582 130226
rect 374154 130046 374210 130102
rect 374278 130046 374334 130102
rect 374402 130046 374458 130102
rect 374526 130046 374582 130102
rect 374154 129922 374210 129978
rect 374278 129922 374334 129978
rect 374402 129922 374458 129978
rect 374526 129922 374582 129978
rect 373884 120842 373940 120898
rect 374154 112294 374210 112350
rect 374278 112294 374334 112350
rect 374402 112294 374458 112350
rect 374526 112294 374582 112350
rect 374154 112170 374210 112226
rect 374278 112170 374334 112226
rect 374402 112170 374458 112226
rect 374526 112170 374582 112226
rect 374154 112046 374210 112102
rect 374278 112046 374334 112102
rect 374402 112046 374458 112102
rect 374526 112046 374582 112102
rect 374154 111922 374210 111978
rect 374278 111922 374334 111978
rect 374402 111922 374458 111978
rect 374526 111922 374582 111978
rect 374154 94294 374210 94350
rect 374278 94294 374334 94350
rect 374402 94294 374458 94350
rect 374526 94294 374582 94350
rect 374154 94170 374210 94226
rect 374278 94170 374334 94226
rect 374402 94170 374458 94226
rect 374526 94170 374582 94226
rect 374154 94046 374210 94102
rect 374278 94046 374334 94102
rect 374402 94046 374458 94102
rect 374526 94046 374582 94102
rect 374154 93922 374210 93978
rect 374278 93922 374334 93978
rect 374402 93922 374458 93978
rect 374526 93922 374582 93978
rect 374154 76294 374210 76350
rect 374278 76294 374334 76350
rect 374402 76294 374458 76350
rect 374526 76294 374582 76350
rect 374154 76170 374210 76226
rect 374278 76170 374334 76226
rect 374402 76170 374458 76226
rect 374526 76170 374582 76226
rect 374154 76046 374210 76102
rect 374278 76046 374334 76102
rect 374402 76046 374458 76102
rect 374526 76046 374582 76102
rect 374154 75922 374210 75978
rect 374278 75922 374334 75978
rect 374402 75922 374458 75978
rect 374526 75922 374582 75978
rect 374154 58294 374210 58350
rect 374278 58294 374334 58350
rect 374402 58294 374458 58350
rect 374526 58294 374582 58350
rect 374154 58170 374210 58226
rect 374278 58170 374334 58226
rect 374402 58170 374458 58226
rect 374526 58170 374582 58226
rect 374154 58046 374210 58102
rect 374278 58046 374334 58102
rect 374402 58046 374458 58102
rect 374526 58046 374582 58102
rect 374154 57922 374210 57978
rect 374278 57922 374334 57978
rect 374402 57922 374458 57978
rect 374526 57922 374582 57978
rect 347154 46294 347210 46350
rect 347278 46294 347334 46350
rect 347402 46294 347458 46350
rect 347526 46294 347582 46350
rect 347154 46170 347210 46226
rect 347278 46170 347334 46226
rect 347402 46170 347458 46226
rect 347526 46170 347582 46226
rect 347154 46046 347210 46102
rect 347278 46046 347334 46102
rect 347402 46046 347458 46102
rect 347526 46046 347582 46102
rect 347154 45922 347210 45978
rect 347278 45922 347334 45978
rect 347402 45922 347458 45978
rect 347526 45922 347582 45978
rect 347154 28294 347210 28350
rect 347278 28294 347334 28350
rect 347402 28294 347458 28350
rect 347526 28294 347582 28350
rect 347154 28170 347210 28226
rect 347278 28170 347334 28226
rect 347402 28170 347458 28226
rect 347526 28170 347582 28226
rect 347154 28046 347210 28102
rect 347278 28046 347334 28102
rect 347402 28046 347458 28102
rect 347526 28046 347582 28102
rect 347154 27922 347210 27978
rect 347278 27922 347334 27978
rect 347402 27922 347458 27978
rect 347526 27922 347582 27978
rect 343434 22294 343490 22350
rect 343558 22294 343614 22350
rect 343682 22294 343738 22350
rect 343806 22294 343862 22350
rect 343434 22170 343490 22226
rect 343558 22170 343614 22226
rect 343682 22170 343738 22226
rect 343806 22170 343862 22226
rect 343434 22046 343490 22102
rect 343558 22046 343614 22102
rect 343682 22046 343738 22102
rect 343806 22046 343862 22102
rect 343434 21922 343490 21978
rect 343558 21922 343614 21978
rect 343682 21922 343738 21978
rect 343806 21922 343862 21978
rect 344514 22294 344570 22350
rect 344638 22294 344694 22350
rect 344514 22170 344570 22226
rect 344638 22170 344694 22226
rect 344514 22046 344570 22102
rect 344638 22046 344694 22102
rect 344514 21922 344570 21978
rect 344638 21922 344694 21978
rect 343434 4294 343490 4350
rect 343558 4294 343614 4350
rect 343682 4294 343738 4350
rect 343806 4294 343862 4350
rect 343434 4170 343490 4226
rect 343558 4170 343614 4226
rect 343682 4170 343738 4226
rect 343806 4170 343862 4226
rect 343434 4046 343490 4102
rect 343558 4046 343614 4102
rect 343682 4046 343738 4102
rect 343806 4046 343862 4102
rect 343434 3922 343490 3978
rect 343558 3922 343614 3978
rect 343682 3922 343738 3978
rect 343806 3922 343862 3978
rect 343434 -216 343490 -160
rect 343558 -216 343614 -160
rect 343682 -216 343738 -160
rect 343806 -216 343862 -160
rect 343434 -340 343490 -284
rect 343558 -340 343614 -284
rect 343682 -340 343738 -284
rect 343806 -340 343862 -284
rect 343434 -464 343490 -408
rect 343558 -464 343614 -408
rect 343682 -464 343738 -408
rect 343806 -464 343862 -408
rect 343434 -588 343490 -532
rect 343558 -588 343614 -532
rect 343682 -588 343738 -532
rect 343806 -588 343862 -532
rect 347154 10294 347210 10350
rect 347278 10294 347334 10350
rect 347402 10294 347458 10350
rect 347526 10294 347582 10350
rect 347154 10170 347210 10226
rect 347278 10170 347334 10226
rect 347402 10170 347458 10226
rect 347526 10170 347582 10226
rect 347154 10046 347210 10102
rect 347278 10046 347334 10102
rect 347402 10046 347458 10102
rect 347526 10046 347582 10102
rect 347154 9922 347210 9978
rect 347278 9922 347334 9978
rect 347402 9922 347458 9978
rect 347526 9922 347582 9978
rect 347154 -1176 347210 -1120
rect 347278 -1176 347334 -1120
rect 347402 -1176 347458 -1120
rect 347526 -1176 347582 -1120
rect 347154 -1300 347210 -1244
rect 347278 -1300 347334 -1244
rect 347402 -1300 347458 -1244
rect 347526 -1300 347582 -1244
rect 347154 -1424 347210 -1368
rect 347278 -1424 347334 -1368
rect 347402 -1424 347458 -1368
rect 347526 -1424 347582 -1368
rect 347154 -1548 347210 -1492
rect 347278 -1548 347334 -1492
rect 347402 -1548 347458 -1492
rect 347526 -1548 347582 -1492
rect 375676 212102 375732 212158
rect 377132 260342 377188 260398
rect 377874 316294 377930 316350
rect 377998 316294 378054 316350
rect 378122 316294 378178 316350
rect 378246 316294 378302 316350
rect 377874 316170 377930 316226
rect 377998 316170 378054 316226
rect 378122 316170 378178 316226
rect 378246 316170 378302 316226
rect 377874 316046 377930 316102
rect 377998 316046 378054 316102
rect 378122 316046 378178 316102
rect 378246 316046 378302 316102
rect 377874 315922 377930 315978
rect 377998 315922 378054 315978
rect 378122 315922 378178 315978
rect 378246 315922 378302 315978
rect 377874 298294 377930 298350
rect 377998 298294 378054 298350
rect 378122 298294 378178 298350
rect 378246 298294 378302 298350
rect 377874 298170 377930 298226
rect 377998 298170 378054 298226
rect 378122 298170 378178 298226
rect 378246 298170 378302 298226
rect 377874 298046 377930 298102
rect 377998 298046 378054 298102
rect 378122 298046 378178 298102
rect 378246 298046 378302 298102
rect 377874 297922 377930 297978
rect 377998 297922 378054 297978
rect 378122 297922 378178 297978
rect 378246 297922 378302 297978
rect 377874 280294 377930 280350
rect 377998 280294 378054 280350
rect 378122 280294 378178 280350
rect 378246 280294 378302 280350
rect 377874 280170 377930 280226
rect 377998 280170 378054 280226
rect 378122 280170 378178 280226
rect 378246 280170 378302 280226
rect 377874 280046 377930 280102
rect 377998 280046 378054 280102
rect 378122 280046 378178 280102
rect 378246 280046 378302 280102
rect 377874 279922 377930 279978
rect 377998 279922 378054 279978
rect 378122 279922 378178 279978
rect 378246 279922 378302 279978
rect 377874 262294 377930 262350
rect 377998 262294 378054 262350
rect 378122 262294 378178 262350
rect 378246 262294 378302 262350
rect 377874 262170 377930 262226
rect 377998 262170 378054 262226
rect 378122 262170 378178 262226
rect 378246 262170 378302 262226
rect 377874 262046 377930 262102
rect 377998 262046 378054 262102
rect 378122 262046 378178 262102
rect 378246 262046 378302 262102
rect 377874 261922 377930 261978
rect 377998 261922 378054 261978
rect 378122 261922 378178 261978
rect 378246 261922 378302 261978
rect 377580 261602 377636 261658
rect 377874 244294 377930 244350
rect 377998 244294 378054 244350
rect 378122 244294 378178 244350
rect 378246 244294 378302 244350
rect 377874 244170 377930 244226
rect 377998 244170 378054 244226
rect 378122 244170 378178 244226
rect 378246 244170 378302 244226
rect 377874 244046 377930 244102
rect 377998 244046 378054 244102
rect 378122 244046 378178 244102
rect 378246 244046 378302 244102
rect 377874 243922 377930 243978
rect 377998 243922 378054 243978
rect 378122 243922 378178 243978
rect 378246 243922 378302 243978
rect 376124 216962 376180 217018
rect 376124 105722 376180 105778
rect 376124 91502 376180 91558
rect 377356 156302 377412 156358
rect 376908 133622 376964 133678
rect 378812 267182 378868 267238
rect 377874 226294 377930 226350
rect 377998 226294 378054 226350
rect 378122 226294 378178 226350
rect 378246 226294 378302 226350
rect 377874 226170 377930 226226
rect 377998 226170 378054 226226
rect 378122 226170 378178 226226
rect 378246 226170 378302 226226
rect 377874 226046 377930 226102
rect 377998 226046 378054 226102
rect 378122 226046 378178 226102
rect 378246 226046 378302 226102
rect 377874 225922 377930 225978
rect 377998 225922 378054 225978
rect 378122 225922 378178 225978
rect 378246 225922 378302 225978
rect 377874 208294 377930 208350
rect 377998 208294 378054 208350
rect 378122 208294 378178 208350
rect 378246 208294 378302 208350
rect 377874 208170 377930 208226
rect 377998 208170 378054 208226
rect 378122 208170 378178 208226
rect 378246 208170 378302 208226
rect 377874 208046 377930 208102
rect 377998 208046 378054 208102
rect 378122 208046 378178 208102
rect 378246 208046 378302 208102
rect 377874 207922 377930 207978
rect 377998 207922 378054 207978
rect 378122 207922 378178 207978
rect 378246 207922 378302 207978
rect 377874 190294 377930 190350
rect 377998 190294 378054 190350
rect 378122 190294 378178 190350
rect 378246 190294 378302 190350
rect 377874 190170 377930 190226
rect 377998 190170 378054 190226
rect 378122 190170 378178 190226
rect 378246 190170 378302 190226
rect 377874 190046 377930 190102
rect 377998 190046 378054 190102
rect 378122 190046 378178 190102
rect 378246 190046 378302 190102
rect 377874 189922 377930 189978
rect 377998 189922 378054 189978
rect 378122 189922 378178 189978
rect 378246 189922 378302 189978
rect 377874 172294 377930 172350
rect 377998 172294 378054 172350
rect 378122 172294 378178 172350
rect 378246 172294 378302 172350
rect 377874 172170 377930 172226
rect 377998 172170 378054 172226
rect 378122 172170 378178 172226
rect 378246 172170 378302 172226
rect 377874 172046 377930 172102
rect 377998 172046 378054 172102
rect 378122 172046 378178 172102
rect 378246 172046 378302 172102
rect 377874 171922 377930 171978
rect 377998 171922 378054 171978
rect 378122 171922 378178 171978
rect 378246 171922 378302 171978
rect 377874 154294 377930 154350
rect 377998 154294 378054 154350
rect 378122 154294 378178 154350
rect 378246 154294 378302 154350
rect 377874 154170 377930 154226
rect 377998 154170 378054 154226
rect 378122 154170 378178 154226
rect 378246 154170 378302 154226
rect 377874 154046 377930 154102
rect 377998 154046 378054 154102
rect 378122 154046 378178 154102
rect 378246 154046 378302 154102
rect 377874 153922 377930 153978
rect 377998 153922 378054 153978
rect 378122 153922 378178 153978
rect 378246 153922 378302 153978
rect 377874 136294 377930 136350
rect 377998 136294 378054 136350
rect 378122 136294 378178 136350
rect 378246 136294 378302 136350
rect 377874 136170 377930 136226
rect 377998 136170 378054 136226
rect 378122 136170 378178 136226
rect 378246 136170 378302 136226
rect 377874 136046 377930 136102
rect 377998 136046 378054 136102
rect 378122 136046 378178 136102
rect 378246 136046 378302 136102
rect 377874 135922 377930 135978
rect 377998 135922 378054 135978
rect 378122 135922 378178 135978
rect 378246 135922 378302 135978
rect 378700 214082 378756 214138
rect 379260 215572 379316 215578
rect 379260 215522 379316 215572
rect 378924 211022 378980 211078
rect 379484 264482 379540 264538
rect 379596 261242 379652 261298
rect 379484 217142 379540 217198
rect 379484 216422 379540 216478
rect 379484 215342 379540 215398
rect 377874 118294 377930 118350
rect 377998 118294 378054 118350
rect 378122 118294 378178 118350
rect 378246 118294 378302 118350
rect 377874 118170 377930 118226
rect 377998 118170 378054 118226
rect 378122 118170 378178 118226
rect 378246 118170 378302 118226
rect 377874 118046 377930 118102
rect 377998 118046 378054 118102
rect 378122 118046 378178 118102
rect 378246 118046 378302 118102
rect 377874 117922 377930 117978
rect 377998 117922 378054 117978
rect 378122 117922 378178 117978
rect 378246 117922 378302 117978
rect 377580 101582 377636 101638
rect 377874 100294 377930 100350
rect 377998 100294 378054 100350
rect 378122 100294 378178 100350
rect 378246 100294 378302 100350
rect 377874 100170 377930 100226
rect 377998 100170 378054 100226
rect 378122 100170 378178 100226
rect 378246 100170 378302 100226
rect 377874 100046 377930 100102
rect 377998 100046 378054 100102
rect 378122 100046 378178 100102
rect 378246 100046 378302 100102
rect 377874 99922 377930 99978
rect 377998 99922 378054 99978
rect 378122 99922 378178 99978
rect 378246 99922 378302 99978
rect 377874 82294 377930 82350
rect 377998 82294 378054 82350
rect 378122 82294 378178 82350
rect 378246 82294 378302 82350
rect 377874 82170 377930 82226
rect 377998 82170 378054 82226
rect 378122 82170 378178 82226
rect 378246 82170 378302 82226
rect 377874 82046 377930 82102
rect 377998 82046 378054 82102
rect 378122 82046 378178 82102
rect 378246 82046 378302 82102
rect 377874 81922 377930 81978
rect 377998 81922 378054 81978
rect 378122 81922 378178 81978
rect 378246 81922 378302 81978
rect 377580 71342 377636 71398
rect 377580 64862 377636 64918
rect 377580 64682 377636 64738
rect 378588 74222 378644 74278
rect 377874 64294 377930 64350
rect 377998 64294 378054 64350
rect 378122 64294 378178 64350
rect 378246 64294 378302 64350
rect 377874 64170 377930 64226
rect 377998 64170 378054 64226
rect 378122 64170 378178 64226
rect 378246 64170 378302 64226
rect 377874 64046 377930 64102
rect 377998 64046 378054 64102
rect 378122 64046 378178 64102
rect 378246 64046 378302 64102
rect 377874 63922 377930 63978
rect 377998 63922 378054 63978
rect 378122 63922 378178 63978
rect 378246 63922 378302 63978
rect 377580 62882 377636 62938
rect 376236 52108 376292 52138
rect 376236 52082 376292 52108
rect 374154 40294 374210 40350
rect 374278 40294 374334 40350
rect 374402 40294 374458 40350
rect 374526 40294 374582 40350
rect 374154 40170 374210 40226
rect 374278 40170 374334 40226
rect 374402 40170 374458 40226
rect 374526 40170 374582 40226
rect 374154 40046 374210 40102
rect 374278 40046 374334 40102
rect 374402 40046 374458 40102
rect 374526 40046 374582 40102
rect 374154 39922 374210 39978
rect 374278 39922 374334 39978
rect 374402 39922 374458 39978
rect 374526 39922 374582 39978
rect 374154 22294 374210 22350
rect 374278 22294 374334 22350
rect 374402 22294 374458 22350
rect 374526 22294 374582 22350
rect 374154 22170 374210 22226
rect 374278 22170 374334 22226
rect 374402 22170 374458 22226
rect 374526 22170 374582 22226
rect 374154 22046 374210 22102
rect 374278 22046 374334 22102
rect 374402 22046 374458 22102
rect 374526 22046 374582 22102
rect 374154 21922 374210 21978
rect 374278 21922 374334 21978
rect 374402 21922 374458 21978
rect 374526 21922 374582 21978
rect 374154 4294 374210 4350
rect 374278 4294 374334 4350
rect 374402 4294 374458 4350
rect 374526 4294 374582 4350
rect 374154 4170 374210 4226
rect 374278 4170 374334 4226
rect 374402 4170 374458 4226
rect 374526 4170 374582 4226
rect 374154 4046 374210 4102
rect 374278 4046 374334 4102
rect 374402 4046 374458 4102
rect 374526 4046 374582 4102
rect 374154 3922 374210 3978
rect 374278 3922 374334 3978
rect 374402 3922 374458 3978
rect 374526 3922 374582 3978
rect 374154 -216 374210 -160
rect 374278 -216 374334 -160
rect 374402 -216 374458 -160
rect 374526 -216 374582 -160
rect 374154 -340 374210 -284
rect 374278 -340 374334 -284
rect 374402 -340 374458 -284
rect 374526 -340 374582 -284
rect 374154 -464 374210 -408
rect 374278 -464 374334 -408
rect 374402 -464 374458 -408
rect 374526 -464 374582 -408
rect 374154 -588 374210 -532
rect 374278 -588 374334 -532
rect 374402 -588 374458 -532
rect 374526 -588 374582 -532
rect 377874 46294 377930 46350
rect 377998 46294 378054 46350
rect 378122 46294 378178 46350
rect 378246 46294 378302 46350
rect 377874 46170 377930 46226
rect 377998 46170 378054 46226
rect 378122 46170 378178 46226
rect 378246 46170 378302 46226
rect 377874 46046 377930 46102
rect 377998 46046 378054 46102
rect 378122 46046 378178 46102
rect 378246 46046 378302 46102
rect 377874 45922 377930 45978
rect 377998 45922 378054 45978
rect 378122 45922 378178 45978
rect 378246 45922 378302 45978
rect 379372 182222 379428 182278
rect 379932 268082 379988 268138
rect 379820 267902 379876 267958
rect 379708 217682 379764 217738
rect 379708 212462 379764 212518
rect 380044 241802 380100 241858
rect 379596 151082 379652 151138
rect 378812 81602 378868 81658
rect 378812 80702 378868 80758
rect 378812 80522 378868 80578
rect 378812 78362 378868 78418
rect 378812 78002 378868 78058
rect 378812 72828 378868 72838
rect 378812 72782 378868 72828
rect 379596 115802 379652 115858
rect 379596 76562 379652 76618
rect 379596 74042 379652 74098
rect 379708 43622 379764 43678
rect 384518 310294 384574 310350
rect 384642 310294 384698 310350
rect 384518 310170 384574 310226
rect 384642 310170 384698 310226
rect 384518 310046 384574 310102
rect 384642 310046 384698 310102
rect 384518 309922 384574 309978
rect 384642 309922 384698 309978
rect 384518 292294 384574 292350
rect 384642 292294 384698 292350
rect 384518 292170 384574 292226
rect 384642 292170 384698 292226
rect 384518 292046 384574 292102
rect 384642 292046 384698 292102
rect 384518 291922 384574 291978
rect 384642 291922 384698 291978
rect 380380 216782 380436 216838
rect 380268 215162 380324 215218
rect 380380 216468 380436 216478
rect 380380 216422 380436 216468
rect 380268 213542 380324 213598
rect 380268 211742 380324 211798
rect 380268 209222 380324 209278
rect 380716 286082 380772 286138
rect 404874 364294 404930 364350
rect 404998 364294 405054 364350
rect 405122 364294 405178 364350
rect 405246 364294 405302 364350
rect 404874 364170 404930 364226
rect 404998 364170 405054 364226
rect 405122 364170 405178 364226
rect 405246 364170 405302 364226
rect 404874 364046 404930 364102
rect 404998 364046 405054 364102
rect 405122 364046 405178 364102
rect 405246 364046 405302 364102
rect 404874 363922 404930 363978
rect 404998 363922 405054 363978
rect 405122 363922 405178 363978
rect 405246 363922 405302 363978
rect 404874 346294 404930 346350
rect 404998 346294 405054 346350
rect 405122 346294 405178 346350
rect 405246 346294 405302 346350
rect 404874 346170 404930 346226
rect 404998 346170 405054 346226
rect 405122 346170 405178 346226
rect 405246 346170 405302 346226
rect 404874 346046 404930 346102
rect 404998 346046 405054 346102
rect 405122 346046 405178 346102
rect 405246 346046 405302 346102
rect 404874 345922 404930 345978
rect 404998 345922 405054 345978
rect 405122 345922 405178 345978
rect 405246 345922 405302 345978
rect 404874 328294 404930 328350
rect 404998 328294 405054 328350
rect 405122 328294 405178 328350
rect 405246 328294 405302 328350
rect 404874 328170 404930 328226
rect 404998 328170 405054 328226
rect 405122 328170 405178 328226
rect 405246 328170 405302 328226
rect 404874 328046 404930 328102
rect 404998 328046 405054 328102
rect 405122 328046 405178 328102
rect 405246 328046 405302 328102
rect 404874 327922 404930 327978
rect 404998 327922 405054 327978
rect 405122 327922 405178 327978
rect 405246 327922 405302 327978
rect 399878 316294 399934 316350
rect 400002 316294 400058 316350
rect 399878 316170 399934 316226
rect 400002 316170 400058 316226
rect 399878 316046 399934 316102
rect 400002 316046 400058 316102
rect 399878 315922 399934 315978
rect 400002 315922 400058 315978
rect 408594 598116 408650 598172
rect 408718 598116 408774 598172
rect 408842 598116 408898 598172
rect 408966 598116 409022 598172
rect 408594 597992 408650 598048
rect 408718 597992 408774 598048
rect 408842 597992 408898 598048
rect 408966 597992 409022 598048
rect 408594 597868 408650 597924
rect 408718 597868 408774 597924
rect 408842 597868 408898 597924
rect 408966 597868 409022 597924
rect 408594 597744 408650 597800
rect 408718 597744 408774 597800
rect 408842 597744 408898 597800
rect 408966 597744 409022 597800
rect 408594 586294 408650 586350
rect 408718 586294 408774 586350
rect 408842 586294 408898 586350
rect 408966 586294 409022 586350
rect 408594 586170 408650 586226
rect 408718 586170 408774 586226
rect 408842 586170 408898 586226
rect 408966 586170 409022 586226
rect 408594 586046 408650 586102
rect 408718 586046 408774 586102
rect 408842 586046 408898 586102
rect 408966 586046 409022 586102
rect 408594 585922 408650 585978
rect 408718 585922 408774 585978
rect 408842 585922 408898 585978
rect 408966 585922 409022 585978
rect 408594 568294 408650 568350
rect 408718 568294 408774 568350
rect 408842 568294 408898 568350
rect 408966 568294 409022 568350
rect 408594 568170 408650 568226
rect 408718 568170 408774 568226
rect 408842 568170 408898 568226
rect 408966 568170 409022 568226
rect 408594 568046 408650 568102
rect 408718 568046 408774 568102
rect 408842 568046 408898 568102
rect 408966 568046 409022 568102
rect 408594 567922 408650 567978
rect 408718 567922 408774 567978
rect 408842 567922 408898 567978
rect 408966 567922 409022 567978
rect 408594 550294 408650 550350
rect 408718 550294 408774 550350
rect 408842 550294 408898 550350
rect 408966 550294 409022 550350
rect 408594 550170 408650 550226
rect 408718 550170 408774 550226
rect 408842 550170 408898 550226
rect 408966 550170 409022 550226
rect 408594 550046 408650 550102
rect 408718 550046 408774 550102
rect 408842 550046 408898 550102
rect 408966 550046 409022 550102
rect 408594 549922 408650 549978
rect 408718 549922 408774 549978
rect 408842 549922 408898 549978
rect 408966 549922 409022 549978
rect 408594 532294 408650 532350
rect 408718 532294 408774 532350
rect 408842 532294 408898 532350
rect 408966 532294 409022 532350
rect 408594 532170 408650 532226
rect 408718 532170 408774 532226
rect 408842 532170 408898 532226
rect 408966 532170 409022 532226
rect 408594 532046 408650 532102
rect 408718 532046 408774 532102
rect 408842 532046 408898 532102
rect 408966 532046 409022 532102
rect 408594 531922 408650 531978
rect 408718 531922 408774 531978
rect 408842 531922 408898 531978
rect 408966 531922 409022 531978
rect 408594 514294 408650 514350
rect 408718 514294 408774 514350
rect 408842 514294 408898 514350
rect 408966 514294 409022 514350
rect 408594 514170 408650 514226
rect 408718 514170 408774 514226
rect 408842 514170 408898 514226
rect 408966 514170 409022 514226
rect 408594 514046 408650 514102
rect 408718 514046 408774 514102
rect 408842 514046 408898 514102
rect 408966 514046 409022 514102
rect 408594 513922 408650 513978
rect 408718 513922 408774 513978
rect 408842 513922 408898 513978
rect 408966 513922 409022 513978
rect 408594 496294 408650 496350
rect 408718 496294 408774 496350
rect 408842 496294 408898 496350
rect 408966 496294 409022 496350
rect 408594 496170 408650 496226
rect 408718 496170 408774 496226
rect 408842 496170 408898 496226
rect 408966 496170 409022 496226
rect 408594 496046 408650 496102
rect 408718 496046 408774 496102
rect 408842 496046 408898 496102
rect 408966 496046 409022 496102
rect 408594 495922 408650 495978
rect 408718 495922 408774 495978
rect 408842 495922 408898 495978
rect 408966 495922 409022 495978
rect 408594 478294 408650 478350
rect 408718 478294 408774 478350
rect 408842 478294 408898 478350
rect 408966 478294 409022 478350
rect 408594 478170 408650 478226
rect 408718 478170 408774 478226
rect 408842 478170 408898 478226
rect 408966 478170 409022 478226
rect 408594 478046 408650 478102
rect 408718 478046 408774 478102
rect 408842 478046 408898 478102
rect 408966 478046 409022 478102
rect 408594 477922 408650 477978
rect 408718 477922 408774 477978
rect 408842 477922 408898 477978
rect 408966 477922 409022 477978
rect 408594 460294 408650 460350
rect 408718 460294 408774 460350
rect 408842 460294 408898 460350
rect 408966 460294 409022 460350
rect 408594 460170 408650 460226
rect 408718 460170 408774 460226
rect 408842 460170 408898 460226
rect 408966 460170 409022 460226
rect 408594 460046 408650 460102
rect 408718 460046 408774 460102
rect 408842 460046 408898 460102
rect 408966 460046 409022 460102
rect 408594 459922 408650 459978
rect 408718 459922 408774 459978
rect 408842 459922 408898 459978
rect 408966 459922 409022 459978
rect 408594 442294 408650 442350
rect 408718 442294 408774 442350
rect 408842 442294 408898 442350
rect 408966 442294 409022 442350
rect 408594 442170 408650 442226
rect 408718 442170 408774 442226
rect 408842 442170 408898 442226
rect 408966 442170 409022 442226
rect 408594 442046 408650 442102
rect 408718 442046 408774 442102
rect 408842 442046 408898 442102
rect 408966 442046 409022 442102
rect 408594 441922 408650 441978
rect 408718 441922 408774 441978
rect 408842 441922 408898 441978
rect 408966 441922 409022 441978
rect 408594 424294 408650 424350
rect 408718 424294 408774 424350
rect 408842 424294 408898 424350
rect 408966 424294 409022 424350
rect 408594 424170 408650 424226
rect 408718 424170 408774 424226
rect 408842 424170 408898 424226
rect 408966 424170 409022 424226
rect 408594 424046 408650 424102
rect 408718 424046 408774 424102
rect 408842 424046 408898 424102
rect 408966 424046 409022 424102
rect 408594 423922 408650 423978
rect 408718 423922 408774 423978
rect 408842 423922 408898 423978
rect 408966 423922 409022 423978
rect 408594 406294 408650 406350
rect 408718 406294 408774 406350
rect 408842 406294 408898 406350
rect 408966 406294 409022 406350
rect 408594 406170 408650 406226
rect 408718 406170 408774 406226
rect 408842 406170 408898 406226
rect 408966 406170 409022 406226
rect 408594 406046 408650 406102
rect 408718 406046 408774 406102
rect 408842 406046 408898 406102
rect 408966 406046 409022 406102
rect 408594 405922 408650 405978
rect 408718 405922 408774 405978
rect 408842 405922 408898 405978
rect 408966 405922 409022 405978
rect 408594 388294 408650 388350
rect 408718 388294 408774 388350
rect 408842 388294 408898 388350
rect 408966 388294 409022 388350
rect 408594 388170 408650 388226
rect 408718 388170 408774 388226
rect 408842 388170 408898 388226
rect 408966 388170 409022 388226
rect 408594 388046 408650 388102
rect 408718 388046 408774 388102
rect 408842 388046 408898 388102
rect 408966 388046 409022 388102
rect 408594 387922 408650 387978
rect 408718 387922 408774 387978
rect 408842 387922 408898 387978
rect 408966 387922 409022 387978
rect 408594 370294 408650 370350
rect 408718 370294 408774 370350
rect 408842 370294 408898 370350
rect 408966 370294 409022 370350
rect 408594 370170 408650 370226
rect 408718 370170 408774 370226
rect 408842 370170 408898 370226
rect 408966 370170 409022 370226
rect 408594 370046 408650 370102
rect 408718 370046 408774 370102
rect 408842 370046 408898 370102
rect 408966 370046 409022 370102
rect 408594 369922 408650 369978
rect 408718 369922 408774 369978
rect 408842 369922 408898 369978
rect 408966 369922 409022 369978
rect 408594 352294 408650 352350
rect 408718 352294 408774 352350
rect 408842 352294 408898 352350
rect 408966 352294 409022 352350
rect 408594 352170 408650 352226
rect 408718 352170 408774 352226
rect 408842 352170 408898 352226
rect 408966 352170 409022 352226
rect 408594 352046 408650 352102
rect 408718 352046 408774 352102
rect 408842 352046 408898 352102
rect 408966 352046 409022 352102
rect 408594 351922 408650 351978
rect 408718 351922 408774 351978
rect 408842 351922 408898 351978
rect 408966 351922 409022 351978
rect 408594 334294 408650 334350
rect 408718 334294 408774 334350
rect 408842 334294 408898 334350
rect 408966 334294 409022 334350
rect 408594 334170 408650 334226
rect 408718 334170 408774 334226
rect 408842 334170 408898 334226
rect 408966 334170 409022 334226
rect 408594 334046 408650 334102
rect 408718 334046 408774 334102
rect 408842 334046 408898 334102
rect 408966 334046 409022 334102
rect 408594 333922 408650 333978
rect 408718 333922 408774 333978
rect 408842 333922 408898 333978
rect 408966 333922 409022 333978
rect 435594 597156 435650 597212
rect 435718 597156 435774 597212
rect 435842 597156 435898 597212
rect 435966 597156 436022 597212
rect 435594 597032 435650 597088
rect 435718 597032 435774 597088
rect 435842 597032 435898 597088
rect 435966 597032 436022 597088
rect 435594 596908 435650 596964
rect 435718 596908 435774 596964
rect 435842 596908 435898 596964
rect 435966 596908 436022 596964
rect 435594 596784 435650 596840
rect 435718 596784 435774 596840
rect 435842 596784 435898 596840
rect 435966 596784 436022 596840
rect 435594 580294 435650 580350
rect 435718 580294 435774 580350
rect 435842 580294 435898 580350
rect 435966 580294 436022 580350
rect 435594 580170 435650 580226
rect 435718 580170 435774 580226
rect 435842 580170 435898 580226
rect 435966 580170 436022 580226
rect 435594 580046 435650 580102
rect 435718 580046 435774 580102
rect 435842 580046 435898 580102
rect 435966 580046 436022 580102
rect 435594 579922 435650 579978
rect 435718 579922 435774 579978
rect 435842 579922 435898 579978
rect 435966 579922 436022 579978
rect 435594 562294 435650 562350
rect 435718 562294 435774 562350
rect 435842 562294 435898 562350
rect 435966 562294 436022 562350
rect 435594 562170 435650 562226
rect 435718 562170 435774 562226
rect 435842 562170 435898 562226
rect 435966 562170 436022 562226
rect 435594 562046 435650 562102
rect 435718 562046 435774 562102
rect 435842 562046 435898 562102
rect 435966 562046 436022 562102
rect 435594 561922 435650 561978
rect 435718 561922 435774 561978
rect 435842 561922 435898 561978
rect 435966 561922 436022 561978
rect 435594 544294 435650 544350
rect 435718 544294 435774 544350
rect 435842 544294 435898 544350
rect 435966 544294 436022 544350
rect 435594 544170 435650 544226
rect 435718 544170 435774 544226
rect 435842 544170 435898 544226
rect 435966 544170 436022 544226
rect 435594 544046 435650 544102
rect 435718 544046 435774 544102
rect 435842 544046 435898 544102
rect 435966 544046 436022 544102
rect 435594 543922 435650 543978
rect 435718 543922 435774 543978
rect 435842 543922 435898 543978
rect 435966 543922 436022 543978
rect 435594 526294 435650 526350
rect 435718 526294 435774 526350
rect 435842 526294 435898 526350
rect 435966 526294 436022 526350
rect 435594 526170 435650 526226
rect 435718 526170 435774 526226
rect 435842 526170 435898 526226
rect 435966 526170 436022 526226
rect 435594 526046 435650 526102
rect 435718 526046 435774 526102
rect 435842 526046 435898 526102
rect 435966 526046 436022 526102
rect 435594 525922 435650 525978
rect 435718 525922 435774 525978
rect 435842 525922 435898 525978
rect 435966 525922 436022 525978
rect 435594 508294 435650 508350
rect 435718 508294 435774 508350
rect 435842 508294 435898 508350
rect 435966 508294 436022 508350
rect 435594 508170 435650 508226
rect 435718 508170 435774 508226
rect 435842 508170 435898 508226
rect 435966 508170 436022 508226
rect 435594 508046 435650 508102
rect 435718 508046 435774 508102
rect 435842 508046 435898 508102
rect 435966 508046 436022 508102
rect 435594 507922 435650 507978
rect 435718 507922 435774 507978
rect 435842 507922 435898 507978
rect 435966 507922 436022 507978
rect 435594 490294 435650 490350
rect 435718 490294 435774 490350
rect 435842 490294 435898 490350
rect 435966 490294 436022 490350
rect 435594 490170 435650 490226
rect 435718 490170 435774 490226
rect 435842 490170 435898 490226
rect 435966 490170 436022 490226
rect 435594 490046 435650 490102
rect 435718 490046 435774 490102
rect 435842 490046 435898 490102
rect 435966 490046 436022 490102
rect 435594 489922 435650 489978
rect 435718 489922 435774 489978
rect 435842 489922 435898 489978
rect 435966 489922 436022 489978
rect 435594 472294 435650 472350
rect 435718 472294 435774 472350
rect 435842 472294 435898 472350
rect 435966 472294 436022 472350
rect 435594 472170 435650 472226
rect 435718 472170 435774 472226
rect 435842 472170 435898 472226
rect 435966 472170 436022 472226
rect 435594 472046 435650 472102
rect 435718 472046 435774 472102
rect 435842 472046 435898 472102
rect 435966 472046 436022 472102
rect 435594 471922 435650 471978
rect 435718 471922 435774 471978
rect 435842 471922 435898 471978
rect 435966 471922 436022 471978
rect 435594 454294 435650 454350
rect 435718 454294 435774 454350
rect 435842 454294 435898 454350
rect 435966 454294 436022 454350
rect 435594 454170 435650 454226
rect 435718 454170 435774 454226
rect 435842 454170 435898 454226
rect 435966 454170 436022 454226
rect 435594 454046 435650 454102
rect 435718 454046 435774 454102
rect 435842 454046 435898 454102
rect 435966 454046 436022 454102
rect 435594 453922 435650 453978
rect 435718 453922 435774 453978
rect 435842 453922 435898 453978
rect 435966 453922 436022 453978
rect 435594 436294 435650 436350
rect 435718 436294 435774 436350
rect 435842 436294 435898 436350
rect 435966 436294 436022 436350
rect 435594 436170 435650 436226
rect 435718 436170 435774 436226
rect 435842 436170 435898 436226
rect 435966 436170 436022 436226
rect 435594 436046 435650 436102
rect 435718 436046 435774 436102
rect 435842 436046 435898 436102
rect 435966 436046 436022 436102
rect 435594 435922 435650 435978
rect 435718 435922 435774 435978
rect 435842 435922 435898 435978
rect 435966 435922 436022 435978
rect 435594 418294 435650 418350
rect 435718 418294 435774 418350
rect 435842 418294 435898 418350
rect 435966 418294 436022 418350
rect 435594 418170 435650 418226
rect 435718 418170 435774 418226
rect 435842 418170 435898 418226
rect 435966 418170 436022 418226
rect 435594 418046 435650 418102
rect 435718 418046 435774 418102
rect 435842 418046 435898 418102
rect 435966 418046 436022 418102
rect 435594 417922 435650 417978
rect 435718 417922 435774 417978
rect 435842 417922 435898 417978
rect 435966 417922 436022 417978
rect 435594 400294 435650 400350
rect 435718 400294 435774 400350
rect 435842 400294 435898 400350
rect 435966 400294 436022 400350
rect 435594 400170 435650 400226
rect 435718 400170 435774 400226
rect 435842 400170 435898 400226
rect 435966 400170 436022 400226
rect 435594 400046 435650 400102
rect 435718 400046 435774 400102
rect 435842 400046 435898 400102
rect 435966 400046 436022 400102
rect 435594 399922 435650 399978
rect 435718 399922 435774 399978
rect 435842 399922 435898 399978
rect 435966 399922 436022 399978
rect 435594 382294 435650 382350
rect 435718 382294 435774 382350
rect 435842 382294 435898 382350
rect 435966 382294 436022 382350
rect 435594 382170 435650 382226
rect 435718 382170 435774 382226
rect 435842 382170 435898 382226
rect 435966 382170 436022 382226
rect 435594 382046 435650 382102
rect 435718 382046 435774 382102
rect 435842 382046 435898 382102
rect 435966 382046 436022 382102
rect 435594 381922 435650 381978
rect 435718 381922 435774 381978
rect 435842 381922 435898 381978
rect 435966 381922 436022 381978
rect 435594 364294 435650 364350
rect 435718 364294 435774 364350
rect 435842 364294 435898 364350
rect 435966 364294 436022 364350
rect 435594 364170 435650 364226
rect 435718 364170 435774 364226
rect 435842 364170 435898 364226
rect 435966 364170 436022 364226
rect 435594 364046 435650 364102
rect 435718 364046 435774 364102
rect 435842 364046 435898 364102
rect 435966 364046 436022 364102
rect 435594 363922 435650 363978
rect 435718 363922 435774 363978
rect 435842 363922 435898 363978
rect 435966 363922 436022 363978
rect 435594 346294 435650 346350
rect 435718 346294 435774 346350
rect 435842 346294 435898 346350
rect 435966 346294 436022 346350
rect 435594 346170 435650 346226
rect 435718 346170 435774 346226
rect 435842 346170 435898 346226
rect 435966 346170 436022 346226
rect 435594 346046 435650 346102
rect 435718 346046 435774 346102
rect 435842 346046 435898 346102
rect 435966 346046 436022 346102
rect 435594 345922 435650 345978
rect 435718 345922 435774 345978
rect 435842 345922 435898 345978
rect 435966 345922 436022 345978
rect 435594 328294 435650 328350
rect 435718 328294 435774 328350
rect 435842 328294 435898 328350
rect 435966 328294 436022 328350
rect 435594 328170 435650 328226
rect 435718 328170 435774 328226
rect 435842 328170 435898 328226
rect 435966 328170 436022 328226
rect 408594 316294 408650 316350
rect 408718 316294 408774 316350
rect 408842 316294 408898 316350
rect 408966 316294 409022 316350
rect 408594 316170 408650 316226
rect 408718 316170 408774 316226
rect 408842 316170 408898 316226
rect 408966 316170 409022 316226
rect 408594 316046 408650 316102
rect 408718 316046 408774 316102
rect 408842 316046 408898 316102
rect 408966 316046 409022 316102
rect 408594 315922 408650 315978
rect 408718 315922 408774 315978
rect 408842 315922 408898 315978
rect 408966 315922 409022 315978
rect 411516 312542 411572 312598
rect 415238 310294 415294 310350
rect 415362 310294 415418 310350
rect 415238 310170 415294 310226
rect 415362 310170 415418 310226
rect 415238 310046 415294 310102
rect 415362 310046 415418 310102
rect 415238 309922 415294 309978
rect 415362 309922 415418 309978
rect 399878 298294 399934 298350
rect 400002 298294 400058 298350
rect 399878 298170 399934 298226
rect 400002 298170 400058 298226
rect 399878 298046 399934 298102
rect 400002 298046 400058 298102
rect 399878 297922 399934 297978
rect 400002 297922 400058 297978
rect 415238 292294 415294 292350
rect 415362 292294 415418 292350
rect 415238 292170 415294 292226
rect 415362 292170 415418 292226
rect 415238 292046 415294 292102
rect 415362 292046 415418 292102
rect 415238 291922 415294 291978
rect 415362 291922 415418 291978
rect 387324 286082 387380 286138
rect 399878 280294 399934 280350
rect 400002 280294 400058 280350
rect 399878 280170 399934 280226
rect 400002 280170 400058 280226
rect 399878 280046 399934 280102
rect 400002 280046 400058 280102
rect 399878 279922 399934 279978
rect 400002 279922 400058 279978
rect 385420 270602 385476 270658
rect 387996 268802 388052 268858
rect 387436 261602 387492 261658
rect 408594 262294 408650 262350
rect 408718 262294 408774 262350
rect 408842 262294 408898 262350
rect 408966 262294 409022 262350
rect 408594 262170 408650 262226
rect 408718 262170 408774 262226
rect 408842 262170 408898 262226
rect 408966 262170 409022 262226
rect 408594 262046 408650 262102
rect 408718 262046 408774 262102
rect 408842 262046 408898 262102
rect 408966 262046 409022 262102
rect 408594 261922 408650 261978
rect 408718 261922 408774 261978
rect 408842 261922 408898 261978
rect 408966 261922 409022 261978
rect 413308 264482 413364 264538
rect 416332 268082 416388 268138
rect 418572 312542 418628 312598
rect 435594 328046 435650 328102
rect 435718 328046 435774 328102
rect 435842 328046 435898 328102
rect 435966 328046 436022 328102
rect 424620 267902 424676 267958
rect 420364 267204 420420 267238
rect 420364 267182 420420 267204
rect 430598 316294 430654 316350
rect 430722 316294 430778 316350
rect 430598 316170 430654 316226
rect 430722 316170 430778 316226
rect 430598 316046 430654 316102
rect 430722 316046 430778 316102
rect 430598 315922 430654 315978
rect 430722 315922 430778 315978
rect 430598 298294 430654 298350
rect 430722 298294 430778 298350
rect 430598 298170 430654 298226
rect 430722 298170 430778 298226
rect 430598 298046 430654 298102
rect 430722 298046 430778 298102
rect 430598 297922 430654 297978
rect 430722 297922 430778 297978
rect 430598 280294 430654 280350
rect 430722 280294 430778 280350
rect 430598 280170 430654 280226
rect 430722 280170 430778 280226
rect 430598 280046 430654 280102
rect 430722 280046 430778 280102
rect 430598 279922 430654 279978
rect 430722 279922 430778 279978
rect 435594 327922 435650 327978
rect 435718 327922 435774 327978
rect 435842 327922 435898 327978
rect 435966 327922 436022 327978
rect 403564 261242 403620 261298
rect 383852 260342 383908 260398
rect 384518 256294 384574 256350
rect 384642 256294 384698 256350
rect 384518 256170 384574 256226
rect 384642 256170 384698 256226
rect 384518 256046 384574 256102
rect 384642 256046 384698 256102
rect 384518 255922 384574 255978
rect 384642 255922 384698 255978
rect 415238 256294 415294 256350
rect 415362 256294 415418 256350
rect 415238 256170 415294 256226
rect 415362 256170 415418 256226
rect 415238 256046 415294 256102
rect 415362 256046 415418 256102
rect 415238 255922 415294 255978
rect 415362 255922 415418 255978
rect 399878 244294 399934 244350
rect 400002 244294 400058 244350
rect 399878 244170 399934 244226
rect 400002 244170 400058 244226
rect 399878 244046 399934 244102
rect 400002 244046 400058 244102
rect 399878 243922 399934 243978
rect 400002 243922 400058 243978
rect 381500 241802 381556 241858
rect 384518 238294 384574 238350
rect 384642 238294 384698 238350
rect 384518 238170 384574 238226
rect 384642 238170 384698 238226
rect 384518 238046 384574 238102
rect 384642 238046 384698 238102
rect 384518 237922 384574 237978
rect 384642 237922 384698 237978
rect 415238 238294 415294 238350
rect 415362 238294 415418 238350
rect 415238 238170 415294 238226
rect 415362 238170 415418 238226
rect 415238 238046 415294 238102
rect 415362 238046 415418 238102
rect 415238 237922 415294 237978
rect 415362 237922 415418 237978
rect 399878 226294 399934 226350
rect 400002 226294 400058 226350
rect 399878 226170 399934 226226
rect 400002 226170 400058 226226
rect 399878 226046 399934 226102
rect 400002 226046 400058 226102
rect 399878 225922 399934 225978
rect 400002 225922 400058 225978
rect 384518 220294 384574 220350
rect 384642 220294 384698 220350
rect 384518 220170 384574 220226
rect 384642 220170 384698 220226
rect 384518 220046 384574 220102
rect 384642 220046 384698 220102
rect 384518 219922 384574 219978
rect 384642 219922 384698 219978
rect 415238 220294 415294 220350
rect 415362 220294 415418 220350
rect 415238 220170 415294 220226
rect 415362 220170 415418 220226
rect 415238 220046 415294 220102
rect 415362 220046 415418 220102
rect 415238 219922 415294 219978
rect 415362 219922 415418 219978
rect 381388 218402 381444 218458
rect 383852 217682 383908 217738
rect 381724 216962 381780 217018
rect 381388 215882 381444 215938
rect 381500 216782 381556 216838
rect 381164 209042 381220 209098
rect 380380 166572 380436 166618
rect 380380 166562 380436 166572
rect 380604 149828 380660 149878
rect 380604 149822 380660 149828
rect 380604 144962 380660 145018
rect 380156 117422 380212 117478
rect 379932 72062 379988 72118
rect 381612 215162 381668 215218
rect 382060 215522 382116 215578
rect 381836 215342 381892 215398
rect 381948 213542 382004 213598
rect 381612 156302 381668 156358
rect 381724 166562 381780 166618
rect 381500 149822 381556 149878
rect 381388 72062 381444 72118
rect 381500 74222 381556 74278
rect 381388 71342 381444 71398
rect 382508 213182 382564 213238
rect 383404 211742 383460 211798
rect 382284 144962 382340 145018
rect 382508 151082 382564 151138
rect 384076 217502 384132 217558
rect 395724 214262 395780 214318
rect 386764 212102 386820 212158
rect 386092 210842 386148 210898
rect 392252 211922 392308 211978
rect 389452 211022 389508 211078
rect 389788 198100 389844 198118
rect 389788 198062 389844 198100
rect 384076 187802 384132 187858
rect 384518 184294 384574 184350
rect 384642 184294 384698 184350
rect 384518 184170 384574 184226
rect 384642 184170 384698 184226
rect 384518 184046 384574 184102
rect 384642 184046 384698 184102
rect 384518 183922 384574 183978
rect 384642 183922 384698 183978
rect 399836 208337 399892 208393
rect 399940 208337 399996 208393
rect 400044 208337 400100 208393
rect 399836 208233 399892 208289
rect 399940 208233 399996 208289
rect 400044 208233 400100 208289
rect 399836 208129 399892 208185
rect 399940 208129 399996 208185
rect 400044 208129 400100 208185
rect 402220 204002 402276 204058
rect 408594 208294 408650 208350
rect 408718 208294 408774 208350
rect 408842 208294 408898 208350
rect 408966 208294 409022 208350
rect 408594 208170 408650 208226
rect 408718 208170 408774 208226
rect 408842 208170 408898 208226
rect 408966 208170 409022 208226
rect 408594 208046 408650 208102
rect 408718 208046 408774 208102
rect 408842 208046 408898 208102
rect 408966 208046 409022 208102
rect 408594 207922 408650 207978
rect 408718 207922 408774 207978
rect 408842 207922 408898 207978
rect 408966 207922 409022 207978
rect 404874 202294 404930 202350
rect 404998 202294 405054 202350
rect 405122 202294 405178 202350
rect 405246 202294 405302 202350
rect 404874 202170 404930 202226
rect 404998 202170 405054 202226
rect 405122 202170 405178 202226
rect 405246 202170 405302 202226
rect 404874 202046 404930 202102
rect 404998 202046 405054 202102
rect 405122 202046 405178 202102
rect 405246 202046 405302 202102
rect 404874 201922 404930 201978
rect 404998 201922 405054 201978
rect 405122 201922 405178 201978
rect 405246 201922 405302 201978
rect 399878 190294 399934 190350
rect 400002 190294 400058 190350
rect 399878 190170 399934 190226
rect 400002 190170 400058 190226
rect 399878 190046 399934 190102
rect 400002 190046 400058 190102
rect 399878 189922 399934 189978
rect 400002 189922 400058 189978
rect 404874 184330 404930 184386
rect 404998 184330 405054 184386
rect 405122 184330 405178 184386
rect 405246 184330 405302 184386
rect 404874 184206 404930 184262
rect 404998 184206 405054 184262
rect 405122 184206 405178 184262
rect 405246 184206 405302 184262
rect 404874 184082 404930 184138
rect 404998 184082 405054 184138
rect 405122 184082 405178 184138
rect 405246 184082 405302 184138
rect 418348 213362 418404 213418
rect 430598 244294 430654 244350
rect 430722 244294 430778 244350
rect 430598 244170 430654 244226
rect 430722 244170 430778 244226
rect 430598 244046 430654 244102
rect 430722 244046 430778 244102
rect 430598 243922 430654 243978
rect 430722 243922 430778 243978
rect 431004 242702 431060 242758
rect 430598 226294 430654 226350
rect 430722 226294 430778 226350
rect 430598 226170 430654 226226
rect 430722 226170 430778 226226
rect 430598 226046 430654 226102
rect 430722 226046 430778 226102
rect 430598 225922 430654 225978
rect 430722 225922 430778 225978
rect 430556 208337 430612 208393
rect 430660 208337 430716 208393
rect 430764 208337 430820 208393
rect 430556 208233 430612 208289
rect 430660 208233 430716 208289
rect 430764 208233 430820 208289
rect 430556 208129 430612 208185
rect 430660 208129 430716 208185
rect 430764 208129 430820 208185
rect 430108 198062 430164 198118
rect 408594 190294 408650 190350
rect 408718 190294 408774 190350
rect 408842 190294 408898 190350
rect 408966 190294 409022 190350
rect 408594 190170 408650 190226
rect 408718 190170 408774 190226
rect 408842 190170 408898 190226
rect 408966 190170 409022 190226
rect 408594 190046 408650 190102
rect 408718 190046 408774 190102
rect 408842 190046 408898 190102
rect 408966 190046 409022 190102
rect 408594 189922 408650 189978
rect 408718 189922 408774 189978
rect 408842 189922 408898 189978
rect 408966 189922 409022 189978
rect 430598 190294 430654 190350
rect 430722 190294 430778 190350
rect 430598 190170 430654 190226
rect 430722 190170 430778 190226
rect 430598 190046 430654 190102
rect 430722 190046 430778 190102
rect 430598 189922 430654 189978
rect 430722 189922 430778 189978
rect 431004 187982 431060 188038
rect 415238 184294 415294 184350
rect 415362 184294 415418 184350
rect 415238 184170 415294 184226
rect 415362 184170 415418 184226
rect 415238 184046 415294 184102
rect 415362 184046 415418 184102
rect 415238 183922 415294 183978
rect 415362 183922 415418 183978
rect 395612 182222 395668 182278
rect 399878 172294 399934 172350
rect 400002 172294 400058 172350
rect 399878 172170 399934 172226
rect 400002 172170 400058 172226
rect 399878 172046 399934 172102
rect 400002 172046 400058 172102
rect 399878 171922 399934 171978
rect 400002 171922 400058 171978
rect 430598 172294 430654 172350
rect 430722 172294 430778 172350
rect 430598 172170 430654 172226
rect 430722 172170 430778 172226
rect 430598 172046 430654 172102
rect 430722 172046 430778 172102
rect 430598 171922 430654 171978
rect 430722 171922 430778 171978
rect 384518 166294 384574 166350
rect 384642 166294 384698 166350
rect 384518 166170 384574 166226
rect 384642 166170 384698 166226
rect 384518 166046 384574 166102
rect 384642 166046 384698 166102
rect 384518 165922 384574 165978
rect 384642 165922 384698 165978
rect 415238 166294 415294 166350
rect 415362 166294 415418 166350
rect 415238 166170 415294 166226
rect 415362 166170 415418 166226
rect 415238 166046 415294 166102
rect 415362 166046 415418 166102
rect 415238 165922 415294 165978
rect 415362 165922 415418 165978
rect 399878 154294 399934 154350
rect 400002 154294 400058 154350
rect 399878 154170 399934 154226
rect 400002 154170 400058 154226
rect 399878 154046 399934 154102
rect 400002 154046 400058 154102
rect 399878 153922 399934 153978
rect 400002 153922 400058 153978
rect 430598 154294 430654 154350
rect 430722 154294 430778 154350
rect 430598 154170 430654 154226
rect 430722 154170 430778 154226
rect 430598 154046 430654 154102
rect 430722 154046 430778 154102
rect 430598 153922 430654 153978
rect 430722 153922 430778 153978
rect 384518 148294 384574 148350
rect 384642 148294 384698 148350
rect 384518 148170 384574 148226
rect 384642 148170 384698 148226
rect 384518 148046 384574 148102
rect 384642 148046 384698 148102
rect 384518 147922 384574 147978
rect 384642 147922 384698 147978
rect 415238 148294 415294 148350
rect 415362 148294 415418 148350
rect 415238 148170 415294 148226
rect 415362 148170 415418 148226
rect 415238 148046 415294 148102
rect 415362 148046 415418 148102
rect 415238 147922 415294 147978
rect 415362 147922 415418 147978
rect 384518 112294 384574 112350
rect 384642 112294 384698 112350
rect 384518 112170 384574 112226
rect 384642 112170 384698 112226
rect 384518 112046 384574 112102
rect 384642 112046 384698 112102
rect 384518 111922 384574 111978
rect 384642 111922 384698 111978
rect 384518 94294 384574 94350
rect 384642 94294 384698 94350
rect 384518 94170 384574 94226
rect 384642 94170 384698 94226
rect 384518 94046 384574 94102
rect 384642 94046 384698 94102
rect 384518 93922 384574 93978
rect 384642 93922 384698 93978
rect 381836 72782 381892 72838
rect 383068 76562 383124 76618
rect 384972 78362 385028 78418
rect 384518 76294 384574 76350
rect 384642 76294 384698 76350
rect 384518 76170 384574 76226
rect 384642 76170 384698 76226
rect 384518 76046 384574 76102
rect 384642 76046 384698 76102
rect 384518 75922 384574 75978
rect 384642 75922 384698 75978
rect 383852 74042 383908 74098
rect 384518 58294 384574 58350
rect 384642 58294 384698 58350
rect 384518 58170 384574 58226
rect 384642 58170 384698 58226
rect 384518 58046 384574 58102
rect 384642 58046 384698 58102
rect 384518 57922 384574 57978
rect 384642 57922 384698 57978
rect 385644 80522 385700 80578
rect 386428 80702 386484 80758
rect 385644 78002 385700 78058
rect 386540 81602 386596 81658
rect 388332 71342 388388 71398
rect 388108 64682 388164 64738
rect 388332 64862 388388 64918
rect 389788 62882 389844 62938
rect 389900 80522 389956 80578
rect 390012 78002 390068 78058
rect 391468 100862 391524 100918
rect 392364 105722 392420 105778
rect 392476 100862 392532 100918
rect 393148 74042 393204 74098
rect 394156 91502 394212 91558
rect 394828 52082 394884 52138
rect 396396 115982 396452 116038
rect 408594 136294 408650 136350
rect 408718 136294 408774 136350
rect 408842 136294 408898 136350
rect 408966 136294 409022 136350
rect 408594 136170 408650 136226
rect 408718 136170 408774 136226
rect 408842 136170 408898 136226
rect 408966 136170 409022 136226
rect 408594 136046 408650 136102
rect 408718 136046 408774 136102
rect 408842 136046 408898 136102
rect 408966 136046 409022 136102
rect 408594 135922 408650 135978
rect 408718 135922 408774 135978
rect 408842 135922 408898 135978
rect 408966 135922 409022 135978
rect 399878 118294 399934 118350
rect 400002 118294 400058 118350
rect 399878 118170 399934 118226
rect 400002 118170 400058 118226
rect 399878 118046 399934 118102
rect 400002 118046 400058 118102
rect 399878 117922 399934 117978
rect 400002 117922 400058 117978
rect 439314 598116 439370 598172
rect 439438 598116 439494 598172
rect 439562 598116 439618 598172
rect 439686 598116 439742 598172
rect 439314 597992 439370 598048
rect 439438 597992 439494 598048
rect 439562 597992 439618 598048
rect 439686 597992 439742 598048
rect 439314 597868 439370 597924
rect 439438 597868 439494 597924
rect 439562 597868 439618 597924
rect 439686 597868 439742 597924
rect 439314 597744 439370 597800
rect 439438 597744 439494 597800
rect 439562 597744 439618 597800
rect 439686 597744 439742 597800
rect 439314 586294 439370 586350
rect 439438 586294 439494 586350
rect 439562 586294 439618 586350
rect 439686 586294 439742 586350
rect 439314 586170 439370 586226
rect 439438 586170 439494 586226
rect 439562 586170 439618 586226
rect 439686 586170 439742 586226
rect 439314 586046 439370 586102
rect 439438 586046 439494 586102
rect 439562 586046 439618 586102
rect 439686 586046 439742 586102
rect 439314 585922 439370 585978
rect 439438 585922 439494 585978
rect 439562 585922 439618 585978
rect 439686 585922 439742 585978
rect 439314 568294 439370 568350
rect 439438 568294 439494 568350
rect 439562 568294 439618 568350
rect 439686 568294 439742 568350
rect 439314 568170 439370 568226
rect 439438 568170 439494 568226
rect 439562 568170 439618 568226
rect 439686 568170 439742 568226
rect 439314 568046 439370 568102
rect 439438 568046 439494 568102
rect 439562 568046 439618 568102
rect 439686 568046 439742 568102
rect 439314 567922 439370 567978
rect 439438 567922 439494 567978
rect 439562 567922 439618 567978
rect 439686 567922 439742 567978
rect 439314 550294 439370 550350
rect 439438 550294 439494 550350
rect 439562 550294 439618 550350
rect 439686 550294 439742 550350
rect 439314 550170 439370 550226
rect 439438 550170 439494 550226
rect 439562 550170 439618 550226
rect 439686 550170 439742 550226
rect 439314 550046 439370 550102
rect 439438 550046 439494 550102
rect 439562 550046 439618 550102
rect 439686 550046 439742 550102
rect 439314 549922 439370 549978
rect 439438 549922 439494 549978
rect 439562 549922 439618 549978
rect 439686 549922 439742 549978
rect 439314 532294 439370 532350
rect 439438 532294 439494 532350
rect 439562 532294 439618 532350
rect 439686 532294 439742 532350
rect 439314 532170 439370 532226
rect 439438 532170 439494 532226
rect 439562 532170 439618 532226
rect 439686 532170 439742 532226
rect 439314 532046 439370 532102
rect 439438 532046 439494 532102
rect 439562 532046 439618 532102
rect 439686 532046 439742 532102
rect 439314 531922 439370 531978
rect 439438 531922 439494 531978
rect 439562 531922 439618 531978
rect 439686 531922 439742 531978
rect 439314 514294 439370 514350
rect 439438 514294 439494 514350
rect 439562 514294 439618 514350
rect 439686 514294 439742 514350
rect 439314 514170 439370 514226
rect 439438 514170 439494 514226
rect 439562 514170 439618 514226
rect 439686 514170 439742 514226
rect 439314 514046 439370 514102
rect 439438 514046 439494 514102
rect 439562 514046 439618 514102
rect 439686 514046 439742 514102
rect 439314 513922 439370 513978
rect 439438 513922 439494 513978
rect 439562 513922 439618 513978
rect 439686 513922 439742 513978
rect 439314 496294 439370 496350
rect 439438 496294 439494 496350
rect 439562 496294 439618 496350
rect 439686 496294 439742 496350
rect 439314 496170 439370 496226
rect 439438 496170 439494 496226
rect 439562 496170 439618 496226
rect 439686 496170 439742 496226
rect 439314 496046 439370 496102
rect 439438 496046 439494 496102
rect 439562 496046 439618 496102
rect 439686 496046 439742 496102
rect 439314 495922 439370 495978
rect 439438 495922 439494 495978
rect 439562 495922 439618 495978
rect 439686 495922 439742 495978
rect 439314 478294 439370 478350
rect 439438 478294 439494 478350
rect 439562 478294 439618 478350
rect 439686 478294 439742 478350
rect 439314 478170 439370 478226
rect 439438 478170 439494 478226
rect 439562 478170 439618 478226
rect 439686 478170 439742 478226
rect 439314 478046 439370 478102
rect 439438 478046 439494 478102
rect 439562 478046 439618 478102
rect 439686 478046 439742 478102
rect 439314 477922 439370 477978
rect 439438 477922 439494 477978
rect 439562 477922 439618 477978
rect 439686 477922 439742 477978
rect 439314 460294 439370 460350
rect 439438 460294 439494 460350
rect 439562 460294 439618 460350
rect 439686 460294 439742 460350
rect 439314 460170 439370 460226
rect 439438 460170 439494 460226
rect 439562 460170 439618 460226
rect 439686 460170 439742 460226
rect 439314 460046 439370 460102
rect 439438 460046 439494 460102
rect 439562 460046 439618 460102
rect 439686 460046 439742 460102
rect 439314 459922 439370 459978
rect 439438 459922 439494 459978
rect 439562 459922 439618 459978
rect 439686 459922 439742 459978
rect 439314 442294 439370 442350
rect 439438 442294 439494 442350
rect 439562 442294 439618 442350
rect 439686 442294 439742 442350
rect 439314 442170 439370 442226
rect 439438 442170 439494 442226
rect 439562 442170 439618 442226
rect 439686 442170 439742 442226
rect 439314 442046 439370 442102
rect 439438 442046 439494 442102
rect 439562 442046 439618 442102
rect 439686 442046 439742 442102
rect 439314 441922 439370 441978
rect 439438 441922 439494 441978
rect 439562 441922 439618 441978
rect 439686 441922 439742 441978
rect 439314 424294 439370 424350
rect 439438 424294 439494 424350
rect 439562 424294 439618 424350
rect 439686 424294 439742 424350
rect 439314 424170 439370 424226
rect 439438 424170 439494 424226
rect 439562 424170 439618 424226
rect 439686 424170 439742 424226
rect 439314 424046 439370 424102
rect 439438 424046 439494 424102
rect 439562 424046 439618 424102
rect 439686 424046 439742 424102
rect 439314 423922 439370 423978
rect 439438 423922 439494 423978
rect 439562 423922 439618 423978
rect 439686 423922 439742 423978
rect 439314 406294 439370 406350
rect 439438 406294 439494 406350
rect 439562 406294 439618 406350
rect 439686 406294 439742 406350
rect 439314 406170 439370 406226
rect 439438 406170 439494 406226
rect 439562 406170 439618 406226
rect 439686 406170 439742 406226
rect 439314 406046 439370 406102
rect 439438 406046 439494 406102
rect 439562 406046 439618 406102
rect 439686 406046 439742 406102
rect 439314 405922 439370 405978
rect 439438 405922 439494 405978
rect 439562 405922 439618 405978
rect 439686 405922 439742 405978
rect 439314 388294 439370 388350
rect 439438 388294 439494 388350
rect 439562 388294 439618 388350
rect 439686 388294 439742 388350
rect 439314 388170 439370 388226
rect 439438 388170 439494 388226
rect 439562 388170 439618 388226
rect 439686 388170 439742 388226
rect 439314 388046 439370 388102
rect 439438 388046 439494 388102
rect 439562 388046 439618 388102
rect 439686 388046 439742 388102
rect 439314 387922 439370 387978
rect 439438 387922 439494 387978
rect 439562 387922 439618 387978
rect 439686 387922 439742 387978
rect 439314 370294 439370 370350
rect 439438 370294 439494 370350
rect 439562 370294 439618 370350
rect 439686 370294 439742 370350
rect 439314 370170 439370 370226
rect 439438 370170 439494 370226
rect 439562 370170 439618 370226
rect 439686 370170 439742 370226
rect 439314 370046 439370 370102
rect 439438 370046 439494 370102
rect 439562 370046 439618 370102
rect 439686 370046 439742 370102
rect 439314 369922 439370 369978
rect 439438 369922 439494 369978
rect 439562 369922 439618 369978
rect 439686 369922 439742 369978
rect 439314 352294 439370 352350
rect 439438 352294 439494 352350
rect 439562 352294 439618 352350
rect 439686 352294 439742 352350
rect 439314 352170 439370 352226
rect 439438 352170 439494 352226
rect 439562 352170 439618 352226
rect 439686 352170 439742 352226
rect 439314 352046 439370 352102
rect 439438 352046 439494 352102
rect 439562 352046 439618 352102
rect 439686 352046 439742 352102
rect 439314 351922 439370 351978
rect 439438 351922 439494 351978
rect 439562 351922 439618 351978
rect 439686 351922 439742 351978
rect 439314 334294 439370 334350
rect 439438 334294 439494 334350
rect 439562 334294 439618 334350
rect 439686 334294 439742 334350
rect 439314 334170 439370 334226
rect 439438 334170 439494 334226
rect 439562 334170 439618 334226
rect 439686 334170 439742 334226
rect 439314 334046 439370 334102
rect 439438 334046 439494 334102
rect 439562 334046 439618 334102
rect 439686 334046 439742 334102
rect 439314 333922 439370 333978
rect 439438 333922 439494 333978
rect 439562 333922 439618 333978
rect 439686 333922 439742 333978
rect 435594 310294 435650 310350
rect 435718 310294 435774 310350
rect 435842 310294 435898 310350
rect 435966 310294 436022 310350
rect 435594 310170 435650 310226
rect 435718 310170 435774 310226
rect 435842 310170 435898 310226
rect 435966 310170 436022 310226
rect 435594 310046 435650 310102
rect 435718 310046 435774 310102
rect 435842 310046 435898 310102
rect 435966 310046 436022 310102
rect 435594 309922 435650 309978
rect 435718 309922 435774 309978
rect 435842 309922 435898 309978
rect 435966 309922 436022 309978
rect 435594 292294 435650 292350
rect 435718 292294 435774 292350
rect 435842 292294 435898 292350
rect 435966 292294 436022 292350
rect 435594 292170 435650 292226
rect 435718 292170 435774 292226
rect 435842 292170 435898 292226
rect 435966 292170 436022 292226
rect 435594 292046 435650 292102
rect 435718 292046 435774 292102
rect 435842 292046 435898 292102
rect 435966 292046 436022 292102
rect 435594 291922 435650 291978
rect 435718 291922 435774 291978
rect 435842 291922 435898 291978
rect 435966 291922 436022 291978
rect 432124 204002 432180 204058
rect 435594 274294 435650 274350
rect 435718 274294 435774 274350
rect 435842 274294 435898 274350
rect 435966 274294 436022 274350
rect 435594 274170 435650 274226
rect 435718 274170 435774 274226
rect 435842 274170 435898 274226
rect 435966 274170 436022 274226
rect 435594 274046 435650 274102
rect 435718 274046 435774 274102
rect 435842 274046 435898 274102
rect 435966 274046 436022 274102
rect 435594 273922 435650 273978
rect 435718 273922 435774 273978
rect 435842 273922 435898 273978
rect 435966 273922 436022 273978
rect 434252 240002 434308 240058
rect 435594 256294 435650 256350
rect 435718 256294 435774 256350
rect 435842 256294 435898 256350
rect 435966 256294 436022 256350
rect 435594 256170 435650 256226
rect 435718 256170 435774 256226
rect 435842 256170 435898 256226
rect 435966 256170 436022 256226
rect 435594 256046 435650 256102
rect 435718 256046 435774 256102
rect 435842 256046 435898 256102
rect 435966 256046 436022 256102
rect 435594 255922 435650 255978
rect 435718 255922 435774 255978
rect 435842 255922 435898 255978
rect 435966 255922 436022 255978
rect 436828 242702 436884 242758
rect 466314 597156 466370 597212
rect 466438 597156 466494 597212
rect 466562 597156 466618 597212
rect 466686 597156 466742 597212
rect 466314 597032 466370 597088
rect 466438 597032 466494 597088
rect 466562 597032 466618 597088
rect 466686 597032 466742 597088
rect 466314 596908 466370 596964
rect 466438 596908 466494 596964
rect 466562 596908 466618 596964
rect 466686 596908 466742 596964
rect 466314 596784 466370 596840
rect 466438 596784 466494 596840
rect 466562 596784 466618 596840
rect 466686 596784 466742 596840
rect 466314 580294 466370 580350
rect 466438 580294 466494 580350
rect 466562 580294 466618 580350
rect 466686 580294 466742 580350
rect 466314 580170 466370 580226
rect 466438 580170 466494 580226
rect 466562 580170 466618 580226
rect 466686 580170 466742 580226
rect 466314 580046 466370 580102
rect 466438 580046 466494 580102
rect 466562 580046 466618 580102
rect 466686 580046 466742 580102
rect 466314 579922 466370 579978
rect 466438 579922 466494 579978
rect 466562 579922 466618 579978
rect 466686 579922 466742 579978
rect 466314 562294 466370 562350
rect 466438 562294 466494 562350
rect 466562 562294 466618 562350
rect 466686 562294 466742 562350
rect 466314 562170 466370 562226
rect 466438 562170 466494 562226
rect 466562 562170 466618 562226
rect 466686 562170 466742 562226
rect 466314 562046 466370 562102
rect 466438 562046 466494 562102
rect 466562 562046 466618 562102
rect 466686 562046 466742 562102
rect 466314 561922 466370 561978
rect 466438 561922 466494 561978
rect 466562 561922 466618 561978
rect 466686 561922 466742 561978
rect 466314 544294 466370 544350
rect 466438 544294 466494 544350
rect 466562 544294 466618 544350
rect 466686 544294 466742 544350
rect 466314 544170 466370 544226
rect 466438 544170 466494 544226
rect 466562 544170 466618 544226
rect 466686 544170 466742 544226
rect 466314 544046 466370 544102
rect 466438 544046 466494 544102
rect 466562 544046 466618 544102
rect 466686 544046 466742 544102
rect 466314 543922 466370 543978
rect 466438 543922 466494 543978
rect 466562 543922 466618 543978
rect 466686 543922 466742 543978
rect 466314 526294 466370 526350
rect 466438 526294 466494 526350
rect 466562 526294 466618 526350
rect 466686 526294 466742 526350
rect 466314 526170 466370 526226
rect 466438 526170 466494 526226
rect 466562 526170 466618 526226
rect 466686 526170 466742 526226
rect 466314 526046 466370 526102
rect 466438 526046 466494 526102
rect 466562 526046 466618 526102
rect 466686 526046 466742 526102
rect 466314 525922 466370 525978
rect 466438 525922 466494 525978
rect 466562 525922 466618 525978
rect 466686 525922 466742 525978
rect 466314 508294 466370 508350
rect 466438 508294 466494 508350
rect 466562 508294 466618 508350
rect 466686 508294 466742 508350
rect 466314 508170 466370 508226
rect 466438 508170 466494 508226
rect 466562 508170 466618 508226
rect 466686 508170 466742 508226
rect 466314 508046 466370 508102
rect 466438 508046 466494 508102
rect 466562 508046 466618 508102
rect 466686 508046 466742 508102
rect 466314 507922 466370 507978
rect 466438 507922 466494 507978
rect 466562 507922 466618 507978
rect 466686 507922 466742 507978
rect 466314 490294 466370 490350
rect 466438 490294 466494 490350
rect 466562 490294 466618 490350
rect 466686 490294 466742 490350
rect 466314 490170 466370 490226
rect 466438 490170 466494 490226
rect 466562 490170 466618 490226
rect 466686 490170 466742 490226
rect 466314 490046 466370 490102
rect 466438 490046 466494 490102
rect 466562 490046 466618 490102
rect 466686 490046 466742 490102
rect 466314 489922 466370 489978
rect 466438 489922 466494 489978
rect 466562 489922 466618 489978
rect 466686 489922 466742 489978
rect 466314 472294 466370 472350
rect 466438 472294 466494 472350
rect 466562 472294 466618 472350
rect 466686 472294 466742 472350
rect 466314 472170 466370 472226
rect 466438 472170 466494 472226
rect 466562 472170 466618 472226
rect 466686 472170 466742 472226
rect 466314 472046 466370 472102
rect 466438 472046 466494 472102
rect 466562 472046 466618 472102
rect 466686 472046 466742 472102
rect 466314 471922 466370 471978
rect 466438 471922 466494 471978
rect 466562 471922 466618 471978
rect 466686 471922 466742 471978
rect 466314 454294 466370 454350
rect 466438 454294 466494 454350
rect 466562 454294 466618 454350
rect 466686 454294 466742 454350
rect 466314 454170 466370 454226
rect 466438 454170 466494 454226
rect 466562 454170 466618 454226
rect 466686 454170 466742 454226
rect 466314 454046 466370 454102
rect 466438 454046 466494 454102
rect 466562 454046 466618 454102
rect 466686 454046 466742 454102
rect 466314 453922 466370 453978
rect 466438 453922 466494 453978
rect 466562 453922 466618 453978
rect 466686 453922 466742 453978
rect 466314 436294 466370 436350
rect 466438 436294 466494 436350
rect 466562 436294 466618 436350
rect 466686 436294 466742 436350
rect 466314 436170 466370 436226
rect 466438 436170 466494 436226
rect 466562 436170 466618 436226
rect 466686 436170 466742 436226
rect 466314 436046 466370 436102
rect 466438 436046 466494 436102
rect 466562 436046 466618 436102
rect 466686 436046 466742 436102
rect 466314 435922 466370 435978
rect 466438 435922 466494 435978
rect 466562 435922 466618 435978
rect 466686 435922 466742 435978
rect 466314 418294 466370 418350
rect 466438 418294 466494 418350
rect 466562 418294 466618 418350
rect 466686 418294 466742 418350
rect 466314 418170 466370 418226
rect 466438 418170 466494 418226
rect 466562 418170 466618 418226
rect 466686 418170 466742 418226
rect 466314 418046 466370 418102
rect 466438 418046 466494 418102
rect 466562 418046 466618 418102
rect 466686 418046 466742 418102
rect 466314 417922 466370 417978
rect 466438 417922 466494 417978
rect 466562 417922 466618 417978
rect 466686 417922 466742 417978
rect 466314 400294 466370 400350
rect 466438 400294 466494 400350
rect 466562 400294 466618 400350
rect 466686 400294 466742 400350
rect 466314 400170 466370 400226
rect 466438 400170 466494 400226
rect 466562 400170 466618 400226
rect 466686 400170 466742 400226
rect 466314 400046 466370 400102
rect 466438 400046 466494 400102
rect 466562 400046 466618 400102
rect 466686 400046 466742 400102
rect 466314 399922 466370 399978
rect 466438 399922 466494 399978
rect 466562 399922 466618 399978
rect 466686 399922 466742 399978
rect 466314 382294 466370 382350
rect 466438 382294 466494 382350
rect 466562 382294 466618 382350
rect 466686 382294 466742 382350
rect 466314 382170 466370 382226
rect 466438 382170 466494 382226
rect 466562 382170 466618 382226
rect 466686 382170 466742 382226
rect 466314 382046 466370 382102
rect 466438 382046 466494 382102
rect 466562 382046 466618 382102
rect 466686 382046 466742 382102
rect 466314 381922 466370 381978
rect 466438 381922 466494 381978
rect 466562 381922 466618 381978
rect 466686 381922 466742 381978
rect 466314 364294 466370 364350
rect 466438 364294 466494 364350
rect 466562 364294 466618 364350
rect 466686 364294 466742 364350
rect 466314 364170 466370 364226
rect 466438 364170 466494 364226
rect 466562 364170 466618 364226
rect 466686 364170 466742 364226
rect 466314 364046 466370 364102
rect 466438 364046 466494 364102
rect 466562 364046 466618 364102
rect 466686 364046 466742 364102
rect 466314 363922 466370 363978
rect 466438 363922 466494 363978
rect 466562 363922 466618 363978
rect 466686 363922 466742 363978
rect 466314 346294 466370 346350
rect 466438 346294 466494 346350
rect 466562 346294 466618 346350
rect 466686 346294 466742 346350
rect 466314 346170 466370 346226
rect 466438 346170 466494 346226
rect 466562 346170 466618 346226
rect 466686 346170 466742 346226
rect 466314 346046 466370 346102
rect 466438 346046 466494 346102
rect 466562 346046 466618 346102
rect 466686 346046 466742 346102
rect 466314 345922 466370 345978
rect 466438 345922 466494 345978
rect 466562 345922 466618 345978
rect 466686 345922 466742 345978
rect 466314 328294 466370 328350
rect 466438 328294 466494 328350
rect 466562 328294 466618 328350
rect 466686 328294 466742 328350
rect 466314 328170 466370 328226
rect 466438 328170 466494 328226
rect 466562 328170 466618 328226
rect 466686 328170 466742 328226
rect 466314 328046 466370 328102
rect 466438 328046 466494 328102
rect 466562 328046 466618 328102
rect 466686 328046 466742 328102
rect 466314 327922 466370 327978
rect 466438 327922 466494 327978
rect 466562 327922 466618 327978
rect 466686 327922 466742 327978
rect 439314 316294 439370 316350
rect 439438 316294 439494 316350
rect 439562 316294 439618 316350
rect 439686 316294 439742 316350
rect 439314 316170 439370 316226
rect 439438 316170 439494 316226
rect 439562 316170 439618 316226
rect 439686 316170 439742 316226
rect 439314 316046 439370 316102
rect 439438 316046 439494 316102
rect 439562 316046 439618 316102
rect 439686 316046 439742 316102
rect 439314 315922 439370 315978
rect 439438 315922 439494 315978
rect 439562 315922 439618 315978
rect 439686 315922 439742 315978
rect 439314 298294 439370 298350
rect 439438 298294 439494 298350
rect 439562 298294 439618 298350
rect 439686 298294 439742 298350
rect 439314 298170 439370 298226
rect 439438 298170 439494 298226
rect 439562 298170 439618 298226
rect 439686 298170 439742 298226
rect 439314 298046 439370 298102
rect 439438 298046 439494 298102
rect 439562 298046 439618 298102
rect 439686 298046 439742 298102
rect 439314 297922 439370 297978
rect 439438 297922 439494 297978
rect 439562 297922 439618 297978
rect 439686 297922 439742 297978
rect 440524 310922 440580 310978
rect 439314 280294 439370 280350
rect 439438 280294 439494 280350
rect 439562 280294 439618 280350
rect 439686 280294 439742 280350
rect 439314 280170 439370 280226
rect 439438 280170 439494 280226
rect 439562 280170 439618 280226
rect 439686 280170 439742 280226
rect 439314 280046 439370 280102
rect 439438 280046 439494 280102
rect 439562 280046 439618 280102
rect 439686 280046 439742 280102
rect 439314 279922 439370 279978
rect 439438 279922 439494 279978
rect 439562 279922 439618 279978
rect 439686 279922 439742 279978
rect 439314 262294 439370 262350
rect 439438 262294 439494 262350
rect 439562 262294 439618 262350
rect 439686 262294 439742 262350
rect 439314 262170 439370 262226
rect 439438 262170 439494 262226
rect 439562 262170 439618 262226
rect 439686 262170 439742 262226
rect 439314 262046 439370 262102
rect 439438 262046 439494 262102
rect 439562 262046 439618 262102
rect 439686 262046 439742 262102
rect 439314 261922 439370 261978
rect 439438 261922 439494 261978
rect 439562 261922 439618 261978
rect 439686 261922 439742 261978
rect 439314 244294 439370 244350
rect 439438 244294 439494 244350
rect 439562 244294 439618 244350
rect 439686 244294 439742 244350
rect 439314 244170 439370 244226
rect 439438 244170 439494 244226
rect 439562 244170 439618 244226
rect 439686 244170 439742 244226
rect 439314 244046 439370 244102
rect 439438 244046 439494 244102
rect 439562 244046 439618 244102
rect 439686 244046 439742 244102
rect 439314 243922 439370 243978
rect 439438 243922 439494 243978
rect 439562 243922 439618 243978
rect 439686 243922 439742 243978
rect 435594 238294 435650 238350
rect 435718 238294 435774 238350
rect 435842 238294 435898 238350
rect 435966 238294 436022 238350
rect 435594 238170 435650 238226
rect 435718 238170 435774 238226
rect 435842 238170 435898 238226
rect 435966 238170 436022 238226
rect 435594 238046 435650 238102
rect 435718 238046 435774 238102
rect 435842 238046 435898 238102
rect 435966 238046 436022 238102
rect 435594 237922 435650 237978
rect 435718 237922 435774 237978
rect 435842 237922 435898 237978
rect 435966 237922 436022 237978
rect 435594 220294 435650 220350
rect 435718 220294 435774 220350
rect 435842 220294 435898 220350
rect 435966 220294 436022 220350
rect 435594 220170 435650 220226
rect 435718 220170 435774 220226
rect 435842 220170 435898 220226
rect 435966 220170 436022 220226
rect 435594 220046 435650 220102
rect 435718 220046 435774 220102
rect 435842 220046 435898 220102
rect 435966 220046 436022 220102
rect 435594 219922 435650 219978
rect 435718 219922 435774 219978
rect 435842 219922 435898 219978
rect 435966 219922 436022 219978
rect 435594 202294 435650 202350
rect 435718 202294 435774 202350
rect 435842 202294 435898 202350
rect 435966 202294 436022 202350
rect 435594 202170 435650 202226
rect 435718 202170 435774 202226
rect 435842 202170 435898 202226
rect 435966 202170 436022 202226
rect 435594 202046 435650 202102
rect 435718 202046 435774 202102
rect 435842 202046 435898 202102
rect 435966 202046 436022 202102
rect 435594 201922 435650 201978
rect 435718 201922 435774 201978
rect 435842 201922 435898 201978
rect 435966 201922 436022 201978
rect 440188 242702 440244 242758
rect 439964 240002 440020 240058
rect 439314 226294 439370 226350
rect 439438 226294 439494 226350
rect 439562 226294 439618 226350
rect 439686 226294 439742 226350
rect 439314 226170 439370 226226
rect 439438 226170 439494 226226
rect 439562 226170 439618 226226
rect 439686 226170 439742 226226
rect 439314 226046 439370 226102
rect 439438 226046 439494 226102
rect 439562 226046 439618 226102
rect 439686 226046 439742 226102
rect 439314 225922 439370 225978
rect 439438 225922 439494 225978
rect 439562 225922 439618 225978
rect 439686 225922 439742 225978
rect 443548 216602 443604 216658
rect 466314 310294 466370 310350
rect 466438 310294 466494 310350
rect 466562 310294 466618 310350
rect 466686 310294 466742 310350
rect 466314 310170 466370 310226
rect 466438 310170 466494 310226
rect 466562 310170 466618 310226
rect 466686 310170 466742 310226
rect 466314 310046 466370 310102
rect 466438 310046 466494 310102
rect 466562 310046 466618 310102
rect 466686 310046 466742 310102
rect 466314 309922 466370 309978
rect 466438 309922 466494 309978
rect 466562 309922 466618 309978
rect 466686 309922 466742 309978
rect 445340 217322 445396 217378
rect 466314 292294 466370 292350
rect 466438 292294 466494 292350
rect 466562 292294 466618 292350
rect 466686 292294 466742 292350
rect 466314 292170 466370 292226
rect 466438 292170 466494 292226
rect 466562 292170 466618 292226
rect 466686 292170 466742 292226
rect 466314 292046 466370 292102
rect 466438 292046 466494 292102
rect 466562 292046 466618 292102
rect 466686 292046 466742 292102
rect 466314 291922 466370 291978
rect 466438 291922 466494 291978
rect 466562 291922 466618 291978
rect 466686 291922 466742 291978
rect 466314 274294 466370 274350
rect 466438 274294 466494 274350
rect 466562 274294 466618 274350
rect 466686 274294 466742 274350
rect 466314 274170 466370 274226
rect 466438 274170 466494 274226
rect 466562 274170 466618 274226
rect 466686 274170 466742 274226
rect 466314 274046 466370 274102
rect 466438 274046 466494 274102
rect 466562 274046 466618 274102
rect 466686 274046 466742 274102
rect 466314 273922 466370 273978
rect 466438 273922 466494 273978
rect 466562 273922 466618 273978
rect 466686 273922 466742 273978
rect 466314 256294 466370 256350
rect 466438 256294 466494 256350
rect 466562 256294 466618 256350
rect 466686 256294 466742 256350
rect 466314 256170 466370 256226
rect 466438 256170 466494 256226
rect 466562 256170 466618 256226
rect 466686 256170 466742 256226
rect 466314 256046 466370 256102
rect 466438 256046 466494 256102
rect 466562 256046 466618 256102
rect 466686 256046 466742 256102
rect 466314 255922 466370 255978
rect 466438 255922 466494 255978
rect 466562 255922 466618 255978
rect 466686 255922 466742 255978
rect 466314 238294 466370 238350
rect 466438 238294 466494 238350
rect 466562 238294 466618 238350
rect 466686 238294 466742 238350
rect 466314 238170 466370 238226
rect 466438 238170 466494 238226
rect 466562 238170 466618 238226
rect 466686 238170 466742 238226
rect 466314 238046 466370 238102
rect 466438 238046 466494 238102
rect 466562 238046 466618 238102
rect 466686 238046 466742 238102
rect 466314 237922 466370 237978
rect 466438 237922 466494 237978
rect 466562 237922 466618 237978
rect 466686 237922 466742 237978
rect 466314 220294 466370 220350
rect 466438 220294 466494 220350
rect 466562 220294 466618 220350
rect 466686 220294 466742 220350
rect 466314 220170 466370 220226
rect 466438 220170 466494 220226
rect 466562 220170 466618 220226
rect 466686 220170 466742 220226
rect 466314 220046 466370 220102
rect 466438 220046 466494 220102
rect 466562 220046 466618 220102
rect 466686 220046 466742 220102
rect 466314 219922 466370 219978
rect 466438 219922 466494 219978
rect 466562 219922 466618 219978
rect 466686 219922 466742 219978
rect 445228 216422 445284 216478
rect 439314 208294 439370 208350
rect 439438 208294 439494 208350
rect 439562 208294 439618 208350
rect 439686 208294 439742 208350
rect 439314 208170 439370 208226
rect 439438 208170 439494 208226
rect 439562 208170 439618 208226
rect 439686 208170 439742 208226
rect 439314 208046 439370 208102
rect 439438 208046 439494 208102
rect 439562 208046 439618 208102
rect 439686 208046 439742 208102
rect 439314 207922 439370 207978
rect 439438 207922 439494 207978
rect 439562 207922 439618 207978
rect 439686 207922 439742 207978
rect 435594 184294 435650 184350
rect 435718 184294 435774 184350
rect 435842 184294 435898 184350
rect 435966 184294 436022 184350
rect 435594 184170 435650 184226
rect 435718 184170 435774 184226
rect 435842 184170 435898 184226
rect 435966 184170 436022 184226
rect 435594 184046 435650 184102
rect 435718 184046 435774 184102
rect 435842 184046 435898 184102
rect 435966 184046 436022 184102
rect 435594 183922 435650 183978
rect 435718 183922 435774 183978
rect 435842 183922 435898 183978
rect 435966 183922 436022 183978
rect 435594 166294 435650 166350
rect 435718 166294 435774 166350
rect 435842 166294 435898 166350
rect 435966 166294 436022 166350
rect 435594 166170 435650 166226
rect 435718 166170 435774 166226
rect 435842 166170 435898 166226
rect 435966 166170 436022 166226
rect 435594 166046 435650 166102
rect 435718 166046 435774 166102
rect 435842 166046 435898 166102
rect 435966 166046 436022 166102
rect 435594 165922 435650 165978
rect 435718 165922 435774 165978
rect 435842 165922 435898 165978
rect 435966 165922 436022 165978
rect 435594 148294 435650 148350
rect 435718 148294 435774 148350
rect 435842 148294 435898 148350
rect 435966 148294 436022 148350
rect 435594 148170 435650 148226
rect 435718 148170 435774 148226
rect 435842 148170 435898 148226
rect 435966 148170 436022 148226
rect 435594 148046 435650 148102
rect 435718 148046 435774 148102
rect 435842 148046 435898 148102
rect 435966 148046 436022 148102
rect 435594 147922 435650 147978
rect 435718 147922 435774 147978
rect 435842 147922 435898 147978
rect 435966 147922 436022 147978
rect 442092 215882 442148 215938
rect 439314 190294 439370 190350
rect 439438 190294 439494 190350
rect 439562 190294 439618 190350
rect 439686 190294 439742 190350
rect 439314 190170 439370 190226
rect 439438 190170 439494 190226
rect 439562 190170 439618 190226
rect 439686 190170 439742 190226
rect 439314 190046 439370 190102
rect 439438 190046 439494 190102
rect 439562 190046 439618 190102
rect 439686 190046 439742 190102
rect 439314 189922 439370 189978
rect 439438 189922 439494 189978
rect 439562 189922 439618 189978
rect 439686 189922 439742 189978
rect 439314 172294 439370 172350
rect 439438 172294 439494 172350
rect 439562 172294 439618 172350
rect 439686 172294 439742 172350
rect 439314 172170 439370 172226
rect 439438 172170 439494 172226
rect 439562 172170 439618 172226
rect 439686 172170 439742 172226
rect 439314 172046 439370 172102
rect 439438 172046 439494 172102
rect 439562 172046 439618 172102
rect 439686 172046 439742 172102
rect 439314 171922 439370 171978
rect 439438 171922 439494 171978
rect 439562 171922 439618 171978
rect 439686 171922 439742 171978
rect 439314 154294 439370 154350
rect 439438 154294 439494 154350
rect 439562 154294 439618 154350
rect 439686 154294 439742 154350
rect 439314 154170 439370 154226
rect 439438 154170 439494 154226
rect 439562 154170 439618 154226
rect 439686 154170 439742 154226
rect 439314 154046 439370 154102
rect 439438 154046 439494 154102
rect 439562 154046 439618 154102
rect 439686 154046 439742 154102
rect 439314 153922 439370 153978
rect 439438 153922 439494 153978
rect 439562 153922 439618 153978
rect 439686 153922 439742 153978
rect 439314 136294 439370 136350
rect 439438 136294 439494 136350
rect 439562 136294 439618 136350
rect 439686 136294 439742 136350
rect 439314 136170 439370 136226
rect 439438 136170 439494 136226
rect 439562 136170 439618 136226
rect 439686 136170 439742 136226
rect 439314 136046 439370 136102
rect 439438 136046 439494 136102
rect 439562 136046 439618 136102
rect 439686 136046 439742 136102
rect 439314 135922 439370 135978
rect 439438 135922 439494 135978
rect 439562 135922 439618 135978
rect 439686 135922 439742 135978
rect 408594 118294 408650 118350
rect 408718 118294 408774 118350
rect 408842 118294 408898 118350
rect 408966 118294 409022 118350
rect 408594 118170 408650 118226
rect 408718 118170 408774 118226
rect 408842 118170 408898 118226
rect 408966 118170 409022 118226
rect 408594 118046 408650 118102
rect 408718 118046 408774 118102
rect 408842 118046 408898 118102
rect 408966 118046 409022 118102
rect 408594 117922 408650 117978
rect 408718 117922 408774 117978
rect 408842 117922 408898 117978
rect 408966 117922 409022 117978
rect 435594 130294 435650 130350
rect 435718 130294 435774 130350
rect 435842 130294 435898 130350
rect 435966 130294 436022 130350
rect 435594 130170 435650 130226
rect 435718 130170 435774 130226
rect 435842 130170 435898 130226
rect 435966 130170 436022 130226
rect 435594 130046 435650 130102
rect 435718 130046 435774 130102
rect 435842 130046 435898 130102
rect 435966 130046 436022 130102
rect 435594 129922 435650 129978
rect 435718 129922 435774 129978
rect 435842 129922 435898 129978
rect 435966 129922 436022 129978
rect 398188 115982 398244 116038
rect 415238 112294 415294 112350
rect 415362 112294 415418 112350
rect 415238 112170 415294 112226
rect 415362 112170 415418 112226
rect 415238 112046 415294 112102
rect 415362 112046 415418 112102
rect 415238 111922 415294 111978
rect 415362 111922 415418 111978
rect 399878 100294 399934 100350
rect 400002 100294 400058 100350
rect 399878 100170 399934 100226
rect 400002 100170 400058 100226
rect 399878 100046 399934 100102
rect 400002 100046 400058 100102
rect 399878 99922 399934 99978
rect 400002 99922 400058 99978
rect 415238 94294 415294 94350
rect 415362 94294 415418 94350
rect 415238 94170 415294 94226
rect 415362 94170 415418 94226
rect 415238 94046 415294 94102
rect 415362 94046 415418 94102
rect 415238 93922 415294 93978
rect 415362 93922 415418 93978
rect 399878 82294 399934 82350
rect 400002 82294 400058 82350
rect 399878 82170 399934 82226
rect 400002 82170 400058 82226
rect 399878 82046 399934 82102
rect 400002 82046 400058 82102
rect 399878 81922 399934 81978
rect 400002 81922 400058 81978
rect 415238 76294 415294 76350
rect 415362 76294 415418 76350
rect 415238 76170 415294 76226
rect 415362 76170 415418 76226
rect 415238 76046 415294 76102
rect 415362 76046 415418 76102
rect 415238 75922 415294 75978
rect 415362 75922 415418 75978
rect 399878 64294 399934 64350
rect 400002 64294 400058 64350
rect 399878 64170 399934 64226
rect 400002 64170 400058 64226
rect 399878 64046 399934 64102
rect 400002 64046 400058 64102
rect 399878 63922 399934 63978
rect 400002 63922 400058 63978
rect 415238 58294 415294 58350
rect 415362 58294 415418 58350
rect 415238 58170 415294 58226
rect 415362 58170 415418 58226
rect 415238 58046 415294 58102
rect 415362 58046 415418 58102
rect 415238 57922 415294 57978
rect 415362 57922 415418 57978
rect 404874 40294 404930 40350
rect 404998 40294 405054 40350
rect 405122 40294 405178 40350
rect 405246 40294 405302 40350
rect 377874 28294 377930 28350
rect 377998 28294 378054 28350
rect 378122 28294 378178 28350
rect 378246 28294 378302 28350
rect 377874 28170 377930 28226
rect 377998 28170 378054 28226
rect 378122 28170 378178 28226
rect 378246 28170 378302 28226
rect 377874 28046 377930 28102
rect 377998 28046 378054 28102
rect 378122 28046 378178 28102
rect 378246 28046 378302 28102
rect 377874 27922 377930 27978
rect 377998 27922 378054 27978
rect 378122 27922 378178 27978
rect 378246 27922 378302 27978
rect 377874 10294 377930 10350
rect 377998 10294 378054 10350
rect 378122 10294 378178 10350
rect 378246 10294 378302 10350
rect 377874 10170 377930 10226
rect 377998 10170 378054 10226
rect 378122 10170 378178 10226
rect 378246 10170 378302 10226
rect 377874 10046 377930 10102
rect 377998 10046 378054 10102
rect 378122 10046 378178 10102
rect 378246 10046 378302 10102
rect 377874 9922 377930 9978
rect 377998 9922 378054 9978
rect 378122 9922 378178 9978
rect 378246 9922 378302 9978
rect 377874 -1176 377930 -1120
rect 377998 -1176 378054 -1120
rect 378122 -1176 378178 -1120
rect 378246 -1176 378302 -1120
rect 377874 -1300 377930 -1244
rect 377998 -1300 378054 -1244
rect 378122 -1300 378178 -1244
rect 378246 -1300 378302 -1244
rect 377874 -1424 377930 -1368
rect 377998 -1424 378054 -1368
rect 378122 -1424 378178 -1368
rect 378246 -1424 378302 -1368
rect 377874 -1548 377930 -1492
rect 377998 -1548 378054 -1492
rect 378122 -1548 378178 -1492
rect 378246 -1548 378302 -1492
rect 404874 40170 404930 40226
rect 404998 40170 405054 40226
rect 405122 40170 405178 40226
rect 405246 40170 405302 40226
rect 404874 40046 404930 40102
rect 404998 40046 405054 40102
rect 405122 40046 405178 40102
rect 405246 40046 405302 40102
rect 404874 39922 404930 39978
rect 404998 39922 405054 39978
rect 405122 39922 405178 39978
rect 405246 39922 405302 39978
rect 408594 46142 408650 46198
rect 408718 46142 408774 46198
rect 408842 46142 408898 46198
rect 408966 46142 409022 46198
rect 408594 46018 408650 46074
rect 408718 46018 408774 46074
rect 408842 46018 408898 46074
rect 408966 46018 409022 46074
rect 408594 45894 408650 45950
rect 408718 45894 408774 45950
rect 408842 45894 408898 45950
rect 408966 45894 409022 45950
rect 419692 43652 419748 43678
rect 419692 43622 419748 43652
rect 430598 118294 430654 118350
rect 430722 118294 430778 118350
rect 430598 118170 430654 118226
rect 430722 118170 430778 118226
rect 430598 118046 430654 118102
rect 430722 118046 430778 118102
rect 430598 117922 430654 117978
rect 430722 117922 430778 117978
rect 430598 100294 430654 100350
rect 430722 100294 430778 100350
rect 430598 100170 430654 100226
rect 430722 100170 430778 100226
rect 430598 100046 430654 100102
rect 430722 100046 430778 100102
rect 430598 99922 430654 99978
rect 430722 99922 430778 99978
rect 430598 82294 430654 82350
rect 430722 82294 430778 82350
rect 430598 82170 430654 82226
rect 430722 82170 430778 82226
rect 430598 82046 430654 82102
rect 430722 82046 430778 82102
rect 430598 81922 430654 81978
rect 430722 81922 430778 81978
rect 430598 64294 430654 64350
rect 430722 64294 430778 64350
rect 430598 64170 430654 64226
rect 430722 64170 430778 64226
rect 430598 64046 430654 64102
rect 430722 64046 430778 64102
rect 430598 63922 430654 63978
rect 430722 63922 430778 63978
rect 435594 112294 435650 112350
rect 435718 112294 435774 112350
rect 435842 112294 435898 112350
rect 435966 112294 436022 112350
rect 435594 112170 435650 112226
rect 435718 112170 435774 112226
rect 435842 112170 435898 112226
rect 435966 112170 436022 112226
rect 435594 112046 435650 112102
rect 435718 112046 435774 112102
rect 435842 112046 435898 112102
rect 435966 112046 436022 112102
rect 435594 111922 435650 111978
rect 435718 111922 435774 111978
rect 435842 111922 435898 111978
rect 435966 111922 436022 111978
rect 435594 94294 435650 94350
rect 435718 94294 435774 94350
rect 435842 94294 435898 94350
rect 435966 94294 436022 94350
rect 435594 94170 435650 94226
rect 435718 94170 435774 94226
rect 435842 94170 435898 94226
rect 435966 94170 436022 94226
rect 435594 94046 435650 94102
rect 435718 94046 435774 94102
rect 435842 94046 435898 94102
rect 435966 94046 436022 94102
rect 435594 93922 435650 93978
rect 435718 93922 435774 93978
rect 435842 93922 435898 93978
rect 435966 93922 436022 93978
rect 435594 76294 435650 76350
rect 435718 76294 435774 76350
rect 435842 76294 435898 76350
rect 435966 76294 436022 76350
rect 435594 76170 435650 76226
rect 435718 76170 435774 76226
rect 435842 76170 435898 76226
rect 435966 76170 436022 76226
rect 435594 76046 435650 76102
rect 435718 76046 435774 76102
rect 435842 76046 435898 76102
rect 435966 76046 436022 76102
rect 435594 75922 435650 75978
rect 435718 75922 435774 75978
rect 435842 75922 435898 75978
rect 435966 75922 436022 75978
rect 435594 58294 435650 58350
rect 435718 58294 435774 58350
rect 435842 58294 435898 58350
rect 435966 58294 436022 58350
rect 435594 58170 435650 58226
rect 435718 58170 435774 58226
rect 435842 58170 435898 58226
rect 435966 58170 436022 58226
rect 435594 58046 435650 58102
rect 435718 58046 435774 58102
rect 435842 58046 435898 58102
rect 435966 58046 436022 58102
rect 435594 57922 435650 57978
rect 435718 57922 435774 57978
rect 435842 57922 435898 57978
rect 435966 57922 436022 57978
rect 435594 40294 435650 40350
rect 435718 40294 435774 40350
rect 435842 40294 435898 40350
rect 435966 40294 436022 40350
rect 435594 40170 435650 40226
rect 435718 40170 435774 40226
rect 435842 40170 435898 40226
rect 435966 40170 436022 40226
rect 435594 40046 435650 40102
rect 435718 40046 435774 40102
rect 435842 40046 435898 40102
rect 435966 40046 436022 40102
rect 435594 39922 435650 39978
rect 435718 39922 435774 39978
rect 435842 39922 435898 39978
rect 435966 39922 436022 39978
rect 409166 28294 409222 28350
rect 409290 28294 409346 28350
rect 409166 28170 409222 28226
rect 409290 28170 409346 28226
rect 409166 28046 409222 28102
rect 409290 28046 409346 28102
rect 409166 27922 409222 27978
rect 409290 27922 409346 27978
rect 404874 22294 404930 22350
rect 404998 22294 405054 22350
rect 405122 22294 405178 22350
rect 405246 22294 405302 22350
rect 404874 22170 404930 22226
rect 404998 22170 405054 22226
rect 405122 22170 405178 22226
rect 405246 22170 405302 22226
rect 404874 22046 404930 22102
rect 404998 22046 405054 22102
rect 405122 22046 405178 22102
rect 405246 22046 405302 22102
rect 404874 21922 404930 21978
rect 404998 21922 405054 21978
rect 405122 21922 405178 21978
rect 405246 21922 405302 21978
rect 435594 22294 435650 22350
rect 435718 22294 435774 22350
rect 435842 22294 435898 22350
rect 435966 22294 436022 22350
rect 435594 22170 435650 22226
rect 435718 22170 435774 22226
rect 435842 22170 435898 22226
rect 435966 22170 436022 22226
rect 435594 22046 435650 22102
rect 435718 22046 435774 22102
rect 435842 22046 435898 22102
rect 435966 22046 436022 22102
rect 435594 21922 435650 21978
rect 435718 21922 435774 21978
rect 435842 21922 435898 21978
rect 435966 21922 436022 21978
rect 409166 10294 409222 10350
rect 409290 10294 409346 10350
rect 409166 10170 409222 10226
rect 409290 10170 409346 10226
rect 409166 10046 409222 10102
rect 409290 10046 409346 10102
rect 409166 9922 409222 9978
rect 409290 9922 409346 9978
rect 404874 4294 404930 4350
rect 404998 4294 405054 4350
rect 405122 4294 405178 4350
rect 405246 4294 405302 4350
rect 404874 4170 404930 4226
rect 404998 4170 405054 4226
rect 405122 4170 405178 4226
rect 405246 4170 405302 4226
rect 404874 4046 404930 4102
rect 404998 4046 405054 4102
rect 405122 4046 405178 4102
rect 405246 4046 405302 4102
rect 404874 3922 404930 3978
rect 404998 3922 405054 3978
rect 405122 3922 405178 3978
rect 405246 3922 405302 3978
rect 404874 -216 404930 -160
rect 404998 -216 405054 -160
rect 405122 -216 405178 -160
rect 405246 -216 405302 -160
rect 404874 -340 404930 -284
rect 404998 -340 405054 -284
rect 405122 -340 405178 -284
rect 405246 -340 405302 -284
rect 404874 -464 404930 -408
rect 404998 -464 405054 -408
rect 405122 -464 405178 -408
rect 405246 -464 405302 -408
rect 404874 -588 404930 -532
rect 404998 -588 405054 -532
rect 405122 -588 405178 -532
rect 405246 -588 405302 -532
rect 435594 4294 435650 4350
rect 435718 4294 435774 4350
rect 435842 4294 435898 4350
rect 435966 4294 436022 4350
rect 435594 4170 435650 4226
rect 435718 4170 435774 4226
rect 435842 4170 435898 4226
rect 435966 4170 436022 4226
rect 435594 4046 435650 4102
rect 435718 4046 435774 4102
rect 435842 4046 435898 4102
rect 435966 4046 436022 4102
rect 435594 3922 435650 3978
rect 435718 3922 435774 3978
rect 435842 3922 435898 3978
rect 435966 3922 436022 3978
rect 439314 118294 439370 118350
rect 439438 118294 439494 118350
rect 439562 118294 439618 118350
rect 439686 118294 439742 118350
rect 439314 118170 439370 118226
rect 439438 118170 439494 118226
rect 439562 118170 439618 118226
rect 439686 118170 439742 118226
rect 439314 118046 439370 118102
rect 439438 118046 439494 118102
rect 439562 118046 439618 118102
rect 439686 118046 439742 118102
rect 439314 117922 439370 117978
rect 439438 117922 439494 117978
rect 439562 117922 439618 117978
rect 439686 117922 439742 117978
rect 439314 100294 439370 100350
rect 439438 100294 439494 100350
rect 439562 100294 439618 100350
rect 439686 100294 439742 100350
rect 439314 100170 439370 100226
rect 439438 100170 439494 100226
rect 439562 100170 439618 100226
rect 439686 100170 439742 100226
rect 439314 100046 439370 100102
rect 439438 100046 439494 100102
rect 439562 100046 439618 100102
rect 439686 100046 439742 100102
rect 439314 99922 439370 99978
rect 439438 99922 439494 99978
rect 439562 99922 439618 99978
rect 439686 99922 439742 99978
rect 439314 82294 439370 82350
rect 439438 82294 439494 82350
rect 439562 82294 439618 82350
rect 439686 82294 439742 82350
rect 439314 82170 439370 82226
rect 439438 82170 439494 82226
rect 439562 82170 439618 82226
rect 439686 82170 439742 82226
rect 439314 82046 439370 82102
rect 439438 82046 439494 82102
rect 439562 82046 439618 82102
rect 439686 82046 439742 82102
rect 441980 193202 442036 193258
rect 442540 214082 442596 214138
rect 442652 212462 442708 212518
rect 466314 202294 466370 202350
rect 466438 202294 466494 202350
rect 466562 202294 466618 202350
rect 466686 202294 466742 202350
rect 466314 202170 466370 202226
rect 466438 202170 466494 202226
rect 466562 202170 466618 202226
rect 466686 202170 466742 202226
rect 466314 202046 466370 202102
rect 466438 202046 466494 202102
rect 466562 202046 466618 202102
rect 466686 202046 466742 202102
rect 466314 201922 466370 201978
rect 466438 201922 466494 201978
rect 466562 201922 466618 201978
rect 466686 201922 466742 201978
rect 439314 81922 439370 81978
rect 439438 81922 439494 81978
rect 439562 81922 439618 81978
rect 439686 81922 439742 81978
rect 441868 133622 441924 133678
rect 441980 133442 442036 133498
rect 440636 120842 440692 120898
rect 440524 115802 440580 115858
rect 442092 117422 442148 117478
rect 443660 184922 443716 184978
rect 466314 184294 466370 184350
rect 466438 184294 466494 184350
rect 466562 184294 466618 184350
rect 466686 184294 466742 184350
rect 466314 184170 466370 184226
rect 466438 184170 466494 184226
rect 466562 184170 466618 184226
rect 466686 184170 466742 184226
rect 466314 184046 466370 184102
rect 466438 184046 466494 184102
rect 466562 184046 466618 184102
rect 466686 184046 466742 184102
rect 466314 183922 466370 183978
rect 466438 183922 466494 183978
rect 466562 183922 466618 183978
rect 466686 183922 466742 183978
rect 466314 166294 466370 166350
rect 466438 166294 466494 166350
rect 466562 166294 466618 166350
rect 466686 166294 466742 166350
rect 466314 166170 466370 166226
rect 466438 166170 466494 166226
rect 466562 166170 466618 166226
rect 466686 166170 466742 166226
rect 466314 166046 466370 166102
rect 466438 166046 466494 166102
rect 466562 166046 466618 166102
rect 466686 166046 466742 166102
rect 466314 165922 466370 165978
rect 466438 165922 466494 165978
rect 466562 165922 466618 165978
rect 466686 165922 466742 165978
rect 466314 148294 466370 148350
rect 466438 148294 466494 148350
rect 466562 148294 466618 148350
rect 466686 148294 466742 148350
rect 466314 148170 466370 148226
rect 466438 148170 466494 148226
rect 466562 148170 466618 148226
rect 466686 148170 466742 148226
rect 466314 148046 466370 148102
rect 466438 148046 466494 148102
rect 466562 148046 466618 148102
rect 466686 148046 466742 148102
rect 466314 147922 466370 147978
rect 466438 147922 466494 147978
rect 466562 147922 466618 147978
rect 466686 147922 466742 147978
rect 466314 130294 466370 130350
rect 466438 130294 466494 130350
rect 466562 130294 466618 130350
rect 466686 130294 466742 130350
rect 466314 130170 466370 130226
rect 466438 130170 466494 130226
rect 466562 130170 466618 130226
rect 466686 130170 466742 130226
rect 466314 130046 466370 130102
rect 466438 130046 466494 130102
rect 466562 130046 466618 130102
rect 466686 130046 466742 130102
rect 466314 129922 466370 129978
rect 466438 129922 466494 129978
rect 466562 129922 466618 129978
rect 466686 129922 466742 129978
rect 466314 112294 466370 112350
rect 466438 112294 466494 112350
rect 466562 112294 466618 112350
rect 466686 112294 466742 112350
rect 466314 112170 466370 112226
rect 466438 112170 466494 112226
rect 466562 112170 466618 112226
rect 466686 112170 466742 112226
rect 466314 112046 466370 112102
rect 466438 112046 466494 112102
rect 466562 112046 466618 112102
rect 466686 112046 466742 112102
rect 466314 111922 466370 111978
rect 466438 111922 466494 111978
rect 466562 111922 466618 111978
rect 466686 111922 466742 111978
rect 466314 94294 466370 94350
rect 466438 94294 466494 94350
rect 466562 94294 466618 94350
rect 466686 94294 466742 94350
rect 466314 94170 466370 94226
rect 466438 94170 466494 94226
rect 466562 94170 466618 94226
rect 466686 94170 466742 94226
rect 466314 94046 466370 94102
rect 466438 94046 466494 94102
rect 466562 94046 466618 94102
rect 466686 94046 466742 94102
rect 466314 93922 466370 93978
rect 466438 93922 466494 93978
rect 466562 93922 466618 93978
rect 466686 93922 466742 93978
rect 464518 76294 464574 76350
rect 464642 76294 464698 76350
rect 464518 76170 464574 76226
rect 464642 76170 464698 76226
rect 464518 76046 464574 76102
rect 464642 76046 464698 76102
rect 464518 75922 464574 75978
rect 464642 75922 464698 75978
rect 466314 76294 466370 76350
rect 466438 76294 466494 76350
rect 466562 76294 466618 76350
rect 466686 76294 466742 76350
rect 466314 76170 466370 76226
rect 466438 76170 466494 76226
rect 466562 76170 466618 76226
rect 466686 76170 466742 76226
rect 466314 76046 466370 76102
rect 466438 76046 466494 76102
rect 466562 76046 466618 76102
rect 466686 76046 466742 76102
rect 466314 75922 466370 75978
rect 466438 75922 466494 75978
rect 466562 75922 466618 75978
rect 466686 75922 466742 75978
rect 439314 64294 439370 64350
rect 439438 64294 439494 64350
rect 439562 64294 439618 64350
rect 439686 64294 439742 64350
rect 439314 64170 439370 64226
rect 439438 64170 439494 64226
rect 439562 64170 439618 64226
rect 439686 64170 439742 64226
rect 439314 64046 439370 64102
rect 439438 64046 439494 64102
rect 439562 64046 439618 64102
rect 439686 64046 439742 64102
rect 439314 63922 439370 63978
rect 439438 63922 439494 63978
rect 439562 63922 439618 63978
rect 439686 63922 439742 63978
rect 464518 58294 464574 58350
rect 464642 58294 464698 58350
rect 464518 58170 464574 58226
rect 464642 58170 464698 58226
rect 464518 58046 464574 58102
rect 464642 58046 464698 58102
rect 464518 57922 464574 57978
rect 464642 57922 464698 57978
rect 466314 58294 466370 58350
rect 466438 58294 466494 58350
rect 466562 58294 466618 58350
rect 466686 58294 466742 58350
rect 466314 58170 466370 58226
rect 466438 58170 466494 58226
rect 466562 58170 466618 58226
rect 466686 58170 466742 58226
rect 466314 58046 466370 58102
rect 466438 58046 466494 58102
rect 466562 58046 466618 58102
rect 466686 58046 466742 58102
rect 466314 57922 466370 57978
rect 466438 57922 466494 57978
rect 466562 57922 466618 57978
rect 466686 57922 466742 57978
rect 439314 46294 439370 46350
rect 439438 46294 439494 46350
rect 439562 46294 439618 46350
rect 439686 46294 439742 46350
rect 439314 46170 439370 46226
rect 439438 46170 439494 46226
rect 439562 46170 439618 46226
rect 439686 46170 439742 46226
rect 439314 46046 439370 46102
rect 439438 46046 439494 46102
rect 439562 46046 439618 46102
rect 439686 46046 439742 46102
rect 439314 45922 439370 45978
rect 439438 45922 439494 45978
rect 439562 45922 439618 45978
rect 439686 45922 439742 45978
rect 439314 28294 439370 28350
rect 439438 28294 439494 28350
rect 439562 28294 439618 28350
rect 439686 28294 439742 28350
rect 439314 28170 439370 28226
rect 439438 28170 439494 28226
rect 439562 28170 439618 28226
rect 439686 28170 439742 28226
rect 439314 28046 439370 28102
rect 439438 28046 439494 28102
rect 439562 28046 439618 28102
rect 439686 28046 439742 28102
rect 439314 27922 439370 27978
rect 439438 27922 439494 27978
rect 439562 27922 439618 27978
rect 439686 27922 439742 27978
rect 439314 10294 439370 10350
rect 439438 10294 439494 10350
rect 439562 10294 439618 10350
rect 439686 10294 439742 10350
rect 439314 10170 439370 10226
rect 439438 10170 439494 10226
rect 439562 10170 439618 10226
rect 439686 10170 439742 10226
rect 439314 10046 439370 10102
rect 439438 10046 439494 10102
rect 439562 10046 439618 10102
rect 439686 10046 439742 10102
rect 439314 9922 439370 9978
rect 439438 9922 439494 9978
rect 439562 9922 439618 9978
rect 439686 9922 439742 9978
rect 435594 -216 435650 -160
rect 435718 -216 435774 -160
rect 435842 -216 435898 -160
rect 435966 -216 436022 -160
rect 435594 -340 435650 -284
rect 435718 -340 435774 -284
rect 435842 -340 435898 -284
rect 435966 -340 436022 -284
rect 435594 -464 435650 -408
rect 435718 -464 435774 -408
rect 435842 -464 435898 -408
rect 435966 -464 436022 -408
rect 435594 -588 435650 -532
rect 435718 -588 435774 -532
rect 435842 -588 435898 -532
rect 435966 -588 436022 -532
rect 466314 40294 466370 40350
rect 466438 40294 466494 40350
rect 466562 40294 466618 40350
rect 466686 40294 466742 40350
rect 466314 40170 466370 40226
rect 466438 40170 466494 40226
rect 466562 40170 466618 40226
rect 466686 40170 466742 40226
rect 466314 40046 466370 40102
rect 466438 40046 466494 40102
rect 466562 40046 466618 40102
rect 466686 40046 466742 40102
rect 466314 39922 466370 39978
rect 466438 39922 466494 39978
rect 466562 39922 466618 39978
rect 466686 39922 466742 39978
rect 466314 22294 466370 22350
rect 466438 22294 466494 22350
rect 466562 22294 466618 22350
rect 466686 22294 466742 22350
rect 466314 22170 466370 22226
rect 466438 22170 466494 22226
rect 466562 22170 466618 22226
rect 466686 22170 466742 22226
rect 466314 22046 466370 22102
rect 466438 22046 466494 22102
rect 466562 22046 466618 22102
rect 466686 22046 466742 22102
rect 466314 21922 466370 21978
rect 466438 21922 466494 21978
rect 466562 21922 466618 21978
rect 466686 21922 466742 21978
rect 442988 5124 443044 5158
rect 442988 5102 443044 5124
rect 466314 4294 466370 4350
rect 466438 4294 466494 4350
rect 466562 4294 466618 4350
rect 466686 4294 466742 4350
rect 466314 4170 466370 4226
rect 466438 4170 466494 4226
rect 466562 4170 466618 4226
rect 466686 4170 466742 4226
rect 466314 4046 466370 4102
rect 466438 4046 466494 4102
rect 466562 4046 466618 4102
rect 466686 4046 466742 4102
rect 466314 3922 466370 3978
rect 466438 3922 466494 3978
rect 466562 3922 466618 3978
rect 466686 3922 466742 3978
rect 447692 3332 447748 3358
rect 447692 3302 447748 3332
rect 457100 422 457156 478
rect 439314 -1176 439370 -1120
rect 439438 -1176 439494 -1120
rect 439562 -1176 439618 -1120
rect 439686 -1176 439742 -1120
rect 439314 -1300 439370 -1244
rect 439438 -1300 439494 -1244
rect 439562 -1300 439618 -1244
rect 439686 -1300 439742 -1244
rect 439314 -1424 439370 -1368
rect 439438 -1424 439494 -1368
rect 439562 -1424 439618 -1368
rect 439686 -1424 439742 -1368
rect 439314 -1548 439370 -1492
rect 439438 -1548 439494 -1492
rect 439562 -1548 439618 -1492
rect 439686 -1548 439742 -1492
rect 466314 -216 466370 -160
rect 466438 -216 466494 -160
rect 466562 -216 466618 -160
rect 466686 -216 466742 -160
rect 466314 -340 466370 -284
rect 466438 -340 466494 -284
rect 466562 -340 466618 -284
rect 466686 -340 466742 -284
rect 466314 -464 466370 -408
rect 466438 -464 466494 -408
rect 466562 -464 466618 -408
rect 466686 -464 466742 -408
rect 466314 -588 466370 -532
rect 466438 -588 466494 -532
rect 466562 -588 466618 -532
rect 466686 -588 466742 -532
rect 470034 598116 470090 598172
rect 470158 598116 470214 598172
rect 470282 598116 470338 598172
rect 470406 598116 470462 598172
rect 470034 597992 470090 598048
rect 470158 597992 470214 598048
rect 470282 597992 470338 598048
rect 470406 597992 470462 598048
rect 470034 597868 470090 597924
rect 470158 597868 470214 597924
rect 470282 597868 470338 597924
rect 470406 597868 470462 597924
rect 470034 597744 470090 597800
rect 470158 597744 470214 597800
rect 470282 597744 470338 597800
rect 470406 597744 470462 597800
rect 470034 586294 470090 586350
rect 470158 586294 470214 586350
rect 470282 586294 470338 586350
rect 470406 586294 470462 586350
rect 470034 586170 470090 586226
rect 470158 586170 470214 586226
rect 470282 586170 470338 586226
rect 470406 586170 470462 586226
rect 470034 586046 470090 586102
rect 470158 586046 470214 586102
rect 470282 586046 470338 586102
rect 470406 586046 470462 586102
rect 470034 585922 470090 585978
rect 470158 585922 470214 585978
rect 470282 585922 470338 585978
rect 470406 585922 470462 585978
rect 470034 568294 470090 568350
rect 470158 568294 470214 568350
rect 470282 568294 470338 568350
rect 470406 568294 470462 568350
rect 470034 568170 470090 568226
rect 470158 568170 470214 568226
rect 470282 568170 470338 568226
rect 470406 568170 470462 568226
rect 470034 568046 470090 568102
rect 470158 568046 470214 568102
rect 470282 568046 470338 568102
rect 470406 568046 470462 568102
rect 470034 567922 470090 567978
rect 470158 567922 470214 567978
rect 470282 567922 470338 567978
rect 470406 567922 470462 567978
rect 470034 550294 470090 550350
rect 470158 550294 470214 550350
rect 470282 550294 470338 550350
rect 470406 550294 470462 550350
rect 470034 550170 470090 550226
rect 470158 550170 470214 550226
rect 470282 550170 470338 550226
rect 470406 550170 470462 550226
rect 470034 550046 470090 550102
rect 470158 550046 470214 550102
rect 470282 550046 470338 550102
rect 470406 550046 470462 550102
rect 470034 549922 470090 549978
rect 470158 549922 470214 549978
rect 470282 549922 470338 549978
rect 470406 549922 470462 549978
rect 470034 532294 470090 532350
rect 470158 532294 470214 532350
rect 470282 532294 470338 532350
rect 470406 532294 470462 532350
rect 470034 532170 470090 532226
rect 470158 532170 470214 532226
rect 470282 532170 470338 532226
rect 470406 532170 470462 532226
rect 470034 532046 470090 532102
rect 470158 532046 470214 532102
rect 470282 532046 470338 532102
rect 470406 532046 470462 532102
rect 470034 531922 470090 531978
rect 470158 531922 470214 531978
rect 470282 531922 470338 531978
rect 470406 531922 470462 531978
rect 470034 514294 470090 514350
rect 470158 514294 470214 514350
rect 470282 514294 470338 514350
rect 470406 514294 470462 514350
rect 470034 514170 470090 514226
rect 470158 514170 470214 514226
rect 470282 514170 470338 514226
rect 470406 514170 470462 514226
rect 470034 514046 470090 514102
rect 470158 514046 470214 514102
rect 470282 514046 470338 514102
rect 470406 514046 470462 514102
rect 470034 513922 470090 513978
rect 470158 513922 470214 513978
rect 470282 513922 470338 513978
rect 470406 513922 470462 513978
rect 470034 496294 470090 496350
rect 470158 496294 470214 496350
rect 470282 496294 470338 496350
rect 470406 496294 470462 496350
rect 470034 496170 470090 496226
rect 470158 496170 470214 496226
rect 470282 496170 470338 496226
rect 470406 496170 470462 496226
rect 470034 496046 470090 496102
rect 470158 496046 470214 496102
rect 470282 496046 470338 496102
rect 470406 496046 470462 496102
rect 470034 495922 470090 495978
rect 470158 495922 470214 495978
rect 470282 495922 470338 495978
rect 470406 495922 470462 495978
rect 470034 478294 470090 478350
rect 470158 478294 470214 478350
rect 470282 478294 470338 478350
rect 470406 478294 470462 478350
rect 470034 478170 470090 478226
rect 470158 478170 470214 478226
rect 470282 478170 470338 478226
rect 470406 478170 470462 478226
rect 470034 478046 470090 478102
rect 470158 478046 470214 478102
rect 470282 478046 470338 478102
rect 470406 478046 470462 478102
rect 470034 477922 470090 477978
rect 470158 477922 470214 477978
rect 470282 477922 470338 477978
rect 470406 477922 470462 477978
rect 470034 460294 470090 460350
rect 470158 460294 470214 460350
rect 470282 460294 470338 460350
rect 470406 460294 470462 460350
rect 470034 460170 470090 460226
rect 470158 460170 470214 460226
rect 470282 460170 470338 460226
rect 470406 460170 470462 460226
rect 470034 460046 470090 460102
rect 470158 460046 470214 460102
rect 470282 460046 470338 460102
rect 470406 460046 470462 460102
rect 470034 459922 470090 459978
rect 470158 459922 470214 459978
rect 470282 459922 470338 459978
rect 470406 459922 470462 459978
rect 470034 442294 470090 442350
rect 470158 442294 470214 442350
rect 470282 442294 470338 442350
rect 470406 442294 470462 442350
rect 470034 442170 470090 442226
rect 470158 442170 470214 442226
rect 470282 442170 470338 442226
rect 470406 442170 470462 442226
rect 470034 442046 470090 442102
rect 470158 442046 470214 442102
rect 470282 442046 470338 442102
rect 470406 442046 470462 442102
rect 470034 441922 470090 441978
rect 470158 441922 470214 441978
rect 470282 441922 470338 441978
rect 470406 441922 470462 441978
rect 470034 424294 470090 424350
rect 470158 424294 470214 424350
rect 470282 424294 470338 424350
rect 470406 424294 470462 424350
rect 470034 424170 470090 424226
rect 470158 424170 470214 424226
rect 470282 424170 470338 424226
rect 470406 424170 470462 424226
rect 470034 424046 470090 424102
rect 470158 424046 470214 424102
rect 470282 424046 470338 424102
rect 470406 424046 470462 424102
rect 470034 423922 470090 423978
rect 470158 423922 470214 423978
rect 470282 423922 470338 423978
rect 470406 423922 470462 423978
rect 470034 406294 470090 406350
rect 470158 406294 470214 406350
rect 470282 406294 470338 406350
rect 470406 406294 470462 406350
rect 470034 406170 470090 406226
rect 470158 406170 470214 406226
rect 470282 406170 470338 406226
rect 470406 406170 470462 406226
rect 470034 406046 470090 406102
rect 470158 406046 470214 406102
rect 470282 406046 470338 406102
rect 470406 406046 470462 406102
rect 470034 405922 470090 405978
rect 470158 405922 470214 405978
rect 470282 405922 470338 405978
rect 470406 405922 470462 405978
rect 470034 388294 470090 388350
rect 470158 388294 470214 388350
rect 470282 388294 470338 388350
rect 470406 388294 470462 388350
rect 470034 388170 470090 388226
rect 470158 388170 470214 388226
rect 470282 388170 470338 388226
rect 470406 388170 470462 388226
rect 470034 388046 470090 388102
rect 470158 388046 470214 388102
rect 470282 388046 470338 388102
rect 470406 388046 470462 388102
rect 470034 387922 470090 387978
rect 470158 387922 470214 387978
rect 470282 387922 470338 387978
rect 470406 387922 470462 387978
rect 470034 370294 470090 370350
rect 470158 370294 470214 370350
rect 470282 370294 470338 370350
rect 470406 370294 470462 370350
rect 470034 370170 470090 370226
rect 470158 370170 470214 370226
rect 470282 370170 470338 370226
rect 470406 370170 470462 370226
rect 470034 370046 470090 370102
rect 470158 370046 470214 370102
rect 470282 370046 470338 370102
rect 470406 370046 470462 370102
rect 470034 369922 470090 369978
rect 470158 369922 470214 369978
rect 470282 369922 470338 369978
rect 470406 369922 470462 369978
rect 470034 352294 470090 352350
rect 470158 352294 470214 352350
rect 470282 352294 470338 352350
rect 470406 352294 470462 352350
rect 470034 352170 470090 352226
rect 470158 352170 470214 352226
rect 470282 352170 470338 352226
rect 470406 352170 470462 352226
rect 470034 352046 470090 352102
rect 470158 352046 470214 352102
rect 470282 352046 470338 352102
rect 470406 352046 470462 352102
rect 470034 351922 470090 351978
rect 470158 351922 470214 351978
rect 470282 351922 470338 351978
rect 470406 351922 470462 351978
rect 470034 334294 470090 334350
rect 470158 334294 470214 334350
rect 470282 334294 470338 334350
rect 470406 334294 470462 334350
rect 470034 334170 470090 334226
rect 470158 334170 470214 334226
rect 470282 334170 470338 334226
rect 470406 334170 470462 334226
rect 470034 334046 470090 334102
rect 470158 334046 470214 334102
rect 470282 334046 470338 334102
rect 470406 334046 470462 334102
rect 470034 333922 470090 333978
rect 470158 333922 470214 333978
rect 470282 333922 470338 333978
rect 470406 333922 470462 333978
rect 470034 316294 470090 316350
rect 470158 316294 470214 316350
rect 470282 316294 470338 316350
rect 470406 316294 470462 316350
rect 470034 316170 470090 316226
rect 470158 316170 470214 316226
rect 470282 316170 470338 316226
rect 470406 316170 470462 316226
rect 470034 316046 470090 316102
rect 470158 316046 470214 316102
rect 470282 316046 470338 316102
rect 470406 316046 470462 316102
rect 470034 315922 470090 315978
rect 470158 315922 470214 315978
rect 470282 315922 470338 315978
rect 470406 315922 470462 315978
rect 470034 298294 470090 298350
rect 470158 298294 470214 298350
rect 470282 298294 470338 298350
rect 470406 298294 470462 298350
rect 470034 298170 470090 298226
rect 470158 298170 470214 298226
rect 470282 298170 470338 298226
rect 470406 298170 470462 298226
rect 470034 298046 470090 298102
rect 470158 298046 470214 298102
rect 470282 298046 470338 298102
rect 470406 298046 470462 298102
rect 470034 297922 470090 297978
rect 470158 297922 470214 297978
rect 470282 297922 470338 297978
rect 470406 297922 470462 297978
rect 470034 280294 470090 280350
rect 470158 280294 470214 280350
rect 470282 280294 470338 280350
rect 470406 280294 470462 280350
rect 470034 280170 470090 280226
rect 470158 280170 470214 280226
rect 470282 280170 470338 280226
rect 470406 280170 470462 280226
rect 470034 280046 470090 280102
rect 470158 280046 470214 280102
rect 470282 280046 470338 280102
rect 470406 280046 470462 280102
rect 470034 279922 470090 279978
rect 470158 279922 470214 279978
rect 470282 279922 470338 279978
rect 470406 279922 470462 279978
rect 470034 262294 470090 262350
rect 470158 262294 470214 262350
rect 470282 262294 470338 262350
rect 470406 262294 470462 262350
rect 470034 262170 470090 262226
rect 470158 262170 470214 262226
rect 470282 262170 470338 262226
rect 470406 262170 470462 262226
rect 470034 262046 470090 262102
rect 470158 262046 470214 262102
rect 470282 262046 470338 262102
rect 470406 262046 470462 262102
rect 470034 261922 470090 261978
rect 470158 261922 470214 261978
rect 470282 261922 470338 261978
rect 470406 261922 470462 261978
rect 470034 244294 470090 244350
rect 470158 244294 470214 244350
rect 470282 244294 470338 244350
rect 470406 244294 470462 244350
rect 470034 244170 470090 244226
rect 470158 244170 470214 244226
rect 470282 244170 470338 244226
rect 470406 244170 470462 244226
rect 470034 244046 470090 244102
rect 470158 244046 470214 244102
rect 470282 244046 470338 244102
rect 470406 244046 470462 244102
rect 470034 243922 470090 243978
rect 470158 243922 470214 243978
rect 470282 243922 470338 243978
rect 470406 243922 470462 243978
rect 470034 226294 470090 226350
rect 470158 226294 470214 226350
rect 470282 226294 470338 226350
rect 470406 226294 470462 226350
rect 470034 226170 470090 226226
rect 470158 226170 470214 226226
rect 470282 226170 470338 226226
rect 470406 226170 470462 226226
rect 470034 226046 470090 226102
rect 470158 226046 470214 226102
rect 470282 226046 470338 226102
rect 470406 226046 470462 226102
rect 470034 225922 470090 225978
rect 470158 225922 470214 225978
rect 470282 225922 470338 225978
rect 470406 225922 470462 225978
rect 470034 208294 470090 208350
rect 470158 208294 470214 208350
rect 470282 208294 470338 208350
rect 470406 208294 470462 208350
rect 470034 208170 470090 208226
rect 470158 208170 470214 208226
rect 470282 208170 470338 208226
rect 470406 208170 470462 208226
rect 470034 208046 470090 208102
rect 470158 208046 470214 208102
rect 470282 208046 470338 208102
rect 470406 208046 470462 208102
rect 470034 207922 470090 207978
rect 470158 207922 470214 207978
rect 470282 207922 470338 207978
rect 470406 207922 470462 207978
rect 470034 190294 470090 190350
rect 470158 190294 470214 190350
rect 470282 190294 470338 190350
rect 470406 190294 470462 190350
rect 470034 190170 470090 190226
rect 470158 190170 470214 190226
rect 470282 190170 470338 190226
rect 470406 190170 470462 190226
rect 470034 190046 470090 190102
rect 470158 190046 470214 190102
rect 470282 190046 470338 190102
rect 470406 190046 470462 190102
rect 470034 189922 470090 189978
rect 470158 189922 470214 189978
rect 470282 189922 470338 189978
rect 470406 189922 470462 189978
rect 470034 172294 470090 172350
rect 470158 172294 470214 172350
rect 470282 172294 470338 172350
rect 470406 172294 470462 172350
rect 470034 172170 470090 172226
rect 470158 172170 470214 172226
rect 470282 172170 470338 172226
rect 470406 172170 470462 172226
rect 470034 172046 470090 172102
rect 470158 172046 470214 172102
rect 470282 172046 470338 172102
rect 470406 172046 470462 172102
rect 470034 171922 470090 171978
rect 470158 171922 470214 171978
rect 470282 171922 470338 171978
rect 470406 171922 470462 171978
rect 470034 154294 470090 154350
rect 470158 154294 470214 154350
rect 470282 154294 470338 154350
rect 470406 154294 470462 154350
rect 470034 154170 470090 154226
rect 470158 154170 470214 154226
rect 470282 154170 470338 154226
rect 470406 154170 470462 154226
rect 470034 154046 470090 154102
rect 470158 154046 470214 154102
rect 470282 154046 470338 154102
rect 470406 154046 470462 154102
rect 470034 153922 470090 153978
rect 470158 153922 470214 153978
rect 470282 153922 470338 153978
rect 470406 153922 470462 153978
rect 470034 136294 470090 136350
rect 470158 136294 470214 136350
rect 470282 136294 470338 136350
rect 470406 136294 470462 136350
rect 470034 136170 470090 136226
rect 470158 136170 470214 136226
rect 470282 136170 470338 136226
rect 470406 136170 470462 136226
rect 470034 136046 470090 136102
rect 470158 136046 470214 136102
rect 470282 136046 470338 136102
rect 470406 136046 470462 136102
rect 470034 135922 470090 135978
rect 470158 135922 470214 135978
rect 470282 135922 470338 135978
rect 470406 135922 470462 135978
rect 470034 118294 470090 118350
rect 470158 118294 470214 118350
rect 470282 118294 470338 118350
rect 470406 118294 470462 118350
rect 470034 118170 470090 118226
rect 470158 118170 470214 118226
rect 470282 118170 470338 118226
rect 470406 118170 470462 118226
rect 470034 118046 470090 118102
rect 470158 118046 470214 118102
rect 470282 118046 470338 118102
rect 470406 118046 470462 118102
rect 470034 117922 470090 117978
rect 470158 117922 470214 117978
rect 470282 117922 470338 117978
rect 470406 117922 470462 117978
rect 470034 100294 470090 100350
rect 470158 100294 470214 100350
rect 470282 100294 470338 100350
rect 470406 100294 470462 100350
rect 470034 100170 470090 100226
rect 470158 100170 470214 100226
rect 470282 100170 470338 100226
rect 470406 100170 470462 100226
rect 470034 100046 470090 100102
rect 470158 100046 470214 100102
rect 470282 100046 470338 100102
rect 470406 100046 470462 100102
rect 470034 99922 470090 99978
rect 470158 99922 470214 99978
rect 470282 99922 470338 99978
rect 470406 99922 470462 99978
rect 497034 597156 497090 597212
rect 497158 597156 497214 597212
rect 497282 597156 497338 597212
rect 497406 597156 497462 597212
rect 497034 597032 497090 597088
rect 497158 597032 497214 597088
rect 497282 597032 497338 597088
rect 497406 597032 497462 597088
rect 497034 596908 497090 596964
rect 497158 596908 497214 596964
rect 497282 596908 497338 596964
rect 497406 596908 497462 596964
rect 497034 596784 497090 596840
rect 497158 596784 497214 596840
rect 497282 596784 497338 596840
rect 497406 596784 497462 596840
rect 497034 580294 497090 580350
rect 497158 580294 497214 580350
rect 497282 580294 497338 580350
rect 497406 580294 497462 580350
rect 497034 580170 497090 580226
rect 497158 580170 497214 580226
rect 497282 580170 497338 580226
rect 497406 580170 497462 580226
rect 497034 580046 497090 580102
rect 497158 580046 497214 580102
rect 497282 580046 497338 580102
rect 497406 580046 497462 580102
rect 497034 579922 497090 579978
rect 497158 579922 497214 579978
rect 497282 579922 497338 579978
rect 497406 579922 497462 579978
rect 497034 562294 497090 562350
rect 497158 562294 497214 562350
rect 497282 562294 497338 562350
rect 497406 562294 497462 562350
rect 497034 562170 497090 562226
rect 497158 562170 497214 562226
rect 497282 562170 497338 562226
rect 497406 562170 497462 562226
rect 497034 562046 497090 562102
rect 497158 562046 497214 562102
rect 497282 562046 497338 562102
rect 497406 562046 497462 562102
rect 497034 561922 497090 561978
rect 497158 561922 497214 561978
rect 497282 561922 497338 561978
rect 497406 561922 497462 561978
rect 497034 544294 497090 544350
rect 497158 544294 497214 544350
rect 497282 544294 497338 544350
rect 497406 544294 497462 544350
rect 497034 544170 497090 544226
rect 497158 544170 497214 544226
rect 497282 544170 497338 544226
rect 497406 544170 497462 544226
rect 497034 544046 497090 544102
rect 497158 544046 497214 544102
rect 497282 544046 497338 544102
rect 497406 544046 497462 544102
rect 497034 543922 497090 543978
rect 497158 543922 497214 543978
rect 497282 543922 497338 543978
rect 497406 543922 497462 543978
rect 497034 526294 497090 526350
rect 497158 526294 497214 526350
rect 497282 526294 497338 526350
rect 497406 526294 497462 526350
rect 497034 526170 497090 526226
rect 497158 526170 497214 526226
rect 497282 526170 497338 526226
rect 497406 526170 497462 526226
rect 497034 526046 497090 526102
rect 497158 526046 497214 526102
rect 497282 526046 497338 526102
rect 497406 526046 497462 526102
rect 497034 525922 497090 525978
rect 497158 525922 497214 525978
rect 497282 525922 497338 525978
rect 497406 525922 497462 525978
rect 497034 508294 497090 508350
rect 497158 508294 497214 508350
rect 497282 508294 497338 508350
rect 497406 508294 497462 508350
rect 497034 508170 497090 508226
rect 497158 508170 497214 508226
rect 497282 508170 497338 508226
rect 497406 508170 497462 508226
rect 497034 508046 497090 508102
rect 497158 508046 497214 508102
rect 497282 508046 497338 508102
rect 497406 508046 497462 508102
rect 497034 507922 497090 507978
rect 497158 507922 497214 507978
rect 497282 507922 497338 507978
rect 497406 507922 497462 507978
rect 497034 490294 497090 490350
rect 497158 490294 497214 490350
rect 497282 490294 497338 490350
rect 497406 490294 497462 490350
rect 497034 490170 497090 490226
rect 497158 490170 497214 490226
rect 497282 490170 497338 490226
rect 497406 490170 497462 490226
rect 497034 490046 497090 490102
rect 497158 490046 497214 490102
rect 497282 490046 497338 490102
rect 497406 490046 497462 490102
rect 497034 489922 497090 489978
rect 497158 489922 497214 489978
rect 497282 489922 497338 489978
rect 497406 489922 497462 489978
rect 497034 472294 497090 472350
rect 497158 472294 497214 472350
rect 497282 472294 497338 472350
rect 497406 472294 497462 472350
rect 497034 472170 497090 472226
rect 497158 472170 497214 472226
rect 497282 472170 497338 472226
rect 497406 472170 497462 472226
rect 497034 472046 497090 472102
rect 497158 472046 497214 472102
rect 497282 472046 497338 472102
rect 497406 472046 497462 472102
rect 497034 471922 497090 471978
rect 497158 471922 497214 471978
rect 497282 471922 497338 471978
rect 497406 471922 497462 471978
rect 497034 454294 497090 454350
rect 497158 454294 497214 454350
rect 497282 454294 497338 454350
rect 497406 454294 497462 454350
rect 497034 454170 497090 454226
rect 497158 454170 497214 454226
rect 497282 454170 497338 454226
rect 497406 454170 497462 454226
rect 497034 454046 497090 454102
rect 497158 454046 497214 454102
rect 497282 454046 497338 454102
rect 497406 454046 497462 454102
rect 497034 453922 497090 453978
rect 497158 453922 497214 453978
rect 497282 453922 497338 453978
rect 497406 453922 497462 453978
rect 497034 436294 497090 436350
rect 497158 436294 497214 436350
rect 497282 436294 497338 436350
rect 497406 436294 497462 436350
rect 497034 436170 497090 436226
rect 497158 436170 497214 436226
rect 497282 436170 497338 436226
rect 497406 436170 497462 436226
rect 497034 436046 497090 436102
rect 497158 436046 497214 436102
rect 497282 436046 497338 436102
rect 497406 436046 497462 436102
rect 497034 435922 497090 435978
rect 497158 435922 497214 435978
rect 497282 435922 497338 435978
rect 497406 435922 497462 435978
rect 497034 418294 497090 418350
rect 497158 418294 497214 418350
rect 497282 418294 497338 418350
rect 497406 418294 497462 418350
rect 497034 418170 497090 418226
rect 497158 418170 497214 418226
rect 497282 418170 497338 418226
rect 497406 418170 497462 418226
rect 497034 418046 497090 418102
rect 497158 418046 497214 418102
rect 497282 418046 497338 418102
rect 497406 418046 497462 418102
rect 497034 417922 497090 417978
rect 497158 417922 497214 417978
rect 497282 417922 497338 417978
rect 497406 417922 497462 417978
rect 497034 400294 497090 400350
rect 497158 400294 497214 400350
rect 497282 400294 497338 400350
rect 497406 400294 497462 400350
rect 497034 400170 497090 400226
rect 497158 400170 497214 400226
rect 497282 400170 497338 400226
rect 497406 400170 497462 400226
rect 497034 400046 497090 400102
rect 497158 400046 497214 400102
rect 497282 400046 497338 400102
rect 497406 400046 497462 400102
rect 497034 399922 497090 399978
rect 497158 399922 497214 399978
rect 497282 399922 497338 399978
rect 497406 399922 497462 399978
rect 497034 382294 497090 382350
rect 497158 382294 497214 382350
rect 497282 382294 497338 382350
rect 497406 382294 497462 382350
rect 497034 382170 497090 382226
rect 497158 382170 497214 382226
rect 497282 382170 497338 382226
rect 497406 382170 497462 382226
rect 497034 382046 497090 382102
rect 497158 382046 497214 382102
rect 497282 382046 497338 382102
rect 497406 382046 497462 382102
rect 497034 381922 497090 381978
rect 497158 381922 497214 381978
rect 497282 381922 497338 381978
rect 497406 381922 497462 381978
rect 497034 364294 497090 364350
rect 497158 364294 497214 364350
rect 497282 364294 497338 364350
rect 497406 364294 497462 364350
rect 497034 364170 497090 364226
rect 497158 364170 497214 364226
rect 497282 364170 497338 364226
rect 497406 364170 497462 364226
rect 497034 364046 497090 364102
rect 497158 364046 497214 364102
rect 497282 364046 497338 364102
rect 497406 364046 497462 364102
rect 497034 363922 497090 363978
rect 497158 363922 497214 363978
rect 497282 363922 497338 363978
rect 497406 363922 497462 363978
rect 497034 346294 497090 346350
rect 497158 346294 497214 346350
rect 497282 346294 497338 346350
rect 497406 346294 497462 346350
rect 497034 346170 497090 346226
rect 497158 346170 497214 346226
rect 497282 346170 497338 346226
rect 497406 346170 497462 346226
rect 497034 346046 497090 346102
rect 497158 346046 497214 346102
rect 497282 346046 497338 346102
rect 497406 346046 497462 346102
rect 497034 345922 497090 345978
rect 497158 345922 497214 345978
rect 497282 345922 497338 345978
rect 497406 345922 497462 345978
rect 497034 328294 497090 328350
rect 497158 328294 497214 328350
rect 497282 328294 497338 328350
rect 497406 328294 497462 328350
rect 497034 328170 497090 328226
rect 497158 328170 497214 328226
rect 497282 328170 497338 328226
rect 497406 328170 497462 328226
rect 497034 328046 497090 328102
rect 497158 328046 497214 328102
rect 497282 328046 497338 328102
rect 497406 328046 497462 328102
rect 497034 327922 497090 327978
rect 497158 327922 497214 327978
rect 497282 327922 497338 327978
rect 497406 327922 497462 327978
rect 497034 310294 497090 310350
rect 497158 310294 497214 310350
rect 497282 310294 497338 310350
rect 497406 310294 497462 310350
rect 497034 310170 497090 310226
rect 497158 310170 497214 310226
rect 497282 310170 497338 310226
rect 497406 310170 497462 310226
rect 497034 310046 497090 310102
rect 497158 310046 497214 310102
rect 497282 310046 497338 310102
rect 497406 310046 497462 310102
rect 497034 309922 497090 309978
rect 497158 309922 497214 309978
rect 497282 309922 497338 309978
rect 497406 309922 497462 309978
rect 497034 292294 497090 292350
rect 497158 292294 497214 292350
rect 497282 292294 497338 292350
rect 497406 292294 497462 292350
rect 497034 292170 497090 292226
rect 497158 292170 497214 292226
rect 497282 292170 497338 292226
rect 497406 292170 497462 292226
rect 497034 292046 497090 292102
rect 497158 292046 497214 292102
rect 497282 292046 497338 292102
rect 497406 292046 497462 292102
rect 497034 291922 497090 291978
rect 497158 291922 497214 291978
rect 497282 291922 497338 291978
rect 497406 291922 497462 291978
rect 497034 274294 497090 274350
rect 497158 274294 497214 274350
rect 497282 274294 497338 274350
rect 497406 274294 497462 274350
rect 497034 274170 497090 274226
rect 497158 274170 497214 274226
rect 497282 274170 497338 274226
rect 497406 274170 497462 274226
rect 497034 274046 497090 274102
rect 497158 274046 497214 274102
rect 497282 274046 497338 274102
rect 497406 274046 497462 274102
rect 497034 273922 497090 273978
rect 497158 273922 497214 273978
rect 497282 273922 497338 273978
rect 497406 273922 497462 273978
rect 497034 256294 497090 256350
rect 497158 256294 497214 256350
rect 497282 256294 497338 256350
rect 497406 256294 497462 256350
rect 497034 256170 497090 256226
rect 497158 256170 497214 256226
rect 497282 256170 497338 256226
rect 497406 256170 497462 256226
rect 497034 256046 497090 256102
rect 497158 256046 497214 256102
rect 497282 256046 497338 256102
rect 497406 256046 497462 256102
rect 497034 255922 497090 255978
rect 497158 255922 497214 255978
rect 497282 255922 497338 255978
rect 497406 255922 497462 255978
rect 497034 238294 497090 238350
rect 497158 238294 497214 238350
rect 497282 238294 497338 238350
rect 497406 238294 497462 238350
rect 497034 238170 497090 238226
rect 497158 238170 497214 238226
rect 497282 238170 497338 238226
rect 497406 238170 497462 238226
rect 497034 238046 497090 238102
rect 497158 238046 497214 238102
rect 497282 238046 497338 238102
rect 497406 238046 497462 238102
rect 497034 237922 497090 237978
rect 497158 237922 497214 237978
rect 497282 237922 497338 237978
rect 497406 237922 497462 237978
rect 497034 220294 497090 220350
rect 497158 220294 497214 220350
rect 497282 220294 497338 220350
rect 497406 220294 497462 220350
rect 497034 220170 497090 220226
rect 497158 220170 497214 220226
rect 497282 220170 497338 220226
rect 497406 220170 497462 220226
rect 497034 220046 497090 220102
rect 497158 220046 497214 220102
rect 497282 220046 497338 220102
rect 497406 220046 497462 220102
rect 497034 219922 497090 219978
rect 497158 219922 497214 219978
rect 497282 219922 497338 219978
rect 497406 219922 497462 219978
rect 497034 202294 497090 202350
rect 497158 202294 497214 202350
rect 497282 202294 497338 202350
rect 497406 202294 497462 202350
rect 497034 202170 497090 202226
rect 497158 202170 497214 202226
rect 497282 202170 497338 202226
rect 497406 202170 497462 202226
rect 497034 202046 497090 202102
rect 497158 202046 497214 202102
rect 497282 202046 497338 202102
rect 497406 202046 497462 202102
rect 497034 201922 497090 201978
rect 497158 201922 497214 201978
rect 497282 201922 497338 201978
rect 497406 201922 497462 201978
rect 497034 184294 497090 184350
rect 497158 184294 497214 184350
rect 497282 184294 497338 184350
rect 497406 184294 497462 184350
rect 497034 184170 497090 184226
rect 497158 184170 497214 184226
rect 497282 184170 497338 184226
rect 497406 184170 497462 184226
rect 497034 184046 497090 184102
rect 497158 184046 497214 184102
rect 497282 184046 497338 184102
rect 497406 184046 497462 184102
rect 497034 183922 497090 183978
rect 497158 183922 497214 183978
rect 497282 183922 497338 183978
rect 497406 183922 497462 183978
rect 497034 166294 497090 166350
rect 497158 166294 497214 166350
rect 497282 166294 497338 166350
rect 497406 166294 497462 166350
rect 497034 166170 497090 166226
rect 497158 166170 497214 166226
rect 497282 166170 497338 166226
rect 497406 166170 497462 166226
rect 497034 166046 497090 166102
rect 497158 166046 497214 166102
rect 497282 166046 497338 166102
rect 497406 166046 497462 166102
rect 497034 165922 497090 165978
rect 497158 165922 497214 165978
rect 497282 165922 497338 165978
rect 497406 165922 497462 165978
rect 497034 148294 497090 148350
rect 497158 148294 497214 148350
rect 497282 148294 497338 148350
rect 497406 148294 497462 148350
rect 497034 148170 497090 148226
rect 497158 148170 497214 148226
rect 497282 148170 497338 148226
rect 497406 148170 497462 148226
rect 497034 148046 497090 148102
rect 497158 148046 497214 148102
rect 497282 148046 497338 148102
rect 497406 148046 497462 148102
rect 497034 147922 497090 147978
rect 497158 147922 497214 147978
rect 497282 147922 497338 147978
rect 497406 147922 497462 147978
rect 497034 130294 497090 130350
rect 497158 130294 497214 130350
rect 497282 130294 497338 130350
rect 497406 130294 497462 130350
rect 497034 130170 497090 130226
rect 497158 130170 497214 130226
rect 497282 130170 497338 130226
rect 497406 130170 497462 130226
rect 497034 130046 497090 130102
rect 497158 130046 497214 130102
rect 497282 130046 497338 130102
rect 497406 130046 497462 130102
rect 497034 129922 497090 129978
rect 497158 129922 497214 129978
rect 497282 129922 497338 129978
rect 497406 129922 497462 129978
rect 497034 112294 497090 112350
rect 497158 112294 497214 112350
rect 497282 112294 497338 112350
rect 497406 112294 497462 112350
rect 497034 112170 497090 112226
rect 497158 112170 497214 112226
rect 497282 112170 497338 112226
rect 497406 112170 497462 112226
rect 497034 112046 497090 112102
rect 497158 112046 497214 112102
rect 497282 112046 497338 112102
rect 497406 112046 497462 112102
rect 497034 111922 497090 111978
rect 497158 111922 497214 111978
rect 497282 111922 497338 111978
rect 497406 111922 497462 111978
rect 497034 94294 497090 94350
rect 497158 94294 497214 94350
rect 497282 94294 497338 94350
rect 497406 94294 497462 94350
rect 497034 94170 497090 94226
rect 497158 94170 497214 94226
rect 497282 94170 497338 94226
rect 497406 94170 497462 94226
rect 497034 94046 497090 94102
rect 497158 94046 497214 94102
rect 497282 94046 497338 94102
rect 497406 94046 497462 94102
rect 497034 93922 497090 93978
rect 497158 93922 497214 93978
rect 497282 93922 497338 93978
rect 497406 93922 497462 93978
rect 470034 82294 470090 82350
rect 470158 82294 470214 82350
rect 470282 82294 470338 82350
rect 470406 82294 470462 82350
rect 470034 82170 470090 82226
rect 470158 82170 470214 82226
rect 470282 82170 470338 82226
rect 470406 82170 470462 82226
rect 470034 82046 470090 82102
rect 470158 82046 470214 82102
rect 470282 82046 470338 82102
rect 470406 82046 470462 82102
rect 470034 81922 470090 81978
rect 470158 81922 470214 81978
rect 470282 81922 470338 81978
rect 470406 81922 470462 81978
rect 479878 82294 479934 82350
rect 480002 82294 480058 82350
rect 479878 82170 479934 82226
rect 480002 82170 480058 82226
rect 479878 82046 479934 82102
rect 480002 82046 480058 82102
rect 479878 81922 479934 81978
rect 480002 81922 480058 81978
rect 495238 76294 495294 76350
rect 495362 76294 495418 76350
rect 495238 76170 495294 76226
rect 495362 76170 495418 76226
rect 495238 76046 495294 76102
rect 495362 76046 495418 76102
rect 495238 75922 495294 75978
rect 495362 75922 495418 75978
rect 497034 76294 497090 76350
rect 497158 76294 497214 76350
rect 497282 76294 497338 76350
rect 497406 76294 497462 76350
rect 497034 76170 497090 76226
rect 497158 76170 497214 76226
rect 497282 76170 497338 76226
rect 497406 76170 497462 76226
rect 497034 76046 497090 76102
rect 497158 76046 497214 76102
rect 497282 76046 497338 76102
rect 497406 76046 497462 76102
rect 497034 75922 497090 75978
rect 497158 75922 497214 75978
rect 497282 75922 497338 75978
rect 497406 75922 497462 75978
rect 470034 64294 470090 64350
rect 470158 64294 470214 64350
rect 470282 64294 470338 64350
rect 470406 64294 470462 64350
rect 470034 64170 470090 64226
rect 470158 64170 470214 64226
rect 470282 64170 470338 64226
rect 470406 64170 470462 64226
rect 470034 64046 470090 64102
rect 470158 64046 470214 64102
rect 470282 64046 470338 64102
rect 470406 64046 470462 64102
rect 470034 63922 470090 63978
rect 470158 63922 470214 63978
rect 470282 63922 470338 63978
rect 470406 63922 470462 63978
rect 479878 64294 479934 64350
rect 480002 64294 480058 64350
rect 479878 64170 479934 64226
rect 480002 64170 480058 64226
rect 479878 64046 479934 64102
rect 480002 64046 480058 64102
rect 479878 63922 479934 63978
rect 480002 63922 480058 63978
rect 495238 58294 495294 58350
rect 495362 58294 495418 58350
rect 495238 58170 495294 58226
rect 495362 58170 495418 58226
rect 495238 58046 495294 58102
rect 495362 58046 495418 58102
rect 495238 57922 495294 57978
rect 495362 57922 495418 57978
rect 497034 58294 497090 58350
rect 497158 58294 497214 58350
rect 497282 58294 497338 58350
rect 497406 58294 497462 58350
rect 497034 58170 497090 58226
rect 497158 58170 497214 58226
rect 497282 58170 497338 58226
rect 497406 58170 497462 58226
rect 497034 58046 497090 58102
rect 497158 58046 497214 58102
rect 497282 58046 497338 58102
rect 497406 58046 497462 58102
rect 497034 57922 497090 57978
rect 497158 57922 497214 57978
rect 497282 57922 497338 57978
rect 497406 57922 497462 57978
rect 470034 46294 470090 46350
rect 470158 46294 470214 46350
rect 470282 46294 470338 46350
rect 470406 46294 470462 46350
rect 470034 46170 470090 46226
rect 470158 46170 470214 46226
rect 470282 46170 470338 46226
rect 470406 46170 470462 46226
rect 470034 46046 470090 46102
rect 470158 46046 470214 46102
rect 470282 46046 470338 46102
rect 470406 46046 470462 46102
rect 470034 45922 470090 45978
rect 470158 45922 470214 45978
rect 470282 45922 470338 45978
rect 470406 45922 470462 45978
rect 470034 28294 470090 28350
rect 470158 28294 470214 28350
rect 470282 28294 470338 28350
rect 470406 28294 470462 28350
rect 470034 28170 470090 28226
rect 470158 28170 470214 28226
rect 470282 28170 470338 28226
rect 470406 28170 470462 28226
rect 470034 28046 470090 28102
rect 470158 28046 470214 28102
rect 470282 28046 470338 28102
rect 470406 28046 470462 28102
rect 470034 27922 470090 27978
rect 470158 27922 470214 27978
rect 470282 27922 470338 27978
rect 470406 27922 470462 27978
rect 497034 40294 497090 40350
rect 497158 40294 497214 40350
rect 497282 40294 497338 40350
rect 497406 40294 497462 40350
rect 497034 40170 497090 40226
rect 497158 40170 497214 40226
rect 497282 40170 497338 40226
rect 497406 40170 497462 40226
rect 497034 40046 497090 40102
rect 497158 40046 497214 40102
rect 497282 40046 497338 40102
rect 497406 40046 497462 40102
rect 497034 39922 497090 39978
rect 497158 39922 497214 39978
rect 497282 39922 497338 39978
rect 497406 39922 497462 39978
rect 473818 22294 473874 22350
rect 473942 22294 473998 22350
rect 473818 22170 473874 22226
rect 473942 22170 473998 22226
rect 473818 22046 473874 22102
rect 473942 22046 473998 22102
rect 473818 21922 473874 21978
rect 473942 21922 473998 21978
rect 497034 22294 497090 22350
rect 497158 22294 497214 22350
rect 497282 22294 497338 22350
rect 497406 22294 497462 22350
rect 497034 22170 497090 22226
rect 497158 22170 497214 22226
rect 497282 22170 497338 22226
rect 497406 22170 497462 22226
rect 497034 22046 497090 22102
rect 497158 22046 497214 22102
rect 497282 22046 497338 22102
rect 497406 22046 497462 22102
rect 497034 21922 497090 21978
rect 497158 21922 497214 21978
rect 497282 21922 497338 21978
rect 497406 21922 497462 21978
rect 470034 10294 470090 10350
rect 470158 10294 470214 10350
rect 470282 10294 470338 10350
rect 470406 10294 470462 10350
rect 470034 10170 470090 10226
rect 470158 10170 470214 10226
rect 470282 10170 470338 10226
rect 470406 10170 470462 10226
rect 470034 10046 470090 10102
rect 470158 10046 470214 10102
rect 470282 10046 470338 10102
rect 470406 10046 470462 10102
rect 470034 9922 470090 9978
rect 470158 9922 470214 9978
rect 470282 9922 470338 9978
rect 470406 9922 470462 9978
rect 475468 5282 475524 5338
rect 494956 5102 495012 5158
rect 500754 598116 500810 598172
rect 500878 598116 500934 598172
rect 501002 598116 501058 598172
rect 501126 598116 501182 598172
rect 500754 597992 500810 598048
rect 500878 597992 500934 598048
rect 501002 597992 501058 598048
rect 501126 597992 501182 598048
rect 500754 597868 500810 597924
rect 500878 597868 500934 597924
rect 501002 597868 501058 597924
rect 501126 597868 501182 597924
rect 500754 597744 500810 597800
rect 500878 597744 500934 597800
rect 501002 597744 501058 597800
rect 501126 597744 501182 597800
rect 500754 586294 500810 586350
rect 500878 586294 500934 586350
rect 501002 586294 501058 586350
rect 501126 586294 501182 586350
rect 500754 586170 500810 586226
rect 500878 586170 500934 586226
rect 501002 586170 501058 586226
rect 501126 586170 501182 586226
rect 500754 586046 500810 586102
rect 500878 586046 500934 586102
rect 501002 586046 501058 586102
rect 501126 586046 501182 586102
rect 500754 585922 500810 585978
rect 500878 585922 500934 585978
rect 501002 585922 501058 585978
rect 501126 585922 501182 585978
rect 500754 568294 500810 568350
rect 500878 568294 500934 568350
rect 501002 568294 501058 568350
rect 501126 568294 501182 568350
rect 500754 568170 500810 568226
rect 500878 568170 500934 568226
rect 501002 568170 501058 568226
rect 501126 568170 501182 568226
rect 500754 568046 500810 568102
rect 500878 568046 500934 568102
rect 501002 568046 501058 568102
rect 501126 568046 501182 568102
rect 500754 567922 500810 567978
rect 500878 567922 500934 567978
rect 501002 567922 501058 567978
rect 501126 567922 501182 567978
rect 500754 550294 500810 550350
rect 500878 550294 500934 550350
rect 501002 550294 501058 550350
rect 501126 550294 501182 550350
rect 500754 550170 500810 550226
rect 500878 550170 500934 550226
rect 501002 550170 501058 550226
rect 501126 550170 501182 550226
rect 500754 550046 500810 550102
rect 500878 550046 500934 550102
rect 501002 550046 501058 550102
rect 501126 550046 501182 550102
rect 500754 549922 500810 549978
rect 500878 549922 500934 549978
rect 501002 549922 501058 549978
rect 501126 549922 501182 549978
rect 500754 532294 500810 532350
rect 500878 532294 500934 532350
rect 501002 532294 501058 532350
rect 501126 532294 501182 532350
rect 500754 532170 500810 532226
rect 500878 532170 500934 532226
rect 501002 532170 501058 532226
rect 501126 532170 501182 532226
rect 500754 532046 500810 532102
rect 500878 532046 500934 532102
rect 501002 532046 501058 532102
rect 501126 532046 501182 532102
rect 500754 531922 500810 531978
rect 500878 531922 500934 531978
rect 501002 531922 501058 531978
rect 501126 531922 501182 531978
rect 500754 514294 500810 514350
rect 500878 514294 500934 514350
rect 501002 514294 501058 514350
rect 501126 514294 501182 514350
rect 500754 514170 500810 514226
rect 500878 514170 500934 514226
rect 501002 514170 501058 514226
rect 501126 514170 501182 514226
rect 500754 514046 500810 514102
rect 500878 514046 500934 514102
rect 501002 514046 501058 514102
rect 501126 514046 501182 514102
rect 500754 513922 500810 513978
rect 500878 513922 500934 513978
rect 501002 513922 501058 513978
rect 501126 513922 501182 513978
rect 500754 496294 500810 496350
rect 500878 496294 500934 496350
rect 501002 496294 501058 496350
rect 501126 496294 501182 496350
rect 500754 496170 500810 496226
rect 500878 496170 500934 496226
rect 501002 496170 501058 496226
rect 501126 496170 501182 496226
rect 500754 496046 500810 496102
rect 500878 496046 500934 496102
rect 501002 496046 501058 496102
rect 501126 496046 501182 496102
rect 500754 495922 500810 495978
rect 500878 495922 500934 495978
rect 501002 495922 501058 495978
rect 501126 495922 501182 495978
rect 500754 478294 500810 478350
rect 500878 478294 500934 478350
rect 501002 478294 501058 478350
rect 501126 478294 501182 478350
rect 500754 478170 500810 478226
rect 500878 478170 500934 478226
rect 501002 478170 501058 478226
rect 501126 478170 501182 478226
rect 500754 478046 500810 478102
rect 500878 478046 500934 478102
rect 501002 478046 501058 478102
rect 501126 478046 501182 478102
rect 500754 477922 500810 477978
rect 500878 477922 500934 477978
rect 501002 477922 501058 477978
rect 501126 477922 501182 477978
rect 500754 460294 500810 460350
rect 500878 460294 500934 460350
rect 501002 460294 501058 460350
rect 501126 460294 501182 460350
rect 500754 460170 500810 460226
rect 500878 460170 500934 460226
rect 501002 460170 501058 460226
rect 501126 460170 501182 460226
rect 500754 460046 500810 460102
rect 500878 460046 500934 460102
rect 501002 460046 501058 460102
rect 501126 460046 501182 460102
rect 500754 459922 500810 459978
rect 500878 459922 500934 459978
rect 501002 459922 501058 459978
rect 501126 459922 501182 459978
rect 500754 442294 500810 442350
rect 500878 442294 500934 442350
rect 501002 442294 501058 442350
rect 501126 442294 501182 442350
rect 500754 442170 500810 442226
rect 500878 442170 500934 442226
rect 501002 442170 501058 442226
rect 501126 442170 501182 442226
rect 500754 442046 500810 442102
rect 500878 442046 500934 442102
rect 501002 442046 501058 442102
rect 501126 442046 501182 442102
rect 500754 441922 500810 441978
rect 500878 441922 500934 441978
rect 501002 441922 501058 441978
rect 501126 441922 501182 441978
rect 500754 424294 500810 424350
rect 500878 424294 500934 424350
rect 501002 424294 501058 424350
rect 501126 424294 501182 424350
rect 500754 424170 500810 424226
rect 500878 424170 500934 424226
rect 501002 424170 501058 424226
rect 501126 424170 501182 424226
rect 500754 424046 500810 424102
rect 500878 424046 500934 424102
rect 501002 424046 501058 424102
rect 501126 424046 501182 424102
rect 500754 423922 500810 423978
rect 500878 423922 500934 423978
rect 501002 423922 501058 423978
rect 501126 423922 501182 423978
rect 500754 406294 500810 406350
rect 500878 406294 500934 406350
rect 501002 406294 501058 406350
rect 501126 406294 501182 406350
rect 500754 406170 500810 406226
rect 500878 406170 500934 406226
rect 501002 406170 501058 406226
rect 501126 406170 501182 406226
rect 500754 406046 500810 406102
rect 500878 406046 500934 406102
rect 501002 406046 501058 406102
rect 501126 406046 501182 406102
rect 500754 405922 500810 405978
rect 500878 405922 500934 405978
rect 501002 405922 501058 405978
rect 501126 405922 501182 405978
rect 527754 597156 527810 597212
rect 527878 597156 527934 597212
rect 528002 597156 528058 597212
rect 528126 597156 528182 597212
rect 527754 597032 527810 597088
rect 527878 597032 527934 597088
rect 528002 597032 528058 597088
rect 528126 597032 528182 597088
rect 527754 596908 527810 596964
rect 527878 596908 527934 596964
rect 528002 596908 528058 596964
rect 528126 596908 528182 596964
rect 527754 596784 527810 596840
rect 527878 596784 527934 596840
rect 528002 596784 528058 596840
rect 528126 596784 528182 596840
rect 527754 580294 527810 580350
rect 527878 580294 527934 580350
rect 528002 580294 528058 580350
rect 528126 580294 528182 580350
rect 527754 580170 527810 580226
rect 527878 580170 527934 580226
rect 528002 580170 528058 580226
rect 528126 580170 528182 580226
rect 527754 580046 527810 580102
rect 527878 580046 527934 580102
rect 528002 580046 528058 580102
rect 528126 580046 528182 580102
rect 527754 579922 527810 579978
rect 527878 579922 527934 579978
rect 528002 579922 528058 579978
rect 528126 579922 528182 579978
rect 527754 562294 527810 562350
rect 527878 562294 527934 562350
rect 528002 562294 528058 562350
rect 528126 562294 528182 562350
rect 527754 562170 527810 562226
rect 527878 562170 527934 562226
rect 528002 562170 528058 562226
rect 528126 562170 528182 562226
rect 527754 562046 527810 562102
rect 527878 562046 527934 562102
rect 528002 562046 528058 562102
rect 528126 562046 528182 562102
rect 527754 561922 527810 561978
rect 527878 561922 527934 561978
rect 528002 561922 528058 561978
rect 528126 561922 528182 561978
rect 527754 544294 527810 544350
rect 527878 544294 527934 544350
rect 528002 544294 528058 544350
rect 528126 544294 528182 544350
rect 527754 544170 527810 544226
rect 527878 544170 527934 544226
rect 528002 544170 528058 544226
rect 528126 544170 528182 544226
rect 527754 544046 527810 544102
rect 527878 544046 527934 544102
rect 528002 544046 528058 544102
rect 528126 544046 528182 544102
rect 527754 543922 527810 543978
rect 527878 543922 527934 543978
rect 528002 543922 528058 543978
rect 528126 543922 528182 543978
rect 527754 526294 527810 526350
rect 527878 526294 527934 526350
rect 528002 526294 528058 526350
rect 528126 526294 528182 526350
rect 527754 526170 527810 526226
rect 527878 526170 527934 526226
rect 528002 526170 528058 526226
rect 528126 526170 528182 526226
rect 527754 526046 527810 526102
rect 527878 526046 527934 526102
rect 528002 526046 528058 526102
rect 528126 526046 528182 526102
rect 527754 525922 527810 525978
rect 527878 525922 527934 525978
rect 528002 525922 528058 525978
rect 528126 525922 528182 525978
rect 527754 508294 527810 508350
rect 527878 508294 527934 508350
rect 528002 508294 528058 508350
rect 528126 508294 528182 508350
rect 527754 508170 527810 508226
rect 527878 508170 527934 508226
rect 528002 508170 528058 508226
rect 528126 508170 528182 508226
rect 527754 508046 527810 508102
rect 527878 508046 527934 508102
rect 528002 508046 528058 508102
rect 528126 508046 528182 508102
rect 527754 507922 527810 507978
rect 527878 507922 527934 507978
rect 528002 507922 528058 507978
rect 528126 507922 528182 507978
rect 527754 490294 527810 490350
rect 527878 490294 527934 490350
rect 528002 490294 528058 490350
rect 528126 490294 528182 490350
rect 527754 490170 527810 490226
rect 527878 490170 527934 490226
rect 528002 490170 528058 490226
rect 528126 490170 528182 490226
rect 527754 490046 527810 490102
rect 527878 490046 527934 490102
rect 528002 490046 528058 490102
rect 528126 490046 528182 490102
rect 527754 489922 527810 489978
rect 527878 489922 527934 489978
rect 528002 489922 528058 489978
rect 528126 489922 528182 489978
rect 527754 472294 527810 472350
rect 527878 472294 527934 472350
rect 528002 472294 528058 472350
rect 528126 472294 528182 472350
rect 527754 472170 527810 472226
rect 527878 472170 527934 472226
rect 528002 472170 528058 472226
rect 528126 472170 528182 472226
rect 527754 472046 527810 472102
rect 527878 472046 527934 472102
rect 528002 472046 528058 472102
rect 528126 472046 528182 472102
rect 527754 471922 527810 471978
rect 527878 471922 527934 471978
rect 528002 471922 528058 471978
rect 528126 471922 528182 471978
rect 527754 454294 527810 454350
rect 527878 454294 527934 454350
rect 528002 454294 528058 454350
rect 528126 454294 528182 454350
rect 527754 454170 527810 454226
rect 527878 454170 527934 454226
rect 528002 454170 528058 454226
rect 528126 454170 528182 454226
rect 527754 454046 527810 454102
rect 527878 454046 527934 454102
rect 528002 454046 528058 454102
rect 528126 454046 528182 454102
rect 527754 453922 527810 453978
rect 527878 453922 527934 453978
rect 528002 453922 528058 453978
rect 528126 453922 528182 453978
rect 527754 436294 527810 436350
rect 527878 436294 527934 436350
rect 528002 436294 528058 436350
rect 528126 436294 528182 436350
rect 527754 436170 527810 436226
rect 527878 436170 527934 436226
rect 528002 436170 528058 436226
rect 528126 436170 528182 436226
rect 527754 436046 527810 436102
rect 527878 436046 527934 436102
rect 528002 436046 528058 436102
rect 528126 436046 528182 436102
rect 527754 435922 527810 435978
rect 527878 435922 527934 435978
rect 528002 435922 528058 435978
rect 528126 435922 528182 435978
rect 527754 418294 527810 418350
rect 527878 418294 527934 418350
rect 528002 418294 528058 418350
rect 528126 418294 528182 418350
rect 527754 418170 527810 418226
rect 527878 418170 527934 418226
rect 528002 418170 528058 418226
rect 528126 418170 528182 418226
rect 527754 418046 527810 418102
rect 527878 418046 527934 418102
rect 528002 418046 528058 418102
rect 528126 418046 528182 418102
rect 527754 417922 527810 417978
rect 527878 417922 527934 417978
rect 528002 417922 528058 417978
rect 528126 417922 528182 417978
rect 527754 400294 527810 400350
rect 527878 400294 527934 400350
rect 528002 400294 528058 400350
rect 528126 400294 528182 400350
rect 527754 400170 527810 400226
rect 527878 400170 527934 400226
rect 528002 400170 528058 400226
rect 528126 400170 528182 400226
rect 527754 400046 527810 400102
rect 527878 400046 527934 400102
rect 528002 400046 528058 400102
rect 528126 400046 528182 400102
rect 527754 399922 527810 399978
rect 527878 399922 527934 399978
rect 528002 399922 528058 399978
rect 528126 399922 528182 399978
rect 500754 388294 500810 388350
rect 500878 388294 500934 388350
rect 501002 388294 501058 388350
rect 501126 388294 501182 388350
rect 500754 388170 500810 388226
rect 500878 388170 500934 388226
rect 501002 388170 501058 388226
rect 501126 388170 501182 388226
rect 500754 388046 500810 388102
rect 500878 388046 500934 388102
rect 501002 388046 501058 388102
rect 501126 388046 501182 388102
rect 500754 387922 500810 387978
rect 500878 387922 500934 387978
rect 501002 387922 501058 387978
rect 501126 387922 501182 387978
rect 500754 370294 500810 370350
rect 500878 370294 500934 370350
rect 501002 370294 501058 370350
rect 501126 370294 501182 370350
rect 500754 370170 500810 370226
rect 500878 370170 500934 370226
rect 501002 370170 501058 370226
rect 501126 370170 501182 370226
rect 500754 370046 500810 370102
rect 500878 370046 500934 370102
rect 501002 370046 501058 370102
rect 501126 370046 501182 370102
rect 500754 369922 500810 369978
rect 500878 369922 500934 369978
rect 501002 369922 501058 369978
rect 501126 369922 501182 369978
rect 500754 352294 500810 352350
rect 500878 352294 500934 352350
rect 501002 352294 501058 352350
rect 501126 352294 501182 352350
rect 500754 352170 500810 352226
rect 500878 352170 500934 352226
rect 501002 352170 501058 352226
rect 501126 352170 501182 352226
rect 500754 352046 500810 352102
rect 500878 352046 500934 352102
rect 501002 352046 501058 352102
rect 501126 352046 501182 352102
rect 500754 351922 500810 351978
rect 500878 351922 500934 351978
rect 501002 351922 501058 351978
rect 501126 351922 501182 351978
rect 500754 334294 500810 334350
rect 500878 334294 500934 334350
rect 501002 334294 501058 334350
rect 501126 334294 501182 334350
rect 500754 334170 500810 334226
rect 500878 334170 500934 334226
rect 501002 334170 501058 334226
rect 501126 334170 501182 334226
rect 500754 334046 500810 334102
rect 500878 334046 500934 334102
rect 501002 334046 501058 334102
rect 501126 334046 501182 334102
rect 500754 333922 500810 333978
rect 500878 333922 500934 333978
rect 501002 333922 501058 333978
rect 501126 333922 501182 333978
rect 500754 316294 500810 316350
rect 500878 316294 500934 316350
rect 501002 316294 501058 316350
rect 501126 316294 501182 316350
rect 500754 316170 500810 316226
rect 500878 316170 500934 316226
rect 501002 316170 501058 316226
rect 501126 316170 501182 316226
rect 500754 316046 500810 316102
rect 500878 316046 500934 316102
rect 501002 316046 501058 316102
rect 501126 316046 501182 316102
rect 500754 315922 500810 315978
rect 500878 315922 500934 315978
rect 501002 315922 501058 315978
rect 501126 315922 501182 315978
rect 500754 298294 500810 298350
rect 500878 298294 500934 298350
rect 501002 298294 501058 298350
rect 501126 298294 501182 298350
rect 500754 298170 500810 298226
rect 500878 298170 500934 298226
rect 501002 298170 501058 298226
rect 501126 298170 501182 298226
rect 500754 298046 500810 298102
rect 500878 298046 500934 298102
rect 501002 298046 501058 298102
rect 501126 298046 501182 298102
rect 500754 297922 500810 297978
rect 500878 297922 500934 297978
rect 501002 297922 501058 297978
rect 501126 297922 501182 297978
rect 500754 280294 500810 280350
rect 500878 280294 500934 280350
rect 501002 280294 501058 280350
rect 501126 280294 501182 280350
rect 500754 280170 500810 280226
rect 500878 280170 500934 280226
rect 501002 280170 501058 280226
rect 501126 280170 501182 280226
rect 500754 280046 500810 280102
rect 500878 280046 500934 280102
rect 501002 280046 501058 280102
rect 501126 280046 501182 280102
rect 500754 279922 500810 279978
rect 500878 279922 500934 279978
rect 501002 279922 501058 279978
rect 501126 279922 501182 279978
rect 500754 262294 500810 262350
rect 500878 262294 500934 262350
rect 501002 262294 501058 262350
rect 501126 262294 501182 262350
rect 500754 262170 500810 262226
rect 500878 262170 500934 262226
rect 501002 262170 501058 262226
rect 501126 262170 501182 262226
rect 500754 262046 500810 262102
rect 500878 262046 500934 262102
rect 501002 262046 501058 262102
rect 501126 262046 501182 262102
rect 500754 261922 500810 261978
rect 500878 261922 500934 261978
rect 501002 261922 501058 261978
rect 501126 261922 501182 261978
rect 500754 244294 500810 244350
rect 500878 244294 500934 244350
rect 501002 244294 501058 244350
rect 501126 244294 501182 244350
rect 500754 244170 500810 244226
rect 500878 244170 500934 244226
rect 501002 244170 501058 244226
rect 501126 244170 501182 244226
rect 500754 244046 500810 244102
rect 500878 244046 500934 244102
rect 501002 244046 501058 244102
rect 501126 244046 501182 244102
rect 500754 243922 500810 243978
rect 500878 243922 500934 243978
rect 501002 243922 501058 243978
rect 501126 243922 501182 243978
rect 500754 226294 500810 226350
rect 500878 226294 500934 226350
rect 501002 226294 501058 226350
rect 501126 226294 501182 226350
rect 500754 226170 500810 226226
rect 500878 226170 500934 226226
rect 501002 226170 501058 226226
rect 501126 226170 501182 226226
rect 500754 226046 500810 226102
rect 500878 226046 500934 226102
rect 501002 226046 501058 226102
rect 501126 226046 501182 226102
rect 500754 225922 500810 225978
rect 500878 225922 500934 225978
rect 501002 225922 501058 225978
rect 501126 225922 501182 225978
rect 500754 208294 500810 208350
rect 500878 208294 500934 208350
rect 501002 208294 501058 208350
rect 501126 208294 501182 208350
rect 500754 208170 500810 208226
rect 500878 208170 500934 208226
rect 501002 208170 501058 208226
rect 501126 208170 501182 208226
rect 500754 208046 500810 208102
rect 500878 208046 500934 208102
rect 501002 208046 501058 208102
rect 501126 208046 501182 208102
rect 500754 207922 500810 207978
rect 500878 207922 500934 207978
rect 501002 207922 501058 207978
rect 501126 207922 501182 207978
rect 500754 190294 500810 190350
rect 500878 190294 500934 190350
rect 501002 190294 501058 190350
rect 501126 190294 501182 190350
rect 500754 190170 500810 190226
rect 500878 190170 500934 190226
rect 501002 190170 501058 190226
rect 501126 190170 501182 190226
rect 500754 190046 500810 190102
rect 500878 190046 500934 190102
rect 501002 190046 501058 190102
rect 501126 190046 501182 190102
rect 500754 189922 500810 189978
rect 500878 189922 500934 189978
rect 501002 189922 501058 189978
rect 501126 189922 501182 189978
rect 500754 172294 500810 172350
rect 500878 172294 500934 172350
rect 501002 172294 501058 172350
rect 501126 172294 501182 172350
rect 500754 172170 500810 172226
rect 500878 172170 500934 172226
rect 501002 172170 501058 172226
rect 501126 172170 501182 172226
rect 500754 172046 500810 172102
rect 500878 172046 500934 172102
rect 501002 172046 501058 172102
rect 501126 172046 501182 172102
rect 500754 171922 500810 171978
rect 500878 171922 500934 171978
rect 501002 171922 501058 171978
rect 501126 171922 501182 171978
rect 500754 154294 500810 154350
rect 500878 154294 500934 154350
rect 501002 154294 501058 154350
rect 501126 154294 501182 154350
rect 500754 154170 500810 154226
rect 500878 154170 500934 154226
rect 501002 154170 501058 154226
rect 501126 154170 501182 154226
rect 500754 154046 500810 154102
rect 500878 154046 500934 154102
rect 501002 154046 501058 154102
rect 501126 154046 501182 154102
rect 500754 153922 500810 153978
rect 500878 153922 500934 153978
rect 501002 153922 501058 153978
rect 501126 153922 501182 153978
rect 500754 136294 500810 136350
rect 500878 136294 500934 136350
rect 501002 136294 501058 136350
rect 501126 136294 501182 136350
rect 500754 136170 500810 136226
rect 500878 136170 500934 136226
rect 501002 136170 501058 136226
rect 501126 136170 501182 136226
rect 500754 136046 500810 136102
rect 500878 136046 500934 136102
rect 501002 136046 501058 136102
rect 501126 136046 501182 136102
rect 500754 135922 500810 135978
rect 500878 135922 500934 135978
rect 501002 135922 501058 135978
rect 501126 135922 501182 135978
rect 500754 118294 500810 118350
rect 500878 118294 500934 118350
rect 501002 118294 501058 118350
rect 501126 118294 501182 118350
rect 500754 118170 500810 118226
rect 500878 118170 500934 118226
rect 501002 118170 501058 118226
rect 501126 118170 501182 118226
rect 500754 118046 500810 118102
rect 500878 118046 500934 118102
rect 501002 118046 501058 118102
rect 501126 118046 501182 118102
rect 500754 117922 500810 117978
rect 500878 117922 500934 117978
rect 501002 117922 501058 117978
rect 501126 117922 501182 117978
rect 500754 100294 500810 100350
rect 500878 100294 500934 100350
rect 501002 100294 501058 100350
rect 501126 100294 501182 100350
rect 500754 100170 500810 100226
rect 500878 100170 500934 100226
rect 501002 100170 501058 100226
rect 501126 100170 501182 100226
rect 500754 100046 500810 100102
rect 500878 100046 500934 100102
rect 501002 100046 501058 100102
rect 501126 100046 501182 100102
rect 500754 99922 500810 99978
rect 500878 99922 500934 99978
rect 501002 99922 501058 99978
rect 501126 99922 501182 99978
rect 500754 82294 500810 82350
rect 500878 82294 500934 82350
rect 501002 82294 501058 82350
rect 501126 82294 501182 82350
rect 500754 82170 500810 82226
rect 500878 82170 500934 82226
rect 501002 82170 501058 82226
rect 501126 82170 501182 82226
rect 500754 82046 500810 82102
rect 500878 82046 500934 82102
rect 501002 82046 501058 82102
rect 501126 82046 501182 82102
rect 500754 81922 500810 81978
rect 500878 81922 500934 81978
rect 501002 81922 501058 81978
rect 501126 81922 501182 81978
rect 527754 382294 527810 382350
rect 527878 382294 527934 382350
rect 528002 382294 528058 382350
rect 528126 382294 528182 382350
rect 527754 382170 527810 382226
rect 527878 382170 527934 382226
rect 528002 382170 528058 382226
rect 528126 382170 528182 382226
rect 527754 382046 527810 382102
rect 527878 382046 527934 382102
rect 528002 382046 528058 382102
rect 528126 382046 528182 382102
rect 527754 381922 527810 381978
rect 527878 381922 527934 381978
rect 528002 381922 528058 381978
rect 528126 381922 528182 381978
rect 527754 364294 527810 364350
rect 527878 364294 527934 364350
rect 528002 364294 528058 364350
rect 528126 364294 528182 364350
rect 527754 364170 527810 364226
rect 527878 364170 527934 364226
rect 528002 364170 528058 364226
rect 528126 364170 528182 364226
rect 527754 364046 527810 364102
rect 527878 364046 527934 364102
rect 528002 364046 528058 364102
rect 528126 364046 528182 364102
rect 527754 363922 527810 363978
rect 527878 363922 527934 363978
rect 528002 363922 528058 363978
rect 528126 363922 528182 363978
rect 527754 346294 527810 346350
rect 527878 346294 527934 346350
rect 528002 346294 528058 346350
rect 528126 346294 528182 346350
rect 527754 346170 527810 346226
rect 527878 346170 527934 346226
rect 528002 346170 528058 346226
rect 528126 346170 528182 346226
rect 527754 346046 527810 346102
rect 527878 346046 527934 346102
rect 528002 346046 528058 346102
rect 528126 346046 528182 346102
rect 527754 345922 527810 345978
rect 527878 345922 527934 345978
rect 528002 345922 528058 345978
rect 528126 345922 528182 345978
rect 527754 328294 527810 328350
rect 527878 328294 527934 328350
rect 528002 328294 528058 328350
rect 528126 328294 528182 328350
rect 527754 328170 527810 328226
rect 527878 328170 527934 328226
rect 528002 328170 528058 328226
rect 528126 328170 528182 328226
rect 527754 328046 527810 328102
rect 527878 328046 527934 328102
rect 528002 328046 528058 328102
rect 528126 328046 528182 328102
rect 527754 327922 527810 327978
rect 527878 327922 527934 327978
rect 528002 327922 528058 327978
rect 528126 327922 528182 327978
rect 527754 310294 527810 310350
rect 527878 310294 527934 310350
rect 528002 310294 528058 310350
rect 528126 310294 528182 310350
rect 527754 310170 527810 310226
rect 527878 310170 527934 310226
rect 528002 310170 528058 310226
rect 528126 310170 528182 310226
rect 527754 310046 527810 310102
rect 527878 310046 527934 310102
rect 528002 310046 528058 310102
rect 528126 310046 528182 310102
rect 527754 309922 527810 309978
rect 527878 309922 527934 309978
rect 528002 309922 528058 309978
rect 528126 309922 528182 309978
rect 527754 292294 527810 292350
rect 527878 292294 527934 292350
rect 528002 292294 528058 292350
rect 528126 292294 528182 292350
rect 527754 292170 527810 292226
rect 527878 292170 527934 292226
rect 528002 292170 528058 292226
rect 528126 292170 528182 292226
rect 527754 292046 527810 292102
rect 527878 292046 527934 292102
rect 528002 292046 528058 292102
rect 528126 292046 528182 292102
rect 527754 291922 527810 291978
rect 527878 291922 527934 291978
rect 528002 291922 528058 291978
rect 528126 291922 528182 291978
rect 531474 598116 531530 598172
rect 531598 598116 531654 598172
rect 531722 598116 531778 598172
rect 531846 598116 531902 598172
rect 531474 597992 531530 598048
rect 531598 597992 531654 598048
rect 531722 597992 531778 598048
rect 531846 597992 531902 598048
rect 531474 597868 531530 597924
rect 531598 597868 531654 597924
rect 531722 597868 531778 597924
rect 531846 597868 531902 597924
rect 531474 597744 531530 597800
rect 531598 597744 531654 597800
rect 531722 597744 531778 597800
rect 531846 597744 531902 597800
rect 531474 586294 531530 586350
rect 531598 586294 531654 586350
rect 531722 586294 531778 586350
rect 531846 586294 531902 586350
rect 531474 586170 531530 586226
rect 531598 586170 531654 586226
rect 531722 586170 531778 586226
rect 531846 586170 531902 586226
rect 531474 586046 531530 586102
rect 531598 586046 531654 586102
rect 531722 586046 531778 586102
rect 531846 586046 531902 586102
rect 531474 585922 531530 585978
rect 531598 585922 531654 585978
rect 531722 585922 531778 585978
rect 531846 585922 531902 585978
rect 531474 568294 531530 568350
rect 531598 568294 531654 568350
rect 531722 568294 531778 568350
rect 531846 568294 531902 568350
rect 531474 568170 531530 568226
rect 531598 568170 531654 568226
rect 531722 568170 531778 568226
rect 531846 568170 531902 568226
rect 531474 568046 531530 568102
rect 531598 568046 531654 568102
rect 531722 568046 531778 568102
rect 531846 568046 531902 568102
rect 531474 567922 531530 567978
rect 531598 567922 531654 567978
rect 531722 567922 531778 567978
rect 531846 567922 531902 567978
rect 531474 550294 531530 550350
rect 531598 550294 531654 550350
rect 531722 550294 531778 550350
rect 531846 550294 531902 550350
rect 531474 550170 531530 550226
rect 531598 550170 531654 550226
rect 531722 550170 531778 550226
rect 531846 550170 531902 550226
rect 531474 550046 531530 550102
rect 531598 550046 531654 550102
rect 531722 550046 531778 550102
rect 531846 550046 531902 550102
rect 531474 549922 531530 549978
rect 531598 549922 531654 549978
rect 531722 549922 531778 549978
rect 531846 549922 531902 549978
rect 531474 532294 531530 532350
rect 531598 532294 531654 532350
rect 531722 532294 531778 532350
rect 531846 532294 531902 532350
rect 531474 532170 531530 532226
rect 531598 532170 531654 532226
rect 531722 532170 531778 532226
rect 531846 532170 531902 532226
rect 531474 532046 531530 532102
rect 531598 532046 531654 532102
rect 531722 532046 531778 532102
rect 531846 532046 531902 532102
rect 531474 531922 531530 531978
rect 531598 531922 531654 531978
rect 531722 531922 531778 531978
rect 531846 531922 531902 531978
rect 531474 514294 531530 514350
rect 531598 514294 531654 514350
rect 531722 514294 531778 514350
rect 531846 514294 531902 514350
rect 531474 514170 531530 514226
rect 531598 514170 531654 514226
rect 531722 514170 531778 514226
rect 531846 514170 531902 514226
rect 531474 514046 531530 514102
rect 531598 514046 531654 514102
rect 531722 514046 531778 514102
rect 531846 514046 531902 514102
rect 531474 513922 531530 513978
rect 531598 513922 531654 513978
rect 531722 513922 531778 513978
rect 531846 513922 531902 513978
rect 531474 496294 531530 496350
rect 531598 496294 531654 496350
rect 531722 496294 531778 496350
rect 531846 496294 531902 496350
rect 531474 496170 531530 496226
rect 531598 496170 531654 496226
rect 531722 496170 531778 496226
rect 531846 496170 531902 496226
rect 531474 496046 531530 496102
rect 531598 496046 531654 496102
rect 531722 496046 531778 496102
rect 531846 496046 531902 496102
rect 531474 495922 531530 495978
rect 531598 495922 531654 495978
rect 531722 495922 531778 495978
rect 531846 495922 531902 495978
rect 531474 478294 531530 478350
rect 531598 478294 531654 478350
rect 531722 478294 531778 478350
rect 531846 478294 531902 478350
rect 531474 478170 531530 478226
rect 531598 478170 531654 478226
rect 531722 478170 531778 478226
rect 531846 478170 531902 478226
rect 531474 478046 531530 478102
rect 531598 478046 531654 478102
rect 531722 478046 531778 478102
rect 531846 478046 531902 478102
rect 531474 477922 531530 477978
rect 531598 477922 531654 477978
rect 531722 477922 531778 477978
rect 531846 477922 531902 477978
rect 531474 460294 531530 460350
rect 531598 460294 531654 460350
rect 531722 460294 531778 460350
rect 531846 460294 531902 460350
rect 531474 460170 531530 460226
rect 531598 460170 531654 460226
rect 531722 460170 531778 460226
rect 531846 460170 531902 460226
rect 531474 460046 531530 460102
rect 531598 460046 531654 460102
rect 531722 460046 531778 460102
rect 531846 460046 531902 460102
rect 531474 459922 531530 459978
rect 531598 459922 531654 459978
rect 531722 459922 531778 459978
rect 531846 459922 531902 459978
rect 531474 442294 531530 442350
rect 531598 442294 531654 442350
rect 531722 442294 531778 442350
rect 531846 442294 531902 442350
rect 531474 442170 531530 442226
rect 531598 442170 531654 442226
rect 531722 442170 531778 442226
rect 531846 442170 531902 442226
rect 531474 442046 531530 442102
rect 531598 442046 531654 442102
rect 531722 442046 531778 442102
rect 531846 442046 531902 442102
rect 531474 441922 531530 441978
rect 531598 441922 531654 441978
rect 531722 441922 531778 441978
rect 531846 441922 531902 441978
rect 531474 424294 531530 424350
rect 531598 424294 531654 424350
rect 531722 424294 531778 424350
rect 531846 424294 531902 424350
rect 531474 424170 531530 424226
rect 531598 424170 531654 424226
rect 531722 424170 531778 424226
rect 531846 424170 531902 424226
rect 531474 424046 531530 424102
rect 531598 424046 531654 424102
rect 531722 424046 531778 424102
rect 531846 424046 531902 424102
rect 531474 423922 531530 423978
rect 531598 423922 531654 423978
rect 531722 423922 531778 423978
rect 531846 423922 531902 423978
rect 531474 406294 531530 406350
rect 531598 406294 531654 406350
rect 531722 406294 531778 406350
rect 531846 406294 531902 406350
rect 531474 406170 531530 406226
rect 531598 406170 531654 406226
rect 531722 406170 531778 406226
rect 531846 406170 531902 406226
rect 531474 406046 531530 406102
rect 531598 406046 531654 406102
rect 531722 406046 531778 406102
rect 531846 406046 531902 406102
rect 531474 405922 531530 405978
rect 531598 405922 531654 405978
rect 531722 405922 531778 405978
rect 531846 405922 531902 405978
rect 531474 388294 531530 388350
rect 531598 388294 531654 388350
rect 531722 388294 531778 388350
rect 531846 388294 531902 388350
rect 531474 388170 531530 388226
rect 531598 388170 531654 388226
rect 531722 388170 531778 388226
rect 531846 388170 531902 388226
rect 531474 388046 531530 388102
rect 531598 388046 531654 388102
rect 531722 388046 531778 388102
rect 531846 388046 531902 388102
rect 531474 387922 531530 387978
rect 531598 387922 531654 387978
rect 531722 387922 531778 387978
rect 531846 387922 531902 387978
rect 531474 370294 531530 370350
rect 531598 370294 531654 370350
rect 531722 370294 531778 370350
rect 531846 370294 531902 370350
rect 531474 370170 531530 370226
rect 531598 370170 531654 370226
rect 531722 370170 531778 370226
rect 531846 370170 531902 370226
rect 531474 370046 531530 370102
rect 531598 370046 531654 370102
rect 531722 370046 531778 370102
rect 531846 370046 531902 370102
rect 531474 369922 531530 369978
rect 531598 369922 531654 369978
rect 531722 369922 531778 369978
rect 531846 369922 531902 369978
rect 531474 352294 531530 352350
rect 531598 352294 531654 352350
rect 531722 352294 531778 352350
rect 531846 352294 531902 352350
rect 531474 352170 531530 352226
rect 531598 352170 531654 352226
rect 531722 352170 531778 352226
rect 531846 352170 531902 352226
rect 531474 352046 531530 352102
rect 531598 352046 531654 352102
rect 531722 352046 531778 352102
rect 531846 352046 531902 352102
rect 531474 351922 531530 351978
rect 531598 351922 531654 351978
rect 531722 351922 531778 351978
rect 531846 351922 531902 351978
rect 531474 334294 531530 334350
rect 531598 334294 531654 334350
rect 531722 334294 531778 334350
rect 531846 334294 531902 334350
rect 531474 334170 531530 334226
rect 531598 334170 531654 334226
rect 531722 334170 531778 334226
rect 531846 334170 531902 334226
rect 531474 334046 531530 334102
rect 531598 334046 531654 334102
rect 531722 334046 531778 334102
rect 531846 334046 531902 334102
rect 531474 333922 531530 333978
rect 531598 333922 531654 333978
rect 531722 333922 531778 333978
rect 531846 333922 531902 333978
rect 531474 316294 531530 316350
rect 531598 316294 531654 316350
rect 531722 316294 531778 316350
rect 531846 316294 531902 316350
rect 531474 316170 531530 316226
rect 531598 316170 531654 316226
rect 531722 316170 531778 316226
rect 531846 316170 531902 316226
rect 531474 316046 531530 316102
rect 531598 316046 531654 316102
rect 531722 316046 531778 316102
rect 531846 316046 531902 316102
rect 531474 315922 531530 315978
rect 531598 315922 531654 315978
rect 531722 315922 531778 315978
rect 531846 315922 531902 315978
rect 558474 597156 558530 597212
rect 558598 597156 558654 597212
rect 558722 597156 558778 597212
rect 558846 597156 558902 597212
rect 558474 597032 558530 597088
rect 558598 597032 558654 597088
rect 558722 597032 558778 597088
rect 558846 597032 558902 597088
rect 558474 596908 558530 596964
rect 558598 596908 558654 596964
rect 558722 596908 558778 596964
rect 558846 596908 558902 596964
rect 558474 596784 558530 596840
rect 558598 596784 558654 596840
rect 558722 596784 558778 596840
rect 558846 596784 558902 596840
rect 558474 580294 558530 580350
rect 558598 580294 558654 580350
rect 558722 580294 558778 580350
rect 558846 580294 558902 580350
rect 558474 580170 558530 580226
rect 558598 580170 558654 580226
rect 558722 580170 558778 580226
rect 558846 580170 558902 580226
rect 558474 580046 558530 580102
rect 558598 580046 558654 580102
rect 558722 580046 558778 580102
rect 558846 580046 558902 580102
rect 558474 579922 558530 579978
rect 558598 579922 558654 579978
rect 558722 579922 558778 579978
rect 558846 579922 558902 579978
rect 558474 562294 558530 562350
rect 558598 562294 558654 562350
rect 558722 562294 558778 562350
rect 558846 562294 558902 562350
rect 558474 562170 558530 562226
rect 558598 562170 558654 562226
rect 558722 562170 558778 562226
rect 558846 562170 558902 562226
rect 558474 562046 558530 562102
rect 558598 562046 558654 562102
rect 558722 562046 558778 562102
rect 558846 562046 558902 562102
rect 558474 561922 558530 561978
rect 558598 561922 558654 561978
rect 558722 561922 558778 561978
rect 558846 561922 558902 561978
rect 558474 544294 558530 544350
rect 558598 544294 558654 544350
rect 558722 544294 558778 544350
rect 558846 544294 558902 544350
rect 558474 544170 558530 544226
rect 558598 544170 558654 544226
rect 558722 544170 558778 544226
rect 558846 544170 558902 544226
rect 558474 544046 558530 544102
rect 558598 544046 558654 544102
rect 558722 544046 558778 544102
rect 558846 544046 558902 544102
rect 558474 543922 558530 543978
rect 558598 543922 558654 543978
rect 558722 543922 558778 543978
rect 558846 543922 558902 543978
rect 558474 526294 558530 526350
rect 558598 526294 558654 526350
rect 558722 526294 558778 526350
rect 558846 526294 558902 526350
rect 558474 526170 558530 526226
rect 558598 526170 558654 526226
rect 558722 526170 558778 526226
rect 558846 526170 558902 526226
rect 558474 526046 558530 526102
rect 558598 526046 558654 526102
rect 558722 526046 558778 526102
rect 558846 526046 558902 526102
rect 558474 525922 558530 525978
rect 558598 525922 558654 525978
rect 558722 525922 558778 525978
rect 558846 525922 558902 525978
rect 558474 508294 558530 508350
rect 558598 508294 558654 508350
rect 558722 508294 558778 508350
rect 558846 508294 558902 508350
rect 558474 508170 558530 508226
rect 558598 508170 558654 508226
rect 558722 508170 558778 508226
rect 558846 508170 558902 508226
rect 558474 508046 558530 508102
rect 558598 508046 558654 508102
rect 558722 508046 558778 508102
rect 558846 508046 558902 508102
rect 558474 507922 558530 507978
rect 558598 507922 558654 507978
rect 558722 507922 558778 507978
rect 558846 507922 558902 507978
rect 558474 490294 558530 490350
rect 558598 490294 558654 490350
rect 558722 490294 558778 490350
rect 558846 490294 558902 490350
rect 558474 490170 558530 490226
rect 558598 490170 558654 490226
rect 558722 490170 558778 490226
rect 558846 490170 558902 490226
rect 558474 490046 558530 490102
rect 558598 490046 558654 490102
rect 558722 490046 558778 490102
rect 558846 490046 558902 490102
rect 558474 489922 558530 489978
rect 558598 489922 558654 489978
rect 558722 489922 558778 489978
rect 558846 489922 558902 489978
rect 558474 472294 558530 472350
rect 558598 472294 558654 472350
rect 558722 472294 558778 472350
rect 558846 472294 558902 472350
rect 558474 472170 558530 472226
rect 558598 472170 558654 472226
rect 558722 472170 558778 472226
rect 558846 472170 558902 472226
rect 558474 472046 558530 472102
rect 558598 472046 558654 472102
rect 558722 472046 558778 472102
rect 558846 472046 558902 472102
rect 558474 471922 558530 471978
rect 558598 471922 558654 471978
rect 558722 471922 558778 471978
rect 558846 471922 558902 471978
rect 558474 454294 558530 454350
rect 558598 454294 558654 454350
rect 558722 454294 558778 454350
rect 558846 454294 558902 454350
rect 558474 454170 558530 454226
rect 558598 454170 558654 454226
rect 558722 454170 558778 454226
rect 558846 454170 558902 454226
rect 558474 454046 558530 454102
rect 558598 454046 558654 454102
rect 558722 454046 558778 454102
rect 558846 454046 558902 454102
rect 558474 453922 558530 453978
rect 558598 453922 558654 453978
rect 558722 453922 558778 453978
rect 558846 453922 558902 453978
rect 558474 436294 558530 436350
rect 558598 436294 558654 436350
rect 558722 436294 558778 436350
rect 558846 436294 558902 436350
rect 558474 436170 558530 436226
rect 558598 436170 558654 436226
rect 558722 436170 558778 436226
rect 558846 436170 558902 436226
rect 558474 436046 558530 436102
rect 558598 436046 558654 436102
rect 558722 436046 558778 436102
rect 558846 436046 558902 436102
rect 558474 435922 558530 435978
rect 558598 435922 558654 435978
rect 558722 435922 558778 435978
rect 558846 435922 558902 435978
rect 558474 418294 558530 418350
rect 558598 418294 558654 418350
rect 558722 418294 558778 418350
rect 558846 418294 558902 418350
rect 558474 418170 558530 418226
rect 558598 418170 558654 418226
rect 558722 418170 558778 418226
rect 558846 418170 558902 418226
rect 558474 418046 558530 418102
rect 558598 418046 558654 418102
rect 558722 418046 558778 418102
rect 558846 418046 558902 418102
rect 558474 417922 558530 417978
rect 558598 417922 558654 417978
rect 558722 417922 558778 417978
rect 558846 417922 558902 417978
rect 558474 400294 558530 400350
rect 558598 400294 558654 400350
rect 558722 400294 558778 400350
rect 558846 400294 558902 400350
rect 558474 400170 558530 400226
rect 558598 400170 558654 400226
rect 558722 400170 558778 400226
rect 558846 400170 558902 400226
rect 558474 400046 558530 400102
rect 558598 400046 558654 400102
rect 558722 400046 558778 400102
rect 558846 400046 558902 400102
rect 558474 399922 558530 399978
rect 558598 399922 558654 399978
rect 558722 399922 558778 399978
rect 558846 399922 558902 399978
rect 558474 382294 558530 382350
rect 558598 382294 558654 382350
rect 558722 382294 558778 382350
rect 558846 382294 558902 382350
rect 558474 382170 558530 382226
rect 558598 382170 558654 382226
rect 558722 382170 558778 382226
rect 558846 382170 558902 382226
rect 558474 382046 558530 382102
rect 558598 382046 558654 382102
rect 558722 382046 558778 382102
rect 558846 382046 558902 382102
rect 558474 381922 558530 381978
rect 558598 381922 558654 381978
rect 558722 381922 558778 381978
rect 558846 381922 558902 381978
rect 558474 364294 558530 364350
rect 558598 364294 558654 364350
rect 558722 364294 558778 364350
rect 558846 364294 558902 364350
rect 558474 364170 558530 364226
rect 558598 364170 558654 364226
rect 558722 364170 558778 364226
rect 558846 364170 558902 364226
rect 558474 364046 558530 364102
rect 558598 364046 558654 364102
rect 558722 364046 558778 364102
rect 558846 364046 558902 364102
rect 558474 363922 558530 363978
rect 558598 363922 558654 363978
rect 558722 363922 558778 363978
rect 558846 363922 558902 363978
rect 558474 346294 558530 346350
rect 558598 346294 558654 346350
rect 558722 346294 558778 346350
rect 558846 346294 558902 346350
rect 558474 346170 558530 346226
rect 558598 346170 558654 346226
rect 558722 346170 558778 346226
rect 558846 346170 558902 346226
rect 558474 346046 558530 346102
rect 558598 346046 558654 346102
rect 558722 346046 558778 346102
rect 558846 346046 558902 346102
rect 558474 345922 558530 345978
rect 558598 345922 558654 345978
rect 558722 345922 558778 345978
rect 558846 345922 558902 345978
rect 558474 328294 558530 328350
rect 558598 328294 558654 328350
rect 558722 328294 558778 328350
rect 558846 328294 558902 328350
rect 558474 328170 558530 328226
rect 558598 328170 558654 328226
rect 558722 328170 558778 328226
rect 558846 328170 558902 328226
rect 558474 328046 558530 328102
rect 558598 328046 558654 328102
rect 558722 328046 558778 328102
rect 558846 328046 558902 328102
rect 558474 327922 558530 327978
rect 558598 327922 558654 327978
rect 558722 327922 558778 327978
rect 558846 327922 558902 327978
rect 531474 298294 531530 298350
rect 531598 298294 531654 298350
rect 531722 298294 531778 298350
rect 531846 298294 531902 298350
rect 531474 298170 531530 298226
rect 531598 298170 531654 298226
rect 531722 298170 531778 298226
rect 531846 298170 531902 298226
rect 531474 298046 531530 298102
rect 531598 298046 531654 298102
rect 531722 298046 531778 298102
rect 531846 298046 531902 298102
rect 531474 297922 531530 297978
rect 531598 297922 531654 297978
rect 531722 297922 531778 297978
rect 531846 297922 531902 297978
rect 531474 280294 531530 280350
rect 531598 280294 531654 280350
rect 531722 280294 531778 280350
rect 531846 280294 531902 280350
rect 531474 280170 531530 280226
rect 531598 280170 531654 280226
rect 531722 280170 531778 280226
rect 531846 280170 531902 280226
rect 531474 280046 531530 280102
rect 531598 280046 531654 280102
rect 531722 280046 531778 280102
rect 531846 280046 531902 280102
rect 531474 279922 531530 279978
rect 531598 279922 531654 279978
rect 531722 279922 531778 279978
rect 531846 279922 531902 279978
rect 527754 274294 527810 274350
rect 527878 274294 527934 274350
rect 528002 274294 528058 274350
rect 528126 274294 528182 274350
rect 527754 274170 527810 274226
rect 527878 274170 527934 274226
rect 528002 274170 528058 274226
rect 528126 274170 528182 274226
rect 527754 274046 527810 274102
rect 527878 274046 527934 274102
rect 528002 274046 528058 274102
rect 528126 274046 528182 274102
rect 527754 273922 527810 273978
rect 527878 273922 527934 273978
rect 528002 273922 528058 273978
rect 528126 273922 528182 273978
rect 527754 256294 527810 256350
rect 527878 256294 527934 256350
rect 528002 256294 528058 256350
rect 528126 256294 528182 256350
rect 527754 256170 527810 256226
rect 527878 256170 527934 256226
rect 528002 256170 528058 256226
rect 528126 256170 528182 256226
rect 527754 256046 527810 256102
rect 527878 256046 527934 256102
rect 528002 256046 528058 256102
rect 528126 256046 528182 256102
rect 527754 255922 527810 255978
rect 527878 255922 527934 255978
rect 528002 255922 528058 255978
rect 528126 255922 528182 255978
rect 527754 238294 527810 238350
rect 527878 238294 527934 238350
rect 528002 238294 528058 238350
rect 528126 238294 528182 238350
rect 527754 238170 527810 238226
rect 527878 238170 527934 238226
rect 528002 238170 528058 238226
rect 528126 238170 528182 238226
rect 527754 238046 527810 238102
rect 527878 238046 527934 238102
rect 528002 238046 528058 238102
rect 528126 238046 528182 238102
rect 527754 237922 527810 237978
rect 527878 237922 527934 237978
rect 528002 237922 528058 237978
rect 528126 237922 528182 237978
rect 527754 220294 527810 220350
rect 527878 220294 527934 220350
rect 528002 220294 528058 220350
rect 528126 220294 528182 220350
rect 527754 220170 527810 220226
rect 527878 220170 527934 220226
rect 528002 220170 528058 220226
rect 528126 220170 528182 220226
rect 527754 220046 527810 220102
rect 527878 220046 527934 220102
rect 528002 220046 528058 220102
rect 528126 220046 528182 220102
rect 527754 219922 527810 219978
rect 527878 219922 527934 219978
rect 528002 219922 528058 219978
rect 528126 219922 528182 219978
rect 527754 202294 527810 202350
rect 527878 202294 527934 202350
rect 528002 202294 528058 202350
rect 528126 202294 528182 202350
rect 527754 202170 527810 202226
rect 527878 202170 527934 202226
rect 528002 202170 528058 202226
rect 528126 202170 528182 202226
rect 527754 202046 527810 202102
rect 527878 202046 527934 202102
rect 528002 202046 528058 202102
rect 528126 202046 528182 202102
rect 527754 201922 527810 201978
rect 527878 201922 527934 201978
rect 528002 201922 528058 201978
rect 528126 201922 528182 201978
rect 527754 184294 527810 184350
rect 527878 184294 527934 184350
rect 528002 184294 528058 184350
rect 528126 184294 528182 184350
rect 527754 184170 527810 184226
rect 527878 184170 527934 184226
rect 528002 184170 528058 184226
rect 528126 184170 528182 184226
rect 527754 184046 527810 184102
rect 527878 184046 527934 184102
rect 528002 184046 528058 184102
rect 528126 184046 528182 184102
rect 527754 183922 527810 183978
rect 527878 183922 527934 183978
rect 528002 183922 528058 183978
rect 528126 183922 528182 183978
rect 527754 166294 527810 166350
rect 527878 166294 527934 166350
rect 528002 166294 528058 166350
rect 528126 166294 528182 166350
rect 527754 166170 527810 166226
rect 527878 166170 527934 166226
rect 528002 166170 528058 166226
rect 528126 166170 528182 166226
rect 527754 166046 527810 166102
rect 527878 166046 527934 166102
rect 528002 166046 528058 166102
rect 528126 166046 528182 166102
rect 527754 165922 527810 165978
rect 527878 165922 527934 165978
rect 528002 165922 528058 165978
rect 528126 165922 528182 165978
rect 527754 148294 527810 148350
rect 527878 148294 527934 148350
rect 528002 148294 528058 148350
rect 528126 148294 528182 148350
rect 527754 148170 527810 148226
rect 527878 148170 527934 148226
rect 528002 148170 528058 148226
rect 528126 148170 528182 148226
rect 527754 148046 527810 148102
rect 527878 148046 527934 148102
rect 528002 148046 528058 148102
rect 528126 148046 528182 148102
rect 527754 147922 527810 147978
rect 527878 147922 527934 147978
rect 528002 147922 528058 147978
rect 528126 147922 528182 147978
rect 527754 130294 527810 130350
rect 527878 130294 527934 130350
rect 528002 130294 528058 130350
rect 528126 130294 528182 130350
rect 527754 130170 527810 130226
rect 527878 130170 527934 130226
rect 528002 130170 528058 130226
rect 528126 130170 528182 130226
rect 527754 130046 527810 130102
rect 527878 130046 527934 130102
rect 528002 130046 528058 130102
rect 528126 130046 528182 130102
rect 527754 129922 527810 129978
rect 527878 129922 527934 129978
rect 528002 129922 528058 129978
rect 528126 129922 528182 129978
rect 527754 112294 527810 112350
rect 527878 112294 527934 112350
rect 528002 112294 528058 112350
rect 528126 112294 528182 112350
rect 527754 112170 527810 112226
rect 527878 112170 527934 112226
rect 528002 112170 528058 112226
rect 528126 112170 528182 112226
rect 527754 112046 527810 112102
rect 527878 112046 527934 112102
rect 528002 112046 528058 112102
rect 528126 112046 528182 112102
rect 527754 111922 527810 111978
rect 527878 111922 527934 111978
rect 528002 111922 528058 111978
rect 528126 111922 528182 111978
rect 527754 94294 527810 94350
rect 527878 94294 527934 94350
rect 528002 94294 528058 94350
rect 528126 94294 528182 94350
rect 527754 94170 527810 94226
rect 527878 94170 527934 94226
rect 528002 94170 528058 94226
rect 528126 94170 528182 94226
rect 527754 94046 527810 94102
rect 527878 94046 527934 94102
rect 528002 94046 528058 94102
rect 528126 94046 528182 94102
rect 527754 93922 527810 93978
rect 527878 93922 527934 93978
rect 528002 93922 528058 93978
rect 528126 93922 528182 93978
rect 527754 76294 527810 76350
rect 527878 76294 527934 76350
rect 528002 76294 528058 76350
rect 528126 76294 528182 76350
rect 527754 76170 527810 76226
rect 527878 76170 527934 76226
rect 528002 76170 528058 76226
rect 528126 76170 528182 76226
rect 527754 76046 527810 76102
rect 527878 76046 527934 76102
rect 528002 76046 528058 76102
rect 528126 76046 528182 76102
rect 527754 75922 527810 75978
rect 527878 75922 527934 75978
rect 528002 75922 528058 75978
rect 528126 75922 528182 75978
rect 500754 64294 500810 64350
rect 500878 64294 500934 64350
rect 501002 64294 501058 64350
rect 501126 64294 501182 64350
rect 500754 64170 500810 64226
rect 500878 64170 500934 64226
rect 501002 64170 501058 64226
rect 501126 64170 501182 64226
rect 500754 64046 500810 64102
rect 500878 64046 500934 64102
rect 501002 64046 501058 64102
rect 501126 64046 501182 64102
rect 500754 63922 500810 63978
rect 500878 63922 500934 63978
rect 501002 63922 501058 63978
rect 501126 63922 501182 63978
rect 500754 46294 500810 46350
rect 500878 46294 500934 46350
rect 501002 46294 501058 46350
rect 501126 46294 501182 46350
rect 500754 46170 500810 46226
rect 500878 46170 500934 46226
rect 501002 46170 501058 46226
rect 501126 46170 501182 46226
rect 500754 46046 500810 46102
rect 500878 46046 500934 46102
rect 501002 46046 501058 46102
rect 501126 46046 501182 46102
rect 500754 45922 500810 45978
rect 500878 45922 500934 45978
rect 501002 45922 501058 45978
rect 501126 45922 501182 45978
rect 500754 28294 500810 28350
rect 500878 28294 500934 28350
rect 501002 28294 501058 28350
rect 501126 28294 501182 28350
rect 500754 28170 500810 28226
rect 500878 28170 500934 28226
rect 501002 28170 501058 28226
rect 501126 28170 501182 28226
rect 500754 28046 500810 28102
rect 500878 28046 500934 28102
rect 501002 28046 501058 28102
rect 501126 28046 501182 28102
rect 500754 27922 500810 27978
rect 500878 27922 500934 27978
rect 501002 27922 501058 27978
rect 501126 27922 501182 27978
rect 500754 10294 500810 10350
rect 500878 10294 500934 10350
rect 501002 10294 501058 10350
rect 501126 10294 501182 10350
rect 500754 10170 500810 10226
rect 500878 10170 500934 10226
rect 501002 10170 501058 10226
rect 501126 10170 501182 10226
rect 500754 10046 500810 10102
rect 500878 10046 500934 10102
rect 501002 10046 501058 10102
rect 501126 10046 501182 10102
rect 500754 9922 500810 9978
rect 500878 9922 500934 9978
rect 501002 9922 501058 9978
rect 501126 9922 501182 9978
rect 498988 5124 499044 5158
rect 498988 5102 499044 5124
rect 497034 4294 497090 4350
rect 497158 4294 497214 4350
rect 497282 4294 497338 4350
rect 497406 4294 497462 4350
rect 497034 4170 497090 4226
rect 497158 4170 497214 4226
rect 497282 4170 497338 4226
rect 497406 4170 497462 4226
rect 497034 4046 497090 4102
rect 497158 4046 497214 4102
rect 497282 4046 497338 4102
rect 497406 4046 497462 4102
rect 497034 3922 497090 3978
rect 497158 3922 497214 3978
rect 497282 3922 497338 3978
rect 497406 3922 497462 3978
rect 470034 -1176 470090 -1120
rect 470158 -1176 470214 -1120
rect 470282 -1176 470338 -1120
rect 470406 -1176 470462 -1120
rect 470034 -1300 470090 -1244
rect 470158 -1300 470214 -1244
rect 470282 -1300 470338 -1244
rect 470406 -1300 470462 -1244
rect 470034 -1424 470090 -1368
rect 470158 -1424 470214 -1368
rect 470282 -1424 470338 -1368
rect 470406 -1424 470462 -1368
rect 470034 -1548 470090 -1492
rect 470158 -1548 470214 -1492
rect 470282 -1548 470338 -1492
rect 470406 -1548 470462 -1492
rect 498988 3302 499044 3358
rect 499436 3122 499492 3178
rect 497034 -216 497090 -160
rect 497158 -216 497214 -160
rect 497282 -216 497338 -160
rect 497406 -216 497462 -160
rect 497034 -340 497090 -284
rect 497158 -340 497214 -284
rect 497282 -340 497338 -284
rect 497406 -340 497462 -284
rect 497034 -464 497090 -408
rect 497158 -464 497214 -408
rect 497282 -464 497338 -408
rect 497406 -464 497462 -408
rect 497034 -588 497090 -532
rect 497158 -588 497214 -532
rect 497282 -588 497338 -532
rect 497406 -588 497462 -532
rect 531474 262294 531530 262350
rect 531598 262294 531654 262350
rect 531722 262294 531778 262350
rect 531846 262294 531902 262350
rect 531474 262170 531530 262226
rect 531598 262170 531654 262226
rect 531722 262170 531778 262226
rect 531846 262170 531902 262226
rect 531474 262046 531530 262102
rect 531598 262046 531654 262102
rect 531722 262046 531778 262102
rect 531846 262046 531902 262102
rect 531474 261922 531530 261978
rect 531598 261922 531654 261978
rect 531722 261922 531778 261978
rect 531846 261922 531902 261978
rect 531474 244294 531530 244350
rect 531598 244294 531654 244350
rect 531722 244294 531778 244350
rect 531846 244294 531902 244350
rect 531474 244170 531530 244226
rect 531598 244170 531654 244226
rect 531722 244170 531778 244226
rect 531846 244170 531902 244226
rect 531474 244046 531530 244102
rect 531598 244046 531654 244102
rect 531722 244046 531778 244102
rect 531846 244046 531902 244102
rect 531474 243922 531530 243978
rect 531598 243922 531654 243978
rect 531722 243922 531778 243978
rect 531846 243922 531902 243978
rect 531474 226294 531530 226350
rect 531598 226294 531654 226350
rect 531722 226294 531778 226350
rect 531846 226294 531902 226350
rect 531474 226170 531530 226226
rect 531598 226170 531654 226226
rect 531722 226170 531778 226226
rect 531846 226170 531902 226226
rect 531474 226046 531530 226102
rect 531598 226046 531654 226102
rect 531722 226046 531778 226102
rect 531846 226046 531902 226102
rect 531474 225922 531530 225978
rect 531598 225922 531654 225978
rect 531722 225922 531778 225978
rect 531846 225922 531902 225978
rect 531474 208294 531530 208350
rect 531598 208294 531654 208350
rect 531722 208294 531778 208350
rect 531846 208294 531902 208350
rect 531474 208170 531530 208226
rect 531598 208170 531654 208226
rect 531722 208170 531778 208226
rect 531846 208170 531902 208226
rect 531474 208046 531530 208102
rect 531598 208046 531654 208102
rect 531722 208046 531778 208102
rect 531846 208046 531902 208102
rect 531474 207922 531530 207978
rect 531598 207922 531654 207978
rect 531722 207922 531778 207978
rect 531846 207922 531902 207978
rect 531474 190294 531530 190350
rect 531598 190294 531654 190350
rect 531722 190294 531778 190350
rect 531846 190294 531902 190350
rect 531474 190170 531530 190226
rect 531598 190170 531654 190226
rect 531722 190170 531778 190226
rect 531846 190170 531902 190226
rect 531474 190046 531530 190102
rect 531598 190046 531654 190102
rect 531722 190046 531778 190102
rect 531846 190046 531902 190102
rect 531474 189922 531530 189978
rect 531598 189922 531654 189978
rect 531722 189922 531778 189978
rect 531846 189922 531902 189978
rect 531474 172294 531530 172350
rect 531598 172294 531654 172350
rect 531722 172294 531778 172350
rect 531846 172294 531902 172350
rect 531474 172170 531530 172226
rect 531598 172170 531654 172226
rect 531722 172170 531778 172226
rect 531846 172170 531902 172226
rect 531474 172046 531530 172102
rect 531598 172046 531654 172102
rect 531722 172046 531778 172102
rect 531846 172046 531902 172102
rect 531474 171922 531530 171978
rect 531598 171922 531654 171978
rect 531722 171922 531778 171978
rect 531846 171922 531902 171978
rect 531474 154294 531530 154350
rect 531598 154294 531654 154350
rect 531722 154294 531778 154350
rect 531846 154294 531902 154350
rect 531474 154170 531530 154226
rect 531598 154170 531654 154226
rect 531722 154170 531778 154226
rect 531846 154170 531902 154226
rect 531474 154046 531530 154102
rect 531598 154046 531654 154102
rect 531722 154046 531778 154102
rect 531846 154046 531902 154102
rect 531474 153922 531530 153978
rect 531598 153922 531654 153978
rect 531722 153922 531778 153978
rect 531846 153922 531902 153978
rect 531474 136294 531530 136350
rect 531598 136294 531654 136350
rect 531722 136294 531778 136350
rect 531846 136294 531902 136350
rect 531474 136170 531530 136226
rect 531598 136170 531654 136226
rect 531722 136170 531778 136226
rect 531846 136170 531902 136226
rect 531474 136046 531530 136102
rect 531598 136046 531654 136102
rect 531722 136046 531778 136102
rect 531846 136046 531902 136102
rect 531474 135922 531530 135978
rect 531598 135922 531654 135978
rect 531722 135922 531778 135978
rect 531846 135922 531902 135978
rect 531474 118294 531530 118350
rect 531598 118294 531654 118350
rect 531722 118294 531778 118350
rect 531846 118294 531902 118350
rect 531474 118170 531530 118226
rect 531598 118170 531654 118226
rect 531722 118170 531778 118226
rect 531846 118170 531902 118226
rect 531474 118046 531530 118102
rect 531598 118046 531654 118102
rect 531722 118046 531778 118102
rect 531846 118046 531902 118102
rect 531474 117922 531530 117978
rect 531598 117922 531654 117978
rect 531722 117922 531778 117978
rect 531846 117922 531902 117978
rect 531474 100294 531530 100350
rect 531598 100294 531654 100350
rect 531722 100294 531778 100350
rect 531846 100294 531902 100350
rect 531474 100170 531530 100226
rect 531598 100170 531654 100226
rect 531722 100170 531778 100226
rect 531846 100170 531902 100226
rect 531474 100046 531530 100102
rect 531598 100046 531654 100102
rect 531722 100046 531778 100102
rect 531846 100046 531902 100102
rect 531474 99922 531530 99978
rect 531598 99922 531654 99978
rect 531722 99922 531778 99978
rect 531846 99922 531902 99978
rect 531474 82294 531530 82350
rect 531598 82294 531654 82350
rect 531722 82294 531778 82350
rect 531846 82294 531902 82350
rect 531474 82170 531530 82226
rect 531598 82170 531654 82226
rect 531722 82170 531778 82226
rect 531846 82170 531902 82226
rect 531474 82046 531530 82102
rect 531598 82046 531654 82102
rect 531722 82046 531778 82102
rect 531846 82046 531902 82102
rect 531474 81922 531530 81978
rect 531598 81922 531654 81978
rect 531722 81922 531778 81978
rect 531846 81922 531902 81978
rect 527754 58294 527810 58350
rect 527878 58294 527934 58350
rect 528002 58294 528058 58350
rect 528126 58294 528182 58350
rect 527754 58170 527810 58226
rect 527878 58170 527934 58226
rect 528002 58170 528058 58226
rect 528126 58170 528182 58226
rect 527754 58046 527810 58102
rect 527878 58046 527934 58102
rect 528002 58046 528058 58102
rect 528126 58046 528182 58102
rect 527754 57922 527810 57978
rect 527878 57922 527934 57978
rect 528002 57922 528058 57978
rect 528126 57922 528182 57978
rect 527754 40294 527810 40350
rect 527878 40294 527934 40350
rect 528002 40294 528058 40350
rect 528126 40294 528182 40350
rect 527754 40170 527810 40226
rect 527878 40170 527934 40226
rect 528002 40170 528058 40226
rect 528126 40170 528182 40226
rect 527754 40046 527810 40102
rect 527878 40046 527934 40102
rect 528002 40046 528058 40102
rect 528126 40046 528182 40102
rect 527754 39922 527810 39978
rect 527878 39922 527934 39978
rect 528002 39922 528058 39978
rect 528126 39922 528182 39978
rect 527754 22294 527810 22350
rect 527878 22294 527934 22350
rect 528002 22294 528058 22350
rect 528126 22294 528182 22350
rect 527754 22170 527810 22226
rect 527878 22170 527934 22226
rect 528002 22170 528058 22226
rect 528126 22170 528182 22226
rect 527754 22046 527810 22102
rect 527878 22046 527934 22102
rect 528002 22046 528058 22102
rect 528126 22046 528182 22102
rect 527754 21922 527810 21978
rect 527878 21922 527934 21978
rect 528002 21922 528058 21978
rect 528126 21922 528182 21978
rect 531474 64294 531530 64350
rect 531598 64294 531654 64350
rect 531722 64294 531778 64350
rect 531846 64294 531902 64350
rect 531474 64170 531530 64226
rect 531598 64170 531654 64226
rect 531722 64170 531778 64226
rect 531846 64170 531902 64226
rect 531474 64046 531530 64102
rect 531598 64046 531654 64102
rect 531722 64046 531778 64102
rect 531846 64046 531902 64102
rect 531474 63922 531530 63978
rect 531598 63922 531654 63978
rect 531722 63922 531778 63978
rect 531846 63922 531902 63978
rect 531474 46294 531530 46350
rect 531598 46294 531654 46350
rect 531722 46294 531778 46350
rect 531846 46294 531902 46350
rect 531474 46170 531530 46226
rect 531598 46170 531654 46226
rect 531722 46170 531778 46226
rect 531846 46170 531902 46226
rect 531474 46046 531530 46102
rect 531598 46046 531654 46102
rect 531722 46046 531778 46102
rect 531846 46046 531902 46102
rect 531474 45922 531530 45978
rect 531598 45922 531654 45978
rect 531722 45922 531778 45978
rect 531846 45922 531902 45978
rect 558474 310294 558530 310350
rect 558598 310294 558654 310350
rect 558722 310294 558778 310350
rect 558846 310294 558902 310350
rect 558474 310170 558530 310226
rect 558598 310170 558654 310226
rect 558722 310170 558778 310226
rect 558846 310170 558902 310226
rect 558474 310046 558530 310102
rect 558598 310046 558654 310102
rect 558722 310046 558778 310102
rect 558846 310046 558902 310102
rect 558474 309922 558530 309978
rect 558598 309922 558654 309978
rect 558722 309922 558778 309978
rect 558846 309922 558902 309978
rect 558474 292294 558530 292350
rect 558598 292294 558654 292350
rect 558722 292294 558778 292350
rect 558846 292294 558902 292350
rect 558474 292170 558530 292226
rect 558598 292170 558654 292226
rect 558722 292170 558778 292226
rect 558846 292170 558902 292226
rect 558474 292046 558530 292102
rect 558598 292046 558654 292102
rect 558722 292046 558778 292102
rect 558846 292046 558902 292102
rect 558474 291922 558530 291978
rect 558598 291922 558654 291978
rect 558722 291922 558778 291978
rect 558846 291922 558902 291978
rect 558474 274294 558530 274350
rect 558598 274294 558654 274350
rect 558722 274294 558778 274350
rect 558846 274294 558902 274350
rect 558474 274170 558530 274226
rect 558598 274170 558654 274226
rect 558722 274170 558778 274226
rect 558846 274170 558902 274226
rect 558474 274046 558530 274102
rect 558598 274046 558654 274102
rect 558722 274046 558778 274102
rect 558846 274046 558902 274102
rect 558474 273922 558530 273978
rect 558598 273922 558654 273978
rect 558722 273922 558778 273978
rect 558846 273922 558902 273978
rect 531474 28294 531530 28350
rect 531598 28294 531654 28350
rect 531722 28294 531778 28350
rect 531846 28294 531902 28350
rect 531474 28170 531530 28226
rect 531598 28170 531654 28226
rect 531722 28170 531778 28226
rect 531846 28170 531902 28226
rect 531474 28046 531530 28102
rect 531598 28046 531654 28102
rect 531722 28046 531778 28102
rect 531846 28046 531902 28102
rect 531474 27922 531530 27978
rect 531598 27922 531654 27978
rect 531722 27922 531778 27978
rect 531846 27922 531902 27978
rect 538470 28294 538526 28350
rect 538594 28294 538650 28350
rect 538470 28170 538526 28226
rect 538594 28170 538650 28226
rect 538470 28046 538526 28102
rect 538594 28046 538650 28102
rect 538470 27922 538526 27978
rect 538594 27922 538650 27978
rect 531474 10294 531530 10350
rect 531598 10294 531654 10350
rect 531722 10294 531778 10350
rect 531846 10294 531902 10350
rect 531474 10170 531530 10226
rect 531598 10170 531654 10226
rect 531722 10170 531778 10226
rect 531846 10170 531902 10226
rect 531474 10046 531530 10102
rect 531598 10046 531654 10102
rect 531722 10046 531778 10102
rect 531846 10046 531902 10102
rect 531474 9922 531530 9978
rect 531598 9922 531654 9978
rect 531722 9922 531778 9978
rect 531846 9922 531902 9978
rect 527754 4294 527810 4350
rect 527878 4294 527934 4350
rect 528002 4294 528058 4350
rect 528126 4294 528182 4350
rect 527754 4170 527810 4226
rect 527878 4170 527934 4226
rect 528002 4170 528058 4226
rect 528126 4170 528182 4226
rect 527754 4046 527810 4102
rect 527878 4046 527934 4102
rect 528002 4046 528058 4102
rect 528126 4046 528182 4102
rect 527754 3922 527810 3978
rect 527878 3922 527934 3978
rect 528002 3922 528058 3978
rect 528126 3922 528182 3978
rect 501676 3332 501732 3358
rect 501676 3302 501732 3332
rect 512092 422 512148 478
rect 510748 242 510804 298
rect 504140 62 504196 118
rect 500754 -1176 500810 -1120
rect 500878 -1176 500934 -1120
rect 501002 -1176 501058 -1120
rect 501126 -1176 501182 -1120
rect 500754 -1300 500810 -1244
rect 500878 -1300 500934 -1244
rect 501002 -1300 501058 -1244
rect 501126 -1300 501182 -1244
rect 500754 -1424 500810 -1368
rect 500878 -1424 500934 -1368
rect 501002 -1424 501058 -1368
rect 501126 -1424 501182 -1368
rect 500754 -1548 500810 -1492
rect 500878 -1548 500934 -1492
rect 501002 -1548 501058 -1492
rect 501126 -1548 501182 -1492
rect 529228 5282 529284 5338
rect 527754 -216 527810 -160
rect 527878 -216 527934 -160
rect 528002 -216 528058 -160
rect 528126 -216 528182 -160
rect 527754 -340 527810 -284
rect 527878 -340 527934 -284
rect 528002 -340 528058 -284
rect 528126 -340 528182 -284
rect 527754 -464 527810 -408
rect 527878 -464 527934 -408
rect 528002 -464 528058 -408
rect 528126 -464 528182 -408
rect 527754 -588 527810 -532
rect 527878 -588 527934 -532
rect 528002 -588 528058 -532
rect 528126 -588 528182 -532
rect 538470 10294 538526 10350
rect 538594 10294 538650 10350
rect 538470 10170 538526 10226
rect 538594 10170 538650 10226
rect 538470 10046 538526 10102
rect 538594 10046 538650 10102
rect 538470 9922 538526 9978
rect 538594 9922 538650 9978
rect 558474 256294 558530 256350
rect 558598 256294 558654 256350
rect 558722 256294 558778 256350
rect 558846 256294 558902 256350
rect 558474 256170 558530 256226
rect 558598 256170 558654 256226
rect 558722 256170 558778 256226
rect 558846 256170 558902 256226
rect 558474 256046 558530 256102
rect 558598 256046 558654 256102
rect 558722 256046 558778 256102
rect 558846 256046 558902 256102
rect 558474 255922 558530 255978
rect 558598 255922 558654 255978
rect 558722 255922 558778 255978
rect 558846 255922 558902 255978
rect 558474 238294 558530 238350
rect 558598 238294 558654 238350
rect 558722 238294 558778 238350
rect 558846 238294 558902 238350
rect 558474 238170 558530 238226
rect 558598 238170 558654 238226
rect 558722 238170 558778 238226
rect 558846 238170 558902 238226
rect 558474 238046 558530 238102
rect 558598 238046 558654 238102
rect 558722 238046 558778 238102
rect 558846 238046 558902 238102
rect 558474 237922 558530 237978
rect 558598 237922 558654 237978
rect 558722 237922 558778 237978
rect 558846 237922 558902 237978
rect 558474 220294 558530 220350
rect 558598 220294 558654 220350
rect 558722 220294 558778 220350
rect 558846 220294 558902 220350
rect 558474 220170 558530 220226
rect 558598 220170 558654 220226
rect 558722 220170 558778 220226
rect 558846 220170 558902 220226
rect 558474 220046 558530 220102
rect 558598 220046 558654 220102
rect 558722 220046 558778 220102
rect 558846 220046 558902 220102
rect 558474 219922 558530 219978
rect 558598 219922 558654 219978
rect 558722 219922 558778 219978
rect 558846 219922 558902 219978
rect 562194 598116 562250 598172
rect 562318 598116 562374 598172
rect 562442 598116 562498 598172
rect 562566 598116 562622 598172
rect 562194 597992 562250 598048
rect 562318 597992 562374 598048
rect 562442 597992 562498 598048
rect 562566 597992 562622 598048
rect 562194 597868 562250 597924
rect 562318 597868 562374 597924
rect 562442 597868 562498 597924
rect 562566 597868 562622 597924
rect 562194 597744 562250 597800
rect 562318 597744 562374 597800
rect 562442 597744 562498 597800
rect 562566 597744 562622 597800
rect 589194 597156 589250 597212
rect 589318 597156 589374 597212
rect 589442 597156 589498 597212
rect 589566 597156 589622 597212
rect 589194 597032 589250 597088
rect 589318 597032 589374 597088
rect 589442 597032 589498 597088
rect 589566 597032 589622 597088
rect 589194 596908 589250 596964
rect 589318 596908 589374 596964
rect 589442 596908 589498 596964
rect 589566 596908 589622 596964
rect 589194 596784 589250 596840
rect 589318 596784 589374 596840
rect 589442 596784 589498 596840
rect 589566 596784 589622 596840
rect 562194 586294 562250 586350
rect 562318 586294 562374 586350
rect 562442 586294 562498 586350
rect 562566 586294 562622 586350
rect 562194 586170 562250 586226
rect 562318 586170 562374 586226
rect 562442 586170 562498 586226
rect 562566 586170 562622 586226
rect 562194 586046 562250 586102
rect 562318 586046 562374 586102
rect 562442 586046 562498 586102
rect 562566 586046 562622 586102
rect 562194 585922 562250 585978
rect 562318 585922 562374 585978
rect 562442 585922 562498 585978
rect 562566 585922 562622 585978
rect 562194 568294 562250 568350
rect 562318 568294 562374 568350
rect 562442 568294 562498 568350
rect 562566 568294 562622 568350
rect 562194 568170 562250 568226
rect 562318 568170 562374 568226
rect 562442 568170 562498 568226
rect 562566 568170 562622 568226
rect 562194 568046 562250 568102
rect 562318 568046 562374 568102
rect 562442 568046 562498 568102
rect 562566 568046 562622 568102
rect 562194 567922 562250 567978
rect 562318 567922 562374 567978
rect 562442 567922 562498 567978
rect 562566 567922 562622 567978
rect 562194 550294 562250 550350
rect 562318 550294 562374 550350
rect 562442 550294 562498 550350
rect 562566 550294 562622 550350
rect 562194 550170 562250 550226
rect 562318 550170 562374 550226
rect 562442 550170 562498 550226
rect 562566 550170 562622 550226
rect 562194 550046 562250 550102
rect 562318 550046 562374 550102
rect 562442 550046 562498 550102
rect 562566 550046 562622 550102
rect 562194 549922 562250 549978
rect 562318 549922 562374 549978
rect 562442 549922 562498 549978
rect 562566 549922 562622 549978
rect 562194 532294 562250 532350
rect 562318 532294 562374 532350
rect 562442 532294 562498 532350
rect 562566 532294 562622 532350
rect 562194 532170 562250 532226
rect 562318 532170 562374 532226
rect 562442 532170 562498 532226
rect 562566 532170 562622 532226
rect 562194 532046 562250 532102
rect 562318 532046 562374 532102
rect 562442 532046 562498 532102
rect 562566 532046 562622 532102
rect 562194 531922 562250 531978
rect 562318 531922 562374 531978
rect 562442 531922 562498 531978
rect 562566 531922 562622 531978
rect 562194 514294 562250 514350
rect 562318 514294 562374 514350
rect 562442 514294 562498 514350
rect 562566 514294 562622 514350
rect 562194 514170 562250 514226
rect 562318 514170 562374 514226
rect 562442 514170 562498 514226
rect 562566 514170 562622 514226
rect 562194 514046 562250 514102
rect 562318 514046 562374 514102
rect 562442 514046 562498 514102
rect 562566 514046 562622 514102
rect 562194 513922 562250 513978
rect 562318 513922 562374 513978
rect 562442 513922 562498 513978
rect 562566 513922 562622 513978
rect 562194 496294 562250 496350
rect 562318 496294 562374 496350
rect 562442 496294 562498 496350
rect 562566 496294 562622 496350
rect 562194 496170 562250 496226
rect 562318 496170 562374 496226
rect 562442 496170 562498 496226
rect 562566 496170 562622 496226
rect 562194 496046 562250 496102
rect 562318 496046 562374 496102
rect 562442 496046 562498 496102
rect 562566 496046 562622 496102
rect 562194 495922 562250 495978
rect 562318 495922 562374 495978
rect 562442 495922 562498 495978
rect 562566 495922 562622 495978
rect 562194 478294 562250 478350
rect 562318 478294 562374 478350
rect 562442 478294 562498 478350
rect 562566 478294 562622 478350
rect 562194 478170 562250 478226
rect 562318 478170 562374 478226
rect 562442 478170 562498 478226
rect 562566 478170 562622 478226
rect 562194 478046 562250 478102
rect 562318 478046 562374 478102
rect 562442 478046 562498 478102
rect 562566 478046 562622 478102
rect 562194 477922 562250 477978
rect 562318 477922 562374 477978
rect 562442 477922 562498 477978
rect 562566 477922 562622 477978
rect 562194 460294 562250 460350
rect 562318 460294 562374 460350
rect 562442 460294 562498 460350
rect 562566 460294 562622 460350
rect 562194 460170 562250 460226
rect 562318 460170 562374 460226
rect 562442 460170 562498 460226
rect 562566 460170 562622 460226
rect 562194 460046 562250 460102
rect 562318 460046 562374 460102
rect 562442 460046 562498 460102
rect 562566 460046 562622 460102
rect 562194 459922 562250 459978
rect 562318 459922 562374 459978
rect 562442 459922 562498 459978
rect 562566 459922 562622 459978
rect 562194 442294 562250 442350
rect 562318 442294 562374 442350
rect 562442 442294 562498 442350
rect 562566 442294 562622 442350
rect 562194 442170 562250 442226
rect 562318 442170 562374 442226
rect 562442 442170 562498 442226
rect 562566 442170 562622 442226
rect 562194 442046 562250 442102
rect 562318 442046 562374 442102
rect 562442 442046 562498 442102
rect 562566 442046 562622 442102
rect 562194 441922 562250 441978
rect 562318 441922 562374 441978
rect 562442 441922 562498 441978
rect 562566 441922 562622 441978
rect 562194 424294 562250 424350
rect 562318 424294 562374 424350
rect 562442 424294 562498 424350
rect 562566 424294 562622 424350
rect 562194 424170 562250 424226
rect 562318 424170 562374 424226
rect 562442 424170 562498 424226
rect 562566 424170 562622 424226
rect 562194 424046 562250 424102
rect 562318 424046 562374 424102
rect 562442 424046 562498 424102
rect 562566 424046 562622 424102
rect 562194 423922 562250 423978
rect 562318 423922 562374 423978
rect 562442 423922 562498 423978
rect 562566 423922 562622 423978
rect 562194 406294 562250 406350
rect 562318 406294 562374 406350
rect 562442 406294 562498 406350
rect 562566 406294 562622 406350
rect 562194 406170 562250 406226
rect 562318 406170 562374 406226
rect 562442 406170 562498 406226
rect 562566 406170 562622 406226
rect 562194 406046 562250 406102
rect 562318 406046 562374 406102
rect 562442 406046 562498 406102
rect 562566 406046 562622 406102
rect 562194 405922 562250 405978
rect 562318 405922 562374 405978
rect 562442 405922 562498 405978
rect 562566 405922 562622 405978
rect 562194 388294 562250 388350
rect 562318 388294 562374 388350
rect 562442 388294 562498 388350
rect 562566 388294 562622 388350
rect 562194 388170 562250 388226
rect 562318 388170 562374 388226
rect 562442 388170 562498 388226
rect 562566 388170 562622 388226
rect 562194 388046 562250 388102
rect 562318 388046 562374 388102
rect 562442 388046 562498 388102
rect 562566 388046 562622 388102
rect 562194 387922 562250 387978
rect 562318 387922 562374 387978
rect 562442 387922 562498 387978
rect 562566 387922 562622 387978
rect 562194 370294 562250 370350
rect 562318 370294 562374 370350
rect 562442 370294 562498 370350
rect 562566 370294 562622 370350
rect 562194 370170 562250 370226
rect 562318 370170 562374 370226
rect 562442 370170 562498 370226
rect 562566 370170 562622 370226
rect 562194 370046 562250 370102
rect 562318 370046 562374 370102
rect 562442 370046 562498 370102
rect 562566 370046 562622 370102
rect 562194 369922 562250 369978
rect 562318 369922 562374 369978
rect 562442 369922 562498 369978
rect 562566 369922 562622 369978
rect 584668 368702 584724 368758
rect 592914 598116 592970 598172
rect 593038 598116 593094 598172
rect 593162 598116 593218 598172
rect 593286 598116 593342 598172
rect 592914 597992 592970 598048
rect 593038 597992 593094 598048
rect 593162 597992 593218 598048
rect 593286 597992 593342 598048
rect 592914 597868 592970 597924
rect 593038 597868 593094 597924
rect 593162 597868 593218 597924
rect 593286 597868 593342 597924
rect 592914 597744 592970 597800
rect 593038 597744 593094 597800
rect 593162 597744 593218 597800
rect 593286 597744 593342 597800
rect 589194 580294 589250 580350
rect 589318 580294 589374 580350
rect 589442 580294 589498 580350
rect 589566 580294 589622 580350
rect 589194 580170 589250 580226
rect 589318 580170 589374 580226
rect 589442 580170 589498 580226
rect 589566 580170 589622 580226
rect 589194 580046 589250 580102
rect 589318 580046 589374 580102
rect 589442 580046 589498 580102
rect 589566 580046 589622 580102
rect 589194 579922 589250 579978
rect 589318 579922 589374 579978
rect 589442 579922 589498 579978
rect 589566 579922 589622 579978
rect 589194 562294 589250 562350
rect 589318 562294 589374 562350
rect 589442 562294 589498 562350
rect 589566 562294 589622 562350
rect 589194 562170 589250 562226
rect 589318 562170 589374 562226
rect 589442 562170 589498 562226
rect 589566 562170 589622 562226
rect 589194 562046 589250 562102
rect 589318 562046 589374 562102
rect 589442 562046 589498 562102
rect 589566 562046 589622 562102
rect 589194 561922 589250 561978
rect 589318 561922 589374 561978
rect 589442 561922 589498 561978
rect 589566 561922 589622 561978
rect 589194 544294 589250 544350
rect 589318 544294 589374 544350
rect 589442 544294 589498 544350
rect 589566 544294 589622 544350
rect 589194 544170 589250 544226
rect 589318 544170 589374 544226
rect 589442 544170 589498 544226
rect 589566 544170 589622 544226
rect 589194 544046 589250 544102
rect 589318 544046 589374 544102
rect 589442 544046 589498 544102
rect 589566 544046 589622 544102
rect 589194 543922 589250 543978
rect 589318 543922 589374 543978
rect 589442 543922 589498 543978
rect 589566 543922 589622 543978
rect 589194 526294 589250 526350
rect 589318 526294 589374 526350
rect 589442 526294 589498 526350
rect 589566 526294 589622 526350
rect 589194 526170 589250 526226
rect 589318 526170 589374 526226
rect 589442 526170 589498 526226
rect 589566 526170 589622 526226
rect 589194 526046 589250 526102
rect 589318 526046 589374 526102
rect 589442 526046 589498 526102
rect 589566 526046 589622 526102
rect 589194 525922 589250 525978
rect 589318 525922 589374 525978
rect 589442 525922 589498 525978
rect 589566 525922 589622 525978
rect 589194 508294 589250 508350
rect 589318 508294 589374 508350
rect 589442 508294 589498 508350
rect 589566 508294 589622 508350
rect 589194 508170 589250 508226
rect 589318 508170 589374 508226
rect 589442 508170 589498 508226
rect 589566 508170 589622 508226
rect 589194 508046 589250 508102
rect 589318 508046 589374 508102
rect 589442 508046 589498 508102
rect 589566 508046 589622 508102
rect 589194 507922 589250 507978
rect 589318 507922 589374 507978
rect 589442 507922 589498 507978
rect 589566 507922 589622 507978
rect 589194 490294 589250 490350
rect 589318 490294 589374 490350
rect 589442 490294 589498 490350
rect 589566 490294 589622 490350
rect 589194 490170 589250 490226
rect 589318 490170 589374 490226
rect 589442 490170 589498 490226
rect 589566 490170 589622 490226
rect 589194 490046 589250 490102
rect 589318 490046 589374 490102
rect 589442 490046 589498 490102
rect 589566 490046 589622 490102
rect 589194 489922 589250 489978
rect 589318 489922 589374 489978
rect 589442 489922 589498 489978
rect 589566 489922 589622 489978
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 592914 586294 592970 586350
rect 593038 586294 593094 586350
rect 593162 586294 593218 586350
rect 593286 586294 593342 586350
rect 592914 586170 592970 586226
rect 593038 586170 593094 586226
rect 593162 586170 593218 586226
rect 593286 586170 593342 586226
rect 592914 586046 592970 586102
rect 593038 586046 593094 586102
rect 593162 586046 593218 586102
rect 593286 586046 593342 586102
rect 592914 585922 592970 585978
rect 593038 585922 593094 585978
rect 593162 585922 593218 585978
rect 593286 585922 593342 585978
rect 592914 568294 592970 568350
rect 593038 568294 593094 568350
rect 593162 568294 593218 568350
rect 593286 568294 593342 568350
rect 592914 568170 592970 568226
rect 593038 568170 593094 568226
rect 593162 568170 593218 568226
rect 593286 568170 593342 568226
rect 592914 568046 592970 568102
rect 593038 568046 593094 568102
rect 593162 568046 593218 568102
rect 593286 568046 593342 568102
rect 592914 567922 592970 567978
rect 593038 567922 593094 567978
rect 593162 567922 593218 567978
rect 593286 567922 593342 567978
rect 592914 550294 592970 550350
rect 593038 550294 593094 550350
rect 593162 550294 593218 550350
rect 593286 550294 593342 550350
rect 592914 550170 592970 550226
rect 593038 550170 593094 550226
rect 593162 550170 593218 550226
rect 593286 550170 593342 550226
rect 592914 550046 592970 550102
rect 593038 550046 593094 550102
rect 593162 550046 593218 550102
rect 593286 550046 593342 550102
rect 592914 549922 592970 549978
rect 593038 549922 593094 549978
rect 593162 549922 593218 549978
rect 593286 549922 593342 549978
rect 592914 532294 592970 532350
rect 593038 532294 593094 532350
rect 593162 532294 593218 532350
rect 593286 532294 593342 532350
rect 592914 532170 592970 532226
rect 593038 532170 593094 532226
rect 593162 532170 593218 532226
rect 593286 532170 593342 532226
rect 592914 532046 592970 532102
rect 593038 532046 593094 532102
rect 593162 532046 593218 532102
rect 593286 532046 593342 532102
rect 592914 531922 592970 531978
rect 593038 531922 593094 531978
rect 593162 531922 593218 531978
rect 593286 531922 593342 531978
rect 592914 514294 592970 514350
rect 593038 514294 593094 514350
rect 593162 514294 593218 514350
rect 593286 514294 593342 514350
rect 592914 514170 592970 514226
rect 593038 514170 593094 514226
rect 593162 514170 593218 514226
rect 593286 514170 593342 514226
rect 592914 514046 592970 514102
rect 593038 514046 593094 514102
rect 593162 514046 593218 514102
rect 593286 514046 593342 514102
rect 592914 513922 592970 513978
rect 593038 513922 593094 513978
rect 593162 513922 593218 513978
rect 593286 513922 593342 513978
rect 592914 496294 592970 496350
rect 593038 496294 593094 496350
rect 593162 496294 593218 496350
rect 593286 496294 593342 496350
rect 592914 496170 592970 496226
rect 593038 496170 593094 496226
rect 593162 496170 593218 496226
rect 593286 496170 593342 496226
rect 592914 496046 592970 496102
rect 593038 496046 593094 496102
rect 593162 496046 593218 496102
rect 593286 496046 593342 496102
rect 592914 495922 592970 495978
rect 593038 495922 593094 495978
rect 593162 495922 593218 495978
rect 593286 495922 593342 495978
rect 589194 472294 589250 472350
rect 589318 472294 589374 472350
rect 589442 472294 589498 472350
rect 589566 472294 589622 472350
rect 589194 472170 589250 472226
rect 589318 472170 589374 472226
rect 589442 472170 589498 472226
rect 589566 472170 589622 472226
rect 589194 472046 589250 472102
rect 589318 472046 589374 472102
rect 589442 472046 589498 472102
rect 589566 472046 589622 472102
rect 589194 471922 589250 471978
rect 589318 471922 589374 471978
rect 589442 471922 589498 471978
rect 589566 471922 589622 471978
rect 589194 454294 589250 454350
rect 589318 454294 589374 454350
rect 589442 454294 589498 454350
rect 589566 454294 589622 454350
rect 589194 454170 589250 454226
rect 589318 454170 589374 454226
rect 589442 454170 589498 454226
rect 589566 454170 589622 454226
rect 589194 454046 589250 454102
rect 589318 454046 589374 454102
rect 589442 454046 589498 454102
rect 589566 454046 589622 454102
rect 589194 453922 589250 453978
rect 589318 453922 589374 453978
rect 589442 453922 589498 453978
rect 589566 453922 589622 453978
rect 589194 436294 589250 436350
rect 589318 436294 589374 436350
rect 589442 436294 589498 436350
rect 589566 436294 589622 436350
rect 589194 436170 589250 436226
rect 589318 436170 589374 436226
rect 589442 436170 589498 436226
rect 589566 436170 589622 436226
rect 589194 436046 589250 436102
rect 589318 436046 589374 436102
rect 589442 436046 589498 436102
rect 589566 436046 589622 436102
rect 589194 435922 589250 435978
rect 589318 435922 589374 435978
rect 589442 435922 589498 435978
rect 589566 435922 589622 435978
rect 589194 418294 589250 418350
rect 589318 418294 589374 418350
rect 589442 418294 589498 418350
rect 589566 418294 589622 418350
rect 589194 418170 589250 418226
rect 589318 418170 589374 418226
rect 589442 418170 589498 418226
rect 589566 418170 589622 418226
rect 589194 418046 589250 418102
rect 589318 418046 589374 418102
rect 589442 418046 589498 418102
rect 589566 418046 589622 418102
rect 589194 417922 589250 417978
rect 589318 417922 589374 417978
rect 589442 417922 589498 417978
rect 589566 417922 589622 417978
rect 589194 400294 589250 400350
rect 589318 400294 589374 400350
rect 589442 400294 589498 400350
rect 589566 400294 589622 400350
rect 589194 400170 589250 400226
rect 589318 400170 589374 400226
rect 589442 400170 589498 400226
rect 589566 400170 589622 400226
rect 589194 400046 589250 400102
rect 589318 400046 589374 400102
rect 589442 400046 589498 400102
rect 589566 400046 589622 400102
rect 589194 399922 589250 399978
rect 589318 399922 589374 399978
rect 589442 399922 589498 399978
rect 589566 399922 589622 399978
rect 589194 382294 589250 382350
rect 589318 382294 589374 382350
rect 589442 382294 589498 382350
rect 589566 382294 589622 382350
rect 589194 382170 589250 382226
rect 589318 382170 589374 382226
rect 589442 382170 589498 382226
rect 589566 382170 589622 382226
rect 589194 382046 589250 382102
rect 589318 382046 589374 382102
rect 589442 382046 589498 382102
rect 589566 382046 589622 382102
rect 589194 381922 589250 381978
rect 589318 381922 589374 381978
rect 589442 381922 589498 381978
rect 589566 381922 589622 381978
rect 562194 352294 562250 352350
rect 562318 352294 562374 352350
rect 562442 352294 562498 352350
rect 562566 352294 562622 352350
rect 562194 352170 562250 352226
rect 562318 352170 562374 352226
rect 562442 352170 562498 352226
rect 562566 352170 562622 352226
rect 562194 352046 562250 352102
rect 562318 352046 562374 352102
rect 562442 352046 562498 352102
rect 562566 352046 562622 352102
rect 562194 351922 562250 351978
rect 562318 351922 562374 351978
rect 562442 351922 562498 351978
rect 562566 351922 562622 351978
rect 562194 334294 562250 334350
rect 562318 334294 562374 334350
rect 562442 334294 562498 334350
rect 562566 334294 562622 334350
rect 562194 334170 562250 334226
rect 562318 334170 562374 334226
rect 562442 334170 562498 334226
rect 562566 334170 562622 334226
rect 562194 334046 562250 334102
rect 562318 334046 562374 334102
rect 562442 334046 562498 334102
rect 562566 334046 562622 334102
rect 562194 333922 562250 333978
rect 562318 333922 562374 333978
rect 562442 333922 562498 333978
rect 562566 333922 562622 333978
rect 562194 316294 562250 316350
rect 562318 316294 562374 316350
rect 562442 316294 562498 316350
rect 562566 316294 562622 316350
rect 562194 316170 562250 316226
rect 562318 316170 562374 316226
rect 562442 316170 562498 316226
rect 562566 316170 562622 316226
rect 562194 316046 562250 316102
rect 562318 316046 562374 316102
rect 562442 316046 562498 316102
rect 562566 316046 562622 316102
rect 562194 315922 562250 315978
rect 562318 315922 562374 315978
rect 562442 315922 562498 315978
rect 562566 315922 562622 315978
rect 562194 298294 562250 298350
rect 562318 298294 562374 298350
rect 562442 298294 562498 298350
rect 562566 298294 562622 298350
rect 562194 298170 562250 298226
rect 562318 298170 562374 298226
rect 562442 298170 562498 298226
rect 562566 298170 562622 298226
rect 562194 298046 562250 298102
rect 562318 298046 562374 298102
rect 562442 298046 562498 298102
rect 562566 298046 562622 298102
rect 562194 297922 562250 297978
rect 562318 297922 562374 297978
rect 562442 297922 562498 297978
rect 562566 297922 562622 297978
rect 589194 364294 589250 364350
rect 589318 364294 589374 364350
rect 589442 364294 589498 364350
rect 589566 364294 589622 364350
rect 589194 364170 589250 364226
rect 589318 364170 589374 364226
rect 589442 364170 589498 364226
rect 589566 364170 589622 364226
rect 589194 364046 589250 364102
rect 589318 364046 589374 364102
rect 589442 364046 589498 364102
rect 589566 364046 589622 364102
rect 592914 478294 592970 478350
rect 593038 478294 593094 478350
rect 593162 478294 593218 478350
rect 593286 478294 593342 478350
rect 592914 478170 592970 478226
rect 593038 478170 593094 478226
rect 593162 478170 593218 478226
rect 593286 478170 593342 478226
rect 592914 478046 592970 478102
rect 593038 478046 593094 478102
rect 593162 478046 593218 478102
rect 593286 478046 593342 478102
rect 592914 477922 592970 477978
rect 593038 477922 593094 477978
rect 593162 477922 593218 477978
rect 593286 477922 593342 477978
rect 592914 460294 592970 460350
rect 593038 460294 593094 460350
rect 593162 460294 593218 460350
rect 593286 460294 593342 460350
rect 592914 460170 592970 460226
rect 593038 460170 593094 460226
rect 593162 460170 593218 460226
rect 593286 460170 593342 460226
rect 592914 460046 592970 460102
rect 593038 460046 593094 460102
rect 593162 460046 593218 460102
rect 593286 460046 593342 460102
rect 592914 459922 592970 459978
rect 593038 459922 593094 459978
rect 593162 459922 593218 459978
rect 593286 459922 593342 459978
rect 592914 442294 592970 442350
rect 593038 442294 593094 442350
rect 593162 442294 593218 442350
rect 593286 442294 593342 442350
rect 592914 442170 592970 442226
rect 593038 442170 593094 442226
rect 593162 442170 593218 442226
rect 593286 442170 593342 442226
rect 592914 442046 592970 442102
rect 593038 442046 593094 442102
rect 593162 442046 593218 442102
rect 593286 442046 593342 442102
rect 592914 441922 592970 441978
rect 593038 441922 593094 441978
rect 593162 441922 593218 441978
rect 593286 441922 593342 441978
rect 592914 424294 592970 424350
rect 593038 424294 593094 424350
rect 593162 424294 593218 424350
rect 593286 424294 593342 424350
rect 592914 424170 592970 424226
rect 593038 424170 593094 424226
rect 593162 424170 593218 424226
rect 593286 424170 593342 424226
rect 592914 424046 592970 424102
rect 593038 424046 593094 424102
rect 593162 424046 593218 424102
rect 593286 424046 593342 424102
rect 592914 423922 592970 423978
rect 593038 423922 593094 423978
rect 593162 423922 593218 423978
rect 593286 423922 593342 423978
rect 592914 406294 592970 406350
rect 593038 406294 593094 406350
rect 593162 406294 593218 406350
rect 593286 406294 593342 406350
rect 592914 406170 592970 406226
rect 593038 406170 593094 406226
rect 593162 406170 593218 406226
rect 593286 406170 593342 406226
rect 592914 406046 592970 406102
rect 593038 406046 593094 406102
rect 593162 406046 593218 406102
rect 593286 406046 593342 406102
rect 592914 405922 592970 405978
rect 593038 405922 593094 405978
rect 593162 405922 593218 405978
rect 593286 405922 593342 405978
rect 592914 388294 592970 388350
rect 593038 388294 593094 388350
rect 593162 388294 593218 388350
rect 593286 388294 593342 388350
rect 592914 388170 592970 388226
rect 593038 388170 593094 388226
rect 593162 388170 593218 388226
rect 593286 388170 593342 388226
rect 592914 388046 592970 388102
rect 593038 388046 593094 388102
rect 593162 388046 593218 388102
rect 593286 388046 593342 388102
rect 592914 387922 592970 387978
rect 593038 387922 593094 387978
rect 593162 387922 593218 387978
rect 593286 387922 593342 387978
rect 592914 370294 592970 370350
rect 593038 370294 593094 370350
rect 593162 370294 593218 370350
rect 593286 370294 593342 370350
rect 592914 370170 592970 370226
rect 593038 370170 593094 370226
rect 593162 370170 593218 370226
rect 593286 370170 593342 370226
rect 592914 370046 592970 370102
rect 593038 370046 593094 370102
rect 593162 370046 593218 370102
rect 593286 370046 593342 370102
rect 592914 369922 592970 369978
rect 593038 369922 593094 369978
rect 593162 369922 593218 369978
rect 593286 369922 593342 369978
rect 589194 363922 589250 363978
rect 589318 363922 589374 363978
rect 589442 363922 589498 363978
rect 589566 363922 589622 363978
rect 589194 346294 589250 346350
rect 589318 346294 589374 346350
rect 589442 346294 589498 346350
rect 589566 346294 589622 346350
rect 589194 346170 589250 346226
rect 589318 346170 589374 346226
rect 589442 346170 589498 346226
rect 589566 346170 589622 346226
rect 589194 346046 589250 346102
rect 589318 346046 589374 346102
rect 589442 346046 589498 346102
rect 589566 346046 589622 346102
rect 589194 345922 589250 345978
rect 589318 345922 589374 345978
rect 589442 345922 589498 345978
rect 589566 345922 589622 345978
rect 589194 328294 589250 328350
rect 589318 328294 589374 328350
rect 589442 328294 589498 328350
rect 589566 328294 589622 328350
rect 589194 328170 589250 328226
rect 589318 328170 589374 328226
rect 589442 328170 589498 328226
rect 589566 328170 589622 328226
rect 589194 328046 589250 328102
rect 589318 328046 589374 328102
rect 589442 328046 589498 328102
rect 589566 328046 589622 328102
rect 589194 327922 589250 327978
rect 589318 327922 589374 327978
rect 589442 327922 589498 327978
rect 589566 327922 589622 327978
rect 589194 310294 589250 310350
rect 589318 310294 589374 310350
rect 589442 310294 589498 310350
rect 589566 310294 589622 310350
rect 589194 310170 589250 310226
rect 589318 310170 589374 310226
rect 589442 310170 589498 310226
rect 589566 310170 589622 310226
rect 589194 310046 589250 310102
rect 589318 310046 589374 310102
rect 589442 310046 589498 310102
rect 589566 310046 589622 310102
rect 589194 309922 589250 309978
rect 589318 309922 589374 309978
rect 589442 309922 589498 309978
rect 589566 309922 589622 309978
rect 562194 280294 562250 280350
rect 562318 280294 562374 280350
rect 562442 280294 562498 280350
rect 562566 280294 562622 280350
rect 562194 280170 562250 280226
rect 562318 280170 562374 280226
rect 562442 280170 562498 280226
rect 562566 280170 562622 280226
rect 562194 280046 562250 280102
rect 562318 280046 562374 280102
rect 562442 280046 562498 280102
rect 562566 280046 562622 280102
rect 562194 279922 562250 279978
rect 562318 279922 562374 279978
rect 562442 279922 562498 279978
rect 562566 279922 562622 279978
rect 562194 262294 562250 262350
rect 562318 262294 562374 262350
rect 562442 262294 562498 262350
rect 562566 262294 562622 262350
rect 562194 262170 562250 262226
rect 562318 262170 562374 262226
rect 562442 262170 562498 262226
rect 562566 262170 562622 262226
rect 562194 262046 562250 262102
rect 562318 262046 562374 262102
rect 562442 262046 562498 262102
rect 562566 262046 562622 262102
rect 562194 261922 562250 261978
rect 562318 261922 562374 261978
rect 562442 261922 562498 261978
rect 562566 261922 562622 261978
rect 562194 244294 562250 244350
rect 562318 244294 562374 244350
rect 562442 244294 562498 244350
rect 562566 244294 562622 244350
rect 562194 244170 562250 244226
rect 562318 244170 562374 244226
rect 562442 244170 562498 244226
rect 562566 244170 562622 244226
rect 562194 244046 562250 244102
rect 562318 244046 562374 244102
rect 562442 244046 562498 244102
rect 562566 244046 562622 244102
rect 562194 243922 562250 243978
rect 562318 243922 562374 243978
rect 562442 243922 562498 243978
rect 562566 243922 562622 243978
rect 562194 226294 562250 226350
rect 562318 226294 562374 226350
rect 562442 226294 562498 226350
rect 562566 226294 562622 226350
rect 562194 226170 562250 226226
rect 562318 226170 562374 226226
rect 562442 226170 562498 226226
rect 562566 226170 562622 226226
rect 562194 226046 562250 226102
rect 562318 226046 562374 226102
rect 562442 226046 562498 226102
rect 562566 226046 562622 226102
rect 562194 225922 562250 225978
rect 562318 225922 562374 225978
rect 562442 225922 562498 225978
rect 562566 225922 562622 225978
rect 562194 208294 562250 208350
rect 562318 208294 562374 208350
rect 562442 208294 562498 208350
rect 562566 208294 562622 208350
rect 562194 208170 562250 208226
rect 562318 208170 562374 208226
rect 562442 208170 562498 208226
rect 562566 208170 562622 208226
rect 562194 208046 562250 208102
rect 562318 208046 562374 208102
rect 562442 208046 562498 208102
rect 562566 208046 562622 208102
rect 562194 207922 562250 207978
rect 562318 207922 562374 207978
rect 562442 207922 562498 207978
rect 562566 207922 562622 207978
rect 558474 202294 558530 202350
rect 558598 202294 558654 202350
rect 558722 202294 558778 202350
rect 558846 202294 558902 202350
rect 558474 202170 558530 202226
rect 558598 202170 558654 202226
rect 558722 202170 558778 202226
rect 558846 202170 558902 202226
rect 558474 202046 558530 202102
rect 558598 202046 558654 202102
rect 558722 202046 558778 202102
rect 558846 202046 558902 202102
rect 558474 201922 558530 201978
rect 558598 201922 558654 201978
rect 558722 201922 558778 201978
rect 558846 201922 558902 201978
rect 558474 184294 558530 184350
rect 558598 184294 558654 184350
rect 558722 184294 558778 184350
rect 558846 184294 558902 184350
rect 558474 184170 558530 184226
rect 558598 184170 558654 184226
rect 558722 184170 558778 184226
rect 558846 184170 558902 184226
rect 558474 184046 558530 184102
rect 558598 184046 558654 184102
rect 558722 184046 558778 184102
rect 558846 184046 558902 184102
rect 558474 183922 558530 183978
rect 558598 183922 558654 183978
rect 558722 183922 558778 183978
rect 558846 183922 558902 183978
rect 558474 166294 558530 166350
rect 558598 166294 558654 166350
rect 558722 166294 558778 166350
rect 558846 166294 558902 166350
rect 558474 166170 558530 166226
rect 558598 166170 558654 166226
rect 558722 166170 558778 166226
rect 558846 166170 558902 166226
rect 558474 166046 558530 166102
rect 558598 166046 558654 166102
rect 558722 166046 558778 166102
rect 558846 166046 558902 166102
rect 558474 165922 558530 165978
rect 558598 165922 558654 165978
rect 558722 165922 558778 165978
rect 558846 165922 558902 165978
rect 558474 148294 558530 148350
rect 558598 148294 558654 148350
rect 558722 148294 558778 148350
rect 558846 148294 558902 148350
rect 558474 148170 558530 148226
rect 558598 148170 558654 148226
rect 558722 148170 558778 148226
rect 558846 148170 558902 148226
rect 558474 148046 558530 148102
rect 558598 148046 558654 148102
rect 558722 148046 558778 148102
rect 558846 148046 558902 148102
rect 558474 147922 558530 147978
rect 558598 147922 558654 147978
rect 558722 147922 558778 147978
rect 558846 147922 558902 147978
rect 558474 130294 558530 130350
rect 558598 130294 558654 130350
rect 558722 130294 558778 130350
rect 558846 130294 558902 130350
rect 558474 130170 558530 130226
rect 558598 130170 558654 130226
rect 558722 130170 558778 130226
rect 558846 130170 558902 130226
rect 558474 130046 558530 130102
rect 558598 130046 558654 130102
rect 558722 130046 558778 130102
rect 558846 130046 558902 130102
rect 558474 129922 558530 129978
rect 558598 129922 558654 129978
rect 558722 129922 558778 129978
rect 558846 129922 558902 129978
rect 558474 112294 558530 112350
rect 558598 112294 558654 112350
rect 558722 112294 558778 112350
rect 558846 112294 558902 112350
rect 558474 112170 558530 112226
rect 558598 112170 558654 112226
rect 558722 112170 558778 112226
rect 558846 112170 558902 112226
rect 558474 112046 558530 112102
rect 558598 112046 558654 112102
rect 558722 112046 558778 112102
rect 558846 112046 558902 112102
rect 558474 111922 558530 111978
rect 558598 111922 558654 111978
rect 558722 111922 558778 111978
rect 558846 111922 558902 111978
rect 558474 94294 558530 94350
rect 558598 94294 558654 94350
rect 558722 94294 558778 94350
rect 558846 94294 558902 94350
rect 558474 94170 558530 94226
rect 558598 94170 558654 94226
rect 558722 94170 558778 94226
rect 558846 94170 558902 94226
rect 558474 94046 558530 94102
rect 558598 94046 558654 94102
rect 558722 94046 558778 94102
rect 558846 94046 558902 94102
rect 558474 93922 558530 93978
rect 558598 93922 558654 93978
rect 558722 93922 558778 93978
rect 558846 93922 558902 93978
rect 558474 76294 558530 76350
rect 558598 76294 558654 76350
rect 558722 76294 558778 76350
rect 558846 76294 558902 76350
rect 558474 76170 558530 76226
rect 558598 76170 558654 76226
rect 558722 76170 558778 76226
rect 558846 76170 558902 76226
rect 558474 76046 558530 76102
rect 558598 76046 558654 76102
rect 558722 76046 558778 76102
rect 558846 76046 558902 76102
rect 558474 75922 558530 75978
rect 558598 75922 558654 75978
rect 558722 75922 558778 75978
rect 558846 75922 558902 75978
rect 558474 58294 558530 58350
rect 558598 58294 558654 58350
rect 558722 58294 558778 58350
rect 558846 58294 558902 58350
rect 558474 58170 558530 58226
rect 558598 58170 558654 58226
rect 558722 58170 558778 58226
rect 558846 58170 558902 58226
rect 558474 58046 558530 58102
rect 558598 58046 558654 58102
rect 558722 58046 558778 58102
rect 558846 58046 558902 58102
rect 558474 57922 558530 57978
rect 558598 57922 558654 57978
rect 558722 57922 558778 57978
rect 558846 57922 558902 57978
rect 558474 40294 558530 40350
rect 558598 40294 558654 40350
rect 558722 40294 558778 40350
rect 558846 40294 558902 40350
rect 558474 40170 558530 40226
rect 558598 40170 558654 40226
rect 558722 40170 558778 40226
rect 558846 40170 558902 40226
rect 558474 40046 558530 40102
rect 558598 40046 558654 40102
rect 558722 40046 558778 40102
rect 558846 40046 558902 40102
rect 558474 39922 558530 39978
rect 558598 39922 558654 39978
rect 558722 39922 558778 39978
rect 558846 39922 558902 39978
rect 562194 190294 562250 190350
rect 562318 190294 562374 190350
rect 562442 190294 562498 190350
rect 562566 190294 562622 190350
rect 562194 190170 562250 190226
rect 562318 190170 562374 190226
rect 562442 190170 562498 190226
rect 562566 190170 562622 190226
rect 562194 190046 562250 190102
rect 562318 190046 562374 190102
rect 562442 190046 562498 190102
rect 562566 190046 562622 190102
rect 562194 189922 562250 189978
rect 562318 189922 562374 189978
rect 562442 189922 562498 189978
rect 562566 189922 562622 189978
rect 562194 172294 562250 172350
rect 562318 172294 562374 172350
rect 562442 172294 562498 172350
rect 562566 172294 562622 172350
rect 562194 172170 562250 172226
rect 562318 172170 562374 172226
rect 562442 172170 562498 172226
rect 562566 172170 562622 172226
rect 562194 172046 562250 172102
rect 562318 172046 562374 172102
rect 562442 172046 562498 172102
rect 562566 172046 562622 172102
rect 562194 171922 562250 171978
rect 562318 171922 562374 171978
rect 562442 171922 562498 171978
rect 562566 171922 562622 171978
rect 562194 154294 562250 154350
rect 562318 154294 562374 154350
rect 562442 154294 562498 154350
rect 562566 154294 562622 154350
rect 562194 154170 562250 154226
rect 562318 154170 562374 154226
rect 562442 154170 562498 154226
rect 562566 154170 562622 154226
rect 562194 154046 562250 154102
rect 562318 154046 562374 154102
rect 562442 154046 562498 154102
rect 562566 154046 562622 154102
rect 562194 153922 562250 153978
rect 562318 153922 562374 153978
rect 562442 153922 562498 153978
rect 562566 153922 562622 153978
rect 562194 136294 562250 136350
rect 562318 136294 562374 136350
rect 562442 136294 562498 136350
rect 562566 136294 562622 136350
rect 562194 136170 562250 136226
rect 562318 136170 562374 136226
rect 562442 136170 562498 136226
rect 562566 136170 562622 136226
rect 562194 136046 562250 136102
rect 562318 136046 562374 136102
rect 562442 136046 562498 136102
rect 562566 136046 562622 136102
rect 562194 135922 562250 135978
rect 562318 135922 562374 135978
rect 562442 135922 562498 135978
rect 562566 135922 562622 135978
rect 562194 118294 562250 118350
rect 562318 118294 562374 118350
rect 562442 118294 562498 118350
rect 562566 118294 562622 118350
rect 562194 118170 562250 118226
rect 562318 118170 562374 118226
rect 562442 118170 562498 118226
rect 562566 118170 562622 118226
rect 562194 118046 562250 118102
rect 562318 118046 562374 118102
rect 562442 118046 562498 118102
rect 562566 118046 562622 118102
rect 562194 117922 562250 117978
rect 562318 117922 562374 117978
rect 562442 117922 562498 117978
rect 562566 117922 562622 117978
rect 562194 100294 562250 100350
rect 562318 100294 562374 100350
rect 562442 100294 562498 100350
rect 562566 100294 562622 100350
rect 562194 100170 562250 100226
rect 562318 100170 562374 100226
rect 562442 100170 562498 100226
rect 562566 100170 562622 100226
rect 562194 100046 562250 100102
rect 562318 100046 562374 100102
rect 562442 100046 562498 100102
rect 562566 100046 562622 100102
rect 562194 99922 562250 99978
rect 562318 99922 562374 99978
rect 562442 99922 562498 99978
rect 562566 99922 562622 99978
rect 562194 82294 562250 82350
rect 562318 82294 562374 82350
rect 562442 82294 562498 82350
rect 562566 82294 562622 82350
rect 562194 82170 562250 82226
rect 562318 82170 562374 82226
rect 562442 82170 562498 82226
rect 562566 82170 562622 82226
rect 562194 82046 562250 82102
rect 562318 82046 562374 82102
rect 562442 82046 562498 82102
rect 562566 82046 562622 82102
rect 562194 81922 562250 81978
rect 562318 81922 562374 81978
rect 562442 81922 562498 81978
rect 562566 81922 562622 81978
rect 562194 64294 562250 64350
rect 562318 64294 562374 64350
rect 562442 64294 562498 64350
rect 562566 64294 562622 64350
rect 562194 64170 562250 64226
rect 562318 64170 562374 64226
rect 562442 64170 562498 64226
rect 562566 64170 562622 64226
rect 562194 64046 562250 64102
rect 562318 64046 562374 64102
rect 562442 64046 562498 64102
rect 562566 64046 562622 64102
rect 562194 63922 562250 63978
rect 562318 63922 562374 63978
rect 562442 63922 562498 63978
rect 562566 63922 562622 63978
rect 562194 46294 562250 46350
rect 562318 46294 562374 46350
rect 562442 46294 562498 46350
rect 562566 46294 562622 46350
rect 562194 46170 562250 46226
rect 562318 46170 562374 46226
rect 562442 46170 562498 46226
rect 562566 46170 562622 46226
rect 562194 46046 562250 46102
rect 562318 46046 562374 46102
rect 562442 46046 562498 46102
rect 562566 46046 562622 46102
rect 562194 45922 562250 45978
rect 562318 45922 562374 45978
rect 562442 45922 562498 45978
rect 562566 45922 562622 45978
rect 589194 292294 589250 292350
rect 589318 292294 589374 292350
rect 589442 292294 589498 292350
rect 589566 292294 589622 292350
rect 589194 292170 589250 292226
rect 589318 292170 589374 292226
rect 589442 292170 589498 292226
rect 589566 292170 589622 292226
rect 589194 292046 589250 292102
rect 589318 292046 589374 292102
rect 589442 292046 589498 292102
rect 589566 292046 589622 292102
rect 589194 291922 589250 291978
rect 589318 291922 589374 291978
rect 589442 291922 589498 291978
rect 589566 291922 589622 291978
rect 592914 352294 592970 352350
rect 593038 352294 593094 352350
rect 593162 352294 593218 352350
rect 593286 352294 593342 352350
rect 592914 352170 592970 352226
rect 593038 352170 593094 352226
rect 593162 352170 593218 352226
rect 593286 352170 593342 352226
rect 592914 352046 592970 352102
rect 593038 352046 593094 352102
rect 593162 352046 593218 352102
rect 593286 352046 593342 352102
rect 592914 351922 592970 351978
rect 593038 351922 593094 351978
rect 593162 351922 593218 351978
rect 593286 351922 593342 351978
rect 592914 334294 592970 334350
rect 593038 334294 593094 334350
rect 593162 334294 593218 334350
rect 593286 334294 593342 334350
rect 592914 334170 592970 334226
rect 593038 334170 593094 334226
rect 593162 334170 593218 334226
rect 593286 334170 593342 334226
rect 592914 334046 592970 334102
rect 593038 334046 593094 334102
rect 593162 334046 593218 334102
rect 593286 334046 593342 334102
rect 592914 333922 592970 333978
rect 593038 333922 593094 333978
rect 593162 333922 593218 333978
rect 593286 333922 593342 333978
rect 592914 316294 592970 316350
rect 593038 316294 593094 316350
rect 593162 316294 593218 316350
rect 593286 316294 593342 316350
rect 592914 316170 592970 316226
rect 593038 316170 593094 316226
rect 593162 316170 593218 316226
rect 593286 316170 593342 316226
rect 592914 316046 592970 316102
rect 593038 316046 593094 316102
rect 593162 316046 593218 316102
rect 593286 316046 593342 316102
rect 592914 315922 592970 315978
rect 593038 315922 593094 315978
rect 593162 315922 593218 315978
rect 593286 315922 593342 315978
rect 592914 298294 592970 298350
rect 593038 298294 593094 298350
rect 593162 298294 593218 298350
rect 593286 298294 593342 298350
rect 592914 298170 592970 298226
rect 593038 298170 593094 298226
rect 593162 298170 593218 298226
rect 593286 298170 593342 298226
rect 592914 298046 592970 298102
rect 593038 298046 593094 298102
rect 593162 298046 593218 298102
rect 593286 298046 593342 298102
rect 592914 297922 592970 297978
rect 593038 297922 593094 297978
rect 593162 297922 593218 297978
rect 593286 297922 593342 297978
rect 592914 280294 592970 280350
rect 593038 280294 593094 280350
rect 593162 280294 593218 280350
rect 593286 280294 593342 280350
rect 592914 280170 592970 280226
rect 593038 280170 593094 280226
rect 593162 280170 593218 280226
rect 593286 280170 593342 280226
rect 592914 280046 592970 280102
rect 593038 280046 593094 280102
rect 593162 280046 593218 280102
rect 593286 280046 593342 280102
rect 592914 279922 592970 279978
rect 593038 279922 593094 279978
rect 593162 279922 593218 279978
rect 593286 279922 593342 279978
rect 589194 274294 589250 274350
rect 589318 274294 589374 274350
rect 589442 274294 589498 274350
rect 589566 274294 589622 274350
rect 589194 274170 589250 274226
rect 589318 274170 589374 274226
rect 589442 274170 589498 274226
rect 589566 274170 589622 274226
rect 589194 274046 589250 274102
rect 589318 274046 589374 274102
rect 589442 274046 589498 274102
rect 589566 274046 589622 274102
rect 589194 273922 589250 273978
rect 589318 273922 589374 273978
rect 589442 273922 589498 273978
rect 589566 273922 589622 273978
rect 589194 256294 589250 256350
rect 589318 256294 589374 256350
rect 589442 256294 589498 256350
rect 589566 256294 589622 256350
rect 589194 256170 589250 256226
rect 589318 256170 589374 256226
rect 589442 256170 589498 256226
rect 589566 256170 589622 256226
rect 589194 256046 589250 256102
rect 589318 256046 589374 256102
rect 589442 256046 589498 256102
rect 589566 256046 589622 256102
rect 589194 255922 589250 255978
rect 589318 255922 589374 255978
rect 589442 255922 589498 255978
rect 589566 255922 589622 255978
rect 562194 28294 562250 28350
rect 562318 28294 562374 28350
rect 562442 28294 562498 28350
rect 562566 28294 562622 28350
rect 562194 28170 562250 28226
rect 562318 28170 562374 28226
rect 562442 28170 562498 28226
rect 562566 28170 562622 28226
rect 562194 28046 562250 28102
rect 562318 28046 562374 28102
rect 562442 28046 562498 28102
rect 562566 28046 562622 28102
rect 562194 27922 562250 27978
rect 562318 27922 562374 27978
rect 562442 27922 562498 27978
rect 562566 27922 562622 27978
rect 558474 22294 558530 22350
rect 558598 22294 558654 22350
rect 558722 22294 558778 22350
rect 558846 22294 558902 22350
rect 558474 22170 558530 22226
rect 558598 22170 558654 22226
rect 558722 22170 558778 22226
rect 558846 22170 558902 22226
rect 558474 22046 558530 22102
rect 558598 22046 558654 22102
rect 558722 22046 558778 22102
rect 558846 22046 558902 22102
rect 558474 21922 558530 21978
rect 558598 21922 558654 21978
rect 558722 21922 558778 21978
rect 558846 21922 558902 21978
rect 557788 5102 557844 5158
rect 558474 4294 558530 4350
rect 558598 4294 558654 4350
rect 558722 4294 558778 4350
rect 558846 4294 558902 4350
rect 558474 4170 558530 4226
rect 558598 4170 558654 4226
rect 558722 4170 558778 4226
rect 558846 4170 558902 4226
rect 558474 4046 558530 4102
rect 558598 4046 558654 4102
rect 558722 4046 558778 4102
rect 558846 4046 558902 4102
rect 558474 3922 558530 3978
rect 558598 3922 558654 3978
rect 558722 3922 558778 3978
rect 558846 3922 558902 3978
rect 531474 -1176 531530 -1120
rect 531598 -1176 531654 -1120
rect 531722 -1176 531778 -1120
rect 531846 -1176 531902 -1120
rect 531474 -1300 531530 -1244
rect 531598 -1300 531654 -1244
rect 531722 -1300 531778 -1244
rect 531846 -1300 531902 -1244
rect 531474 -1424 531530 -1368
rect 531598 -1424 531654 -1368
rect 531722 -1424 531778 -1368
rect 531846 -1424 531902 -1368
rect 531474 -1548 531530 -1492
rect 531598 -1548 531654 -1492
rect 531722 -1548 531778 -1492
rect 531846 -1548 531902 -1492
rect 558474 -216 558530 -160
rect 558598 -216 558654 -160
rect 558722 -216 558778 -160
rect 558846 -216 558902 -160
rect 558474 -340 558530 -284
rect 558598 -340 558654 -284
rect 558722 -340 558778 -284
rect 558846 -340 558902 -284
rect 558474 -464 558530 -408
rect 558598 -464 558654 -408
rect 558722 -464 558778 -408
rect 558846 -464 558902 -408
rect 558474 -588 558530 -532
rect 558598 -588 558654 -532
rect 558722 -588 558778 -532
rect 558846 -588 558902 -532
rect 589194 238294 589250 238350
rect 589318 238294 589374 238350
rect 589442 238294 589498 238350
rect 589566 238294 589622 238350
rect 589194 238170 589250 238226
rect 589318 238170 589374 238226
rect 589442 238170 589498 238226
rect 589566 238170 589622 238226
rect 589194 238046 589250 238102
rect 589318 238046 589374 238102
rect 589442 238046 589498 238102
rect 589566 238046 589622 238102
rect 589194 237922 589250 237978
rect 589318 237922 589374 237978
rect 589442 237922 589498 237978
rect 589566 237922 589622 237978
rect 589194 220294 589250 220350
rect 589318 220294 589374 220350
rect 589442 220294 589498 220350
rect 589566 220294 589622 220350
rect 589194 220170 589250 220226
rect 589318 220170 589374 220226
rect 589442 220170 589498 220226
rect 589566 220170 589622 220226
rect 589194 220046 589250 220102
rect 589318 220046 589374 220102
rect 589442 220046 589498 220102
rect 589566 220046 589622 220102
rect 589194 219922 589250 219978
rect 589318 219922 589374 219978
rect 589442 219922 589498 219978
rect 589566 219922 589622 219978
rect 589194 202294 589250 202350
rect 589318 202294 589374 202350
rect 589442 202294 589498 202350
rect 589566 202294 589622 202350
rect 589194 202170 589250 202226
rect 589318 202170 589374 202226
rect 589442 202170 589498 202226
rect 589566 202170 589622 202226
rect 589194 202046 589250 202102
rect 589318 202046 589374 202102
rect 589442 202046 589498 202102
rect 589566 202046 589622 202102
rect 589194 201922 589250 201978
rect 589318 201922 589374 201978
rect 589442 201922 589498 201978
rect 589566 201922 589622 201978
rect 589194 184294 589250 184350
rect 589318 184294 589374 184350
rect 589442 184294 589498 184350
rect 589566 184294 589622 184350
rect 589194 184170 589250 184226
rect 589318 184170 589374 184226
rect 589442 184170 589498 184226
rect 589566 184170 589622 184226
rect 589194 184046 589250 184102
rect 589318 184046 589374 184102
rect 589442 184046 589498 184102
rect 589566 184046 589622 184102
rect 589194 183922 589250 183978
rect 589318 183922 589374 183978
rect 589442 183922 589498 183978
rect 589566 183922 589622 183978
rect 589194 166294 589250 166350
rect 589318 166294 589374 166350
rect 589442 166294 589498 166350
rect 589566 166294 589622 166350
rect 589194 166170 589250 166226
rect 589318 166170 589374 166226
rect 589442 166170 589498 166226
rect 589566 166170 589622 166226
rect 589194 166046 589250 166102
rect 589318 166046 589374 166102
rect 589442 166046 589498 166102
rect 589566 166046 589622 166102
rect 589194 165922 589250 165978
rect 589318 165922 589374 165978
rect 589442 165922 589498 165978
rect 589566 165922 589622 165978
rect 592914 262294 592970 262350
rect 593038 262294 593094 262350
rect 593162 262294 593218 262350
rect 593286 262294 593342 262350
rect 592914 262170 592970 262226
rect 593038 262170 593094 262226
rect 593162 262170 593218 262226
rect 593286 262170 593342 262226
rect 592914 262046 592970 262102
rect 593038 262046 593094 262102
rect 593162 262046 593218 262102
rect 593286 262046 593342 262102
rect 592914 261922 592970 261978
rect 593038 261922 593094 261978
rect 593162 261922 593218 261978
rect 593286 261922 593342 261978
rect 592914 244294 592970 244350
rect 593038 244294 593094 244350
rect 593162 244294 593218 244350
rect 593286 244294 593342 244350
rect 592914 244170 592970 244226
rect 593038 244170 593094 244226
rect 593162 244170 593218 244226
rect 593286 244170 593342 244226
rect 592914 244046 592970 244102
rect 593038 244046 593094 244102
rect 593162 244046 593218 244102
rect 593286 244046 593342 244102
rect 592914 243922 592970 243978
rect 593038 243922 593094 243978
rect 593162 243922 593218 243978
rect 593286 243922 593342 243978
rect 592914 226294 592970 226350
rect 593038 226294 593094 226350
rect 593162 226294 593218 226350
rect 593286 226294 593342 226350
rect 592914 226170 592970 226226
rect 593038 226170 593094 226226
rect 593162 226170 593218 226226
rect 593286 226170 593342 226226
rect 592914 226046 592970 226102
rect 593038 226046 593094 226102
rect 593162 226046 593218 226102
rect 593286 226046 593342 226102
rect 592914 225922 592970 225978
rect 593038 225922 593094 225978
rect 593162 225922 593218 225978
rect 593286 225922 593342 225978
rect 592914 208294 592970 208350
rect 593038 208294 593094 208350
rect 593162 208294 593218 208350
rect 593286 208294 593342 208350
rect 592914 208170 592970 208226
rect 593038 208170 593094 208226
rect 593162 208170 593218 208226
rect 593286 208170 593342 208226
rect 592914 208046 592970 208102
rect 593038 208046 593094 208102
rect 593162 208046 593218 208102
rect 593286 208046 593342 208102
rect 592914 207922 592970 207978
rect 593038 207922 593094 207978
rect 593162 207922 593218 207978
rect 593286 207922 593342 207978
rect 592914 190294 592970 190350
rect 593038 190294 593094 190350
rect 593162 190294 593218 190350
rect 593286 190294 593342 190350
rect 592914 190170 592970 190226
rect 593038 190170 593094 190226
rect 593162 190170 593218 190226
rect 593286 190170 593342 190226
rect 592914 190046 592970 190102
rect 593038 190046 593094 190102
rect 593162 190046 593218 190102
rect 593286 190046 593342 190102
rect 592914 189922 592970 189978
rect 593038 189922 593094 189978
rect 593162 189922 593218 189978
rect 593286 189922 593342 189978
rect 592914 172294 592970 172350
rect 593038 172294 593094 172350
rect 593162 172294 593218 172350
rect 593286 172294 593342 172350
rect 592914 172170 592970 172226
rect 593038 172170 593094 172226
rect 593162 172170 593218 172226
rect 593286 172170 593342 172226
rect 592914 172046 592970 172102
rect 593038 172046 593094 172102
rect 593162 172046 593218 172102
rect 593286 172046 593342 172102
rect 592914 171922 592970 171978
rect 593038 171922 593094 171978
rect 593162 171922 593218 171978
rect 593286 171922 593342 171978
rect 589194 148294 589250 148350
rect 589318 148294 589374 148350
rect 589442 148294 589498 148350
rect 589566 148294 589622 148350
rect 589194 148170 589250 148226
rect 589318 148170 589374 148226
rect 589442 148170 589498 148226
rect 589566 148170 589622 148226
rect 589194 148046 589250 148102
rect 589318 148046 589374 148102
rect 589442 148046 589498 148102
rect 589566 148046 589622 148102
rect 589194 147922 589250 147978
rect 589318 147922 589374 147978
rect 589442 147922 589498 147978
rect 589566 147922 589622 147978
rect 589194 130294 589250 130350
rect 589318 130294 589374 130350
rect 589442 130294 589498 130350
rect 589566 130294 589622 130350
rect 589194 130170 589250 130226
rect 589318 130170 589374 130226
rect 589442 130170 589498 130226
rect 589566 130170 589622 130226
rect 589194 130046 589250 130102
rect 589318 130046 589374 130102
rect 589442 130046 589498 130102
rect 589566 130046 589622 130102
rect 589194 129922 589250 129978
rect 589318 129922 589374 129978
rect 589442 129922 589498 129978
rect 589566 129922 589622 129978
rect 589194 112294 589250 112350
rect 589318 112294 589374 112350
rect 589442 112294 589498 112350
rect 589566 112294 589622 112350
rect 589194 112170 589250 112226
rect 589318 112170 589374 112226
rect 589442 112170 589498 112226
rect 589566 112170 589622 112226
rect 589194 112046 589250 112102
rect 589318 112046 589374 112102
rect 589442 112046 589498 112102
rect 589566 112046 589622 112102
rect 589194 111922 589250 111978
rect 589318 111922 589374 111978
rect 589442 111922 589498 111978
rect 589566 111922 589622 111978
rect 589194 94294 589250 94350
rect 589318 94294 589374 94350
rect 589442 94294 589498 94350
rect 589566 94294 589622 94350
rect 589194 94170 589250 94226
rect 589318 94170 589374 94226
rect 589442 94170 589498 94226
rect 589566 94170 589622 94226
rect 589194 94046 589250 94102
rect 589318 94046 589374 94102
rect 589442 94046 589498 94102
rect 589566 94046 589622 94102
rect 589194 93922 589250 93978
rect 589318 93922 589374 93978
rect 589442 93922 589498 93978
rect 589566 93922 589622 93978
rect 589194 76294 589250 76350
rect 589318 76294 589374 76350
rect 589442 76294 589498 76350
rect 589566 76294 589622 76350
rect 589194 76170 589250 76226
rect 589318 76170 589374 76226
rect 589442 76170 589498 76226
rect 589566 76170 589622 76226
rect 589194 76046 589250 76102
rect 589318 76046 589374 76102
rect 589442 76046 589498 76102
rect 589566 76046 589622 76102
rect 589194 75922 589250 75978
rect 589318 75922 589374 75978
rect 589442 75922 589498 75978
rect 589566 75922 589622 75978
rect 589194 58294 589250 58350
rect 589318 58294 589374 58350
rect 589442 58294 589498 58350
rect 589566 58294 589622 58350
rect 589194 58170 589250 58226
rect 589318 58170 589374 58226
rect 589442 58170 589498 58226
rect 589566 58170 589622 58226
rect 589194 58046 589250 58102
rect 589318 58046 589374 58102
rect 589442 58046 589498 58102
rect 589566 58046 589622 58102
rect 589194 57922 589250 57978
rect 589318 57922 589374 57978
rect 589442 57922 589498 57978
rect 589566 57922 589622 57978
rect 589194 40294 589250 40350
rect 589318 40294 589374 40350
rect 589442 40294 589498 40350
rect 589566 40294 589622 40350
rect 589194 40170 589250 40226
rect 589318 40170 589374 40226
rect 589442 40170 589498 40226
rect 589566 40170 589622 40226
rect 589194 40046 589250 40102
rect 589318 40046 589374 40102
rect 589442 40046 589498 40102
rect 589566 40046 589622 40102
rect 589194 39922 589250 39978
rect 589318 39922 589374 39978
rect 589442 39922 589498 39978
rect 589566 39922 589622 39978
rect 592914 154294 592970 154350
rect 593038 154294 593094 154350
rect 593162 154294 593218 154350
rect 593286 154294 593342 154350
rect 592914 154170 592970 154226
rect 593038 154170 593094 154226
rect 593162 154170 593218 154226
rect 593286 154170 593342 154226
rect 592914 154046 592970 154102
rect 593038 154046 593094 154102
rect 593162 154046 593218 154102
rect 593286 154046 593342 154102
rect 592914 153922 592970 153978
rect 593038 153922 593094 153978
rect 593162 153922 593218 153978
rect 593286 153922 593342 153978
rect 592914 136294 592970 136350
rect 593038 136294 593094 136350
rect 593162 136294 593218 136350
rect 593286 136294 593342 136350
rect 592914 136170 592970 136226
rect 593038 136170 593094 136226
rect 593162 136170 593218 136226
rect 593286 136170 593342 136226
rect 592914 136046 592970 136102
rect 593038 136046 593094 136102
rect 593162 136046 593218 136102
rect 593286 136046 593342 136102
rect 592914 135922 592970 135978
rect 593038 135922 593094 135978
rect 593162 135922 593218 135978
rect 593286 135922 593342 135978
rect 592914 118294 592970 118350
rect 593038 118294 593094 118350
rect 593162 118294 593218 118350
rect 593286 118294 593342 118350
rect 592914 118170 592970 118226
rect 593038 118170 593094 118226
rect 593162 118170 593218 118226
rect 593286 118170 593342 118226
rect 592914 118046 592970 118102
rect 593038 118046 593094 118102
rect 593162 118046 593218 118102
rect 593286 118046 593342 118102
rect 592914 117922 592970 117978
rect 593038 117922 593094 117978
rect 593162 117922 593218 117978
rect 593286 117922 593342 117978
rect 592914 100294 592970 100350
rect 593038 100294 593094 100350
rect 593162 100294 593218 100350
rect 593286 100294 593342 100350
rect 592914 100170 592970 100226
rect 593038 100170 593094 100226
rect 593162 100170 593218 100226
rect 593286 100170 593342 100226
rect 592914 100046 592970 100102
rect 593038 100046 593094 100102
rect 593162 100046 593218 100102
rect 593286 100046 593342 100102
rect 592914 99922 592970 99978
rect 593038 99922 593094 99978
rect 593162 99922 593218 99978
rect 593286 99922 593342 99978
rect 592914 82294 592970 82350
rect 593038 82294 593094 82350
rect 593162 82294 593218 82350
rect 593286 82294 593342 82350
rect 592914 82170 592970 82226
rect 593038 82170 593094 82226
rect 593162 82170 593218 82226
rect 593286 82170 593342 82226
rect 592914 82046 592970 82102
rect 593038 82046 593094 82102
rect 593162 82046 593218 82102
rect 593286 82046 593342 82102
rect 592914 81922 592970 81978
rect 593038 81922 593094 81978
rect 593162 81922 593218 81978
rect 593286 81922 593342 81978
rect 592914 64294 592970 64350
rect 593038 64294 593094 64350
rect 593162 64294 593218 64350
rect 593286 64294 593342 64350
rect 592914 64170 592970 64226
rect 593038 64170 593094 64226
rect 593162 64170 593218 64226
rect 593286 64170 593342 64226
rect 592914 64046 592970 64102
rect 593038 64046 593094 64102
rect 593162 64046 593218 64102
rect 593286 64046 593342 64102
rect 592914 63922 592970 63978
rect 593038 63922 593094 63978
rect 593162 63922 593218 63978
rect 593286 63922 593342 63978
rect 589194 22294 589250 22350
rect 589318 22294 589374 22350
rect 589442 22294 589498 22350
rect 589566 22294 589622 22350
rect 589194 22170 589250 22226
rect 589318 22170 589374 22226
rect 589442 22170 589498 22226
rect 589566 22170 589622 22226
rect 589194 22046 589250 22102
rect 589318 22046 589374 22102
rect 589442 22046 589498 22102
rect 589566 22046 589622 22102
rect 589194 21922 589250 21978
rect 589318 21922 589374 21978
rect 589442 21922 589498 21978
rect 589566 21922 589622 21978
rect 562194 10294 562250 10350
rect 562318 10294 562374 10350
rect 562442 10294 562498 10350
rect 562566 10294 562622 10350
rect 562194 10170 562250 10226
rect 562318 10170 562374 10226
rect 562442 10170 562498 10226
rect 562566 10170 562622 10226
rect 562194 10046 562250 10102
rect 562318 10046 562374 10102
rect 562442 10046 562498 10102
rect 562566 10046 562622 10102
rect 562194 9922 562250 9978
rect 562318 9922 562374 9978
rect 562442 9922 562498 9978
rect 562566 9922 562622 9978
rect 592914 46294 592970 46350
rect 593038 46294 593094 46350
rect 593162 46294 593218 46350
rect 593286 46294 593342 46350
rect 592914 46170 592970 46226
rect 593038 46170 593094 46226
rect 593162 46170 593218 46226
rect 593286 46170 593342 46226
rect 592914 46046 592970 46102
rect 593038 46046 593094 46102
rect 593162 46046 593218 46102
rect 593286 46046 593342 46102
rect 592914 45922 592970 45978
rect 593038 45922 593094 45978
rect 593162 45922 593218 45978
rect 593286 45922 593342 45978
rect 592914 28294 592970 28350
rect 593038 28294 593094 28350
rect 593162 28294 593218 28350
rect 593286 28294 593342 28350
rect 592914 28170 592970 28226
rect 593038 28170 593094 28226
rect 593162 28170 593218 28226
rect 593286 28170 593342 28226
rect 592914 28046 592970 28102
rect 593038 28046 593094 28102
rect 593162 28046 593218 28102
rect 593286 28046 593342 28102
rect 592914 27922 592970 27978
rect 593038 27922 593094 27978
rect 593162 27922 593218 27978
rect 593286 27922 593342 27978
rect 589194 4294 589250 4350
rect 589318 4294 589374 4350
rect 589442 4294 589498 4350
rect 589566 4294 589622 4350
rect 589194 4170 589250 4226
rect 589318 4170 589374 4226
rect 589442 4170 589498 4226
rect 589566 4170 589622 4226
rect 589194 4046 589250 4102
rect 589318 4046 589374 4102
rect 589442 4046 589498 4102
rect 589566 4046 589622 4102
rect 589194 3922 589250 3978
rect 589318 3922 589374 3978
rect 589442 3922 589498 3978
rect 589566 3922 589622 3978
rect 565404 3302 565460 3358
rect 563500 3122 563556 3178
rect 571228 242 571284 298
rect 569212 62 569268 118
rect 562194 -1176 562250 -1120
rect 562318 -1176 562374 -1120
rect 562442 -1176 562498 -1120
rect 562566 -1176 562622 -1120
rect 562194 -1300 562250 -1244
rect 562318 -1300 562374 -1244
rect 562442 -1300 562498 -1244
rect 562566 -1300 562622 -1244
rect 562194 -1424 562250 -1368
rect 562318 -1424 562374 -1368
rect 562442 -1424 562498 -1368
rect 562566 -1424 562622 -1368
rect 562194 -1548 562250 -1492
rect 562318 -1548 562374 -1492
rect 562442 -1548 562498 -1492
rect 562566 -1548 562622 -1492
rect 589194 -216 589250 -160
rect 589318 -216 589374 -160
rect 589442 -216 589498 -160
rect 589566 -216 589622 -160
rect 589194 -340 589250 -284
rect 589318 -340 589374 -284
rect 589442 -340 589498 -284
rect 589566 -340 589622 -284
rect 589194 -464 589250 -408
rect 589318 -464 589374 -408
rect 589442 -464 589498 -408
rect 589566 -464 589622 -408
rect 589194 -588 589250 -532
rect 589318 -588 589374 -532
rect 589442 -588 589498 -532
rect 589566 -588 589622 -532
rect 592914 10294 592970 10350
rect 593038 10294 593094 10350
rect 593162 10294 593218 10350
rect 593286 10294 593342 10350
rect 592914 10170 592970 10226
rect 593038 10170 593094 10226
rect 593162 10170 593218 10226
rect 593286 10170 593342 10226
rect 592914 10046 592970 10102
rect 593038 10046 593094 10102
rect 593162 10046 593218 10102
rect 593286 10046 593342 10102
rect 592914 9922 592970 9978
rect 593038 9922 593094 9978
rect 593162 9922 593218 9978
rect 593286 9922 593342 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 592914 -1176 592970 -1120
rect 593038 -1176 593094 -1120
rect 593162 -1176 593218 -1120
rect 593286 -1176 593342 -1120
rect 592914 -1300 592970 -1244
rect 593038 -1300 593094 -1244
rect 593162 -1300 593218 -1244
rect 593286 -1300 593342 -1244
rect 592914 -1424 592970 -1368
rect 593038 -1424 593094 -1368
rect 593162 -1424 593218 -1368
rect 593286 -1424 593342 -1368
rect 592914 -1548 592970 -1492
rect 593038 -1548 593094 -1492
rect 593162 -1548 593218 -1492
rect 593286 -1548 593342 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 224274 568350
rect 224330 568294 224398 568350
rect 224454 568294 224522 568350
rect 224578 568294 224646 568350
rect 224702 568294 254994 568350
rect 255050 568294 255118 568350
rect 255174 568294 255242 568350
rect 255298 568294 255366 568350
rect 255422 568294 285714 568350
rect 285770 568294 285838 568350
rect 285894 568294 285962 568350
rect 286018 568294 286086 568350
rect 286142 568294 316434 568350
rect 316490 568294 316558 568350
rect 316614 568294 316682 568350
rect 316738 568294 316806 568350
rect 316862 568294 347154 568350
rect 347210 568294 347278 568350
rect 347334 568294 347402 568350
rect 347458 568294 347526 568350
rect 347582 568294 377874 568350
rect 377930 568294 377998 568350
rect 378054 568294 378122 568350
rect 378178 568294 378246 568350
rect 378302 568294 408594 568350
rect 408650 568294 408718 568350
rect 408774 568294 408842 568350
rect 408898 568294 408966 568350
rect 409022 568294 439314 568350
rect 439370 568294 439438 568350
rect 439494 568294 439562 568350
rect 439618 568294 439686 568350
rect 439742 568294 470034 568350
rect 470090 568294 470158 568350
rect 470214 568294 470282 568350
rect 470338 568294 470406 568350
rect 470462 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 224274 568226
rect 224330 568170 224398 568226
rect 224454 568170 224522 568226
rect 224578 568170 224646 568226
rect 224702 568170 254994 568226
rect 255050 568170 255118 568226
rect 255174 568170 255242 568226
rect 255298 568170 255366 568226
rect 255422 568170 285714 568226
rect 285770 568170 285838 568226
rect 285894 568170 285962 568226
rect 286018 568170 286086 568226
rect 286142 568170 316434 568226
rect 316490 568170 316558 568226
rect 316614 568170 316682 568226
rect 316738 568170 316806 568226
rect 316862 568170 347154 568226
rect 347210 568170 347278 568226
rect 347334 568170 347402 568226
rect 347458 568170 347526 568226
rect 347582 568170 377874 568226
rect 377930 568170 377998 568226
rect 378054 568170 378122 568226
rect 378178 568170 378246 568226
rect 378302 568170 408594 568226
rect 408650 568170 408718 568226
rect 408774 568170 408842 568226
rect 408898 568170 408966 568226
rect 409022 568170 439314 568226
rect 439370 568170 439438 568226
rect 439494 568170 439562 568226
rect 439618 568170 439686 568226
rect 439742 568170 470034 568226
rect 470090 568170 470158 568226
rect 470214 568170 470282 568226
rect 470338 568170 470406 568226
rect 470462 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 224274 568102
rect 224330 568046 224398 568102
rect 224454 568046 224522 568102
rect 224578 568046 224646 568102
rect 224702 568046 254994 568102
rect 255050 568046 255118 568102
rect 255174 568046 255242 568102
rect 255298 568046 255366 568102
rect 255422 568046 285714 568102
rect 285770 568046 285838 568102
rect 285894 568046 285962 568102
rect 286018 568046 286086 568102
rect 286142 568046 316434 568102
rect 316490 568046 316558 568102
rect 316614 568046 316682 568102
rect 316738 568046 316806 568102
rect 316862 568046 347154 568102
rect 347210 568046 347278 568102
rect 347334 568046 347402 568102
rect 347458 568046 347526 568102
rect 347582 568046 377874 568102
rect 377930 568046 377998 568102
rect 378054 568046 378122 568102
rect 378178 568046 378246 568102
rect 378302 568046 408594 568102
rect 408650 568046 408718 568102
rect 408774 568046 408842 568102
rect 408898 568046 408966 568102
rect 409022 568046 439314 568102
rect 439370 568046 439438 568102
rect 439494 568046 439562 568102
rect 439618 568046 439686 568102
rect 439742 568046 470034 568102
rect 470090 568046 470158 568102
rect 470214 568046 470282 568102
rect 470338 568046 470406 568102
rect 470462 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 224274 567978
rect 224330 567922 224398 567978
rect 224454 567922 224522 567978
rect 224578 567922 224646 567978
rect 224702 567922 254994 567978
rect 255050 567922 255118 567978
rect 255174 567922 255242 567978
rect 255298 567922 255366 567978
rect 255422 567922 285714 567978
rect 285770 567922 285838 567978
rect 285894 567922 285962 567978
rect 286018 567922 286086 567978
rect 286142 567922 316434 567978
rect 316490 567922 316558 567978
rect 316614 567922 316682 567978
rect 316738 567922 316806 567978
rect 316862 567922 347154 567978
rect 347210 567922 347278 567978
rect 347334 567922 347402 567978
rect 347458 567922 347526 567978
rect 347582 567922 377874 567978
rect 377930 567922 377998 567978
rect 378054 567922 378122 567978
rect 378178 567922 378246 567978
rect 378302 567922 408594 567978
rect 408650 567922 408718 567978
rect 408774 567922 408842 567978
rect 408898 567922 408966 567978
rect 409022 567922 439314 567978
rect 439370 567922 439438 567978
rect 439494 567922 439562 567978
rect 439618 567922 439686 567978
rect 439742 567922 470034 567978
rect 470090 567922 470158 567978
rect 470214 567922 470282 567978
rect 470338 567922 470406 567978
rect 470462 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 220554 562350
rect 220610 562294 220678 562350
rect 220734 562294 220802 562350
rect 220858 562294 220926 562350
rect 220982 562294 251274 562350
rect 251330 562294 251398 562350
rect 251454 562294 251522 562350
rect 251578 562294 251646 562350
rect 251702 562294 281994 562350
rect 282050 562294 282118 562350
rect 282174 562294 282242 562350
rect 282298 562294 282366 562350
rect 282422 562294 312714 562350
rect 312770 562294 312838 562350
rect 312894 562294 312962 562350
rect 313018 562294 313086 562350
rect 313142 562294 343434 562350
rect 343490 562294 343558 562350
rect 343614 562294 343682 562350
rect 343738 562294 343806 562350
rect 343862 562294 374154 562350
rect 374210 562294 374278 562350
rect 374334 562294 374402 562350
rect 374458 562294 374526 562350
rect 374582 562294 404874 562350
rect 404930 562294 404998 562350
rect 405054 562294 405122 562350
rect 405178 562294 405246 562350
rect 405302 562294 435594 562350
rect 435650 562294 435718 562350
rect 435774 562294 435842 562350
rect 435898 562294 435966 562350
rect 436022 562294 466314 562350
rect 466370 562294 466438 562350
rect 466494 562294 466562 562350
rect 466618 562294 466686 562350
rect 466742 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 220554 562226
rect 220610 562170 220678 562226
rect 220734 562170 220802 562226
rect 220858 562170 220926 562226
rect 220982 562170 251274 562226
rect 251330 562170 251398 562226
rect 251454 562170 251522 562226
rect 251578 562170 251646 562226
rect 251702 562170 281994 562226
rect 282050 562170 282118 562226
rect 282174 562170 282242 562226
rect 282298 562170 282366 562226
rect 282422 562170 312714 562226
rect 312770 562170 312838 562226
rect 312894 562170 312962 562226
rect 313018 562170 313086 562226
rect 313142 562170 343434 562226
rect 343490 562170 343558 562226
rect 343614 562170 343682 562226
rect 343738 562170 343806 562226
rect 343862 562170 374154 562226
rect 374210 562170 374278 562226
rect 374334 562170 374402 562226
rect 374458 562170 374526 562226
rect 374582 562170 404874 562226
rect 404930 562170 404998 562226
rect 405054 562170 405122 562226
rect 405178 562170 405246 562226
rect 405302 562170 435594 562226
rect 435650 562170 435718 562226
rect 435774 562170 435842 562226
rect 435898 562170 435966 562226
rect 436022 562170 466314 562226
rect 466370 562170 466438 562226
rect 466494 562170 466562 562226
rect 466618 562170 466686 562226
rect 466742 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 220554 562102
rect 220610 562046 220678 562102
rect 220734 562046 220802 562102
rect 220858 562046 220926 562102
rect 220982 562046 251274 562102
rect 251330 562046 251398 562102
rect 251454 562046 251522 562102
rect 251578 562046 251646 562102
rect 251702 562046 281994 562102
rect 282050 562046 282118 562102
rect 282174 562046 282242 562102
rect 282298 562046 282366 562102
rect 282422 562046 312714 562102
rect 312770 562046 312838 562102
rect 312894 562046 312962 562102
rect 313018 562046 313086 562102
rect 313142 562046 343434 562102
rect 343490 562046 343558 562102
rect 343614 562046 343682 562102
rect 343738 562046 343806 562102
rect 343862 562046 374154 562102
rect 374210 562046 374278 562102
rect 374334 562046 374402 562102
rect 374458 562046 374526 562102
rect 374582 562046 404874 562102
rect 404930 562046 404998 562102
rect 405054 562046 405122 562102
rect 405178 562046 405246 562102
rect 405302 562046 435594 562102
rect 435650 562046 435718 562102
rect 435774 562046 435842 562102
rect 435898 562046 435966 562102
rect 436022 562046 466314 562102
rect 466370 562046 466438 562102
rect 466494 562046 466562 562102
rect 466618 562046 466686 562102
rect 466742 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 128394 561978
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 220554 561978
rect 220610 561922 220678 561978
rect 220734 561922 220802 561978
rect 220858 561922 220926 561978
rect 220982 561922 251274 561978
rect 251330 561922 251398 561978
rect 251454 561922 251522 561978
rect 251578 561922 251646 561978
rect 251702 561922 281994 561978
rect 282050 561922 282118 561978
rect 282174 561922 282242 561978
rect 282298 561922 282366 561978
rect 282422 561922 312714 561978
rect 312770 561922 312838 561978
rect 312894 561922 312962 561978
rect 313018 561922 313086 561978
rect 313142 561922 343434 561978
rect 343490 561922 343558 561978
rect 343614 561922 343682 561978
rect 343738 561922 343806 561978
rect 343862 561922 374154 561978
rect 374210 561922 374278 561978
rect 374334 561922 374402 561978
rect 374458 561922 374526 561978
rect 374582 561922 404874 561978
rect 404930 561922 404998 561978
rect 405054 561922 405122 561978
rect 405178 561922 405246 561978
rect 405302 561922 435594 561978
rect 435650 561922 435718 561978
rect 435774 561922 435842 561978
rect 435898 561922 435966 561978
rect 436022 561922 466314 561978
rect 466370 561922 466438 561978
rect 466494 561922 466562 561978
rect 466618 561922 466686 561978
rect 466742 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 224274 550350
rect 224330 550294 224398 550350
rect 224454 550294 224522 550350
rect 224578 550294 224646 550350
rect 224702 550294 254994 550350
rect 255050 550294 255118 550350
rect 255174 550294 255242 550350
rect 255298 550294 255366 550350
rect 255422 550294 285714 550350
rect 285770 550294 285838 550350
rect 285894 550294 285962 550350
rect 286018 550294 286086 550350
rect 286142 550294 316434 550350
rect 316490 550294 316558 550350
rect 316614 550294 316682 550350
rect 316738 550294 316806 550350
rect 316862 550294 347154 550350
rect 347210 550294 347278 550350
rect 347334 550294 347402 550350
rect 347458 550294 347526 550350
rect 347582 550294 377874 550350
rect 377930 550294 377998 550350
rect 378054 550294 378122 550350
rect 378178 550294 378246 550350
rect 378302 550294 408594 550350
rect 408650 550294 408718 550350
rect 408774 550294 408842 550350
rect 408898 550294 408966 550350
rect 409022 550294 439314 550350
rect 439370 550294 439438 550350
rect 439494 550294 439562 550350
rect 439618 550294 439686 550350
rect 439742 550294 470034 550350
rect 470090 550294 470158 550350
rect 470214 550294 470282 550350
rect 470338 550294 470406 550350
rect 470462 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 224274 550226
rect 224330 550170 224398 550226
rect 224454 550170 224522 550226
rect 224578 550170 224646 550226
rect 224702 550170 254994 550226
rect 255050 550170 255118 550226
rect 255174 550170 255242 550226
rect 255298 550170 255366 550226
rect 255422 550170 285714 550226
rect 285770 550170 285838 550226
rect 285894 550170 285962 550226
rect 286018 550170 286086 550226
rect 286142 550170 316434 550226
rect 316490 550170 316558 550226
rect 316614 550170 316682 550226
rect 316738 550170 316806 550226
rect 316862 550170 347154 550226
rect 347210 550170 347278 550226
rect 347334 550170 347402 550226
rect 347458 550170 347526 550226
rect 347582 550170 377874 550226
rect 377930 550170 377998 550226
rect 378054 550170 378122 550226
rect 378178 550170 378246 550226
rect 378302 550170 408594 550226
rect 408650 550170 408718 550226
rect 408774 550170 408842 550226
rect 408898 550170 408966 550226
rect 409022 550170 439314 550226
rect 439370 550170 439438 550226
rect 439494 550170 439562 550226
rect 439618 550170 439686 550226
rect 439742 550170 470034 550226
rect 470090 550170 470158 550226
rect 470214 550170 470282 550226
rect 470338 550170 470406 550226
rect 470462 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 224274 550102
rect 224330 550046 224398 550102
rect 224454 550046 224522 550102
rect 224578 550046 224646 550102
rect 224702 550046 254994 550102
rect 255050 550046 255118 550102
rect 255174 550046 255242 550102
rect 255298 550046 255366 550102
rect 255422 550046 285714 550102
rect 285770 550046 285838 550102
rect 285894 550046 285962 550102
rect 286018 550046 286086 550102
rect 286142 550046 316434 550102
rect 316490 550046 316558 550102
rect 316614 550046 316682 550102
rect 316738 550046 316806 550102
rect 316862 550046 347154 550102
rect 347210 550046 347278 550102
rect 347334 550046 347402 550102
rect 347458 550046 347526 550102
rect 347582 550046 377874 550102
rect 377930 550046 377998 550102
rect 378054 550046 378122 550102
rect 378178 550046 378246 550102
rect 378302 550046 408594 550102
rect 408650 550046 408718 550102
rect 408774 550046 408842 550102
rect 408898 550046 408966 550102
rect 409022 550046 439314 550102
rect 439370 550046 439438 550102
rect 439494 550046 439562 550102
rect 439618 550046 439686 550102
rect 439742 550046 470034 550102
rect 470090 550046 470158 550102
rect 470214 550046 470282 550102
rect 470338 550046 470406 550102
rect 470462 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 224274 549978
rect 224330 549922 224398 549978
rect 224454 549922 224522 549978
rect 224578 549922 224646 549978
rect 224702 549922 254994 549978
rect 255050 549922 255118 549978
rect 255174 549922 255242 549978
rect 255298 549922 255366 549978
rect 255422 549922 285714 549978
rect 285770 549922 285838 549978
rect 285894 549922 285962 549978
rect 286018 549922 286086 549978
rect 286142 549922 316434 549978
rect 316490 549922 316558 549978
rect 316614 549922 316682 549978
rect 316738 549922 316806 549978
rect 316862 549922 347154 549978
rect 347210 549922 347278 549978
rect 347334 549922 347402 549978
rect 347458 549922 347526 549978
rect 347582 549922 377874 549978
rect 377930 549922 377998 549978
rect 378054 549922 378122 549978
rect 378178 549922 378246 549978
rect 378302 549922 408594 549978
rect 408650 549922 408718 549978
rect 408774 549922 408842 549978
rect 408898 549922 408966 549978
rect 409022 549922 439314 549978
rect 439370 549922 439438 549978
rect 439494 549922 439562 549978
rect 439618 549922 439686 549978
rect 439742 549922 470034 549978
rect 470090 549922 470158 549978
rect 470214 549922 470282 549978
rect 470338 549922 470406 549978
rect 470462 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 97674 544350
rect 97730 544294 97798 544350
rect 97854 544294 97922 544350
rect 97978 544294 98046 544350
rect 98102 544294 128394 544350
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 220554 544350
rect 220610 544294 220678 544350
rect 220734 544294 220802 544350
rect 220858 544294 220926 544350
rect 220982 544294 251274 544350
rect 251330 544294 251398 544350
rect 251454 544294 251522 544350
rect 251578 544294 251646 544350
rect 251702 544294 281994 544350
rect 282050 544294 282118 544350
rect 282174 544294 282242 544350
rect 282298 544294 282366 544350
rect 282422 544294 312714 544350
rect 312770 544294 312838 544350
rect 312894 544294 312962 544350
rect 313018 544294 313086 544350
rect 313142 544294 343434 544350
rect 343490 544294 343558 544350
rect 343614 544294 343682 544350
rect 343738 544294 343806 544350
rect 343862 544294 374154 544350
rect 374210 544294 374278 544350
rect 374334 544294 374402 544350
rect 374458 544294 374526 544350
rect 374582 544294 404874 544350
rect 404930 544294 404998 544350
rect 405054 544294 405122 544350
rect 405178 544294 405246 544350
rect 405302 544294 435594 544350
rect 435650 544294 435718 544350
rect 435774 544294 435842 544350
rect 435898 544294 435966 544350
rect 436022 544294 466314 544350
rect 466370 544294 466438 544350
rect 466494 544294 466562 544350
rect 466618 544294 466686 544350
rect 466742 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 97674 544226
rect 97730 544170 97798 544226
rect 97854 544170 97922 544226
rect 97978 544170 98046 544226
rect 98102 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 220554 544226
rect 220610 544170 220678 544226
rect 220734 544170 220802 544226
rect 220858 544170 220926 544226
rect 220982 544170 251274 544226
rect 251330 544170 251398 544226
rect 251454 544170 251522 544226
rect 251578 544170 251646 544226
rect 251702 544170 281994 544226
rect 282050 544170 282118 544226
rect 282174 544170 282242 544226
rect 282298 544170 282366 544226
rect 282422 544170 312714 544226
rect 312770 544170 312838 544226
rect 312894 544170 312962 544226
rect 313018 544170 313086 544226
rect 313142 544170 343434 544226
rect 343490 544170 343558 544226
rect 343614 544170 343682 544226
rect 343738 544170 343806 544226
rect 343862 544170 374154 544226
rect 374210 544170 374278 544226
rect 374334 544170 374402 544226
rect 374458 544170 374526 544226
rect 374582 544170 404874 544226
rect 404930 544170 404998 544226
rect 405054 544170 405122 544226
rect 405178 544170 405246 544226
rect 405302 544170 435594 544226
rect 435650 544170 435718 544226
rect 435774 544170 435842 544226
rect 435898 544170 435966 544226
rect 436022 544170 466314 544226
rect 466370 544170 466438 544226
rect 466494 544170 466562 544226
rect 466618 544170 466686 544226
rect 466742 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 97674 544102
rect 97730 544046 97798 544102
rect 97854 544046 97922 544102
rect 97978 544046 98046 544102
rect 98102 544046 128394 544102
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 220554 544102
rect 220610 544046 220678 544102
rect 220734 544046 220802 544102
rect 220858 544046 220926 544102
rect 220982 544046 251274 544102
rect 251330 544046 251398 544102
rect 251454 544046 251522 544102
rect 251578 544046 251646 544102
rect 251702 544046 281994 544102
rect 282050 544046 282118 544102
rect 282174 544046 282242 544102
rect 282298 544046 282366 544102
rect 282422 544046 312714 544102
rect 312770 544046 312838 544102
rect 312894 544046 312962 544102
rect 313018 544046 313086 544102
rect 313142 544046 343434 544102
rect 343490 544046 343558 544102
rect 343614 544046 343682 544102
rect 343738 544046 343806 544102
rect 343862 544046 374154 544102
rect 374210 544046 374278 544102
rect 374334 544046 374402 544102
rect 374458 544046 374526 544102
rect 374582 544046 404874 544102
rect 404930 544046 404998 544102
rect 405054 544046 405122 544102
rect 405178 544046 405246 544102
rect 405302 544046 435594 544102
rect 435650 544046 435718 544102
rect 435774 544046 435842 544102
rect 435898 544046 435966 544102
rect 436022 544046 466314 544102
rect 466370 544046 466438 544102
rect 466494 544046 466562 544102
rect 466618 544046 466686 544102
rect 466742 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 97674 543978
rect 97730 543922 97798 543978
rect 97854 543922 97922 543978
rect 97978 543922 98046 543978
rect 98102 543922 128394 543978
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 220554 543978
rect 220610 543922 220678 543978
rect 220734 543922 220802 543978
rect 220858 543922 220926 543978
rect 220982 543922 251274 543978
rect 251330 543922 251398 543978
rect 251454 543922 251522 543978
rect 251578 543922 251646 543978
rect 251702 543922 281994 543978
rect 282050 543922 282118 543978
rect 282174 543922 282242 543978
rect 282298 543922 282366 543978
rect 282422 543922 312714 543978
rect 312770 543922 312838 543978
rect 312894 543922 312962 543978
rect 313018 543922 313086 543978
rect 313142 543922 343434 543978
rect 343490 543922 343558 543978
rect 343614 543922 343682 543978
rect 343738 543922 343806 543978
rect 343862 543922 374154 543978
rect 374210 543922 374278 543978
rect 374334 543922 374402 543978
rect 374458 543922 374526 543978
rect 374582 543922 404874 543978
rect 404930 543922 404998 543978
rect 405054 543922 405122 543978
rect 405178 543922 405246 543978
rect 405302 543922 435594 543978
rect 435650 543922 435718 543978
rect 435774 543922 435842 543978
rect 435898 543922 435966 543978
rect 436022 543922 466314 543978
rect 466370 543922 466438 543978
rect 466494 543922 466562 543978
rect 466618 543922 466686 543978
rect 466742 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532294 70674 532350
rect 70730 532294 70798 532350
rect 70854 532294 70922 532350
rect 70978 532294 71046 532350
rect 71102 532294 101394 532350
rect 101450 532294 101518 532350
rect 101574 532294 101642 532350
rect 101698 532294 101766 532350
rect 101822 532294 132114 532350
rect 132170 532294 132238 532350
rect 132294 532294 132362 532350
rect 132418 532294 132486 532350
rect 132542 532294 162834 532350
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 193554 532350
rect 193610 532294 193678 532350
rect 193734 532294 193802 532350
rect 193858 532294 193926 532350
rect 193982 532294 224274 532350
rect 224330 532294 224398 532350
rect 224454 532294 224522 532350
rect 224578 532294 224646 532350
rect 224702 532294 254994 532350
rect 255050 532294 255118 532350
rect 255174 532294 255242 532350
rect 255298 532294 255366 532350
rect 255422 532294 285714 532350
rect 285770 532294 285838 532350
rect 285894 532294 285962 532350
rect 286018 532294 286086 532350
rect 286142 532294 316434 532350
rect 316490 532294 316558 532350
rect 316614 532294 316682 532350
rect 316738 532294 316806 532350
rect 316862 532294 347154 532350
rect 347210 532294 347278 532350
rect 347334 532294 347402 532350
rect 347458 532294 347526 532350
rect 347582 532294 377874 532350
rect 377930 532294 377998 532350
rect 378054 532294 378122 532350
rect 378178 532294 378246 532350
rect 378302 532294 408594 532350
rect 408650 532294 408718 532350
rect 408774 532294 408842 532350
rect 408898 532294 408966 532350
rect 409022 532294 439314 532350
rect 439370 532294 439438 532350
rect 439494 532294 439562 532350
rect 439618 532294 439686 532350
rect 439742 532294 470034 532350
rect 470090 532294 470158 532350
rect 470214 532294 470282 532350
rect 470338 532294 470406 532350
rect 470462 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 70674 532226
rect 70730 532170 70798 532226
rect 70854 532170 70922 532226
rect 70978 532170 71046 532226
rect 71102 532170 101394 532226
rect 101450 532170 101518 532226
rect 101574 532170 101642 532226
rect 101698 532170 101766 532226
rect 101822 532170 132114 532226
rect 132170 532170 132238 532226
rect 132294 532170 132362 532226
rect 132418 532170 132486 532226
rect 132542 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 193554 532226
rect 193610 532170 193678 532226
rect 193734 532170 193802 532226
rect 193858 532170 193926 532226
rect 193982 532170 224274 532226
rect 224330 532170 224398 532226
rect 224454 532170 224522 532226
rect 224578 532170 224646 532226
rect 224702 532170 254994 532226
rect 255050 532170 255118 532226
rect 255174 532170 255242 532226
rect 255298 532170 255366 532226
rect 255422 532170 285714 532226
rect 285770 532170 285838 532226
rect 285894 532170 285962 532226
rect 286018 532170 286086 532226
rect 286142 532170 316434 532226
rect 316490 532170 316558 532226
rect 316614 532170 316682 532226
rect 316738 532170 316806 532226
rect 316862 532170 347154 532226
rect 347210 532170 347278 532226
rect 347334 532170 347402 532226
rect 347458 532170 347526 532226
rect 347582 532170 377874 532226
rect 377930 532170 377998 532226
rect 378054 532170 378122 532226
rect 378178 532170 378246 532226
rect 378302 532170 408594 532226
rect 408650 532170 408718 532226
rect 408774 532170 408842 532226
rect 408898 532170 408966 532226
rect 409022 532170 439314 532226
rect 439370 532170 439438 532226
rect 439494 532170 439562 532226
rect 439618 532170 439686 532226
rect 439742 532170 470034 532226
rect 470090 532170 470158 532226
rect 470214 532170 470282 532226
rect 470338 532170 470406 532226
rect 470462 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 70674 532102
rect 70730 532046 70798 532102
rect 70854 532046 70922 532102
rect 70978 532046 71046 532102
rect 71102 532046 101394 532102
rect 101450 532046 101518 532102
rect 101574 532046 101642 532102
rect 101698 532046 101766 532102
rect 101822 532046 132114 532102
rect 132170 532046 132238 532102
rect 132294 532046 132362 532102
rect 132418 532046 132486 532102
rect 132542 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 193554 532102
rect 193610 532046 193678 532102
rect 193734 532046 193802 532102
rect 193858 532046 193926 532102
rect 193982 532046 224274 532102
rect 224330 532046 224398 532102
rect 224454 532046 224522 532102
rect 224578 532046 224646 532102
rect 224702 532046 254994 532102
rect 255050 532046 255118 532102
rect 255174 532046 255242 532102
rect 255298 532046 255366 532102
rect 255422 532046 285714 532102
rect 285770 532046 285838 532102
rect 285894 532046 285962 532102
rect 286018 532046 286086 532102
rect 286142 532046 316434 532102
rect 316490 532046 316558 532102
rect 316614 532046 316682 532102
rect 316738 532046 316806 532102
rect 316862 532046 347154 532102
rect 347210 532046 347278 532102
rect 347334 532046 347402 532102
rect 347458 532046 347526 532102
rect 347582 532046 377874 532102
rect 377930 532046 377998 532102
rect 378054 532046 378122 532102
rect 378178 532046 378246 532102
rect 378302 532046 408594 532102
rect 408650 532046 408718 532102
rect 408774 532046 408842 532102
rect 408898 532046 408966 532102
rect 409022 532046 439314 532102
rect 439370 532046 439438 532102
rect 439494 532046 439562 532102
rect 439618 532046 439686 532102
rect 439742 532046 470034 532102
rect 470090 532046 470158 532102
rect 470214 532046 470282 532102
rect 470338 532046 470406 532102
rect 470462 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531922 70674 531978
rect 70730 531922 70798 531978
rect 70854 531922 70922 531978
rect 70978 531922 71046 531978
rect 71102 531922 101394 531978
rect 101450 531922 101518 531978
rect 101574 531922 101642 531978
rect 101698 531922 101766 531978
rect 101822 531922 132114 531978
rect 132170 531922 132238 531978
rect 132294 531922 132362 531978
rect 132418 531922 132486 531978
rect 132542 531922 162834 531978
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 193554 531978
rect 193610 531922 193678 531978
rect 193734 531922 193802 531978
rect 193858 531922 193926 531978
rect 193982 531922 224274 531978
rect 224330 531922 224398 531978
rect 224454 531922 224522 531978
rect 224578 531922 224646 531978
rect 224702 531922 254994 531978
rect 255050 531922 255118 531978
rect 255174 531922 255242 531978
rect 255298 531922 255366 531978
rect 255422 531922 285714 531978
rect 285770 531922 285838 531978
rect 285894 531922 285962 531978
rect 286018 531922 286086 531978
rect 286142 531922 316434 531978
rect 316490 531922 316558 531978
rect 316614 531922 316682 531978
rect 316738 531922 316806 531978
rect 316862 531922 347154 531978
rect 347210 531922 347278 531978
rect 347334 531922 347402 531978
rect 347458 531922 347526 531978
rect 347582 531922 377874 531978
rect 377930 531922 377998 531978
rect 378054 531922 378122 531978
rect 378178 531922 378246 531978
rect 378302 531922 408594 531978
rect 408650 531922 408718 531978
rect 408774 531922 408842 531978
rect 408898 531922 408966 531978
rect 409022 531922 439314 531978
rect 439370 531922 439438 531978
rect 439494 531922 439562 531978
rect 439618 531922 439686 531978
rect 439742 531922 470034 531978
rect 470090 531922 470158 531978
rect 470214 531922 470282 531978
rect 470338 531922 470406 531978
rect 470462 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 66954 526350
rect 67010 526294 67078 526350
rect 67134 526294 67202 526350
rect 67258 526294 67326 526350
rect 67382 526294 97674 526350
rect 97730 526294 97798 526350
rect 97854 526294 97922 526350
rect 97978 526294 98046 526350
rect 98102 526294 128394 526350
rect 128450 526294 128518 526350
rect 128574 526294 128642 526350
rect 128698 526294 128766 526350
rect 128822 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 220554 526350
rect 220610 526294 220678 526350
rect 220734 526294 220802 526350
rect 220858 526294 220926 526350
rect 220982 526294 251274 526350
rect 251330 526294 251398 526350
rect 251454 526294 251522 526350
rect 251578 526294 251646 526350
rect 251702 526294 281994 526350
rect 282050 526294 282118 526350
rect 282174 526294 282242 526350
rect 282298 526294 282366 526350
rect 282422 526294 312714 526350
rect 312770 526294 312838 526350
rect 312894 526294 312962 526350
rect 313018 526294 313086 526350
rect 313142 526294 343434 526350
rect 343490 526294 343558 526350
rect 343614 526294 343682 526350
rect 343738 526294 343806 526350
rect 343862 526294 374154 526350
rect 374210 526294 374278 526350
rect 374334 526294 374402 526350
rect 374458 526294 374526 526350
rect 374582 526294 404874 526350
rect 404930 526294 404998 526350
rect 405054 526294 405122 526350
rect 405178 526294 405246 526350
rect 405302 526294 435594 526350
rect 435650 526294 435718 526350
rect 435774 526294 435842 526350
rect 435898 526294 435966 526350
rect 436022 526294 466314 526350
rect 466370 526294 466438 526350
rect 466494 526294 466562 526350
rect 466618 526294 466686 526350
rect 466742 526294 497034 526350
rect 497090 526294 497158 526350
rect 497214 526294 497282 526350
rect 497338 526294 497406 526350
rect 497462 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 66954 526226
rect 67010 526170 67078 526226
rect 67134 526170 67202 526226
rect 67258 526170 67326 526226
rect 67382 526170 97674 526226
rect 97730 526170 97798 526226
rect 97854 526170 97922 526226
rect 97978 526170 98046 526226
rect 98102 526170 128394 526226
rect 128450 526170 128518 526226
rect 128574 526170 128642 526226
rect 128698 526170 128766 526226
rect 128822 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 220554 526226
rect 220610 526170 220678 526226
rect 220734 526170 220802 526226
rect 220858 526170 220926 526226
rect 220982 526170 251274 526226
rect 251330 526170 251398 526226
rect 251454 526170 251522 526226
rect 251578 526170 251646 526226
rect 251702 526170 281994 526226
rect 282050 526170 282118 526226
rect 282174 526170 282242 526226
rect 282298 526170 282366 526226
rect 282422 526170 312714 526226
rect 312770 526170 312838 526226
rect 312894 526170 312962 526226
rect 313018 526170 313086 526226
rect 313142 526170 343434 526226
rect 343490 526170 343558 526226
rect 343614 526170 343682 526226
rect 343738 526170 343806 526226
rect 343862 526170 374154 526226
rect 374210 526170 374278 526226
rect 374334 526170 374402 526226
rect 374458 526170 374526 526226
rect 374582 526170 404874 526226
rect 404930 526170 404998 526226
rect 405054 526170 405122 526226
rect 405178 526170 405246 526226
rect 405302 526170 435594 526226
rect 435650 526170 435718 526226
rect 435774 526170 435842 526226
rect 435898 526170 435966 526226
rect 436022 526170 466314 526226
rect 466370 526170 466438 526226
rect 466494 526170 466562 526226
rect 466618 526170 466686 526226
rect 466742 526170 497034 526226
rect 497090 526170 497158 526226
rect 497214 526170 497282 526226
rect 497338 526170 497406 526226
rect 497462 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 66954 526102
rect 67010 526046 67078 526102
rect 67134 526046 67202 526102
rect 67258 526046 67326 526102
rect 67382 526046 97674 526102
rect 97730 526046 97798 526102
rect 97854 526046 97922 526102
rect 97978 526046 98046 526102
rect 98102 526046 128394 526102
rect 128450 526046 128518 526102
rect 128574 526046 128642 526102
rect 128698 526046 128766 526102
rect 128822 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 220554 526102
rect 220610 526046 220678 526102
rect 220734 526046 220802 526102
rect 220858 526046 220926 526102
rect 220982 526046 251274 526102
rect 251330 526046 251398 526102
rect 251454 526046 251522 526102
rect 251578 526046 251646 526102
rect 251702 526046 281994 526102
rect 282050 526046 282118 526102
rect 282174 526046 282242 526102
rect 282298 526046 282366 526102
rect 282422 526046 312714 526102
rect 312770 526046 312838 526102
rect 312894 526046 312962 526102
rect 313018 526046 313086 526102
rect 313142 526046 343434 526102
rect 343490 526046 343558 526102
rect 343614 526046 343682 526102
rect 343738 526046 343806 526102
rect 343862 526046 374154 526102
rect 374210 526046 374278 526102
rect 374334 526046 374402 526102
rect 374458 526046 374526 526102
rect 374582 526046 404874 526102
rect 404930 526046 404998 526102
rect 405054 526046 405122 526102
rect 405178 526046 405246 526102
rect 405302 526046 435594 526102
rect 435650 526046 435718 526102
rect 435774 526046 435842 526102
rect 435898 526046 435966 526102
rect 436022 526046 466314 526102
rect 466370 526046 466438 526102
rect 466494 526046 466562 526102
rect 466618 526046 466686 526102
rect 466742 526046 497034 526102
rect 497090 526046 497158 526102
rect 497214 526046 497282 526102
rect 497338 526046 497406 526102
rect 497462 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 66954 525978
rect 67010 525922 67078 525978
rect 67134 525922 67202 525978
rect 67258 525922 67326 525978
rect 67382 525922 97674 525978
rect 97730 525922 97798 525978
rect 97854 525922 97922 525978
rect 97978 525922 98046 525978
rect 98102 525922 128394 525978
rect 128450 525922 128518 525978
rect 128574 525922 128642 525978
rect 128698 525922 128766 525978
rect 128822 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 220554 525978
rect 220610 525922 220678 525978
rect 220734 525922 220802 525978
rect 220858 525922 220926 525978
rect 220982 525922 251274 525978
rect 251330 525922 251398 525978
rect 251454 525922 251522 525978
rect 251578 525922 251646 525978
rect 251702 525922 281994 525978
rect 282050 525922 282118 525978
rect 282174 525922 282242 525978
rect 282298 525922 282366 525978
rect 282422 525922 312714 525978
rect 312770 525922 312838 525978
rect 312894 525922 312962 525978
rect 313018 525922 313086 525978
rect 313142 525922 343434 525978
rect 343490 525922 343558 525978
rect 343614 525922 343682 525978
rect 343738 525922 343806 525978
rect 343862 525922 374154 525978
rect 374210 525922 374278 525978
rect 374334 525922 374402 525978
rect 374458 525922 374526 525978
rect 374582 525922 404874 525978
rect 404930 525922 404998 525978
rect 405054 525922 405122 525978
rect 405178 525922 405246 525978
rect 405302 525922 435594 525978
rect 435650 525922 435718 525978
rect 435774 525922 435842 525978
rect 435898 525922 435966 525978
rect 436022 525922 466314 525978
rect 466370 525922 466438 525978
rect 466494 525922 466562 525978
rect 466618 525922 466686 525978
rect 466742 525922 497034 525978
rect 497090 525922 497158 525978
rect 497214 525922 497282 525978
rect 497338 525922 497406 525978
rect 497462 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 70674 514350
rect 70730 514294 70798 514350
rect 70854 514294 70922 514350
rect 70978 514294 71046 514350
rect 71102 514294 101394 514350
rect 101450 514294 101518 514350
rect 101574 514294 101642 514350
rect 101698 514294 101766 514350
rect 101822 514294 132114 514350
rect 132170 514294 132238 514350
rect 132294 514294 132362 514350
rect 132418 514294 132486 514350
rect 132542 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 193554 514350
rect 193610 514294 193678 514350
rect 193734 514294 193802 514350
rect 193858 514294 193926 514350
rect 193982 514294 224274 514350
rect 224330 514294 224398 514350
rect 224454 514294 224522 514350
rect 224578 514294 224646 514350
rect 224702 514294 254994 514350
rect 255050 514294 255118 514350
rect 255174 514294 255242 514350
rect 255298 514294 255366 514350
rect 255422 514294 285714 514350
rect 285770 514294 285838 514350
rect 285894 514294 285962 514350
rect 286018 514294 286086 514350
rect 286142 514294 316434 514350
rect 316490 514294 316558 514350
rect 316614 514294 316682 514350
rect 316738 514294 316806 514350
rect 316862 514294 347154 514350
rect 347210 514294 347278 514350
rect 347334 514294 347402 514350
rect 347458 514294 347526 514350
rect 347582 514294 377874 514350
rect 377930 514294 377998 514350
rect 378054 514294 378122 514350
rect 378178 514294 378246 514350
rect 378302 514294 408594 514350
rect 408650 514294 408718 514350
rect 408774 514294 408842 514350
rect 408898 514294 408966 514350
rect 409022 514294 439314 514350
rect 439370 514294 439438 514350
rect 439494 514294 439562 514350
rect 439618 514294 439686 514350
rect 439742 514294 470034 514350
rect 470090 514294 470158 514350
rect 470214 514294 470282 514350
rect 470338 514294 470406 514350
rect 470462 514294 500754 514350
rect 500810 514294 500878 514350
rect 500934 514294 501002 514350
rect 501058 514294 501126 514350
rect 501182 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 70674 514226
rect 70730 514170 70798 514226
rect 70854 514170 70922 514226
rect 70978 514170 71046 514226
rect 71102 514170 101394 514226
rect 101450 514170 101518 514226
rect 101574 514170 101642 514226
rect 101698 514170 101766 514226
rect 101822 514170 132114 514226
rect 132170 514170 132238 514226
rect 132294 514170 132362 514226
rect 132418 514170 132486 514226
rect 132542 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 193554 514226
rect 193610 514170 193678 514226
rect 193734 514170 193802 514226
rect 193858 514170 193926 514226
rect 193982 514170 224274 514226
rect 224330 514170 224398 514226
rect 224454 514170 224522 514226
rect 224578 514170 224646 514226
rect 224702 514170 254994 514226
rect 255050 514170 255118 514226
rect 255174 514170 255242 514226
rect 255298 514170 255366 514226
rect 255422 514170 285714 514226
rect 285770 514170 285838 514226
rect 285894 514170 285962 514226
rect 286018 514170 286086 514226
rect 286142 514170 316434 514226
rect 316490 514170 316558 514226
rect 316614 514170 316682 514226
rect 316738 514170 316806 514226
rect 316862 514170 347154 514226
rect 347210 514170 347278 514226
rect 347334 514170 347402 514226
rect 347458 514170 347526 514226
rect 347582 514170 377874 514226
rect 377930 514170 377998 514226
rect 378054 514170 378122 514226
rect 378178 514170 378246 514226
rect 378302 514170 408594 514226
rect 408650 514170 408718 514226
rect 408774 514170 408842 514226
rect 408898 514170 408966 514226
rect 409022 514170 439314 514226
rect 439370 514170 439438 514226
rect 439494 514170 439562 514226
rect 439618 514170 439686 514226
rect 439742 514170 470034 514226
rect 470090 514170 470158 514226
rect 470214 514170 470282 514226
rect 470338 514170 470406 514226
rect 470462 514170 500754 514226
rect 500810 514170 500878 514226
rect 500934 514170 501002 514226
rect 501058 514170 501126 514226
rect 501182 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 70674 514102
rect 70730 514046 70798 514102
rect 70854 514046 70922 514102
rect 70978 514046 71046 514102
rect 71102 514046 101394 514102
rect 101450 514046 101518 514102
rect 101574 514046 101642 514102
rect 101698 514046 101766 514102
rect 101822 514046 132114 514102
rect 132170 514046 132238 514102
rect 132294 514046 132362 514102
rect 132418 514046 132486 514102
rect 132542 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 193554 514102
rect 193610 514046 193678 514102
rect 193734 514046 193802 514102
rect 193858 514046 193926 514102
rect 193982 514046 224274 514102
rect 224330 514046 224398 514102
rect 224454 514046 224522 514102
rect 224578 514046 224646 514102
rect 224702 514046 254994 514102
rect 255050 514046 255118 514102
rect 255174 514046 255242 514102
rect 255298 514046 255366 514102
rect 255422 514046 285714 514102
rect 285770 514046 285838 514102
rect 285894 514046 285962 514102
rect 286018 514046 286086 514102
rect 286142 514046 316434 514102
rect 316490 514046 316558 514102
rect 316614 514046 316682 514102
rect 316738 514046 316806 514102
rect 316862 514046 347154 514102
rect 347210 514046 347278 514102
rect 347334 514046 347402 514102
rect 347458 514046 347526 514102
rect 347582 514046 377874 514102
rect 377930 514046 377998 514102
rect 378054 514046 378122 514102
rect 378178 514046 378246 514102
rect 378302 514046 408594 514102
rect 408650 514046 408718 514102
rect 408774 514046 408842 514102
rect 408898 514046 408966 514102
rect 409022 514046 439314 514102
rect 439370 514046 439438 514102
rect 439494 514046 439562 514102
rect 439618 514046 439686 514102
rect 439742 514046 470034 514102
rect 470090 514046 470158 514102
rect 470214 514046 470282 514102
rect 470338 514046 470406 514102
rect 470462 514046 500754 514102
rect 500810 514046 500878 514102
rect 500934 514046 501002 514102
rect 501058 514046 501126 514102
rect 501182 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 70674 513978
rect 70730 513922 70798 513978
rect 70854 513922 70922 513978
rect 70978 513922 71046 513978
rect 71102 513922 101394 513978
rect 101450 513922 101518 513978
rect 101574 513922 101642 513978
rect 101698 513922 101766 513978
rect 101822 513922 132114 513978
rect 132170 513922 132238 513978
rect 132294 513922 132362 513978
rect 132418 513922 132486 513978
rect 132542 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 193554 513978
rect 193610 513922 193678 513978
rect 193734 513922 193802 513978
rect 193858 513922 193926 513978
rect 193982 513922 224274 513978
rect 224330 513922 224398 513978
rect 224454 513922 224522 513978
rect 224578 513922 224646 513978
rect 224702 513922 254994 513978
rect 255050 513922 255118 513978
rect 255174 513922 255242 513978
rect 255298 513922 255366 513978
rect 255422 513922 285714 513978
rect 285770 513922 285838 513978
rect 285894 513922 285962 513978
rect 286018 513922 286086 513978
rect 286142 513922 316434 513978
rect 316490 513922 316558 513978
rect 316614 513922 316682 513978
rect 316738 513922 316806 513978
rect 316862 513922 347154 513978
rect 347210 513922 347278 513978
rect 347334 513922 347402 513978
rect 347458 513922 347526 513978
rect 347582 513922 377874 513978
rect 377930 513922 377998 513978
rect 378054 513922 378122 513978
rect 378178 513922 378246 513978
rect 378302 513922 408594 513978
rect 408650 513922 408718 513978
rect 408774 513922 408842 513978
rect 408898 513922 408966 513978
rect 409022 513922 439314 513978
rect 439370 513922 439438 513978
rect 439494 513922 439562 513978
rect 439618 513922 439686 513978
rect 439742 513922 470034 513978
rect 470090 513922 470158 513978
rect 470214 513922 470282 513978
rect 470338 513922 470406 513978
rect 470462 513922 500754 513978
rect 500810 513922 500878 513978
rect 500934 513922 501002 513978
rect 501058 513922 501126 513978
rect 501182 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 66954 508350
rect 67010 508294 67078 508350
rect 67134 508294 67202 508350
rect 67258 508294 67326 508350
rect 67382 508294 97674 508350
rect 97730 508294 97798 508350
rect 97854 508294 97922 508350
rect 97978 508294 98046 508350
rect 98102 508294 128394 508350
rect 128450 508294 128518 508350
rect 128574 508294 128642 508350
rect 128698 508294 128766 508350
rect 128822 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 220554 508350
rect 220610 508294 220678 508350
rect 220734 508294 220802 508350
rect 220858 508294 220926 508350
rect 220982 508294 251274 508350
rect 251330 508294 251398 508350
rect 251454 508294 251522 508350
rect 251578 508294 251646 508350
rect 251702 508294 281994 508350
rect 282050 508294 282118 508350
rect 282174 508294 282242 508350
rect 282298 508294 282366 508350
rect 282422 508294 312714 508350
rect 312770 508294 312838 508350
rect 312894 508294 312962 508350
rect 313018 508294 313086 508350
rect 313142 508294 343434 508350
rect 343490 508294 343558 508350
rect 343614 508294 343682 508350
rect 343738 508294 343806 508350
rect 343862 508294 374154 508350
rect 374210 508294 374278 508350
rect 374334 508294 374402 508350
rect 374458 508294 374526 508350
rect 374582 508294 404874 508350
rect 404930 508294 404998 508350
rect 405054 508294 405122 508350
rect 405178 508294 405246 508350
rect 405302 508294 435594 508350
rect 435650 508294 435718 508350
rect 435774 508294 435842 508350
rect 435898 508294 435966 508350
rect 436022 508294 466314 508350
rect 466370 508294 466438 508350
rect 466494 508294 466562 508350
rect 466618 508294 466686 508350
rect 466742 508294 497034 508350
rect 497090 508294 497158 508350
rect 497214 508294 497282 508350
rect 497338 508294 497406 508350
rect 497462 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 66954 508226
rect 67010 508170 67078 508226
rect 67134 508170 67202 508226
rect 67258 508170 67326 508226
rect 67382 508170 97674 508226
rect 97730 508170 97798 508226
rect 97854 508170 97922 508226
rect 97978 508170 98046 508226
rect 98102 508170 128394 508226
rect 128450 508170 128518 508226
rect 128574 508170 128642 508226
rect 128698 508170 128766 508226
rect 128822 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 220554 508226
rect 220610 508170 220678 508226
rect 220734 508170 220802 508226
rect 220858 508170 220926 508226
rect 220982 508170 251274 508226
rect 251330 508170 251398 508226
rect 251454 508170 251522 508226
rect 251578 508170 251646 508226
rect 251702 508170 281994 508226
rect 282050 508170 282118 508226
rect 282174 508170 282242 508226
rect 282298 508170 282366 508226
rect 282422 508170 312714 508226
rect 312770 508170 312838 508226
rect 312894 508170 312962 508226
rect 313018 508170 313086 508226
rect 313142 508170 343434 508226
rect 343490 508170 343558 508226
rect 343614 508170 343682 508226
rect 343738 508170 343806 508226
rect 343862 508170 374154 508226
rect 374210 508170 374278 508226
rect 374334 508170 374402 508226
rect 374458 508170 374526 508226
rect 374582 508170 404874 508226
rect 404930 508170 404998 508226
rect 405054 508170 405122 508226
rect 405178 508170 405246 508226
rect 405302 508170 435594 508226
rect 435650 508170 435718 508226
rect 435774 508170 435842 508226
rect 435898 508170 435966 508226
rect 436022 508170 466314 508226
rect 466370 508170 466438 508226
rect 466494 508170 466562 508226
rect 466618 508170 466686 508226
rect 466742 508170 497034 508226
rect 497090 508170 497158 508226
rect 497214 508170 497282 508226
rect 497338 508170 497406 508226
rect 497462 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 66954 508102
rect 67010 508046 67078 508102
rect 67134 508046 67202 508102
rect 67258 508046 67326 508102
rect 67382 508046 97674 508102
rect 97730 508046 97798 508102
rect 97854 508046 97922 508102
rect 97978 508046 98046 508102
rect 98102 508046 128394 508102
rect 128450 508046 128518 508102
rect 128574 508046 128642 508102
rect 128698 508046 128766 508102
rect 128822 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 220554 508102
rect 220610 508046 220678 508102
rect 220734 508046 220802 508102
rect 220858 508046 220926 508102
rect 220982 508046 251274 508102
rect 251330 508046 251398 508102
rect 251454 508046 251522 508102
rect 251578 508046 251646 508102
rect 251702 508046 281994 508102
rect 282050 508046 282118 508102
rect 282174 508046 282242 508102
rect 282298 508046 282366 508102
rect 282422 508046 312714 508102
rect 312770 508046 312838 508102
rect 312894 508046 312962 508102
rect 313018 508046 313086 508102
rect 313142 508046 343434 508102
rect 343490 508046 343558 508102
rect 343614 508046 343682 508102
rect 343738 508046 343806 508102
rect 343862 508046 374154 508102
rect 374210 508046 374278 508102
rect 374334 508046 374402 508102
rect 374458 508046 374526 508102
rect 374582 508046 404874 508102
rect 404930 508046 404998 508102
rect 405054 508046 405122 508102
rect 405178 508046 405246 508102
rect 405302 508046 435594 508102
rect 435650 508046 435718 508102
rect 435774 508046 435842 508102
rect 435898 508046 435966 508102
rect 436022 508046 466314 508102
rect 466370 508046 466438 508102
rect 466494 508046 466562 508102
rect 466618 508046 466686 508102
rect 466742 508046 497034 508102
rect 497090 508046 497158 508102
rect 497214 508046 497282 508102
rect 497338 508046 497406 508102
rect 497462 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 66954 507978
rect 67010 507922 67078 507978
rect 67134 507922 67202 507978
rect 67258 507922 67326 507978
rect 67382 507922 97674 507978
rect 97730 507922 97798 507978
rect 97854 507922 97922 507978
rect 97978 507922 98046 507978
rect 98102 507922 128394 507978
rect 128450 507922 128518 507978
rect 128574 507922 128642 507978
rect 128698 507922 128766 507978
rect 128822 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 220554 507978
rect 220610 507922 220678 507978
rect 220734 507922 220802 507978
rect 220858 507922 220926 507978
rect 220982 507922 251274 507978
rect 251330 507922 251398 507978
rect 251454 507922 251522 507978
rect 251578 507922 251646 507978
rect 251702 507922 281994 507978
rect 282050 507922 282118 507978
rect 282174 507922 282242 507978
rect 282298 507922 282366 507978
rect 282422 507922 312714 507978
rect 312770 507922 312838 507978
rect 312894 507922 312962 507978
rect 313018 507922 313086 507978
rect 313142 507922 343434 507978
rect 343490 507922 343558 507978
rect 343614 507922 343682 507978
rect 343738 507922 343806 507978
rect 343862 507922 374154 507978
rect 374210 507922 374278 507978
rect 374334 507922 374402 507978
rect 374458 507922 374526 507978
rect 374582 507922 404874 507978
rect 404930 507922 404998 507978
rect 405054 507922 405122 507978
rect 405178 507922 405246 507978
rect 405302 507922 435594 507978
rect 435650 507922 435718 507978
rect 435774 507922 435842 507978
rect 435898 507922 435966 507978
rect 436022 507922 466314 507978
rect 466370 507922 466438 507978
rect 466494 507922 466562 507978
rect 466618 507922 466686 507978
rect 466742 507922 497034 507978
rect 497090 507922 497158 507978
rect 497214 507922 497282 507978
rect 497338 507922 497406 507978
rect 497462 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 70674 496350
rect 70730 496294 70798 496350
rect 70854 496294 70922 496350
rect 70978 496294 71046 496350
rect 71102 496294 101394 496350
rect 101450 496294 101518 496350
rect 101574 496294 101642 496350
rect 101698 496294 101766 496350
rect 101822 496294 132114 496350
rect 132170 496294 132238 496350
rect 132294 496294 132362 496350
rect 132418 496294 132486 496350
rect 132542 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 224274 496350
rect 224330 496294 224398 496350
rect 224454 496294 224522 496350
rect 224578 496294 224646 496350
rect 224702 496294 254994 496350
rect 255050 496294 255118 496350
rect 255174 496294 255242 496350
rect 255298 496294 255366 496350
rect 255422 496294 285714 496350
rect 285770 496294 285838 496350
rect 285894 496294 285962 496350
rect 286018 496294 286086 496350
rect 286142 496294 316434 496350
rect 316490 496294 316558 496350
rect 316614 496294 316682 496350
rect 316738 496294 316806 496350
rect 316862 496294 347154 496350
rect 347210 496294 347278 496350
rect 347334 496294 347402 496350
rect 347458 496294 347526 496350
rect 347582 496294 377874 496350
rect 377930 496294 377998 496350
rect 378054 496294 378122 496350
rect 378178 496294 378246 496350
rect 378302 496294 408594 496350
rect 408650 496294 408718 496350
rect 408774 496294 408842 496350
rect 408898 496294 408966 496350
rect 409022 496294 439314 496350
rect 439370 496294 439438 496350
rect 439494 496294 439562 496350
rect 439618 496294 439686 496350
rect 439742 496294 470034 496350
rect 470090 496294 470158 496350
rect 470214 496294 470282 496350
rect 470338 496294 470406 496350
rect 470462 496294 500754 496350
rect 500810 496294 500878 496350
rect 500934 496294 501002 496350
rect 501058 496294 501126 496350
rect 501182 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 70674 496226
rect 70730 496170 70798 496226
rect 70854 496170 70922 496226
rect 70978 496170 71046 496226
rect 71102 496170 101394 496226
rect 101450 496170 101518 496226
rect 101574 496170 101642 496226
rect 101698 496170 101766 496226
rect 101822 496170 132114 496226
rect 132170 496170 132238 496226
rect 132294 496170 132362 496226
rect 132418 496170 132486 496226
rect 132542 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 224274 496226
rect 224330 496170 224398 496226
rect 224454 496170 224522 496226
rect 224578 496170 224646 496226
rect 224702 496170 254994 496226
rect 255050 496170 255118 496226
rect 255174 496170 255242 496226
rect 255298 496170 255366 496226
rect 255422 496170 285714 496226
rect 285770 496170 285838 496226
rect 285894 496170 285962 496226
rect 286018 496170 286086 496226
rect 286142 496170 316434 496226
rect 316490 496170 316558 496226
rect 316614 496170 316682 496226
rect 316738 496170 316806 496226
rect 316862 496170 347154 496226
rect 347210 496170 347278 496226
rect 347334 496170 347402 496226
rect 347458 496170 347526 496226
rect 347582 496170 377874 496226
rect 377930 496170 377998 496226
rect 378054 496170 378122 496226
rect 378178 496170 378246 496226
rect 378302 496170 408594 496226
rect 408650 496170 408718 496226
rect 408774 496170 408842 496226
rect 408898 496170 408966 496226
rect 409022 496170 439314 496226
rect 439370 496170 439438 496226
rect 439494 496170 439562 496226
rect 439618 496170 439686 496226
rect 439742 496170 470034 496226
rect 470090 496170 470158 496226
rect 470214 496170 470282 496226
rect 470338 496170 470406 496226
rect 470462 496170 500754 496226
rect 500810 496170 500878 496226
rect 500934 496170 501002 496226
rect 501058 496170 501126 496226
rect 501182 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496046 70674 496102
rect 70730 496046 70798 496102
rect 70854 496046 70922 496102
rect 70978 496046 71046 496102
rect 71102 496046 101394 496102
rect 101450 496046 101518 496102
rect 101574 496046 101642 496102
rect 101698 496046 101766 496102
rect 101822 496046 132114 496102
rect 132170 496046 132238 496102
rect 132294 496046 132362 496102
rect 132418 496046 132486 496102
rect 132542 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 224274 496102
rect 224330 496046 224398 496102
rect 224454 496046 224522 496102
rect 224578 496046 224646 496102
rect 224702 496046 254994 496102
rect 255050 496046 255118 496102
rect 255174 496046 255242 496102
rect 255298 496046 255366 496102
rect 255422 496046 285714 496102
rect 285770 496046 285838 496102
rect 285894 496046 285962 496102
rect 286018 496046 286086 496102
rect 286142 496046 316434 496102
rect 316490 496046 316558 496102
rect 316614 496046 316682 496102
rect 316738 496046 316806 496102
rect 316862 496046 347154 496102
rect 347210 496046 347278 496102
rect 347334 496046 347402 496102
rect 347458 496046 347526 496102
rect 347582 496046 377874 496102
rect 377930 496046 377998 496102
rect 378054 496046 378122 496102
rect 378178 496046 378246 496102
rect 378302 496046 408594 496102
rect 408650 496046 408718 496102
rect 408774 496046 408842 496102
rect 408898 496046 408966 496102
rect 409022 496046 439314 496102
rect 439370 496046 439438 496102
rect 439494 496046 439562 496102
rect 439618 496046 439686 496102
rect 439742 496046 470034 496102
rect 470090 496046 470158 496102
rect 470214 496046 470282 496102
rect 470338 496046 470406 496102
rect 470462 496046 500754 496102
rect 500810 496046 500878 496102
rect 500934 496046 501002 496102
rect 501058 496046 501126 496102
rect 501182 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 495978 597980 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495922 70674 495978
rect 70730 495922 70798 495978
rect 70854 495922 70922 495978
rect 70978 495922 71046 495978
rect 71102 495922 101394 495978
rect 101450 495922 101518 495978
rect 101574 495922 101642 495978
rect 101698 495922 101766 495978
rect 101822 495922 132114 495978
rect 132170 495922 132238 495978
rect 132294 495922 132362 495978
rect 132418 495922 132486 495978
rect 132542 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 224274 495978
rect 224330 495922 224398 495978
rect 224454 495922 224522 495978
rect 224578 495922 224646 495978
rect 224702 495922 254994 495978
rect 255050 495922 255118 495978
rect 255174 495922 255242 495978
rect 255298 495922 255366 495978
rect 255422 495922 285714 495978
rect 285770 495922 285838 495978
rect 285894 495922 285962 495978
rect 286018 495922 286086 495978
rect 286142 495922 316434 495978
rect 316490 495922 316558 495978
rect 316614 495922 316682 495978
rect 316738 495922 316806 495978
rect 316862 495922 347154 495978
rect 347210 495922 347278 495978
rect 347334 495922 347402 495978
rect 347458 495922 347526 495978
rect 347582 495922 377874 495978
rect 377930 495922 377998 495978
rect 378054 495922 378122 495978
rect 378178 495922 378246 495978
rect 378302 495922 408594 495978
rect 408650 495922 408718 495978
rect 408774 495922 408842 495978
rect 408898 495922 408966 495978
rect 409022 495922 439314 495978
rect 439370 495922 439438 495978
rect 439494 495922 439562 495978
rect 439618 495922 439686 495978
rect 439742 495922 470034 495978
rect 470090 495922 470158 495978
rect 470214 495922 470282 495978
rect 470338 495922 470406 495978
rect 470462 495922 500754 495978
rect 500810 495922 500878 495978
rect 500934 495922 501002 495978
rect 501058 495922 501126 495978
rect 501182 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 66954 490350
rect 67010 490294 67078 490350
rect 67134 490294 67202 490350
rect 67258 490294 67326 490350
rect 67382 490294 97674 490350
rect 97730 490294 97798 490350
rect 97854 490294 97922 490350
rect 97978 490294 98046 490350
rect 98102 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 220554 490350
rect 220610 490294 220678 490350
rect 220734 490294 220802 490350
rect 220858 490294 220926 490350
rect 220982 490294 251274 490350
rect 251330 490294 251398 490350
rect 251454 490294 251522 490350
rect 251578 490294 251646 490350
rect 251702 490294 281994 490350
rect 282050 490294 282118 490350
rect 282174 490294 282242 490350
rect 282298 490294 282366 490350
rect 282422 490294 312714 490350
rect 312770 490294 312838 490350
rect 312894 490294 312962 490350
rect 313018 490294 313086 490350
rect 313142 490294 343434 490350
rect 343490 490294 343558 490350
rect 343614 490294 343682 490350
rect 343738 490294 343806 490350
rect 343862 490294 374154 490350
rect 374210 490294 374278 490350
rect 374334 490294 374402 490350
rect 374458 490294 374526 490350
rect 374582 490294 404874 490350
rect 404930 490294 404998 490350
rect 405054 490294 405122 490350
rect 405178 490294 405246 490350
rect 405302 490294 435594 490350
rect 435650 490294 435718 490350
rect 435774 490294 435842 490350
rect 435898 490294 435966 490350
rect 436022 490294 466314 490350
rect 466370 490294 466438 490350
rect 466494 490294 466562 490350
rect 466618 490294 466686 490350
rect 466742 490294 497034 490350
rect 497090 490294 497158 490350
rect 497214 490294 497282 490350
rect 497338 490294 497406 490350
rect 497462 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 66954 490226
rect 67010 490170 67078 490226
rect 67134 490170 67202 490226
rect 67258 490170 67326 490226
rect 67382 490170 97674 490226
rect 97730 490170 97798 490226
rect 97854 490170 97922 490226
rect 97978 490170 98046 490226
rect 98102 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 220554 490226
rect 220610 490170 220678 490226
rect 220734 490170 220802 490226
rect 220858 490170 220926 490226
rect 220982 490170 251274 490226
rect 251330 490170 251398 490226
rect 251454 490170 251522 490226
rect 251578 490170 251646 490226
rect 251702 490170 281994 490226
rect 282050 490170 282118 490226
rect 282174 490170 282242 490226
rect 282298 490170 282366 490226
rect 282422 490170 312714 490226
rect 312770 490170 312838 490226
rect 312894 490170 312962 490226
rect 313018 490170 313086 490226
rect 313142 490170 343434 490226
rect 343490 490170 343558 490226
rect 343614 490170 343682 490226
rect 343738 490170 343806 490226
rect 343862 490170 374154 490226
rect 374210 490170 374278 490226
rect 374334 490170 374402 490226
rect 374458 490170 374526 490226
rect 374582 490170 404874 490226
rect 404930 490170 404998 490226
rect 405054 490170 405122 490226
rect 405178 490170 405246 490226
rect 405302 490170 435594 490226
rect 435650 490170 435718 490226
rect 435774 490170 435842 490226
rect 435898 490170 435966 490226
rect 436022 490170 466314 490226
rect 466370 490170 466438 490226
rect 466494 490170 466562 490226
rect 466618 490170 466686 490226
rect 466742 490170 497034 490226
rect 497090 490170 497158 490226
rect 497214 490170 497282 490226
rect 497338 490170 497406 490226
rect 497462 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 66954 490102
rect 67010 490046 67078 490102
rect 67134 490046 67202 490102
rect 67258 490046 67326 490102
rect 67382 490046 97674 490102
rect 97730 490046 97798 490102
rect 97854 490046 97922 490102
rect 97978 490046 98046 490102
rect 98102 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 220554 490102
rect 220610 490046 220678 490102
rect 220734 490046 220802 490102
rect 220858 490046 220926 490102
rect 220982 490046 251274 490102
rect 251330 490046 251398 490102
rect 251454 490046 251522 490102
rect 251578 490046 251646 490102
rect 251702 490046 281994 490102
rect 282050 490046 282118 490102
rect 282174 490046 282242 490102
rect 282298 490046 282366 490102
rect 282422 490046 312714 490102
rect 312770 490046 312838 490102
rect 312894 490046 312962 490102
rect 313018 490046 313086 490102
rect 313142 490046 343434 490102
rect 343490 490046 343558 490102
rect 343614 490046 343682 490102
rect 343738 490046 343806 490102
rect 343862 490046 374154 490102
rect 374210 490046 374278 490102
rect 374334 490046 374402 490102
rect 374458 490046 374526 490102
rect 374582 490046 404874 490102
rect 404930 490046 404998 490102
rect 405054 490046 405122 490102
rect 405178 490046 405246 490102
rect 405302 490046 435594 490102
rect 435650 490046 435718 490102
rect 435774 490046 435842 490102
rect 435898 490046 435966 490102
rect 436022 490046 466314 490102
rect 466370 490046 466438 490102
rect 466494 490046 466562 490102
rect 466618 490046 466686 490102
rect 466742 490046 497034 490102
rect 497090 490046 497158 490102
rect 497214 490046 497282 490102
rect 497338 490046 497406 490102
rect 497462 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 66954 489978
rect 67010 489922 67078 489978
rect 67134 489922 67202 489978
rect 67258 489922 67326 489978
rect 67382 489922 97674 489978
rect 97730 489922 97798 489978
rect 97854 489922 97922 489978
rect 97978 489922 98046 489978
rect 98102 489922 128394 489978
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 220554 489978
rect 220610 489922 220678 489978
rect 220734 489922 220802 489978
rect 220858 489922 220926 489978
rect 220982 489922 251274 489978
rect 251330 489922 251398 489978
rect 251454 489922 251522 489978
rect 251578 489922 251646 489978
rect 251702 489922 281994 489978
rect 282050 489922 282118 489978
rect 282174 489922 282242 489978
rect 282298 489922 282366 489978
rect 282422 489922 312714 489978
rect 312770 489922 312838 489978
rect 312894 489922 312962 489978
rect 313018 489922 313086 489978
rect 313142 489922 343434 489978
rect 343490 489922 343558 489978
rect 343614 489922 343682 489978
rect 343738 489922 343806 489978
rect 343862 489922 374154 489978
rect 374210 489922 374278 489978
rect 374334 489922 374402 489978
rect 374458 489922 374526 489978
rect 374582 489922 404874 489978
rect 404930 489922 404998 489978
rect 405054 489922 405122 489978
rect 405178 489922 405246 489978
rect 405302 489922 435594 489978
rect 435650 489922 435718 489978
rect 435774 489922 435842 489978
rect 435898 489922 435966 489978
rect 436022 489922 466314 489978
rect 466370 489922 466438 489978
rect 466494 489922 466562 489978
rect 466618 489922 466686 489978
rect 466742 489922 497034 489978
rect 497090 489922 497158 489978
rect 497214 489922 497282 489978
rect 497338 489922 497406 489978
rect 497462 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 101394 478350
rect 101450 478294 101518 478350
rect 101574 478294 101642 478350
rect 101698 478294 101766 478350
rect 101822 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 224274 478350
rect 224330 478294 224398 478350
rect 224454 478294 224522 478350
rect 224578 478294 224646 478350
rect 224702 478294 254994 478350
rect 255050 478294 255118 478350
rect 255174 478294 255242 478350
rect 255298 478294 255366 478350
rect 255422 478294 285714 478350
rect 285770 478294 285838 478350
rect 285894 478294 285962 478350
rect 286018 478294 286086 478350
rect 286142 478294 316434 478350
rect 316490 478294 316558 478350
rect 316614 478294 316682 478350
rect 316738 478294 316806 478350
rect 316862 478294 347154 478350
rect 347210 478294 347278 478350
rect 347334 478294 347402 478350
rect 347458 478294 347526 478350
rect 347582 478294 377874 478350
rect 377930 478294 377998 478350
rect 378054 478294 378122 478350
rect 378178 478294 378246 478350
rect 378302 478294 408594 478350
rect 408650 478294 408718 478350
rect 408774 478294 408842 478350
rect 408898 478294 408966 478350
rect 409022 478294 439314 478350
rect 439370 478294 439438 478350
rect 439494 478294 439562 478350
rect 439618 478294 439686 478350
rect 439742 478294 470034 478350
rect 470090 478294 470158 478350
rect 470214 478294 470282 478350
rect 470338 478294 470406 478350
rect 470462 478294 500754 478350
rect 500810 478294 500878 478350
rect 500934 478294 501002 478350
rect 501058 478294 501126 478350
rect 501182 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 101394 478226
rect 101450 478170 101518 478226
rect 101574 478170 101642 478226
rect 101698 478170 101766 478226
rect 101822 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 224274 478226
rect 224330 478170 224398 478226
rect 224454 478170 224522 478226
rect 224578 478170 224646 478226
rect 224702 478170 254994 478226
rect 255050 478170 255118 478226
rect 255174 478170 255242 478226
rect 255298 478170 255366 478226
rect 255422 478170 285714 478226
rect 285770 478170 285838 478226
rect 285894 478170 285962 478226
rect 286018 478170 286086 478226
rect 286142 478170 316434 478226
rect 316490 478170 316558 478226
rect 316614 478170 316682 478226
rect 316738 478170 316806 478226
rect 316862 478170 347154 478226
rect 347210 478170 347278 478226
rect 347334 478170 347402 478226
rect 347458 478170 347526 478226
rect 347582 478170 377874 478226
rect 377930 478170 377998 478226
rect 378054 478170 378122 478226
rect 378178 478170 378246 478226
rect 378302 478170 408594 478226
rect 408650 478170 408718 478226
rect 408774 478170 408842 478226
rect 408898 478170 408966 478226
rect 409022 478170 439314 478226
rect 439370 478170 439438 478226
rect 439494 478170 439562 478226
rect 439618 478170 439686 478226
rect 439742 478170 470034 478226
rect 470090 478170 470158 478226
rect 470214 478170 470282 478226
rect 470338 478170 470406 478226
rect 470462 478170 500754 478226
rect 500810 478170 500878 478226
rect 500934 478170 501002 478226
rect 501058 478170 501126 478226
rect 501182 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 101394 478102
rect 101450 478046 101518 478102
rect 101574 478046 101642 478102
rect 101698 478046 101766 478102
rect 101822 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 224274 478102
rect 224330 478046 224398 478102
rect 224454 478046 224522 478102
rect 224578 478046 224646 478102
rect 224702 478046 254994 478102
rect 255050 478046 255118 478102
rect 255174 478046 255242 478102
rect 255298 478046 255366 478102
rect 255422 478046 285714 478102
rect 285770 478046 285838 478102
rect 285894 478046 285962 478102
rect 286018 478046 286086 478102
rect 286142 478046 316434 478102
rect 316490 478046 316558 478102
rect 316614 478046 316682 478102
rect 316738 478046 316806 478102
rect 316862 478046 347154 478102
rect 347210 478046 347278 478102
rect 347334 478046 347402 478102
rect 347458 478046 347526 478102
rect 347582 478046 377874 478102
rect 377930 478046 377998 478102
rect 378054 478046 378122 478102
rect 378178 478046 378246 478102
rect 378302 478046 408594 478102
rect 408650 478046 408718 478102
rect 408774 478046 408842 478102
rect 408898 478046 408966 478102
rect 409022 478046 439314 478102
rect 439370 478046 439438 478102
rect 439494 478046 439562 478102
rect 439618 478046 439686 478102
rect 439742 478046 470034 478102
rect 470090 478046 470158 478102
rect 470214 478046 470282 478102
rect 470338 478046 470406 478102
rect 470462 478046 500754 478102
rect 500810 478046 500878 478102
rect 500934 478046 501002 478102
rect 501058 478046 501126 478102
rect 501182 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 101394 477978
rect 101450 477922 101518 477978
rect 101574 477922 101642 477978
rect 101698 477922 101766 477978
rect 101822 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 224274 477978
rect 224330 477922 224398 477978
rect 224454 477922 224522 477978
rect 224578 477922 224646 477978
rect 224702 477922 254994 477978
rect 255050 477922 255118 477978
rect 255174 477922 255242 477978
rect 255298 477922 255366 477978
rect 255422 477922 285714 477978
rect 285770 477922 285838 477978
rect 285894 477922 285962 477978
rect 286018 477922 286086 477978
rect 286142 477922 316434 477978
rect 316490 477922 316558 477978
rect 316614 477922 316682 477978
rect 316738 477922 316806 477978
rect 316862 477922 347154 477978
rect 347210 477922 347278 477978
rect 347334 477922 347402 477978
rect 347458 477922 347526 477978
rect 347582 477922 377874 477978
rect 377930 477922 377998 477978
rect 378054 477922 378122 477978
rect 378178 477922 378246 477978
rect 378302 477922 408594 477978
rect 408650 477922 408718 477978
rect 408774 477922 408842 477978
rect 408898 477922 408966 477978
rect 409022 477922 439314 477978
rect 439370 477922 439438 477978
rect 439494 477922 439562 477978
rect 439618 477922 439686 477978
rect 439742 477922 470034 477978
rect 470090 477922 470158 477978
rect 470214 477922 470282 477978
rect 470338 477922 470406 477978
rect 470462 477922 500754 477978
rect 500810 477922 500878 477978
rect 500934 477922 501002 477978
rect 501058 477922 501126 477978
rect 501182 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 220554 472350
rect 220610 472294 220678 472350
rect 220734 472294 220802 472350
rect 220858 472294 220926 472350
rect 220982 472294 251274 472350
rect 251330 472294 251398 472350
rect 251454 472294 251522 472350
rect 251578 472294 251646 472350
rect 251702 472294 281994 472350
rect 282050 472294 282118 472350
rect 282174 472294 282242 472350
rect 282298 472294 282366 472350
rect 282422 472294 312714 472350
rect 312770 472294 312838 472350
rect 312894 472294 312962 472350
rect 313018 472294 313086 472350
rect 313142 472294 343434 472350
rect 343490 472294 343558 472350
rect 343614 472294 343682 472350
rect 343738 472294 343806 472350
rect 343862 472294 374154 472350
rect 374210 472294 374278 472350
rect 374334 472294 374402 472350
rect 374458 472294 374526 472350
rect 374582 472294 404874 472350
rect 404930 472294 404998 472350
rect 405054 472294 405122 472350
rect 405178 472294 405246 472350
rect 405302 472294 435594 472350
rect 435650 472294 435718 472350
rect 435774 472294 435842 472350
rect 435898 472294 435966 472350
rect 436022 472294 466314 472350
rect 466370 472294 466438 472350
rect 466494 472294 466562 472350
rect 466618 472294 466686 472350
rect 466742 472294 497034 472350
rect 497090 472294 497158 472350
rect 497214 472294 497282 472350
rect 497338 472294 497406 472350
rect 497462 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 220554 472226
rect 220610 472170 220678 472226
rect 220734 472170 220802 472226
rect 220858 472170 220926 472226
rect 220982 472170 251274 472226
rect 251330 472170 251398 472226
rect 251454 472170 251522 472226
rect 251578 472170 251646 472226
rect 251702 472170 281994 472226
rect 282050 472170 282118 472226
rect 282174 472170 282242 472226
rect 282298 472170 282366 472226
rect 282422 472170 312714 472226
rect 312770 472170 312838 472226
rect 312894 472170 312962 472226
rect 313018 472170 313086 472226
rect 313142 472170 343434 472226
rect 343490 472170 343558 472226
rect 343614 472170 343682 472226
rect 343738 472170 343806 472226
rect 343862 472170 374154 472226
rect 374210 472170 374278 472226
rect 374334 472170 374402 472226
rect 374458 472170 374526 472226
rect 374582 472170 404874 472226
rect 404930 472170 404998 472226
rect 405054 472170 405122 472226
rect 405178 472170 405246 472226
rect 405302 472170 435594 472226
rect 435650 472170 435718 472226
rect 435774 472170 435842 472226
rect 435898 472170 435966 472226
rect 436022 472170 466314 472226
rect 466370 472170 466438 472226
rect 466494 472170 466562 472226
rect 466618 472170 466686 472226
rect 466742 472170 497034 472226
rect 497090 472170 497158 472226
rect 497214 472170 497282 472226
rect 497338 472170 497406 472226
rect 497462 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 220554 472102
rect 220610 472046 220678 472102
rect 220734 472046 220802 472102
rect 220858 472046 220926 472102
rect 220982 472046 251274 472102
rect 251330 472046 251398 472102
rect 251454 472046 251522 472102
rect 251578 472046 251646 472102
rect 251702 472046 281994 472102
rect 282050 472046 282118 472102
rect 282174 472046 282242 472102
rect 282298 472046 282366 472102
rect 282422 472046 312714 472102
rect 312770 472046 312838 472102
rect 312894 472046 312962 472102
rect 313018 472046 313086 472102
rect 313142 472046 343434 472102
rect 343490 472046 343558 472102
rect 343614 472046 343682 472102
rect 343738 472046 343806 472102
rect 343862 472046 374154 472102
rect 374210 472046 374278 472102
rect 374334 472046 374402 472102
rect 374458 472046 374526 472102
rect 374582 472046 404874 472102
rect 404930 472046 404998 472102
rect 405054 472046 405122 472102
rect 405178 472046 405246 472102
rect 405302 472046 435594 472102
rect 435650 472046 435718 472102
rect 435774 472046 435842 472102
rect 435898 472046 435966 472102
rect 436022 472046 466314 472102
rect 466370 472046 466438 472102
rect 466494 472046 466562 472102
rect 466618 472046 466686 472102
rect 466742 472046 497034 472102
rect 497090 472046 497158 472102
rect 497214 472046 497282 472102
rect 497338 472046 497406 472102
rect 497462 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 220554 471978
rect 220610 471922 220678 471978
rect 220734 471922 220802 471978
rect 220858 471922 220926 471978
rect 220982 471922 251274 471978
rect 251330 471922 251398 471978
rect 251454 471922 251522 471978
rect 251578 471922 251646 471978
rect 251702 471922 281994 471978
rect 282050 471922 282118 471978
rect 282174 471922 282242 471978
rect 282298 471922 282366 471978
rect 282422 471922 312714 471978
rect 312770 471922 312838 471978
rect 312894 471922 312962 471978
rect 313018 471922 313086 471978
rect 313142 471922 343434 471978
rect 343490 471922 343558 471978
rect 343614 471922 343682 471978
rect 343738 471922 343806 471978
rect 343862 471922 374154 471978
rect 374210 471922 374278 471978
rect 374334 471922 374402 471978
rect 374458 471922 374526 471978
rect 374582 471922 404874 471978
rect 404930 471922 404998 471978
rect 405054 471922 405122 471978
rect 405178 471922 405246 471978
rect 405302 471922 435594 471978
rect 435650 471922 435718 471978
rect 435774 471922 435842 471978
rect 435898 471922 435966 471978
rect 436022 471922 466314 471978
rect 466370 471922 466438 471978
rect 466494 471922 466562 471978
rect 466618 471922 466686 471978
rect 466742 471922 497034 471978
rect 497090 471922 497158 471978
rect 497214 471922 497282 471978
rect 497338 471922 497406 471978
rect 497462 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 224274 460350
rect 224330 460294 224398 460350
rect 224454 460294 224522 460350
rect 224578 460294 224646 460350
rect 224702 460294 254994 460350
rect 255050 460294 255118 460350
rect 255174 460294 255242 460350
rect 255298 460294 255366 460350
rect 255422 460294 285714 460350
rect 285770 460294 285838 460350
rect 285894 460294 285962 460350
rect 286018 460294 286086 460350
rect 286142 460294 316434 460350
rect 316490 460294 316558 460350
rect 316614 460294 316682 460350
rect 316738 460294 316806 460350
rect 316862 460294 347154 460350
rect 347210 460294 347278 460350
rect 347334 460294 347402 460350
rect 347458 460294 347526 460350
rect 347582 460294 377874 460350
rect 377930 460294 377998 460350
rect 378054 460294 378122 460350
rect 378178 460294 378246 460350
rect 378302 460294 408594 460350
rect 408650 460294 408718 460350
rect 408774 460294 408842 460350
rect 408898 460294 408966 460350
rect 409022 460294 439314 460350
rect 439370 460294 439438 460350
rect 439494 460294 439562 460350
rect 439618 460294 439686 460350
rect 439742 460294 470034 460350
rect 470090 460294 470158 460350
rect 470214 460294 470282 460350
rect 470338 460294 470406 460350
rect 470462 460294 500754 460350
rect 500810 460294 500878 460350
rect 500934 460294 501002 460350
rect 501058 460294 501126 460350
rect 501182 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 224274 460226
rect 224330 460170 224398 460226
rect 224454 460170 224522 460226
rect 224578 460170 224646 460226
rect 224702 460170 254994 460226
rect 255050 460170 255118 460226
rect 255174 460170 255242 460226
rect 255298 460170 255366 460226
rect 255422 460170 285714 460226
rect 285770 460170 285838 460226
rect 285894 460170 285962 460226
rect 286018 460170 286086 460226
rect 286142 460170 316434 460226
rect 316490 460170 316558 460226
rect 316614 460170 316682 460226
rect 316738 460170 316806 460226
rect 316862 460170 347154 460226
rect 347210 460170 347278 460226
rect 347334 460170 347402 460226
rect 347458 460170 347526 460226
rect 347582 460170 377874 460226
rect 377930 460170 377998 460226
rect 378054 460170 378122 460226
rect 378178 460170 378246 460226
rect 378302 460170 408594 460226
rect 408650 460170 408718 460226
rect 408774 460170 408842 460226
rect 408898 460170 408966 460226
rect 409022 460170 439314 460226
rect 439370 460170 439438 460226
rect 439494 460170 439562 460226
rect 439618 460170 439686 460226
rect 439742 460170 470034 460226
rect 470090 460170 470158 460226
rect 470214 460170 470282 460226
rect 470338 460170 470406 460226
rect 470462 460170 500754 460226
rect 500810 460170 500878 460226
rect 500934 460170 501002 460226
rect 501058 460170 501126 460226
rect 501182 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 224274 460102
rect 224330 460046 224398 460102
rect 224454 460046 224522 460102
rect 224578 460046 224646 460102
rect 224702 460046 254994 460102
rect 255050 460046 255118 460102
rect 255174 460046 255242 460102
rect 255298 460046 255366 460102
rect 255422 460046 285714 460102
rect 285770 460046 285838 460102
rect 285894 460046 285962 460102
rect 286018 460046 286086 460102
rect 286142 460046 316434 460102
rect 316490 460046 316558 460102
rect 316614 460046 316682 460102
rect 316738 460046 316806 460102
rect 316862 460046 347154 460102
rect 347210 460046 347278 460102
rect 347334 460046 347402 460102
rect 347458 460046 347526 460102
rect 347582 460046 377874 460102
rect 377930 460046 377998 460102
rect 378054 460046 378122 460102
rect 378178 460046 378246 460102
rect 378302 460046 408594 460102
rect 408650 460046 408718 460102
rect 408774 460046 408842 460102
rect 408898 460046 408966 460102
rect 409022 460046 439314 460102
rect 439370 460046 439438 460102
rect 439494 460046 439562 460102
rect 439618 460046 439686 460102
rect 439742 460046 470034 460102
rect 470090 460046 470158 460102
rect 470214 460046 470282 460102
rect 470338 460046 470406 460102
rect 470462 460046 500754 460102
rect 500810 460046 500878 460102
rect 500934 460046 501002 460102
rect 501058 460046 501126 460102
rect 501182 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 224274 459978
rect 224330 459922 224398 459978
rect 224454 459922 224522 459978
rect 224578 459922 224646 459978
rect 224702 459922 254994 459978
rect 255050 459922 255118 459978
rect 255174 459922 255242 459978
rect 255298 459922 255366 459978
rect 255422 459922 285714 459978
rect 285770 459922 285838 459978
rect 285894 459922 285962 459978
rect 286018 459922 286086 459978
rect 286142 459922 316434 459978
rect 316490 459922 316558 459978
rect 316614 459922 316682 459978
rect 316738 459922 316806 459978
rect 316862 459922 347154 459978
rect 347210 459922 347278 459978
rect 347334 459922 347402 459978
rect 347458 459922 347526 459978
rect 347582 459922 377874 459978
rect 377930 459922 377998 459978
rect 378054 459922 378122 459978
rect 378178 459922 378246 459978
rect 378302 459922 408594 459978
rect 408650 459922 408718 459978
rect 408774 459922 408842 459978
rect 408898 459922 408966 459978
rect 409022 459922 439314 459978
rect 439370 459922 439438 459978
rect 439494 459922 439562 459978
rect 439618 459922 439686 459978
rect 439742 459922 470034 459978
rect 470090 459922 470158 459978
rect 470214 459922 470282 459978
rect 470338 459922 470406 459978
rect 470462 459922 500754 459978
rect 500810 459922 500878 459978
rect 500934 459922 501002 459978
rect 501058 459922 501126 459978
rect 501182 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 220554 454350
rect 220610 454294 220678 454350
rect 220734 454294 220802 454350
rect 220858 454294 220926 454350
rect 220982 454294 251274 454350
rect 251330 454294 251398 454350
rect 251454 454294 251522 454350
rect 251578 454294 251646 454350
rect 251702 454294 281994 454350
rect 282050 454294 282118 454350
rect 282174 454294 282242 454350
rect 282298 454294 282366 454350
rect 282422 454294 312714 454350
rect 312770 454294 312838 454350
rect 312894 454294 312962 454350
rect 313018 454294 313086 454350
rect 313142 454294 343434 454350
rect 343490 454294 343558 454350
rect 343614 454294 343682 454350
rect 343738 454294 343806 454350
rect 343862 454294 374154 454350
rect 374210 454294 374278 454350
rect 374334 454294 374402 454350
rect 374458 454294 374526 454350
rect 374582 454294 404874 454350
rect 404930 454294 404998 454350
rect 405054 454294 405122 454350
rect 405178 454294 405246 454350
rect 405302 454294 435594 454350
rect 435650 454294 435718 454350
rect 435774 454294 435842 454350
rect 435898 454294 435966 454350
rect 436022 454294 466314 454350
rect 466370 454294 466438 454350
rect 466494 454294 466562 454350
rect 466618 454294 466686 454350
rect 466742 454294 497034 454350
rect 497090 454294 497158 454350
rect 497214 454294 497282 454350
rect 497338 454294 497406 454350
rect 497462 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 220554 454226
rect 220610 454170 220678 454226
rect 220734 454170 220802 454226
rect 220858 454170 220926 454226
rect 220982 454170 251274 454226
rect 251330 454170 251398 454226
rect 251454 454170 251522 454226
rect 251578 454170 251646 454226
rect 251702 454170 281994 454226
rect 282050 454170 282118 454226
rect 282174 454170 282242 454226
rect 282298 454170 282366 454226
rect 282422 454170 312714 454226
rect 312770 454170 312838 454226
rect 312894 454170 312962 454226
rect 313018 454170 313086 454226
rect 313142 454170 343434 454226
rect 343490 454170 343558 454226
rect 343614 454170 343682 454226
rect 343738 454170 343806 454226
rect 343862 454170 374154 454226
rect 374210 454170 374278 454226
rect 374334 454170 374402 454226
rect 374458 454170 374526 454226
rect 374582 454170 404874 454226
rect 404930 454170 404998 454226
rect 405054 454170 405122 454226
rect 405178 454170 405246 454226
rect 405302 454170 435594 454226
rect 435650 454170 435718 454226
rect 435774 454170 435842 454226
rect 435898 454170 435966 454226
rect 436022 454170 466314 454226
rect 466370 454170 466438 454226
rect 466494 454170 466562 454226
rect 466618 454170 466686 454226
rect 466742 454170 497034 454226
rect 497090 454170 497158 454226
rect 497214 454170 497282 454226
rect 497338 454170 497406 454226
rect 497462 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 220554 454102
rect 220610 454046 220678 454102
rect 220734 454046 220802 454102
rect 220858 454046 220926 454102
rect 220982 454046 251274 454102
rect 251330 454046 251398 454102
rect 251454 454046 251522 454102
rect 251578 454046 251646 454102
rect 251702 454046 281994 454102
rect 282050 454046 282118 454102
rect 282174 454046 282242 454102
rect 282298 454046 282366 454102
rect 282422 454046 312714 454102
rect 312770 454046 312838 454102
rect 312894 454046 312962 454102
rect 313018 454046 313086 454102
rect 313142 454046 343434 454102
rect 343490 454046 343558 454102
rect 343614 454046 343682 454102
rect 343738 454046 343806 454102
rect 343862 454046 374154 454102
rect 374210 454046 374278 454102
rect 374334 454046 374402 454102
rect 374458 454046 374526 454102
rect 374582 454046 404874 454102
rect 404930 454046 404998 454102
rect 405054 454046 405122 454102
rect 405178 454046 405246 454102
rect 405302 454046 435594 454102
rect 435650 454046 435718 454102
rect 435774 454046 435842 454102
rect 435898 454046 435966 454102
rect 436022 454046 466314 454102
rect 466370 454046 466438 454102
rect 466494 454046 466562 454102
rect 466618 454046 466686 454102
rect 466742 454046 497034 454102
rect 497090 454046 497158 454102
rect 497214 454046 497282 454102
rect 497338 454046 497406 454102
rect 497462 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 220554 453978
rect 220610 453922 220678 453978
rect 220734 453922 220802 453978
rect 220858 453922 220926 453978
rect 220982 453922 251274 453978
rect 251330 453922 251398 453978
rect 251454 453922 251522 453978
rect 251578 453922 251646 453978
rect 251702 453922 281994 453978
rect 282050 453922 282118 453978
rect 282174 453922 282242 453978
rect 282298 453922 282366 453978
rect 282422 453922 312714 453978
rect 312770 453922 312838 453978
rect 312894 453922 312962 453978
rect 313018 453922 313086 453978
rect 313142 453922 343434 453978
rect 343490 453922 343558 453978
rect 343614 453922 343682 453978
rect 343738 453922 343806 453978
rect 343862 453922 374154 453978
rect 374210 453922 374278 453978
rect 374334 453922 374402 453978
rect 374458 453922 374526 453978
rect 374582 453922 404874 453978
rect 404930 453922 404998 453978
rect 405054 453922 405122 453978
rect 405178 453922 405246 453978
rect 405302 453922 435594 453978
rect 435650 453922 435718 453978
rect 435774 453922 435842 453978
rect 435898 453922 435966 453978
rect 436022 453922 466314 453978
rect 466370 453922 466438 453978
rect 466494 453922 466562 453978
rect 466618 453922 466686 453978
rect 466742 453922 497034 453978
rect 497090 453922 497158 453978
rect 497214 453922 497282 453978
rect 497338 453922 497406 453978
rect 497462 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 224274 442350
rect 224330 442294 224398 442350
rect 224454 442294 224522 442350
rect 224578 442294 224646 442350
rect 224702 442294 254994 442350
rect 255050 442294 255118 442350
rect 255174 442294 255242 442350
rect 255298 442294 255366 442350
rect 255422 442294 285714 442350
rect 285770 442294 285838 442350
rect 285894 442294 285962 442350
rect 286018 442294 286086 442350
rect 286142 442294 316434 442350
rect 316490 442294 316558 442350
rect 316614 442294 316682 442350
rect 316738 442294 316806 442350
rect 316862 442294 347154 442350
rect 347210 442294 347278 442350
rect 347334 442294 347402 442350
rect 347458 442294 347526 442350
rect 347582 442294 377874 442350
rect 377930 442294 377998 442350
rect 378054 442294 378122 442350
rect 378178 442294 378246 442350
rect 378302 442294 408594 442350
rect 408650 442294 408718 442350
rect 408774 442294 408842 442350
rect 408898 442294 408966 442350
rect 409022 442294 439314 442350
rect 439370 442294 439438 442350
rect 439494 442294 439562 442350
rect 439618 442294 439686 442350
rect 439742 442294 470034 442350
rect 470090 442294 470158 442350
rect 470214 442294 470282 442350
rect 470338 442294 470406 442350
rect 470462 442294 500754 442350
rect 500810 442294 500878 442350
rect 500934 442294 501002 442350
rect 501058 442294 501126 442350
rect 501182 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 224274 442226
rect 224330 442170 224398 442226
rect 224454 442170 224522 442226
rect 224578 442170 224646 442226
rect 224702 442170 254994 442226
rect 255050 442170 255118 442226
rect 255174 442170 255242 442226
rect 255298 442170 255366 442226
rect 255422 442170 285714 442226
rect 285770 442170 285838 442226
rect 285894 442170 285962 442226
rect 286018 442170 286086 442226
rect 286142 442170 316434 442226
rect 316490 442170 316558 442226
rect 316614 442170 316682 442226
rect 316738 442170 316806 442226
rect 316862 442170 347154 442226
rect 347210 442170 347278 442226
rect 347334 442170 347402 442226
rect 347458 442170 347526 442226
rect 347582 442170 377874 442226
rect 377930 442170 377998 442226
rect 378054 442170 378122 442226
rect 378178 442170 378246 442226
rect 378302 442170 408594 442226
rect 408650 442170 408718 442226
rect 408774 442170 408842 442226
rect 408898 442170 408966 442226
rect 409022 442170 439314 442226
rect 439370 442170 439438 442226
rect 439494 442170 439562 442226
rect 439618 442170 439686 442226
rect 439742 442170 470034 442226
rect 470090 442170 470158 442226
rect 470214 442170 470282 442226
rect 470338 442170 470406 442226
rect 470462 442170 500754 442226
rect 500810 442170 500878 442226
rect 500934 442170 501002 442226
rect 501058 442170 501126 442226
rect 501182 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 224274 442102
rect 224330 442046 224398 442102
rect 224454 442046 224522 442102
rect 224578 442046 224646 442102
rect 224702 442046 254994 442102
rect 255050 442046 255118 442102
rect 255174 442046 255242 442102
rect 255298 442046 255366 442102
rect 255422 442046 285714 442102
rect 285770 442046 285838 442102
rect 285894 442046 285962 442102
rect 286018 442046 286086 442102
rect 286142 442046 316434 442102
rect 316490 442046 316558 442102
rect 316614 442046 316682 442102
rect 316738 442046 316806 442102
rect 316862 442046 347154 442102
rect 347210 442046 347278 442102
rect 347334 442046 347402 442102
rect 347458 442046 347526 442102
rect 347582 442046 377874 442102
rect 377930 442046 377998 442102
rect 378054 442046 378122 442102
rect 378178 442046 378246 442102
rect 378302 442046 408594 442102
rect 408650 442046 408718 442102
rect 408774 442046 408842 442102
rect 408898 442046 408966 442102
rect 409022 442046 439314 442102
rect 439370 442046 439438 442102
rect 439494 442046 439562 442102
rect 439618 442046 439686 442102
rect 439742 442046 470034 442102
rect 470090 442046 470158 442102
rect 470214 442046 470282 442102
rect 470338 442046 470406 442102
rect 470462 442046 500754 442102
rect 500810 442046 500878 442102
rect 500934 442046 501002 442102
rect 501058 442046 501126 442102
rect 501182 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 224274 441978
rect 224330 441922 224398 441978
rect 224454 441922 224522 441978
rect 224578 441922 224646 441978
rect 224702 441922 254994 441978
rect 255050 441922 255118 441978
rect 255174 441922 255242 441978
rect 255298 441922 255366 441978
rect 255422 441922 285714 441978
rect 285770 441922 285838 441978
rect 285894 441922 285962 441978
rect 286018 441922 286086 441978
rect 286142 441922 316434 441978
rect 316490 441922 316558 441978
rect 316614 441922 316682 441978
rect 316738 441922 316806 441978
rect 316862 441922 347154 441978
rect 347210 441922 347278 441978
rect 347334 441922 347402 441978
rect 347458 441922 347526 441978
rect 347582 441922 377874 441978
rect 377930 441922 377998 441978
rect 378054 441922 378122 441978
rect 378178 441922 378246 441978
rect 378302 441922 408594 441978
rect 408650 441922 408718 441978
rect 408774 441922 408842 441978
rect 408898 441922 408966 441978
rect 409022 441922 439314 441978
rect 439370 441922 439438 441978
rect 439494 441922 439562 441978
rect 439618 441922 439686 441978
rect 439742 441922 470034 441978
rect 470090 441922 470158 441978
rect 470214 441922 470282 441978
rect 470338 441922 470406 441978
rect 470462 441922 500754 441978
rect 500810 441922 500878 441978
rect 500934 441922 501002 441978
rect 501058 441922 501126 441978
rect 501182 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 220554 436350
rect 220610 436294 220678 436350
rect 220734 436294 220802 436350
rect 220858 436294 220926 436350
rect 220982 436294 251274 436350
rect 251330 436294 251398 436350
rect 251454 436294 251522 436350
rect 251578 436294 251646 436350
rect 251702 436294 281994 436350
rect 282050 436294 282118 436350
rect 282174 436294 282242 436350
rect 282298 436294 282366 436350
rect 282422 436294 312714 436350
rect 312770 436294 312838 436350
rect 312894 436294 312962 436350
rect 313018 436294 313086 436350
rect 313142 436294 343434 436350
rect 343490 436294 343558 436350
rect 343614 436294 343682 436350
rect 343738 436294 343806 436350
rect 343862 436294 374154 436350
rect 374210 436294 374278 436350
rect 374334 436294 374402 436350
rect 374458 436294 374526 436350
rect 374582 436294 404874 436350
rect 404930 436294 404998 436350
rect 405054 436294 405122 436350
rect 405178 436294 405246 436350
rect 405302 436294 435594 436350
rect 435650 436294 435718 436350
rect 435774 436294 435842 436350
rect 435898 436294 435966 436350
rect 436022 436294 466314 436350
rect 466370 436294 466438 436350
rect 466494 436294 466562 436350
rect 466618 436294 466686 436350
rect 466742 436294 497034 436350
rect 497090 436294 497158 436350
rect 497214 436294 497282 436350
rect 497338 436294 497406 436350
rect 497462 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 220554 436226
rect 220610 436170 220678 436226
rect 220734 436170 220802 436226
rect 220858 436170 220926 436226
rect 220982 436170 251274 436226
rect 251330 436170 251398 436226
rect 251454 436170 251522 436226
rect 251578 436170 251646 436226
rect 251702 436170 281994 436226
rect 282050 436170 282118 436226
rect 282174 436170 282242 436226
rect 282298 436170 282366 436226
rect 282422 436170 312714 436226
rect 312770 436170 312838 436226
rect 312894 436170 312962 436226
rect 313018 436170 313086 436226
rect 313142 436170 343434 436226
rect 343490 436170 343558 436226
rect 343614 436170 343682 436226
rect 343738 436170 343806 436226
rect 343862 436170 374154 436226
rect 374210 436170 374278 436226
rect 374334 436170 374402 436226
rect 374458 436170 374526 436226
rect 374582 436170 404874 436226
rect 404930 436170 404998 436226
rect 405054 436170 405122 436226
rect 405178 436170 405246 436226
rect 405302 436170 435594 436226
rect 435650 436170 435718 436226
rect 435774 436170 435842 436226
rect 435898 436170 435966 436226
rect 436022 436170 466314 436226
rect 466370 436170 466438 436226
rect 466494 436170 466562 436226
rect 466618 436170 466686 436226
rect 466742 436170 497034 436226
rect 497090 436170 497158 436226
rect 497214 436170 497282 436226
rect 497338 436170 497406 436226
rect 497462 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 220554 436102
rect 220610 436046 220678 436102
rect 220734 436046 220802 436102
rect 220858 436046 220926 436102
rect 220982 436046 251274 436102
rect 251330 436046 251398 436102
rect 251454 436046 251522 436102
rect 251578 436046 251646 436102
rect 251702 436046 281994 436102
rect 282050 436046 282118 436102
rect 282174 436046 282242 436102
rect 282298 436046 282366 436102
rect 282422 436046 312714 436102
rect 312770 436046 312838 436102
rect 312894 436046 312962 436102
rect 313018 436046 313086 436102
rect 313142 436046 343434 436102
rect 343490 436046 343558 436102
rect 343614 436046 343682 436102
rect 343738 436046 343806 436102
rect 343862 436046 374154 436102
rect 374210 436046 374278 436102
rect 374334 436046 374402 436102
rect 374458 436046 374526 436102
rect 374582 436046 404874 436102
rect 404930 436046 404998 436102
rect 405054 436046 405122 436102
rect 405178 436046 405246 436102
rect 405302 436046 435594 436102
rect 435650 436046 435718 436102
rect 435774 436046 435842 436102
rect 435898 436046 435966 436102
rect 436022 436046 466314 436102
rect 466370 436046 466438 436102
rect 466494 436046 466562 436102
rect 466618 436046 466686 436102
rect 466742 436046 497034 436102
rect 497090 436046 497158 436102
rect 497214 436046 497282 436102
rect 497338 436046 497406 436102
rect 497462 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 220554 435978
rect 220610 435922 220678 435978
rect 220734 435922 220802 435978
rect 220858 435922 220926 435978
rect 220982 435922 251274 435978
rect 251330 435922 251398 435978
rect 251454 435922 251522 435978
rect 251578 435922 251646 435978
rect 251702 435922 281994 435978
rect 282050 435922 282118 435978
rect 282174 435922 282242 435978
rect 282298 435922 282366 435978
rect 282422 435922 312714 435978
rect 312770 435922 312838 435978
rect 312894 435922 312962 435978
rect 313018 435922 313086 435978
rect 313142 435922 343434 435978
rect 343490 435922 343558 435978
rect 343614 435922 343682 435978
rect 343738 435922 343806 435978
rect 343862 435922 374154 435978
rect 374210 435922 374278 435978
rect 374334 435922 374402 435978
rect 374458 435922 374526 435978
rect 374582 435922 404874 435978
rect 404930 435922 404998 435978
rect 405054 435922 405122 435978
rect 405178 435922 405246 435978
rect 405302 435922 435594 435978
rect 435650 435922 435718 435978
rect 435774 435922 435842 435978
rect 435898 435922 435966 435978
rect 436022 435922 466314 435978
rect 466370 435922 466438 435978
rect 466494 435922 466562 435978
rect 466618 435922 466686 435978
rect 466742 435922 497034 435978
rect 497090 435922 497158 435978
rect 497214 435922 497282 435978
rect 497338 435922 497406 435978
rect 497462 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 193554 424350
rect 193610 424294 193678 424350
rect 193734 424294 193802 424350
rect 193858 424294 193926 424350
rect 193982 424294 224274 424350
rect 224330 424294 224398 424350
rect 224454 424294 224522 424350
rect 224578 424294 224646 424350
rect 224702 424294 254994 424350
rect 255050 424294 255118 424350
rect 255174 424294 255242 424350
rect 255298 424294 255366 424350
rect 255422 424294 285714 424350
rect 285770 424294 285838 424350
rect 285894 424294 285962 424350
rect 286018 424294 286086 424350
rect 286142 424294 316434 424350
rect 316490 424294 316558 424350
rect 316614 424294 316682 424350
rect 316738 424294 316806 424350
rect 316862 424294 347154 424350
rect 347210 424294 347278 424350
rect 347334 424294 347402 424350
rect 347458 424294 347526 424350
rect 347582 424294 377874 424350
rect 377930 424294 377998 424350
rect 378054 424294 378122 424350
rect 378178 424294 378246 424350
rect 378302 424294 408594 424350
rect 408650 424294 408718 424350
rect 408774 424294 408842 424350
rect 408898 424294 408966 424350
rect 409022 424294 439314 424350
rect 439370 424294 439438 424350
rect 439494 424294 439562 424350
rect 439618 424294 439686 424350
rect 439742 424294 470034 424350
rect 470090 424294 470158 424350
rect 470214 424294 470282 424350
rect 470338 424294 470406 424350
rect 470462 424294 500754 424350
rect 500810 424294 500878 424350
rect 500934 424294 501002 424350
rect 501058 424294 501126 424350
rect 501182 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 193554 424226
rect 193610 424170 193678 424226
rect 193734 424170 193802 424226
rect 193858 424170 193926 424226
rect 193982 424170 224274 424226
rect 224330 424170 224398 424226
rect 224454 424170 224522 424226
rect 224578 424170 224646 424226
rect 224702 424170 254994 424226
rect 255050 424170 255118 424226
rect 255174 424170 255242 424226
rect 255298 424170 255366 424226
rect 255422 424170 285714 424226
rect 285770 424170 285838 424226
rect 285894 424170 285962 424226
rect 286018 424170 286086 424226
rect 286142 424170 316434 424226
rect 316490 424170 316558 424226
rect 316614 424170 316682 424226
rect 316738 424170 316806 424226
rect 316862 424170 347154 424226
rect 347210 424170 347278 424226
rect 347334 424170 347402 424226
rect 347458 424170 347526 424226
rect 347582 424170 377874 424226
rect 377930 424170 377998 424226
rect 378054 424170 378122 424226
rect 378178 424170 378246 424226
rect 378302 424170 408594 424226
rect 408650 424170 408718 424226
rect 408774 424170 408842 424226
rect 408898 424170 408966 424226
rect 409022 424170 439314 424226
rect 439370 424170 439438 424226
rect 439494 424170 439562 424226
rect 439618 424170 439686 424226
rect 439742 424170 470034 424226
rect 470090 424170 470158 424226
rect 470214 424170 470282 424226
rect 470338 424170 470406 424226
rect 470462 424170 500754 424226
rect 500810 424170 500878 424226
rect 500934 424170 501002 424226
rect 501058 424170 501126 424226
rect 501182 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 193554 424102
rect 193610 424046 193678 424102
rect 193734 424046 193802 424102
rect 193858 424046 193926 424102
rect 193982 424046 224274 424102
rect 224330 424046 224398 424102
rect 224454 424046 224522 424102
rect 224578 424046 224646 424102
rect 224702 424046 254994 424102
rect 255050 424046 255118 424102
rect 255174 424046 255242 424102
rect 255298 424046 255366 424102
rect 255422 424046 285714 424102
rect 285770 424046 285838 424102
rect 285894 424046 285962 424102
rect 286018 424046 286086 424102
rect 286142 424046 316434 424102
rect 316490 424046 316558 424102
rect 316614 424046 316682 424102
rect 316738 424046 316806 424102
rect 316862 424046 347154 424102
rect 347210 424046 347278 424102
rect 347334 424046 347402 424102
rect 347458 424046 347526 424102
rect 347582 424046 377874 424102
rect 377930 424046 377998 424102
rect 378054 424046 378122 424102
rect 378178 424046 378246 424102
rect 378302 424046 408594 424102
rect 408650 424046 408718 424102
rect 408774 424046 408842 424102
rect 408898 424046 408966 424102
rect 409022 424046 439314 424102
rect 439370 424046 439438 424102
rect 439494 424046 439562 424102
rect 439618 424046 439686 424102
rect 439742 424046 470034 424102
rect 470090 424046 470158 424102
rect 470214 424046 470282 424102
rect 470338 424046 470406 424102
rect 470462 424046 500754 424102
rect 500810 424046 500878 424102
rect 500934 424046 501002 424102
rect 501058 424046 501126 424102
rect 501182 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 193554 423978
rect 193610 423922 193678 423978
rect 193734 423922 193802 423978
rect 193858 423922 193926 423978
rect 193982 423922 224274 423978
rect 224330 423922 224398 423978
rect 224454 423922 224522 423978
rect 224578 423922 224646 423978
rect 224702 423922 254994 423978
rect 255050 423922 255118 423978
rect 255174 423922 255242 423978
rect 255298 423922 255366 423978
rect 255422 423922 285714 423978
rect 285770 423922 285838 423978
rect 285894 423922 285962 423978
rect 286018 423922 286086 423978
rect 286142 423922 316434 423978
rect 316490 423922 316558 423978
rect 316614 423922 316682 423978
rect 316738 423922 316806 423978
rect 316862 423922 347154 423978
rect 347210 423922 347278 423978
rect 347334 423922 347402 423978
rect 347458 423922 347526 423978
rect 347582 423922 377874 423978
rect 377930 423922 377998 423978
rect 378054 423922 378122 423978
rect 378178 423922 378246 423978
rect 378302 423922 408594 423978
rect 408650 423922 408718 423978
rect 408774 423922 408842 423978
rect 408898 423922 408966 423978
rect 409022 423922 439314 423978
rect 439370 423922 439438 423978
rect 439494 423922 439562 423978
rect 439618 423922 439686 423978
rect 439742 423922 470034 423978
rect 470090 423922 470158 423978
rect 470214 423922 470282 423978
rect 470338 423922 470406 423978
rect 470462 423922 500754 423978
rect 500810 423922 500878 423978
rect 500934 423922 501002 423978
rect 501058 423922 501126 423978
rect 501182 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 220554 418350
rect 220610 418294 220678 418350
rect 220734 418294 220802 418350
rect 220858 418294 220926 418350
rect 220982 418294 251274 418350
rect 251330 418294 251398 418350
rect 251454 418294 251522 418350
rect 251578 418294 251646 418350
rect 251702 418294 281994 418350
rect 282050 418294 282118 418350
rect 282174 418294 282242 418350
rect 282298 418294 282366 418350
rect 282422 418294 312714 418350
rect 312770 418294 312838 418350
rect 312894 418294 312962 418350
rect 313018 418294 313086 418350
rect 313142 418294 343434 418350
rect 343490 418294 343558 418350
rect 343614 418294 343682 418350
rect 343738 418294 343806 418350
rect 343862 418294 374154 418350
rect 374210 418294 374278 418350
rect 374334 418294 374402 418350
rect 374458 418294 374526 418350
rect 374582 418294 404874 418350
rect 404930 418294 404998 418350
rect 405054 418294 405122 418350
rect 405178 418294 405246 418350
rect 405302 418294 435594 418350
rect 435650 418294 435718 418350
rect 435774 418294 435842 418350
rect 435898 418294 435966 418350
rect 436022 418294 466314 418350
rect 466370 418294 466438 418350
rect 466494 418294 466562 418350
rect 466618 418294 466686 418350
rect 466742 418294 497034 418350
rect 497090 418294 497158 418350
rect 497214 418294 497282 418350
rect 497338 418294 497406 418350
rect 497462 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 220554 418226
rect 220610 418170 220678 418226
rect 220734 418170 220802 418226
rect 220858 418170 220926 418226
rect 220982 418170 251274 418226
rect 251330 418170 251398 418226
rect 251454 418170 251522 418226
rect 251578 418170 251646 418226
rect 251702 418170 281994 418226
rect 282050 418170 282118 418226
rect 282174 418170 282242 418226
rect 282298 418170 282366 418226
rect 282422 418170 312714 418226
rect 312770 418170 312838 418226
rect 312894 418170 312962 418226
rect 313018 418170 313086 418226
rect 313142 418170 343434 418226
rect 343490 418170 343558 418226
rect 343614 418170 343682 418226
rect 343738 418170 343806 418226
rect 343862 418170 374154 418226
rect 374210 418170 374278 418226
rect 374334 418170 374402 418226
rect 374458 418170 374526 418226
rect 374582 418170 404874 418226
rect 404930 418170 404998 418226
rect 405054 418170 405122 418226
rect 405178 418170 405246 418226
rect 405302 418170 435594 418226
rect 435650 418170 435718 418226
rect 435774 418170 435842 418226
rect 435898 418170 435966 418226
rect 436022 418170 466314 418226
rect 466370 418170 466438 418226
rect 466494 418170 466562 418226
rect 466618 418170 466686 418226
rect 466742 418170 497034 418226
rect 497090 418170 497158 418226
rect 497214 418170 497282 418226
rect 497338 418170 497406 418226
rect 497462 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 220554 418102
rect 220610 418046 220678 418102
rect 220734 418046 220802 418102
rect 220858 418046 220926 418102
rect 220982 418046 251274 418102
rect 251330 418046 251398 418102
rect 251454 418046 251522 418102
rect 251578 418046 251646 418102
rect 251702 418046 281994 418102
rect 282050 418046 282118 418102
rect 282174 418046 282242 418102
rect 282298 418046 282366 418102
rect 282422 418046 312714 418102
rect 312770 418046 312838 418102
rect 312894 418046 312962 418102
rect 313018 418046 313086 418102
rect 313142 418046 343434 418102
rect 343490 418046 343558 418102
rect 343614 418046 343682 418102
rect 343738 418046 343806 418102
rect 343862 418046 374154 418102
rect 374210 418046 374278 418102
rect 374334 418046 374402 418102
rect 374458 418046 374526 418102
rect 374582 418046 404874 418102
rect 404930 418046 404998 418102
rect 405054 418046 405122 418102
rect 405178 418046 405246 418102
rect 405302 418046 435594 418102
rect 435650 418046 435718 418102
rect 435774 418046 435842 418102
rect 435898 418046 435966 418102
rect 436022 418046 466314 418102
rect 466370 418046 466438 418102
rect 466494 418046 466562 418102
rect 466618 418046 466686 418102
rect 466742 418046 497034 418102
rect 497090 418046 497158 418102
rect 497214 418046 497282 418102
rect 497338 418046 497406 418102
rect 497462 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 220554 417978
rect 220610 417922 220678 417978
rect 220734 417922 220802 417978
rect 220858 417922 220926 417978
rect 220982 417922 251274 417978
rect 251330 417922 251398 417978
rect 251454 417922 251522 417978
rect 251578 417922 251646 417978
rect 251702 417922 281994 417978
rect 282050 417922 282118 417978
rect 282174 417922 282242 417978
rect 282298 417922 282366 417978
rect 282422 417922 312714 417978
rect 312770 417922 312838 417978
rect 312894 417922 312962 417978
rect 313018 417922 313086 417978
rect 313142 417922 343434 417978
rect 343490 417922 343558 417978
rect 343614 417922 343682 417978
rect 343738 417922 343806 417978
rect 343862 417922 374154 417978
rect 374210 417922 374278 417978
rect 374334 417922 374402 417978
rect 374458 417922 374526 417978
rect 374582 417922 404874 417978
rect 404930 417922 404998 417978
rect 405054 417922 405122 417978
rect 405178 417922 405246 417978
rect 405302 417922 435594 417978
rect 435650 417922 435718 417978
rect 435774 417922 435842 417978
rect 435898 417922 435966 417978
rect 436022 417922 466314 417978
rect 466370 417922 466438 417978
rect 466494 417922 466562 417978
rect 466618 417922 466686 417978
rect 466742 417922 497034 417978
rect 497090 417922 497158 417978
rect 497214 417922 497282 417978
rect 497338 417922 497406 417978
rect 497462 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 377874 406350
rect 377930 406294 377998 406350
rect 378054 406294 378122 406350
rect 378178 406294 378246 406350
rect 378302 406294 408594 406350
rect 408650 406294 408718 406350
rect 408774 406294 408842 406350
rect 408898 406294 408966 406350
rect 409022 406294 439314 406350
rect 439370 406294 439438 406350
rect 439494 406294 439562 406350
rect 439618 406294 439686 406350
rect 439742 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 500754 406350
rect 500810 406294 500878 406350
rect 500934 406294 501002 406350
rect 501058 406294 501126 406350
rect 501182 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 377874 406226
rect 377930 406170 377998 406226
rect 378054 406170 378122 406226
rect 378178 406170 378246 406226
rect 378302 406170 408594 406226
rect 408650 406170 408718 406226
rect 408774 406170 408842 406226
rect 408898 406170 408966 406226
rect 409022 406170 439314 406226
rect 439370 406170 439438 406226
rect 439494 406170 439562 406226
rect 439618 406170 439686 406226
rect 439742 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 500754 406226
rect 500810 406170 500878 406226
rect 500934 406170 501002 406226
rect 501058 406170 501126 406226
rect 501182 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 377874 406102
rect 377930 406046 377998 406102
rect 378054 406046 378122 406102
rect 378178 406046 378246 406102
rect 378302 406046 408594 406102
rect 408650 406046 408718 406102
rect 408774 406046 408842 406102
rect 408898 406046 408966 406102
rect 409022 406046 439314 406102
rect 439370 406046 439438 406102
rect 439494 406046 439562 406102
rect 439618 406046 439686 406102
rect 439742 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 500754 406102
rect 500810 406046 500878 406102
rect 500934 406046 501002 406102
rect 501058 406046 501126 406102
rect 501182 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 377874 405978
rect 377930 405922 377998 405978
rect 378054 405922 378122 405978
rect 378178 405922 378246 405978
rect 378302 405922 408594 405978
rect 408650 405922 408718 405978
rect 408774 405922 408842 405978
rect 408898 405922 408966 405978
rect 409022 405922 439314 405978
rect 439370 405922 439438 405978
rect 439494 405922 439562 405978
rect 439618 405922 439686 405978
rect 439742 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 500754 405978
rect 500810 405922 500878 405978
rect 500934 405922 501002 405978
rect 501058 405922 501126 405978
rect 501182 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 374154 400350
rect 374210 400294 374278 400350
rect 374334 400294 374402 400350
rect 374458 400294 374526 400350
rect 374582 400294 404874 400350
rect 404930 400294 404998 400350
rect 405054 400294 405122 400350
rect 405178 400294 405246 400350
rect 405302 400294 435594 400350
rect 435650 400294 435718 400350
rect 435774 400294 435842 400350
rect 435898 400294 435966 400350
rect 436022 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 497034 400350
rect 497090 400294 497158 400350
rect 497214 400294 497282 400350
rect 497338 400294 497406 400350
rect 497462 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 374154 400226
rect 374210 400170 374278 400226
rect 374334 400170 374402 400226
rect 374458 400170 374526 400226
rect 374582 400170 404874 400226
rect 404930 400170 404998 400226
rect 405054 400170 405122 400226
rect 405178 400170 405246 400226
rect 405302 400170 435594 400226
rect 435650 400170 435718 400226
rect 435774 400170 435842 400226
rect 435898 400170 435966 400226
rect 436022 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 497034 400226
rect 497090 400170 497158 400226
rect 497214 400170 497282 400226
rect 497338 400170 497406 400226
rect 497462 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 374154 400102
rect 374210 400046 374278 400102
rect 374334 400046 374402 400102
rect 374458 400046 374526 400102
rect 374582 400046 404874 400102
rect 404930 400046 404998 400102
rect 405054 400046 405122 400102
rect 405178 400046 405246 400102
rect 405302 400046 435594 400102
rect 435650 400046 435718 400102
rect 435774 400046 435842 400102
rect 435898 400046 435966 400102
rect 436022 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 497034 400102
rect 497090 400046 497158 400102
rect 497214 400046 497282 400102
rect 497338 400046 497406 400102
rect 497462 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 374154 399978
rect 374210 399922 374278 399978
rect 374334 399922 374402 399978
rect 374458 399922 374526 399978
rect 374582 399922 404874 399978
rect 404930 399922 404998 399978
rect 405054 399922 405122 399978
rect 405178 399922 405246 399978
rect 405302 399922 435594 399978
rect 435650 399922 435718 399978
rect 435774 399922 435842 399978
rect 435898 399922 435966 399978
rect 436022 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 497034 399978
rect 497090 399922 497158 399978
rect 497214 399922 497282 399978
rect 497338 399922 497406 399978
rect 497462 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 377874 388350
rect 377930 388294 377998 388350
rect 378054 388294 378122 388350
rect 378178 388294 378246 388350
rect 378302 388294 408594 388350
rect 408650 388294 408718 388350
rect 408774 388294 408842 388350
rect 408898 388294 408966 388350
rect 409022 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 470034 388350
rect 470090 388294 470158 388350
rect 470214 388294 470282 388350
rect 470338 388294 470406 388350
rect 470462 388294 500754 388350
rect 500810 388294 500878 388350
rect 500934 388294 501002 388350
rect 501058 388294 501126 388350
rect 501182 388294 531474 388350
rect 531530 388294 531598 388350
rect 531654 388294 531722 388350
rect 531778 388294 531846 388350
rect 531902 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 377874 388226
rect 377930 388170 377998 388226
rect 378054 388170 378122 388226
rect 378178 388170 378246 388226
rect 378302 388170 408594 388226
rect 408650 388170 408718 388226
rect 408774 388170 408842 388226
rect 408898 388170 408966 388226
rect 409022 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 470034 388226
rect 470090 388170 470158 388226
rect 470214 388170 470282 388226
rect 470338 388170 470406 388226
rect 470462 388170 500754 388226
rect 500810 388170 500878 388226
rect 500934 388170 501002 388226
rect 501058 388170 501126 388226
rect 501182 388170 531474 388226
rect 531530 388170 531598 388226
rect 531654 388170 531722 388226
rect 531778 388170 531846 388226
rect 531902 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 377874 388102
rect 377930 388046 377998 388102
rect 378054 388046 378122 388102
rect 378178 388046 378246 388102
rect 378302 388046 408594 388102
rect 408650 388046 408718 388102
rect 408774 388046 408842 388102
rect 408898 388046 408966 388102
rect 409022 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 470034 388102
rect 470090 388046 470158 388102
rect 470214 388046 470282 388102
rect 470338 388046 470406 388102
rect 470462 388046 500754 388102
rect 500810 388046 500878 388102
rect 500934 388046 501002 388102
rect 501058 388046 501126 388102
rect 501182 388046 531474 388102
rect 531530 388046 531598 388102
rect 531654 388046 531722 388102
rect 531778 388046 531846 388102
rect 531902 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 377874 387978
rect 377930 387922 377998 387978
rect 378054 387922 378122 387978
rect 378178 387922 378246 387978
rect 378302 387922 408594 387978
rect 408650 387922 408718 387978
rect 408774 387922 408842 387978
rect 408898 387922 408966 387978
rect 409022 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 470034 387978
rect 470090 387922 470158 387978
rect 470214 387922 470282 387978
rect 470338 387922 470406 387978
rect 470462 387922 500754 387978
rect 500810 387922 500878 387978
rect 500934 387922 501002 387978
rect 501058 387922 501126 387978
rect 501182 387922 531474 387978
rect 531530 387922 531598 387978
rect 531654 387922 531722 387978
rect 531778 387922 531846 387978
rect 531902 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 374154 382350
rect 374210 382294 374278 382350
rect 374334 382294 374402 382350
rect 374458 382294 374526 382350
rect 374582 382294 404874 382350
rect 404930 382294 404998 382350
rect 405054 382294 405122 382350
rect 405178 382294 405246 382350
rect 405302 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 466314 382350
rect 466370 382294 466438 382350
rect 466494 382294 466562 382350
rect 466618 382294 466686 382350
rect 466742 382294 497034 382350
rect 497090 382294 497158 382350
rect 497214 382294 497282 382350
rect 497338 382294 497406 382350
rect 497462 382294 527754 382350
rect 527810 382294 527878 382350
rect 527934 382294 528002 382350
rect 528058 382294 528126 382350
rect 528182 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 374154 382226
rect 374210 382170 374278 382226
rect 374334 382170 374402 382226
rect 374458 382170 374526 382226
rect 374582 382170 404874 382226
rect 404930 382170 404998 382226
rect 405054 382170 405122 382226
rect 405178 382170 405246 382226
rect 405302 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 466314 382226
rect 466370 382170 466438 382226
rect 466494 382170 466562 382226
rect 466618 382170 466686 382226
rect 466742 382170 497034 382226
rect 497090 382170 497158 382226
rect 497214 382170 497282 382226
rect 497338 382170 497406 382226
rect 497462 382170 527754 382226
rect 527810 382170 527878 382226
rect 527934 382170 528002 382226
rect 528058 382170 528126 382226
rect 528182 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 374154 382102
rect 374210 382046 374278 382102
rect 374334 382046 374402 382102
rect 374458 382046 374526 382102
rect 374582 382046 404874 382102
rect 404930 382046 404998 382102
rect 405054 382046 405122 382102
rect 405178 382046 405246 382102
rect 405302 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 466314 382102
rect 466370 382046 466438 382102
rect 466494 382046 466562 382102
rect 466618 382046 466686 382102
rect 466742 382046 497034 382102
rect 497090 382046 497158 382102
rect 497214 382046 497282 382102
rect 497338 382046 497406 382102
rect 497462 382046 527754 382102
rect 527810 382046 527878 382102
rect 527934 382046 528002 382102
rect 528058 382046 528126 382102
rect 528182 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 374154 381978
rect 374210 381922 374278 381978
rect 374334 381922 374402 381978
rect 374458 381922 374526 381978
rect 374582 381922 404874 381978
rect 404930 381922 404998 381978
rect 405054 381922 405122 381978
rect 405178 381922 405246 381978
rect 405302 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 466314 381978
rect 466370 381922 466438 381978
rect 466494 381922 466562 381978
rect 466618 381922 466686 381978
rect 466742 381922 497034 381978
rect 497090 381922 497158 381978
rect 497214 381922 497282 381978
rect 497338 381922 497406 381978
rect 497462 381922 527754 381978
rect 527810 381922 527878 381978
rect 527934 381922 528002 381978
rect 528058 381922 528126 381978
rect 528182 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 254994 370350
rect 255050 370294 255118 370350
rect 255174 370294 255242 370350
rect 255298 370294 255366 370350
rect 255422 370294 285714 370350
rect 285770 370294 285838 370350
rect 285894 370294 285962 370350
rect 286018 370294 286086 370350
rect 286142 370294 316434 370350
rect 316490 370294 316558 370350
rect 316614 370294 316682 370350
rect 316738 370294 316806 370350
rect 316862 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 377874 370350
rect 377930 370294 377998 370350
rect 378054 370294 378122 370350
rect 378178 370294 378246 370350
rect 378302 370294 408594 370350
rect 408650 370294 408718 370350
rect 408774 370294 408842 370350
rect 408898 370294 408966 370350
rect 409022 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 470034 370350
rect 470090 370294 470158 370350
rect 470214 370294 470282 370350
rect 470338 370294 470406 370350
rect 470462 370294 500754 370350
rect 500810 370294 500878 370350
rect 500934 370294 501002 370350
rect 501058 370294 501126 370350
rect 501182 370294 531474 370350
rect 531530 370294 531598 370350
rect 531654 370294 531722 370350
rect 531778 370294 531846 370350
rect 531902 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 254994 370226
rect 255050 370170 255118 370226
rect 255174 370170 255242 370226
rect 255298 370170 255366 370226
rect 255422 370170 285714 370226
rect 285770 370170 285838 370226
rect 285894 370170 285962 370226
rect 286018 370170 286086 370226
rect 286142 370170 316434 370226
rect 316490 370170 316558 370226
rect 316614 370170 316682 370226
rect 316738 370170 316806 370226
rect 316862 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 377874 370226
rect 377930 370170 377998 370226
rect 378054 370170 378122 370226
rect 378178 370170 378246 370226
rect 378302 370170 408594 370226
rect 408650 370170 408718 370226
rect 408774 370170 408842 370226
rect 408898 370170 408966 370226
rect 409022 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 470034 370226
rect 470090 370170 470158 370226
rect 470214 370170 470282 370226
rect 470338 370170 470406 370226
rect 470462 370170 500754 370226
rect 500810 370170 500878 370226
rect 500934 370170 501002 370226
rect 501058 370170 501126 370226
rect 501182 370170 531474 370226
rect 531530 370170 531598 370226
rect 531654 370170 531722 370226
rect 531778 370170 531846 370226
rect 531902 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 254994 370102
rect 255050 370046 255118 370102
rect 255174 370046 255242 370102
rect 255298 370046 255366 370102
rect 255422 370046 285714 370102
rect 285770 370046 285838 370102
rect 285894 370046 285962 370102
rect 286018 370046 286086 370102
rect 286142 370046 316434 370102
rect 316490 370046 316558 370102
rect 316614 370046 316682 370102
rect 316738 370046 316806 370102
rect 316862 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 377874 370102
rect 377930 370046 377998 370102
rect 378054 370046 378122 370102
rect 378178 370046 378246 370102
rect 378302 370046 408594 370102
rect 408650 370046 408718 370102
rect 408774 370046 408842 370102
rect 408898 370046 408966 370102
rect 409022 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 470034 370102
rect 470090 370046 470158 370102
rect 470214 370046 470282 370102
rect 470338 370046 470406 370102
rect 470462 370046 500754 370102
rect 500810 370046 500878 370102
rect 500934 370046 501002 370102
rect 501058 370046 501126 370102
rect 501182 370046 531474 370102
rect 531530 370046 531598 370102
rect 531654 370046 531722 370102
rect 531778 370046 531846 370102
rect 531902 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 254994 369978
rect 255050 369922 255118 369978
rect 255174 369922 255242 369978
rect 255298 369922 255366 369978
rect 255422 369922 285714 369978
rect 285770 369922 285838 369978
rect 285894 369922 285962 369978
rect 286018 369922 286086 369978
rect 286142 369922 316434 369978
rect 316490 369922 316558 369978
rect 316614 369922 316682 369978
rect 316738 369922 316806 369978
rect 316862 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 377874 369978
rect 377930 369922 377998 369978
rect 378054 369922 378122 369978
rect 378178 369922 378246 369978
rect 378302 369922 408594 369978
rect 408650 369922 408718 369978
rect 408774 369922 408842 369978
rect 408898 369922 408966 369978
rect 409022 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 470034 369978
rect 470090 369922 470158 369978
rect 470214 369922 470282 369978
rect 470338 369922 470406 369978
rect 470462 369922 500754 369978
rect 500810 369922 500878 369978
rect 500934 369922 501002 369978
rect 501058 369922 501126 369978
rect 501182 369922 531474 369978
rect 531530 369922 531598 369978
rect 531654 369922 531722 369978
rect 531778 369922 531846 369978
rect 531902 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect 59708 368758 584740 368774
rect 59708 368702 59724 368758
rect 59780 368702 584668 368758
rect 584724 368702 584740 368758
rect 59708 368686 584740 368702
rect 171260 366778 202484 366794
rect 171260 366722 171276 366778
rect 171332 366722 202412 366778
rect 202468 366722 202484 366778
rect 171260 366706 202484 366722
rect 110108 366598 202148 366614
rect 110108 366542 110124 366598
rect 110180 366542 202076 366598
rect 202132 366542 202148 366598
rect 110108 366526 202148 366542
rect 2924 366418 201924 366434
rect 2924 366362 2940 366418
rect 2996 366362 201852 366418
rect 201908 366362 201924 366418
rect 2924 366346 201924 366362
rect 109100 365158 160820 365174
rect 109100 365102 109116 365158
rect 109172 365102 160748 365158
rect 160804 365102 160820 365158
rect 109100 365086 160820 365102
rect 119180 364978 164740 364994
rect 119180 364922 119196 364978
rect 119252 364922 164668 364978
rect 164724 364922 164740 364978
rect 119180 364906 164740 364922
rect 156140 364798 204164 364814
rect 156140 364742 156156 364798
rect 156212 364742 204092 364798
rect 204148 364742 204164 364798
rect 156140 364726 204164 364742
rect 157820 364618 205956 364634
rect 157820 364562 157836 364618
rect 157892 364562 205884 364618
rect 205940 364562 205956 364618
rect 157820 364546 205956 364562
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 220554 364350
rect 220610 364294 220678 364350
rect 220734 364294 220802 364350
rect 220858 364294 220926 364350
rect 220982 364294 251274 364350
rect 251330 364294 251398 364350
rect 251454 364294 251522 364350
rect 251578 364294 251646 364350
rect 251702 364294 281994 364350
rect 282050 364294 282118 364350
rect 282174 364294 282242 364350
rect 282298 364294 282366 364350
rect 282422 364294 312714 364350
rect 312770 364294 312838 364350
rect 312894 364294 312962 364350
rect 313018 364294 313086 364350
rect 313142 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 374154 364350
rect 374210 364294 374278 364350
rect 374334 364294 374402 364350
rect 374458 364294 374526 364350
rect 374582 364294 404874 364350
rect 404930 364294 404998 364350
rect 405054 364294 405122 364350
rect 405178 364294 405246 364350
rect 405302 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 466314 364350
rect 466370 364294 466438 364350
rect 466494 364294 466562 364350
rect 466618 364294 466686 364350
rect 466742 364294 497034 364350
rect 497090 364294 497158 364350
rect 497214 364294 497282 364350
rect 497338 364294 497406 364350
rect 497462 364294 527754 364350
rect 527810 364294 527878 364350
rect 527934 364294 528002 364350
rect 528058 364294 528126 364350
rect 528182 364294 558474 364350
rect 558530 364294 558598 364350
rect 558654 364294 558722 364350
rect 558778 364294 558846 364350
rect 558902 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 220554 364226
rect 220610 364170 220678 364226
rect 220734 364170 220802 364226
rect 220858 364170 220926 364226
rect 220982 364170 251274 364226
rect 251330 364170 251398 364226
rect 251454 364170 251522 364226
rect 251578 364170 251646 364226
rect 251702 364170 281994 364226
rect 282050 364170 282118 364226
rect 282174 364170 282242 364226
rect 282298 364170 282366 364226
rect 282422 364170 312714 364226
rect 312770 364170 312838 364226
rect 312894 364170 312962 364226
rect 313018 364170 313086 364226
rect 313142 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 374154 364226
rect 374210 364170 374278 364226
rect 374334 364170 374402 364226
rect 374458 364170 374526 364226
rect 374582 364170 404874 364226
rect 404930 364170 404998 364226
rect 405054 364170 405122 364226
rect 405178 364170 405246 364226
rect 405302 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 466314 364226
rect 466370 364170 466438 364226
rect 466494 364170 466562 364226
rect 466618 364170 466686 364226
rect 466742 364170 497034 364226
rect 497090 364170 497158 364226
rect 497214 364170 497282 364226
rect 497338 364170 497406 364226
rect 497462 364170 527754 364226
rect 527810 364170 527878 364226
rect 527934 364170 528002 364226
rect 528058 364170 528126 364226
rect 528182 364170 558474 364226
rect 558530 364170 558598 364226
rect 558654 364170 558722 364226
rect 558778 364170 558846 364226
rect 558902 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 220554 364102
rect 220610 364046 220678 364102
rect 220734 364046 220802 364102
rect 220858 364046 220926 364102
rect 220982 364046 251274 364102
rect 251330 364046 251398 364102
rect 251454 364046 251522 364102
rect 251578 364046 251646 364102
rect 251702 364046 281994 364102
rect 282050 364046 282118 364102
rect 282174 364046 282242 364102
rect 282298 364046 282366 364102
rect 282422 364046 312714 364102
rect 312770 364046 312838 364102
rect 312894 364046 312962 364102
rect 313018 364046 313086 364102
rect 313142 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 374154 364102
rect 374210 364046 374278 364102
rect 374334 364046 374402 364102
rect 374458 364046 374526 364102
rect 374582 364046 404874 364102
rect 404930 364046 404998 364102
rect 405054 364046 405122 364102
rect 405178 364046 405246 364102
rect 405302 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 466314 364102
rect 466370 364046 466438 364102
rect 466494 364046 466562 364102
rect 466618 364046 466686 364102
rect 466742 364046 497034 364102
rect 497090 364046 497158 364102
rect 497214 364046 497282 364102
rect 497338 364046 497406 364102
rect 497462 364046 527754 364102
rect 527810 364046 527878 364102
rect 527934 364046 528002 364102
rect 528058 364046 528126 364102
rect 528182 364046 558474 364102
rect 558530 364046 558598 364102
rect 558654 364046 558722 364102
rect 558778 364046 558846 364102
rect 558902 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 220554 363978
rect 220610 363922 220678 363978
rect 220734 363922 220802 363978
rect 220858 363922 220926 363978
rect 220982 363922 251274 363978
rect 251330 363922 251398 363978
rect 251454 363922 251522 363978
rect 251578 363922 251646 363978
rect 251702 363922 281994 363978
rect 282050 363922 282118 363978
rect 282174 363922 282242 363978
rect 282298 363922 282366 363978
rect 282422 363922 312714 363978
rect 312770 363922 312838 363978
rect 312894 363922 312962 363978
rect 313018 363922 313086 363978
rect 313142 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 374154 363978
rect 374210 363922 374278 363978
rect 374334 363922 374402 363978
rect 374458 363922 374526 363978
rect 374582 363922 404874 363978
rect 404930 363922 404998 363978
rect 405054 363922 405122 363978
rect 405178 363922 405246 363978
rect 405302 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 466314 363978
rect 466370 363922 466438 363978
rect 466494 363922 466562 363978
rect 466618 363922 466686 363978
rect 466742 363922 497034 363978
rect 497090 363922 497158 363978
rect 497214 363922 497282 363978
rect 497338 363922 497406 363978
rect 497462 363922 527754 363978
rect 527810 363922 527878 363978
rect 527934 363922 528002 363978
rect 528058 363922 528126 363978
rect 528182 363922 558474 363978
rect 558530 363922 558598 363978
rect 558654 363922 558722 363978
rect 558778 363922 558846 363978
rect 558902 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect 151324 363178 206180 363194
rect 151324 363122 151340 363178
rect 151396 363122 206108 363178
rect 206164 363122 206180 363178
rect 151324 363106 206180 363122
rect 151996 362998 212340 363014
rect 151996 362942 152012 362998
rect 152068 362942 212268 362998
rect 212324 362942 212340 362998
rect 151996 362926 212340 362942
rect 117500 362278 163508 362294
rect 117500 362222 117516 362278
rect 117572 362222 163436 362278
rect 163492 362222 163508 362278
rect 117500 362206 163508 362222
rect 150652 362098 207524 362114
rect 150652 362042 150668 362098
rect 150724 362042 207452 362098
rect 207508 362042 207524 362098
rect 150652 362026 207524 362042
rect 161404 361558 209204 361574
rect 161404 361502 161420 361558
rect 161476 361502 209132 361558
rect 209188 361502 209204 361558
rect 161404 361486 209204 361502
rect 1580 361378 202036 361394
rect 1580 361322 1596 361378
rect 1652 361322 201964 361378
rect 202020 361322 202036 361378
rect 1580 361306 202036 361322
rect 173500 360298 194868 360314
rect 173500 360242 173516 360298
rect 173572 360242 194796 360298
rect 194852 360242 194868 360298
rect 173500 360226 194868 360242
rect 110220 360118 199348 360134
rect 110220 360062 110236 360118
rect 110292 360062 199348 360118
rect 110220 360046 199348 360062
rect 112348 359938 199124 359954
rect 112348 359882 112364 359938
rect 112420 359882 199124 359938
rect 112348 359866 199124 359882
rect 190972 359758 195988 359774
rect 190972 359702 190988 359758
rect 191044 359702 195916 359758
rect 195972 359702 195988 359758
rect 190972 359686 195988 359702
rect 190748 359578 196548 359594
rect 190748 359522 190764 359578
rect 190820 359522 196476 359578
rect 196532 359522 196548 359578
rect 190748 359506 196548 359522
rect 199036 359414 199124 359866
rect 199260 359578 199348 360046
rect 199260 359522 199276 359578
rect 199332 359522 199348 359578
rect 199260 359506 199348 359522
rect 199484 359578 202260 359594
rect 199484 359522 202188 359578
rect 202244 359522 202260 359578
rect 199484 359506 202260 359522
rect 199484 359414 199572 359506
rect 199036 359326 199572 359414
rect 182236 359038 205172 359054
rect 182236 358982 182252 359038
rect 182308 358982 205100 359038
rect 205156 358982 205172 359038
rect 182236 358966 205172 358982
rect 189516 358858 212116 358874
rect 189516 358802 189532 358858
rect 189588 358802 212044 358858
rect 212100 358802 212116 358858
rect 189516 358786 212116 358802
rect 166108 358678 205844 358694
rect 166108 358622 166124 358678
rect 166180 358622 205772 358678
rect 205828 358622 205844 358678
rect 166108 358606 205844 358622
rect 110332 357958 199460 357974
rect 110332 357902 110348 357958
rect 110404 357902 199388 357958
rect 199444 357902 199460 357958
rect 110332 357886 199460 357902
rect 108428 357598 191564 357614
rect 108428 357542 108444 357598
rect 108500 357542 191564 357598
rect 108428 357526 191564 357542
rect 196460 357598 203324 357614
rect 196460 357542 196476 357598
rect 196532 357542 203324 357598
rect 196460 357526 203324 357542
rect 191476 357254 191564 357526
rect 203236 357434 203324 357526
rect 192988 357418 199572 357434
rect 192988 357362 193004 357418
rect 193060 357362 199572 357418
rect 192988 357346 199572 357362
rect 203236 357418 205060 357434
rect 203236 357362 204988 357418
rect 205044 357362 205060 357418
rect 203236 357346 205060 357362
rect 199484 357254 199572 357346
rect 191476 357238 199348 357254
rect 191476 357182 199276 357238
rect 199332 357182 199348 357238
rect 191476 357166 199348 357182
rect 199484 357238 208420 357254
rect 199484 357182 208348 357238
rect 208404 357182 208420 357238
rect 199484 357166 208420 357182
rect 186940 357058 208532 357074
rect 186940 357002 186956 357058
rect 187012 357002 208460 357058
rect 208516 357002 208532 357058
rect 186940 356986 208532 357002
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 149222 352350
rect 149278 352294 149346 352350
rect 149402 352294 179942 352350
rect 179998 352294 180066 352350
rect 180122 352294 224274 352350
rect 224330 352294 224398 352350
rect 224454 352294 224522 352350
rect 224578 352294 224646 352350
rect 224702 352294 254994 352350
rect 255050 352294 255118 352350
rect 255174 352294 255242 352350
rect 255298 352294 255366 352350
rect 255422 352294 285714 352350
rect 285770 352294 285838 352350
rect 285894 352294 285962 352350
rect 286018 352294 286086 352350
rect 286142 352294 316434 352350
rect 316490 352294 316558 352350
rect 316614 352294 316682 352350
rect 316738 352294 316806 352350
rect 316862 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 377874 352350
rect 377930 352294 377998 352350
rect 378054 352294 378122 352350
rect 378178 352294 378246 352350
rect 378302 352294 408594 352350
rect 408650 352294 408718 352350
rect 408774 352294 408842 352350
rect 408898 352294 408966 352350
rect 409022 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 470034 352350
rect 470090 352294 470158 352350
rect 470214 352294 470282 352350
rect 470338 352294 470406 352350
rect 470462 352294 500754 352350
rect 500810 352294 500878 352350
rect 500934 352294 501002 352350
rect 501058 352294 501126 352350
rect 501182 352294 531474 352350
rect 531530 352294 531598 352350
rect 531654 352294 531722 352350
rect 531778 352294 531846 352350
rect 531902 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 149222 352226
rect 149278 352170 149346 352226
rect 149402 352170 179942 352226
rect 179998 352170 180066 352226
rect 180122 352170 224274 352226
rect 224330 352170 224398 352226
rect 224454 352170 224522 352226
rect 224578 352170 224646 352226
rect 224702 352170 254994 352226
rect 255050 352170 255118 352226
rect 255174 352170 255242 352226
rect 255298 352170 255366 352226
rect 255422 352170 285714 352226
rect 285770 352170 285838 352226
rect 285894 352170 285962 352226
rect 286018 352170 286086 352226
rect 286142 352170 316434 352226
rect 316490 352170 316558 352226
rect 316614 352170 316682 352226
rect 316738 352170 316806 352226
rect 316862 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 377874 352226
rect 377930 352170 377998 352226
rect 378054 352170 378122 352226
rect 378178 352170 378246 352226
rect 378302 352170 408594 352226
rect 408650 352170 408718 352226
rect 408774 352170 408842 352226
rect 408898 352170 408966 352226
rect 409022 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 470034 352226
rect 470090 352170 470158 352226
rect 470214 352170 470282 352226
rect 470338 352170 470406 352226
rect 470462 352170 500754 352226
rect 500810 352170 500878 352226
rect 500934 352170 501002 352226
rect 501058 352170 501126 352226
rect 501182 352170 531474 352226
rect 531530 352170 531598 352226
rect 531654 352170 531722 352226
rect 531778 352170 531846 352226
rect 531902 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 149222 352102
rect 149278 352046 149346 352102
rect 149402 352046 179942 352102
rect 179998 352046 180066 352102
rect 180122 352046 224274 352102
rect 224330 352046 224398 352102
rect 224454 352046 224522 352102
rect 224578 352046 224646 352102
rect 224702 352046 254994 352102
rect 255050 352046 255118 352102
rect 255174 352046 255242 352102
rect 255298 352046 255366 352102
rect 255422 352046 285714 352102
rect 285770 352046 285838 352102
rect 285894 352046 285962 352102
rect 286018 352046 286086 352102
rect 286142 352046 316434 352102
rect 316490 352046 316558 352102
rect 316614 352046 316682 352102
rect 316738 352046 316806 352102
rect 316862 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 377874 352102
rect 377930 352046 377998 352102
rect 378054 352046 378122 352102
rect 378178 352046 378246 352102
rect 378302 352046 408594 352102
rect 408650 352046 408718 352102
rect 408774 352046 408842 352102
rect 408898 352046 408966 352102
rect 409022 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 470034 352102
rect 470090 352046 470158 352102
rect 470214 352046 470282 352102
rect 470338 352046 470406 352102
rect 470462 352046 500754 352102
rect 500810 352046 500878 352102
rect 500934 352046 501002 352102
rect 501058 352046 501126 352102
rect 501182 352046 531474 352102
rect 531530 352046 531598 352102
rect 531654 352046 531722 352102
rect 531778 352046 531846 352102
rect 531902 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 149222 351978
rect 149278 351922 149346 351978
rect 149402 351922 179942 351978
rect 179998 351922 180066 351978
rect 180122 351922 224274 351978
rect 224330 351922 224398 351978
rect 224454 351922 224522 351978
rect 224578 351922 224646 351978
rect 224702 351922 254994 351978
rect 255050 351922 255118 351978
rect 255174 351922 255242 351978
rect 255298 351922 255366 351978
rect 255422 351922 285714 351978
rect 285770 351922 285838 351978
rect 285894 351922 285962 351978
rect 286018 351922 286086 351978
rect 286142 351922 316434 351978
rect 316490 351922 316558 351978
rect 316614 351922 316682 351978
rect 316738 351922 316806 351978
rect 316862 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 377874 351978
rect 377930 351922 377998 351978
rect 378054 351922 378122 351978
rect 378178 351922 378246 351978
rect 378302 351922 408594 351978
rect 408650 351922 408718 351978
rect 408774 351922 408842 351978
rect 408898 351922 408966 351978
rect 409022 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 470034 351978
rect 470090 351922 470158 351978
rect 470214 351922 470282 351978
rect 470338 351922 470406 351978
rect 470462 351922 500754 351978
rect 500810 351922 500878 351978
rect 500934 351922 501002 351978
rect 501058 351922 501126 351978
rect 501182 351922 531474 351978
rect 531530 351922 531598 351978
rect 531654 351922 531722 351978
rect 531778 351922 531846 351978
rect 531902 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 133862 346350
rect 133918 346294 133986 346350
rect 134042 346294 164582 346350
rect 164638 346294 164706 346350
rect 164762 346294 195302 346350
rect 195358 346294 195426 346350
rect 195482 346294 220554 346350
rect 220610 346294 220678 346350
rect 220734 346294 220802 346350
rect 220858 346294 220926 346350
rect 220982 346294 251274 346350
rect 251330 346294 251398 346350
rect 251454 346294 251522 346350
rect 251578 346294 251646 346350
rect 251702 346294 281994 346350
rect 282050 346294 282118 346350
rect 282174 346294 282242 346350
rect 282298 346294 282366 346350
rect 282422 346294 312714 346350
rect 312770 346294 312838 346350
rect 312894 346294 312962 346350
rect 313018 346294 313086 346350
rect 313142 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 374154 346350
rect 374210 346294 374278 346350
rect 374334 346294 374402 346350
rect 374458 346294 374526 346350
rect 374582 346294 404874 346350
rect 404930 346294 404998 346350
rect 405054 346294 405122 346350
rect 405178 346294 405246 346350
rect 405302 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 466314 346350
rect 466370 346294 466438 346350
rect 466494 346294 466562 346350
rect 466618 346294 466686 346350
rect 466742 346294 497034 346350
rect 497090 346294 497158 346350
rect 497214 346294 497282 346350
rect 497338 346294 497406 346350
rect 497462 346294 527754 346350
rect 527810 346294 527878 346350
rect 527934 346294 528002 346350
rect 528058 346294 528126 346350
rect 528182 346294 558474 346350
rect 558530 346294 558598 346350
rect 558654 346294 558722 346350
rect 558778 346294 558846 346350
rect 558902 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 133862 346226
rect 133918 346170 133986 346226
rect 134042 346170 164582 346226
rect 164638 346170 164706 346226
rect 164762 346170 195302 346226
rect 195358 346170 195426 346226
rect 195482 346170 220554 346226
rect 220610 346170 220678 346226
rect 220734 346170 220802 346226
rect 220858 346170 220926 346226
rect 220982 346170 251274 346226
rect 251330 346170 251398 346226
rect 251454 346170 251522 346226
rect 251578 346170 251646 346226
rect 251702 346170 281994 346226
rect 282050 346170 282118 346226
rect 282174 346170 282242 346226
rect 282298 346170 282366 346226
rect 282422 346170 312714 346226
rect 312770 346170 312838 346226
rect 312894 346170 312962 346226
rect 313018 346170 313086 346226
rect 313142 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 374154 346226
rect 374210 346170 374278 346226
rect 374334 346170 374402 346226
rect 374458 346170 374526 346226
rect 374582 346170 404874 346226
rect 404930 346170 404998 346226
rect 405054 346170 405122 346226
rect 405178 346170 405246 346226
rect 405302 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 466314 346226
rect 466370 346170 466438 346226
rect 466494 346170 466562 346226
rect 466618 346170 466686 346226
rect 466742 346170 497034 346226
rect 497090 346170 497158 346226
rect 497214 346170 497282 346226
rect 497338 346170 497406 346226
rect 497462 346170 527754 346226
rect 527810 346170 527878 346226
rect 527934 346170 528002 346226
rect 528058 346170 528126 346226
rect 528182 346170 558474 346226
rect 558530 346170 558598 346226
rect 558654 346170 558722 346226
rect 558778 346170 558846 346226
rect 558902 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 133862 346102
rect 133918 346046 133986 346102
rect 134042 346046 164582 346102
rect 164638 346046 164706 346102
rect 164762 346046 195302 346102
rect 195358 346046 195426 346102
rect 195482 346046 220554 346102
rect 220610 346046 220678 346102
rect 220734 346046 220802 346102
rect 220858 346046 220926 346102
rect 220982 346046 251274 346102
rect 251330 346046 251398 346102
rect 251454 346046 251522 346102
rect 251578 346046 251646 346102
rect 251702 346046 281994 346102
rect 282050 346046 282118 346102
rect 282174 346046 282242 346102
rect 282298 346046 282366 346102
rect 282422 346046 312714 346102
rect 312770 346046 312838 346102
rect 312894 346046 312962 346102
rect 313018 346046 313086 346102
rect 313142 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 374154 346102
rect 374210 346046 374278 346102
rect 374334 346046 374402 346102
rect 374458 346046 374526 346102
rect 374582 346046 404874 346102
rect 404930 346046 404998 346102
rect 405054 346046 405122 346102
rect 405178 346046 405246 346102
rect 405302 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 466314 346102
rect 466370 346046 466438 346102
rect 466494 346046 466562 346102
rect 466618 346046 466686 346102
rect 466742 346046 497034 346102
rect 497090 346046 497158 346102
rect 497214 346046 497282 346102
rect 497338 346046 497406 346102
rect 497462 346046 527754 346102
rect 527810 346046 527878 346102
rect 527934 346046 528002 346102
rect 528058 346046 528126 346102
rect 528182 346046 558474 346102
rect 558530 346046 558598 346102
rect 558654 346046 558722 346102
rect 558778 346046 558846 346102
rect 558902 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 133862 345978
rect 133918 345922 133986 345978
rect 134042 345922 164582 345978
rect 164638 345922 164706 345978
rect 164762 345922 195302 345978
rect 195358 345922 195426 345978
rect 195482 345922 220554 345978
rect 220610 345922 220678 345978
rect 220734 345922 220802 345978
rect 220858 345922 220926 345978
rect 220982 345922 251274 345978
rect 251330 345922 251398 345978
rect 251454 345922 251522 345978
rect 251578 345922 251646 345978
rect 251702 345922 281994 345978
rect 282050 345922 282118 345978
rect 282174 345922 282242 345978
rect 282298 345922 282366 345978
rect 282422 345922 312714 345978
rect 312770 345922 312838 345978
rect 312894 345922 312962 345978
rect 313018 345922 313086 345978
rect 313142 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 374154 345978
rect 374210 345922 374278 345978
rect 374334 345922 374402 345978
rect 374458 345922 374526 345978
rect 374582 345922 404874 345978
rect 404930 345922 404998 345978
rect 405054 345922 405122 345978
rect 405178 345922 405246 345978
rect 405302 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 466314 345978
rect 466370 345922 466438 345978
rect 466494 345922 466562 345978
rect 466618 345922 466686 345978
rect 466742 345922 497034 345978
rect 497090 345922 497158 345978
rect 497214 345922 497282 345978
rect 497338 345922 497406 345978
rect 497462 345922 527754 345978
rect 527810 345922 527878 345978
rect 527934 345922 528002 345978
rect 528058 345922 528126 345978
rect 528182 345922 558474 345978
rect 558530 345922 558598 345978
rect 558654 345922 558722 345978
rect 558778 345922 558846 345978
rect 558902 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect 197356 336358 199348 336374
rect 197356 336302 197372 336358
rect 197428 336302 199276 336358
rect 199332 336302 199348 336358
rect 197356 336286 199348 336302
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 149222 334350
rect 149278 334294 149346 334350
rect 149402 334294 179942 334350
rect 179998 334294 180066 334350
rect 180122 334294 224274 334350
rect 224330 334294 224398 334350
rect 224454 334294 224522 334350
rect 224578 334294 224646 334350
rect 224702 334294 254994 334350
rect 255050 334294 255118 334350
rect 255174 334294 255242 334350
rect 255298 334294 255366 334350
rect 255422 334294 285714 334350
rect 285770 334294 285838 334350
rect 285894 334294 285962 334350
rect 286018 334294 286086 334350
rect 286142 334294 316434 334350
rect 316490 334294 316558 334350
rect 316614 334294 316682 334350
rect 316738 334294 316806 334350
rect 316862 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 377874 334350
rect 377930 334294 377998 334350
rect 378054 334294 378122 334350
rect 378178 334294 378246 334350
rect 378302 334294 408594 334350
rect 408650 334294 408718 334350
rect 408774 334294 408842 334350
rect 408898 334294 408966 334350
rect 409022 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 470034 334350
rect 470090 334294 470158 334350
rect 470214 334294 470282 334350
rect 470338 334294 470406 334350
rect 470462 334294 500754 334350
rect 500810 334294 500878 334350
rect 500934 334294 501002 334350
rect 501058 334294 501126 334350
rect 501182 334294 531474 334350
rect 531530 334294 531598 334350
rect 531654 334294 531722 334350
rect 531778 334294 531846 334350
rect 531902 334294 562194 334350
rect 562250 334294 562318 334350
rect 562374 334294 562442 334350
rect 562498 334294 562566 334350
rect 562622 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 149222 334226
rect 149278 334170 149346 334226
rect 149402 334170 179942 334226
rect 179998 334170 180066 334226
rect 180122 334170 224274 334226
rect 224330 334170 224398 334226
rect 224454 334170 224522 334226
rect 224578 334170 224646 334226
rect 224702 334170 254994 334226
rect 255050 334170 255118 334226
rect 255174 334170 255242 334226
rect 255298 334170 255366 334226
rect 255422 334170 285714 334226
rect 285770 334170 285838 334226
rect 285894 334170 285962 334226
rect 286018 334170 286086 334226
rect 286142 334170 316434 334226
rect 316490 334170 316558 334226
rect 316614 334170 316682 334226
rect 316738 334170 316806 334226
rect 316862 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 377874 334226
rect 377930 334170 377998 334226
rect 378054 334170 378122 334226
rect 378178 334170 378246 334226
rect 378302 334170 408594 334226
rect 408650 334170 408718 334226
rect 408774 334170 408842 334226
rect 408898 334170 408966 334226
rect 409022 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 470034 334226
rect 470090 334170 470158 334226
rect 470214 334170 470282 334226
rect 470338 334170 470406 334226
rect 470462 334170 500754 334226
rect 500810 334170 500878 334226
rect 500934 334170 501002 334226
rect 501058 334170 501126 334226
rect 501182 334170 531474 334226
rect 531530 334170 531598 334226
rect 531654 334170 531722 334226
rect 531778 334170 531846 334226
rect 531902 334170 562194 334226
rect 562250 334170 562318 334226
rect 562374 334170 562442 334226
rect 562498 334170 562566 334226
rect 562622 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 149222 334102
rect 149278 334046 149346 334102
rect 149402 334046 179942 334102
rect 179998 334046 180066 334102
rect 180122 334046 224274 334102
rect 224330 334046 224398 334102
rect 224454 334046 224522 334102
rect 224578 334046 224646 334102
rect 224702 334046 254994 334102
rect 255050 334046 255118 334102
rect 255174 334046 255242 334102
rect 255298 334046 255366 334102
rect 255422 334046 285714 334102
rect 285770 334046 285838 334102
rect 285894 334046 285962 334102
rect 286018 334046 286086 334102
rect 286142 334046 316434 334102
rect 316490 334046 316558 334102
rect 316614 334046 316682 334102
rect 316738 334046 316806 334102
rect 316862 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 377874 334102
rect 377930 334046 377998 334102
rect 378054 334046 378122 334102
rect 378178 334046 378246 334102
rect 378302 334046 408594 334102
rect 408650 334046 408718 334102
rect 408774 334046 408842 334102
rect 408898 334046 408966 334102
rect 409022 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 470034 334102
rect 470090 334046 470158 334102
rect 470214 334046 470282 334102
rect 470338 334046 470406 334102
rect 470462 334046 500754 334102
rect 500810 334046 500878 334102
rect 500934 334046 501002 334102
rect 501058 334046 501126 334102
rect 501182 334046 531474 334102
rect 531530 334046 531598 334102
rect 531654 334046 531722 334102
rect 531778 334046 531846 334102
rect 531902 334046 562194 334102
rect 562250 334046 562318 334102
rect 562374 334046 562442 334102
rect 562498 334046 562566 334102
rect 562622 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 149222 333978
rect 149278 333922 149346 333978
rect 149402 333922 179942 333978
rect 179998 333922 180066 333978
rect 180122 333922 224274 333978
rect 224330 333922 224398 333978
rect 224454 333922 224522 333978
rect 224578 333922 224646 333978
rect 224702 333922 254994 333978
rect 255050 333922 255118 333978
rect 255174 333922 255242 333978
rect 255298 333922 255366 333978
rect 255422 333922 285714 333978
rect 285770 333922 285838 333978
rect 285894 333922 285962 333978
rect 286018 333922 286086 333978
rect 286142 333922 316434 333978
rect 316490 333922 316558 333978
rect 316614 333922 316682 333978
rect 316738 333922 316806 333978
rect 316862 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 377874 333978
rect 377930 333922 377998 333978
rect 378054 333922 378122 333978
rect 378178 333922 378246 333978
rect 378302 333922 408594 333978
rect 408650 333922 408718 333978
rect 408774 333922 408842 333978
rect 408898 333922 408966 333978
rect 409022 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 470034 333978
rect 470090 333922 470158 333978
rect 470214 333922 470282 333978
rect 470338 333922 470406 333978
rect 470462 333922 500754 333978
rect 500810 333922 500878 333978
rect 500934 333922 501002 333978
rect 501058 333922 501126 333978
rect 501182 333922 531474 333978
rect 531530 333922 531598 333978
rect 531654 333922 531722 333978
rect 531778 333922 531846 333978
rect 531902 333922 562194 333978
rect 562250 333922 562318 333978
rect 562374 333922 562442 333978
rect 562498 333922 562566 333978
rect 562622 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect 3036 332038 114228 332054
rect 3036 331982 3052 332038
rect 3108 331982 114156 332038
rect 114212 331982 114228 332038
rect 3036 331966 114228 331982
rect 5052 331858 117588 331874
rect 5052 331802 5068 331858
rect 5124 331802 117516 331858
rect 117572 331802 117588 331858
rect 5052 331786 117588 331802
rect 197468 330238 199348 330254
rect 197468 330182 197484 330238
rect 197540 330182 199276 330238
rect 199332 330182 199348 330238
rect 197468 330166 199348 330182
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 133862 328350
rect 133918 328294 133986 328350
rect 134042 328294 164582 328350
rect 164638 328294 164706 328350
rect 164762 328294 195302 328350
rect 195358 328294 195426 328350
rect 195482 328294 220554 328350
rect 220610 328294 220678 328350
rect 220734 328294 220802 328350
rect 220858 328294 220926 328350
rect 220982 328294 251274 328350
rect 251330 328294 251398 328350
rect 251454 328294 251522 328350
rect 251578 328294 251646 328350
rect 251702 328294 281994 328350
rect 282050 328294 282118 328350
rect 282174 328294 282242 328350
rect 282298 328294 282366 328350
rect 282422 328294 312714 328350
rect 312770 328294 312838 328350
rect 312894 328294 312962 328350
rect 313018 328294 313086 328350
rect 313142 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 374154 328350
rect 374210 328294 374278 328350
rect 374334 328294 374402 328350
rect 374458 328294 374526 328350
rect 374582 328294 404874 328350
rect 404930 328294 404998 328350
rect 405054 328294 405122 328350
rect 405178 328294 405246 328350
rect 405302 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 466314 328350
rect 466370 328294 466438 328350
rect 466494 328294 466562 328350
rect 466618 328294 466686 328350
rect 466742 328294 497034 328350
rect 497090 328294 497158 328350
rect 497214 328294 497282 328350
rect 497338 328294 497406 328350
rect 497462 328294 527754 328350
rect 527810 328294 527878 328350
rect 527934 328294 528002 328350
rect 528058 328294 528126 328350
rect 528182 328294 558474 328350
rect 558530 328294 558598 328350
rect 558654 328294 558722 328350
rect 558778 328294 558846 328350
rect 558902 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 133862 328226
rect 133918 328170 133986 328226
rect 134042 328170 164582 328226
rect 164638 328170 164706 328226
rect 164762 328170 195302 328226
rect 195358 328170 195426 328226
rect 195482 328170 220554 328226
rect 220610 328170 220678 328226
rect 220734 328170 220802 328226
rect 220858 328170 220926 328226
rect 220982 328170 251274 328226
rect 251330 328170 251398 328226
rect 251454 328170 251522 328226
rect 251578 328170 251646 328226
rect 251702 328170 281994 328226
rect 282050 328170 282118 328226
rect 282174 328170 282242 328226
rect 282298 328170 282366 328226
rect 282422 328170 312714 328226
rect 312770 328170 312838 328226
rect 312894 328170 312962 328226
rect 313018 328170 313086 328226
rect 313142 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 374154 328226
rect 374210 328170 374278 328226
rect 374334 328170 374402 328226
rect 374458 328170 374526 328226
rect 374582 328170 404874 328226
rect 404930 328170 404998 328226
rect 405054 328170 405122 328226
rect 405178 328170 405246 328226
rect 405302 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 466314 328226
rect 466370 328170 466438 328226
rect 466494 328170 466562 328226
rect 466618 328170 466686 328226
rect 466742 328170 497034 328226
rect 497090 328170 497158 328226
rect 497214 328170 497282 328226
rect 497338 328170 497406 328226
rect 497462 328170 527754 328226
rect 527810 328170 527878 328226
rect 527934 328170 528002 328226
rect 528058 328170 528126 328226
rect 528182 328170 558474 328226
rect 558530 328170 558598 328226
rect 558654 328170 558722 328226
rect 558778 328170 558846 328226
rect 558902 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 133862 328102
rect 133918 328046 133986 328102
rect 134042 328046 164582 328102
rect 164638 328046 164706 328102
rect 164762 328046 195302 328102
rect 195358 328046 195426 328102
rect 195482 328046 220554 328102
rect 220610 328046 220678 328102
rect 220734 328046 220802 328102
rect 220858 328046 220926 328102
rect 220982 328046 251274 328102
rect 251330 328046 251398 328102
rect 251454 328046 251522 328102
rect 251578 328046 251646 328102
rect 251702 328046 281994 328102
rect 282050 328046 282118 328102
rect 282174 328046 282242 328102
rect 282298 328046 282366 328102
rect 282422 328046 312714 328102
rect 312770 328046 312838 328102
rect 312894 328046 312962 328102
rect 313018 328046 313086 328102
rect 313142 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 374154 328102
rect 374210 328046 374278 328102
rect 374334 328046 374402 328102
rect 374458 328046 374526 328102
rect 374582 328046 404874 328102
rect 404930 328046 404998 328102
rect 405054 328046 405122 328102
rect 405178 328046 405246 328102
rect 405302 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 466314 328102
rect 466370 328046 466438 328102
rect 466494 328046 466562 328102
rect 466618 328046 466686 328102
rect 466742 328046 497034 328102
rect 497090 328046 497158 328102
rect 497214 328046 497282 328102
rect 497338 328046 497406 328102
rect 497462 328046 527754 328102
rect 527810 328046 527878 328102
rect 527934 328046 528002 328102
rect 528058 328046 528126 328102
rect 528182 328046 558474 328102
rect 558530 328046 558598 328102
rect 558654 328046 558722 328102
rect 558778 328046 558846 328102
rect 558902 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 133862 327978
rect 133918 327922 133986 327978
rect 134042 327922 164582 327978
rect 164638 327922 164706 327978
rect 164762 327922 195302 327978
rect 195358 327922 195426 327978
rect 195482 327922 220554 327978
rect 220610 327922 220678 327978
rect 220734 327922 220802 327978
rect 220858 327922 220926 327978
rect 220982 327922 251274 327978
rect 251330 327922 251398 327978
rect 251454 327922 251522 327978
rect 251578 327922 251646 327978
rect 251702 327922 281994 327978
rect 282050 327922 282118 327978
rect 282174 327922 282242 327978
rect 282298 327922 282366 327978
rect 282422 327922 312714 327978
rect 312770 327922 312838 327978
rect 312894 327922 312962 327978
rect 313018 327922 313086 327978
rect 313142 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 374154 327978
rect 374210 327922 374278 327978
rect 374334 327922 374402 327978
rect 374458 327922 374526 327978
rect 374582 327922 404874 327978
rect 404930 327922 404998 327978
rect 405054 327922 405122 327978
rect 405178 327922 405246 327978
rect 405302 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 466314 327978
rect 466370 327922 466438 327978
rect 466494 327922 466562 327978
rect 466618 327922 466686 327978
rect 466742 327922 497034 327978
rect 497090 327922 497158 327978
rect 497214 327922 497282 327978
rect 497338 327922 497406 327978
rect 497462 327922 527754 327978
rect 527810 327922 527878 327978
rect 527934 327922 528002 327978
rect 528058 327922 528126 327978
rect 528182 327922 558474 327978
rect 558530 327922 558598 327978
rect 558654 327922 558722 327978
rect 558778 327922 558846 327978
rect 558902 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect 106748 326098 116020 326114
rect 106748 326042 106764 326098
rect 106820 326042 115948 326098
rect 116004 326042 116020 326098
rect 106748 326026 116020 326042
rect 5276 325018 57108 325034
rect 5276 324962 5292 325018
rect 5348 324962 57036 325018
rect 57092 324962 57108 325018
rect 5276 324946 57108 324962
rect 60156 321058 61364 321074
rect 60156 321002 60172 321058
rect 60228 321002 61292 321058
rect 61348 321002 61364 321058
rect 60156 320986 61364 321002
rect 118396 319078 121844 319094
rect 118396 319022 118412 319078
rect 118468 319022 121772 319078
rect 121828 319022 121844 319078
rect 118396 319006 121844 319022
rect 197580 317818 199348 317834
rect 197580 317762 197596 317818
rect 197652 317762 199276 317818
rect 199332 317762 199348 317818
rect 197580 317746 199348 317762
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 24878 316350
rect 24934 316294 25002 316350
rect 25058 316294 79878 316350
rect 79934 316294 80002 316350
rect 80058 316294 149222 316350
rect 149278 316294 149346 316350
rect 149402 316294 179942 316350
rect 179998 316294 180066 316350
rect 180122 316294 229878 316350
rect 229934 316294 230002 316350
rect 230058 316294 260598 316350
rect 260654 316294 260722 316350
rect 260778 316294 291318 316350
rect 291374 316294 291442 316350
rect 291498 316294 322038 316350
rect 322094 316294 322162 316350
rect 322218 316294 352758 316350
rect 352814 316294 352882 316350
rect 352938 316294 377874 316350
rect 377930 316294 377998 316350
rect 378054 316294 378122 316350
rect 378178 316294 378246 316350
rect 378302 316294 399878 316350
rect 399934 316294 400002 316350
rect 400058 316294 408594 316350
rect 408650 316294 408718 316350
rect 408774 316294 408842 316350
rect 408898 316294 408966 316350
rect 409022 316294 430598 316350
rect 430654 316294 430722 316350
rect 430778 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 470034 316350
rect 470090 316294 470158 316350
rect 470214 316294 470282 316350
rect 470338 316294 470406 316350
rect 470462 316294 500754 316350
rect 500810 316294 500878 316350
rect 500934 316294 501002 316350
rect 501058 316294 501126 316350
rect 501182 316294 531474 316350
rect 531530 316294 531598 316350
rect 531654 316294 531722 316350
rect 531778 316294 531846 316350
rect 531902 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 24878 316226
rect 24934 316170 25002 316226
rect 25058 316170 79878 316226
rect 79934 316170 80002 316226
rect 80058 316170 149222 316226
rect 149278 316170 149346 316226
rect 149402 316170 179942 316226
rect 179998 316170 180066 316226
rect 180122 316170 229878 316226
rect 229934 316170 230002 316226
rect 230058 316170 260598 316226
rect 260654 316170 260722 316226
rect 260778 316170 291318 316226
rect 291374 316170 291442 316226
rect 291498 316170 322038 316226
rect 322094 316170 322162 316226
rect 322218 316170 352758 316226
rect 352814 316170 352882 316226
rect 352938 316170 377874 316226
rect 377930 316170 377998 316226
rect 378054 316170 378122 316226
rect 378178 316170 378246 316226
rect 378302 316170 399878 316226
rect 399934 316170 400002 316226
rect 400058 316170 408594 316226
rect 408650 316170 408718 316226
rect 408774 316170 408842 316226
rect 408898 316170 408966 316226
rect 409022 316170 430598 316226
rect 430654 316170 430722 316226
rect 430778 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 470034 316226
rect 470090 316170 470158 316226
rect 470214 316170 470282 316226
rect 470338 316170 470406 316226
rect 470462 316170 500754 316226
rect 500810 316170 500878 316226
rect 500934 316170 501002 316226
rect 501058 316170 501126 316226
rect 501182 316170 531474 316226
rect 531530 316170 531598 316226
rect 531654 316170 531722 316226
rect 531778 316170 531846 316226
rect 531902 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 24878 316102
rect 24934 316046 25002 316102
rect 25058 316046 79878 316102
rect 79934 316046 80002 316102
rect 80058 316046 149222 316102
rect 149278 316046 149346 316102
rect 149402 316046 179942 316102
rect 179998 316046 180066 316102
rect 180122 316046 229878 316102
rect 229934 316046 230002 316102
rect 230058 316046 260598 316102
rect 260654 316046 260722 316102
rect 260778 316046 291318 316102
rect 291374 316046 291442 316102
rect 291498 316046 322038 316102
rect 322094 316046 322162 316102
rect 322218 316046 352758 316102
rect 352814 316046 352882 316102
rect 352938 316046 377874 316102
rect 377930 316046 377998 316102
rect 378054 316046 378122 316102
rect 378178 316046 378246 316102
rect 378302 316046 399878 316102
rect 399934 316046 400002 316102
rect 400058 316046 408594 316102
rect 408650 316046 408718 316102
rect 408774 316046 408842 316102
rect 408898 316046 408966 316102
rect 409022 316046 430598 316102
rect 430654 316046 430722 316102
rect 430778 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 470034 316102
rect 470090 316046 470158 316102
rect 470214 316046 470282 316102
rect 470338 316046 470406 316102
rect 470462 316046 500754 316102
rect 500810 316046 500878 316102
rect 500934 316046 501002 316102
rect 501058 316046 501126 316102
rect 501182 316046 531474 316102
rect 531530 316046 531598 316102
rect 531654 316046 531722 316102
rect 531778 316046 531846 316102
rect 531902 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 24878 315978
rect 24934 315922 25002 315978
rect 25058 315922 79878 315978
rect 79934 315922 80002 315978
rect 80058 315922 149222 315978
rect 149278 315922 149346 315978
rect 149402 315922 179942 315978
rect 179998 315922 180066 315978
rect 180122 315922 229878 315978
rect 229934 315922 230002 315978
rect 230058 315922 260598 315978
rect 260654 315922 260722 315978
rect 260778 315922 291318 315978
rect 291374 315922 291442 315978
rect 291498 315922 322038 315978
rect 322094 315922 322162 315978
rect 322218 315922 352758 315978
rect 352814 315922 352882 315978
rect 352938 315922 377874 315978
rect 377930 315922 377998 315978
rect 378054 315922 378122 315978
rect 378178 315922 378246 315978
rect 378302 315922 399878 315978
rect 399934 315922 400002 315978
rect 400058 315922 408594 315978
rect 408650 315922 408718 315978
rect 408774 315922 408842 315978
rect 408898 315922 408966 315978
rect 409022 315922 430598 315978
rect 430654 315922 430722 315978
rect 430778 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 470034 315978
rect 470090 315922 470158 315978
rect 470214 315922 470282 315978
rect 470338 315922 470406 315978
rect 470462 315922 500754 315978
rect 500810 315922 500878 315978
rect 500934 315922 501002 315978
rect 501058 315922 501126 315978
rect 501182 315922 531474 315978
rect 531530 315922 531598 315978
rect 531654 315922 531722 315978
rect 531778 315922 531846 315978
rect 531902 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect 113020 312598 117476 312614
rect 113020 312542 113036 312598
rect 113092 312542 117404 312598
rect 117460 312542 117476 312598
rect 113020 312526 117476 312542
rect 411500 312598 418644 312614
rect 411500 312542 411516 312598
rect 411572 312542 418572 312598
rect 418628 312542 418644 312598
rect 411500 312526 418644 312542
rect 114252 310978 121732 310994
rect 114252 310922 114268 310978
rect 114324 310922 121660 310978
rect 121716 310922 121732 310978
rect 114252 310906 121732 310922
rect 373756 310978 440596 310994
rect 373756 310922 373772 310978
rect 373828 310922 440524 310978
rect 440580 310922 440596 310978
rect 373756 310906 440596 310922
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 9518 310350
rect 9574 310294 9642 310350
rect 9698 310294 40238 310350
rect 40294 310294 40362 310350
rect 40418 310294 64518 310350
rect 64574 310294 64642 310350
rect 64698 310294 95238 310350
rect 95294 310294 95362 310350
rect 95418 310294 133862 310350
rect 133918 310294 133986 310350
rect 134042 310294 164582 310350
rect 164638 310294 164706 310350
rect 164762 310294 195302 310350
rect 195358 310294 195426 310350
rect 195482 310294 214518 310350
rect 214574 310294 214642 310350
rect 214698 310294 245238 310350
rect 245294 310294 245362 310350
rect 245418 310294 275958 310350
rect 276014 310294 276082 310350
rect 276138 310294 306678 310350
rect 306734 310294 306802 310350
rect 306858 310294 337398 310350
rect 337454 310294 337522 310350
rect 337578 310294 368118 310350
rect 368174 310294 368242 310350
rect 368298 310294 374154 310350
rect 374210 310294 374278 310350
rect 374334 310294 374402 310350
rect 374458 310294 374526 310350
rect 374582 310294 384518 310350
rect 384574 310294 384642 310350
rect 384698 310294 415238 310350
rect 415294 310294 415362 310350
rect 415418 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 466314 310350
rect 466370 310294 466438 310350
rect 466494 310294 466562 310350
rect 466618 310294 466686 310350
rect 466742 310294 497034 310350
rect 497090 310294 497158 310350
rect 497214 310294 497282 310350
rect 497338 310294 497406 310350
rect 497462 310294 527754 310350
rect 527810 310294 527878 310350
rect 527934 310294 528002 310350
rect 528058 310294 528126 310350
rect 528182 310294 558474 310350
rect 558530 310294 558598 310350
rect 558654 310294 558722 310350
rect 558778 310294 558846 310350
rect 558902 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 9518 310226
rect 9574 310170 9642 310226
rect 9698 310170 40238 310226
rect 40294 310170 40362 310226
rect 40418 310170 64518 310226
rect 64574 310170 64642 310226
rect 64698 310170 95238 310226
rect 95294 310170 95362 310226
rect 95418 310170 133862 310226
rect 133918 310170 133986 310226
rect 134042 310170 164582 310226
rect 164638 310170 164706 310226
rect 164762 310170 195302 310226
rect 195358 310170 195426 310226
rect 195482 310170 214518 310226
rect 214574 310170 214642 310226
rect 214698 310170 245238 310226
rect 245294 310170 245362 310226
rect 245418 310170 275958 310226
rect 276014 310170 276082 310226
rect 276138 310170 306678 310226
rect 306734 310170 306802 310226
rect 306858 310170 337398 310226
rect 337454 310170 337522 310226
rect 337578 310170 368118 310226
rect 368174 310170 368242 310226
rect 368298 310170 374154 310226
rect 374210 310170 374278 310226
rect 374334 310170 374402 310226
rect 374458 310170 374526 310226
rect 374582 310170 384518 310226
rect 384574 310170 384642 310226
rect 384698 310170 415238 310226
rect 415294 310170 415362 310226
rect 415418 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 466314 310226
rect 466370 310170 466438 310226
rect 466494 310170 466562 310226
rect 466618 310170 466686 310226
rect 466742 310170 497034 310226
rect 497090 310170 497158 310226
rect 497214 310170 497282 310226
rect 497338 310170 497406 310226
rect 497462 310170 527754 310226
rect 527810 310170 527878 310226
rect 527934 310170 528002 310226
rect 528058 310170 528126 310226
rect 528182 310170 558474 310226
rect 558530 310170 558598 310226
rect 558654 310170 558722 310226
rect 558778 310170 558846 310226
rect 558902 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 9518 310102
rect 9574 310046 9642 310102
rect 9698 310046 40238 310102
rect 40294 310046 40362 310102
rect 40418 310046 64518 310102
rect 64574 310046 64642 310102
rect 64698 310046 95238 310102
rect 95294 310046 95362 310102
rect 95418 310046 133862 310102
rect 133918 310046 133986 310102
rect 134042 310046 164582 310102
rect 164638 310046 164706 310102
rect 164762 310046 195302 310102
rect 195358 310046 195426 310102
rect 195482 310046 214518 310102
rect 214574 310046 214642 310102
rect 214698 310046 245238 310102
rect 245294 310046 245362 310102
rect 245418 310046 275958 310102
rect 276014 310046 276082 310102
rect 276138 310046 306678 310102
rect 306734 310046 306802 310102
rect 306858 310046 337398 310102
rect 337454 310046 337522 310102
rect 337578 310046 368118 310102
rect 368174 310046 368242 310102
rect 368298 310046 374154 310102
rect 374210 310046 374278 310102
rect 374334 310046 374402 310102
rect 374458 310046 374526 310102
rect 374582 310046 384518 310102
rect 384574 310046 384642 310102
rect 384698 310046 415238 310102
rect 415294 310046 415362 310102
rect 415418 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 466314 310102
rect 466370 310046 466438 310102
rect 466494 310046 466562 310102
rect 466618 310046 466686 310102
rect 466742 310046 497034 310102
rect 497090 310046 497158 310102
rect 497214 310046 497282 310102
rect 497338 310046 497406 310102
rect 497462 310046 527754 310102
rect 527810 310046 527878 310102
rect 527934 310046 528002 310102
rect 528058 310046 528126 310102
rect 528182 310046 558474 310102
rect 558530 310046 558598 310102
rect 558654 310046 558722 310102
rect 558778 310046 558846 310102
rect 558902 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 9518 309978
rect 9574 309922 9642 309978
rect 9698 309922 40238 309978
rect 40294 309922 40362 309978
rect 40418 309922 64518 309978
rect 64574 309922 64642 309978
rect 64698 309922 95238 309978
rect 95294 309922 95362 309978
rect 95418 309922 133862 309978
rect 133918 309922 133986 309978
rect 134042 309922 164582 309978
rect 164638 309922 164706 309978
rect 164762 309922 195302 309978
rect 195358 309922 195426 309978
rect 195482 309922 214518 309978
rect 214574 309922 214642 309978
rect 214698 309922 245238 309978
rect 245294 309922 245362 309978
rect 245418 309922 275958 309978
rect 276014 309922 276082 309978
rect 276138 309922 306678 309978
rect 306734 309922 306802 309978
rect 306858 309922 337398 309978
rect 337454 309922 337522 309978
rect 337578 309922 368118 309978
rect 368174 309922 368242 309978
rect 368298 309922 374154 309978
rect 374210 309922 374278 309978
rect 374334 309922 374402 309978
rect 374458 309922 374526 309978
rect 374582 309922 384518 309978
rect 384574 309922 384642 309978
rect 384698 309922 415238 309978
rect 415294 309922 415362 309978
rect 415418 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 466314 309978
rect 466370 309922 466438 309978
rect 466494 309922 466562 309978
rect 466618 309922 466686 309978
rect 466742 309922 497034 309978
rect 497090 309922 497158 309978
rect 497214 309922 497282 309978
rect 497338 309922 497406 309978
rect 497462 309922 527754 309978
rect 527810 309922 527878 309978
rect 527934 309922 528002 309978
rect 528058 309922 528126 309978
rect 528182 309922 558474 309978
rect 558530 309922 558598 309978
rect 558654 309922 558722 309978
rect 558778 309922 558846 309978
rect 558902 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect 5276 308998 7604 309014
rect 5276 308942 5292 308998
rect 5348 308942 7532 308998
rect 7588 308942 7604 308998
rect 5276 308926 7604 308942
rect 58700 307558 63044 307574
rect 58700 307502 58716 307558
rect 58772 307502 62972 307558
rect 63028 307502 63044 307558
rect 58700 307486 63044 307502
rect 204860 306658 212228 306674
rect 204860 306602 204876 306658
rect 204932 306602 212156 306658
rect 212212 306602 212228 306658
rect 204860 306586 212228 306602
rect 198140 305758 199908 305774
rect 198140 305702 198156 305758
rect 198212 305702 199836 305758
rect 199892 305702 199908 305758
rect 198140 305686 199908 305702
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 24878 298350
rect 24934 298294 25002 298350
rect 25058 298294 79878 298350
rect 79934 298294 80002 298350
rect 80058 298294 149222 298350
rect 149278 298294 149346 298350
rect 149402 298294 179942 298350
rect 179998 298294 180066 298350
rect 180122 298294 229878 298350
rect 229934 298294 230002 298350
rect 230058 298294 260598 298350
rect 260654 298294 260722 298350
rect 260778 298294 291318 298350
rect 291374 298294 291442 298350
rect 291498 298294 322038 298350
rect 322094 298294 322162 298350
rect 322218 298294 352758 298350
rect 352814 298294 352882 298350
rect 352938 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 399878 298350
rect 399934 298294 400002 298350
rect 400058 298294 430598 298350
rect 430654 298294 430722 298350
rect 430778 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 470034 298350
rect 470090 298294 470158 298350
rect 470214 298294 470282 298350
rect 470338 298294 470406 298350
rect 470462 298294 500754 298350
rect 500810 298294 500878 298350
rect 500934 298294 501002 298350
rect 501058 298294 501126 298350
rect 501182 298294 531474 298350
rect 531530 298294 531598 298350
rect 531654 298294 531722 298350
rect 531778 298294 531846 298350
rect 531902 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 24878 298226
rect 24934 298170 25002 298226
rect 25058 298170 79878 298226
rect 79934 298170 80002 298226
rect 80058 298170 149222 298226
rect 149278 298170 149346 298226
rect 149402 298170 179942 298226
rect 179998 298170 180066 298226
rect 180122 298170 229878 298226
rect 229934 298170 230002 298226
rect 230058 298170 260598 298226
rect 260654 298170 260722 298226
rect 260778 298170 291318 298226
rect 291374 298170 291442 298226
rect 291498 298170 322038 298226
rect 322094 298170 322162 298226
rect 322218 298170 352758 298226
rect 352814 298170 352882 298226
rect 352938 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 399878 298226
rect 399934 298170 400002 298226
rect 400058 298170 430598 298226
rect 430654 298170 430722 298226
rect 430778 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 470034 298226
rect 470090 298170 470158 298226
rect 470214 298170 470282 298226
rect 470338 298170 470406 298226
rect 470462 298170 500754 298226
rect 500810 298170 500878 298226
rect 500934 298170 501002 298226
rect 501058 298170 501126 298226
rect 501182 298170 531474 298226
rect 531530 298170 531598 298226
rect 531654 298170 531722 298226
rect 531778 298170 531846 298226
rect 531902 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 24878 298102
rect 24934 298046 25002 298102
rect 25058 298046 79878 298102
rect 79934 298046 80002 298102
rect 80058 298046 149222 298102
rect 149278 298046 149346 298102
rect 149402 298046 179942 298102
rect 179998 298046 180066 298102
rect 180122 298046 229878 298102
rect 229934 298046 230002 298102
rect 230058 298046 260598 298102
rect 260654 298046 260722 298102
rect 260778 298046 291318 298102
rect 291374 298046 291442 298102
rect 291498 298046 322038 298102
rect 322094 298046 322162 298102
rect 322218 298046 352758 298102
rect 352814 298046 352882 298102
rect 352938 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 399878 298102
rect 399934 298046 400002 298102
rect 400058 298046 430598 298102
rect 430654 298046 430722 298102
rect 430778 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 470034 298102
rect 470090 298046 470158 298102
rect 470214 298046 470282 298102
rect 470338 298046 470406 298102
rect 470462 298046 500754 298102
rect 500810 298046 500878 298102
rect 500934 298046 501002 298102
rect 501058 298046 501126 298102
rect 501182 298046 531474 298102
rect 531530 298046 531598 298102
rect 531654 298046 531722 298102
rect 531778 298046 531846 298102
rect 531902 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 24878 297978
rect 24934 297922 25002 297978
rect 25058 297922 79878 297978
rect 79934 297922 80002 297978
rect 80058 297922 149222 297978
rect 149278 297922 149346 297978
rect 149402 297922 179942 297978
rect 179998 297922 180066 297978
rect 180122 297922 229878 297978
rect 229934 297922 230002 297978
rect 230058 297922 260598 297978
rect 260654 297922 260722 297978
rect 260778 297922 291318 297978
rect 291374 297922 291442 297978
rect 291498 297922 322038 297978
rect 322094 297922 322162 297978
rect 322218 297922 352758 297978
rect 352814 297922 352882 297978
rect 352938 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 399878 297978
rect 399934 297922 400002 297978
rect 400058 297922 430598 297978
rect 430654 297922 430722 297978
rect 430778 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 470034 297978
rect 470090 297922 470158 297978
rect 470214 297922 470282 297978
rect 470338 297922 470406 297978
rect 470462 297922 500754 297978
rect 500810 297922 500878 297978
rect 500934 297922 501002 297978
rect 501058 297922 501126 297978
rect 501182 297922 531474 297978
rect 531530 297922 531598 297978
rect 531654 297922 531722 297978
rect 531778 297922 531846 297978
rect 531902 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect 194332 296758 199348 296774
rect 194332 296702 194348 296758
rect 194404 296702 199276 296758
rect 199332 296702 199348 296758
rect 194332 296686 199348 296702
rect 195788 296398 201924 296414
rect 195788 296342 195804 296398
rect 195860 296342 201852 296398
rect 201908 296342 201924 296398
rect 195788 296326 201924 296342
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 9518 292350
rect 9574 292294 9642 292350
rect 9698 292294 40238 292350
rect 40294 292294 40362 292350
rect 40418 292294 64518 292350
rect 64574 292294 64642 292350
rect 64698 292294 95238 292350
rect 95294 292294 95362 292350
rect 95418 292294 133862 292350
rect 133918 292294 133986 292350
rect 134042 292294 164582 292350
rect 164638 292294 164706 292350
rect 164762 292294 195302 292350
rect 195358 292294 195426 292350
rect 195482 292294 214518 292350
rect 214574 292294 214642 292350
rect 214698 292294 245238 292350
rect 245294 292294 245362 292350
rect 245418 292294 275958 292350
rect 276014 292294 276082 292350
rect 276138 292294 306678 292350
rect 306734 292294 306802 292350
rect 306858 292294 337398 292350
rect 337454 292294 337522 292350
rect 337578 292294 368118 292350
rect 368174 292294 368242 292350
rect 368298 292294 374154 292350
rect 374210 292294 374278 292350
rect 374334 292294 374402 292350
rect 374458 292294 374526 292350
rect 374582 292294 384518 292350
rect 384574 292294 384642 292350
rect 384698 292294 415238 292350
rect 415294 292294 415362 292350
rect 415418 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 466314 292350
rect 466370 292294 466438 292350
rect 466494 292294 466562 292350
rect 466618 292294 466686 292350
rect 466742 292294 497034 292350
rect 497090 292294 497158 292350
rect 497214 292294 497282 292350
rect 497338 292294 497406 292350
rect 497462 292294 527754 292350
rect 527810 292294 527878 292350
rect 527934 292294 528002 292350
rect 528058 292294 528126 292350
rect 528182 292294 558474 292350
rect 558530 292294 558598 292350
rect 558654 292294 558722 292350
rect 558778 292294 558846 292350
rect 558902 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 9518 292226
rect 9574 292170 9642 292226
rect 9698 292170 40238 292226
rect 40294 292170 40362 292226
rect 40418 292170 64518 292226
rect 64574 292170 64642 292226
rect 64698 292170 95238 292226
rect 95294 292170 95362 292226
rect 95418 292170 133862 292226
rect 133918 292170 133986 292226
rect 134042 292170 164582 292226
rect 164638 292170 164706 292226
rect 164762 292170 195302 292226
rect 195358 292170 195426 292226
rect 195482 292170 214518 292226
rect 214574 292170 214642 292226
rect 214698 292170 245238 292226
rect 245294 292170 245362 292226
rect 245418 292170 275958 292226
rect 276014 292170 276082 292226
rect 276138 292170 306678 292226
rect 306734 292170 306802 292226
rect 306858 292170 337398 292226
rect 337454 292170 337522 292226
rect 337578 292170 368118 292226
rect 368174 292170 368242 292226
rect 368298 292170 374154 292226
rect 374210 292170 374278 292226
rect 374334 292170 374402 292226
rect 374458 292170 374526 292226
rect 374582 292170 384518 292226
rect 384574 292170 384642 292226
rect 384698 292170 415238 292226
rect 415294 292170 415362 292226
rect 415418 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 466314 292226
rect 466370 292170 466438 292226
rect 466494 292170 466562 292226
rect 466618 292170 466686 292226
rect 466742 292170 497034 292226
rect 497090 292170 497158 292226
rect 497214 292170 497282 292226
rect 497338 292170 497406 292226
rect 497462 292170 527754 292226
rect 527810 292170 527878 292226
rect 527934 292170 528002 292226
rect 528058 292170 528126 292226
rect 528182 292170 558474 292226
rect 558530 292170 558598 292226
rect 558654 292170 558722 292226
rect 558778 292170 558846 292226
rect 558902 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 9518 292102
rect 9574 292046 9642 292102
rect 9698 292046 40238 292102
rect 40294 292046 40362 292102
rect 40418 292046 64518 292102
rect 64574 292046 64642 292102
rect 64698 292046 95238 292102
rect 95294 292046 95362 292102
rect 95418 292046 133862 292102
rect 133918 292046 133986 292102
rect 134042 292046 164582 292102
rect 164638 292046 164706 292102
rect 164762 292046 195302 292102
rect 195358 292046 195426 292102
rect 195482 292046 214518 292102
rect 214574 292046 214642 292102
rect 214698 292046 245238 292102
rect 245294 292046 245362 292102
rect 245418 292046 275958 292102
rect 276014 292046 276082 292102
rect 276138 292046 306678 292102
rect 306734 292046 306802 292102
rect 306858 292046 337398 292102
rect 337454 292046 337522 292102
rect 337578 292046 368118 292102
rect 368174 292046 368242 292102
rect 368298 292046 374154 292102
rect 374210 292046 374278 292102
rect 374334 292046 374402 292102
rect 374458 292046 374526 292102
rect 374582 292046 384518 292102
rect 384574 292046 384642 292102
rect 384698 292046 415238 292102
rect 415294 292046 415362 292102
rect 415418 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 466314 292102
rect 466370 292046 466438 292102
rect 466494 292046 466562 292102
rect 466618 292046 466686 292102
rect 466742 292046 497034 292102
rect 497090 292046 497158 292102
rect 497214 292046 497282 292102
rect 497338 292046 497406 292102
rect 497462 292046 527754 292102
rect 527810 292046 527878 292102
rect 527934 292046 528002 292102
rect 528058 292046 528126 292102
rect 528182 292046 558474 292102
rect 558530 292046 558598 292102
rect 558654 292046 558722 292102
rect 558778 292046 558846 292102
rect 558902 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 9518 291978
rect 9574 291922 9642 291978
rect 9698 291922 40238 291978
rect 40294 291922 40362 291978
rect 40418 291922 64518 291978
rect 64574 291922 64642 291978
rect 64698 291922 95238 291978
rect 95294 291922 95362 291978
rect 95418 291922 133862 291978
rect 133918 291922 133986 291978
rect 134042 291922 164582 291978
rect 164638 291922 164706 291978
rect 164762 291922 195302 291978
rect 195358 291922 195426 291978
rect 195482 291922 214518 291978
rect 214574 291922 214642 291978
rect 214698 291922 245238 291978
rect 245294 291922 245362 291978
rect 245418 291922 275958 291978
rect 276014 291922 276082 291978
rect 276138 291922 306678 291978
rect 306734 291922 306802 291978
rect 306858 291922 337398 291978
rect 337454 291922 337522 291978
rect 337578 291922 368118 291978
rect 368174 291922 368242 291978
rect 368298 291922 374154 291978
rect 374210 291922 374278 291978
rect 374334 291922 374402 291978
rect 374458 291922 374526 291978
rect 374582 291922 384518 291978
rect 384574 291922 384642 291978
rect 384698 291922 415238 291978
rect 415294 291922 415362 291978
rect 415418 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 466314 291978
rect 466370 291922 466438 291978
rect 466494 291922 466562 291978
rect 466618 291922 466686 291978
rect 466742 291922 497034 291978
rect 497090 291922 497158 291978
rect 497214 291922 497282 291978
rect 497338 291922 497406 291978
rect 497462 291922 527754 291978
rect 527810 291922 527878 291978
rect 527934 291922 528002 291978
rect 528058 291922 528126 291978
rect 528182 291922 558474 291978
rect 558530 291922 558598 291978
rect 558654 291922 558722 291978
rect 558778 291922 558846 291978
rect 558902 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect 4716 290818 7716 290834
rect 4716 290762 4732 290818
rect 4788 290762 7644 290818
rect 7700 290762 7716 290818
rect 4716 290746 7716 290762
rect 197804 287578 199348 287594
rect 197804 287522 197820 287578
rect 197876 287522 199276 287578
rect 199332 287522 199348 287578
rect 197804 287506 199348 287522
rect 58700 287398 68868 287414
rect 58700 287342 58716 287398
rect 58772 287342 68796 287398
rect 68852 287342 68868 287398
rect 58700 287326 68868 287342
rect 77516 286678 106724 286694
rect 77516 286622 77532 286678
rect 77588 286622 106652 286678
rect 106708 286622 106724 286678
rect 77516 286606 106724 286622
rect 58364 286498 120052 286514
rect 58364 286442 58380 286498
rect 58436 286442 119980 286498
rect 120036 286442 120052 286498
rect 58364 286426 120052 286442
rect 380700 286138 387396 286154
rect 380700 286082 380716 286138
rect 380772 286082 387324 286138
rect 387380 286082 387396 286138
rect 380700 286066 387396 286082
rect 58140 284698 121956 284714
rect 58140 284642 58156 284698
rect 58212 284642 121884 284698
rect 121940 284642 121956 284698
rect 58140 284626 121956 284642
rect 58700 283978 119380 283994
rect 58700 283922 58716 283978
rect 58772 283922 119308 283978
rect 119364 283922 119380 283978
rect 58700 283906 119380 283922
rect 57916 283438 121508 283454
rect 57916 283382 57932 283438
rect 57988 283382 121436 283438
rect 121492 283382 121508 283438
rect 57916 283366 121508 283382
rect 58476 283258 141108 283274
rect 58476 283202 58492 283258
rect 58548 283202 141036 283258
rect 141092 283202 141108 283258
rect 58476 283186 141108 283202
rect 56460 283078 139764 283094
rect 56460 283022 56476 283078
rect 56532 283022 139692 283078
rect 139748 283022 139764 283078
rect 56460 283006 139764 283022
rect 58700 282358 122404 282374
rect 58700 282302 58716 282358
rect 58772 282302 122332 282358
rect 122388 282302 122404 282358
rect 58700 282286 122404 282302
rect 58252 282178 146484 282194
rect 58252 282122 58268 282178
rect 58324 282122 146412 282178
rect 146468 282122 146484 282178
rect 58252 282106 146484 282122
rect 193100 282178 194756 282194
rect 193100 282122 193116 282178
rect 193172 282122 194684 282178
rect 194740 282122 194756 282178
rect 193100 282106 194756 282122
rect 56348 281998 163732 282014
rect 56348 281942 56364 281998
rect 56420 281942 163660 281998
rect 163716 281942 163732 281998
rect 56348 281926 163732 281942
rect 5276 281818 121620 281834
rect 5276 281762 5292 281818
rect 5348 281762 121548 281818
rect 121604 281762 121620 281818
rect 5276 281746 121620 281762
rect 3036 281638 127780 281654
rect 3036 281582 3052 281638
rect 3108 281582 127708 281638
rect 127764 281582 127780 281638
rect 3036 281566 127780 281582
rect 5276 281458 133716 281474
rect 5276 281402 5292 281458
rect 5348 281402 133644 281458
rect 133700 281402 133716 281458
rect 5276 281386 133716 281402
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 70674 280350
rect 70730 280294 70798 280350
rect 70854 280294 70922 280350
rect 70978 280294 71046 280350
rect 71102 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 229878 280350
rect 229934 280294 230002 280350
rect 230058 280294 260598 280350
rect 260654 280294 260722 280350
rect 260778 280294 291318 280350
rect 291374 280294 291442 280350
rect 291498 280294 322038 280350
rect 322094 280294 322162 280350
rect 322218 280294 352758 280350
rect 352814 280294 352882 280350
rect 352938 280294 377874 280350
rect 377930 280294 377998 280350
rect 378054 280294 378122 280350
rect 378178 280294 378246 280350
rect 378302 280294 399878 280350
rect 399934 280294 400002 280350
rect 400058 280294 430598 280350
rect 430654 280294 430722 280350
rect 430778 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 470034 280350
rect 470090 280294 470158 280350
rect 470214 280294 470282 280350
rect 470338 280294 470406 280350
rect 470462 280294 500754 280350
rect 500810 280294 500878 280350
rect 500934 280294 501002 280350
rect 501058 280294 501126 280350
rect 501182 280294 531474 280350
rect 531530 280294 531598 280350
rect 531654 280294 531722 280350
rect 531778 280294 531846 280350
rect 531902 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 70674 280226
rect 70730 280170 70798 280226
rect 70854 280170 70922 280226
rect 70978 280170 71046 280226
rect 71102 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 229878 280226
rect 229934 280170 230002 280226
rect 230058 280170 260598 280226
rect 260654 280170 260722 280226
rect 260778 280170 291318 280226
rect 291374 280170 291442 280226
rect 291498 280170 322038 280226
rect 322094 280170 322162 280226
rect 322218 280170 352758 280226
rect 352814 280170 352882 280226
rect 352938 280170 377874 280226
rect 377930 280170 377998 280226
rect 378054 280170 378122 280226
rect 378178 280170 378246 280226
rect 378302 280170 399878 280226
rect 399934 280170 400002 280226
rect 400058 280170 430598 280226
rect 430654 280170 430722 280226
rect 430778 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 470034 280226
rect 470090 280170 470158 280226
rect 470214 280170 470282 280226
rect 470338 280170 470406 280226
rect 470462 280170 500754 280226
rect 500810 280170 500878 280226
rect 500934 280170 501002 280226
rect 501058 280170 501126 280226
rect 501182 280170 531474 280226
rect 531530 280170 531598 280226
rect 531654 280170 531722 280226
rect 531778 280170 531846 280226
rect 531902 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 70674 280102
rect 70730 280046 70798 280102
rect 70854 280046 70922 280102
rect 70978 280046 71046 280102
rect 71102 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 229878 280102
rect 229934 280046 230002 280102
rect 230058 280046 260598 280102
rect 260654 280046 260722 280102
rect 260778 280046 291318 280102
rect 291374 280046 291442 280102
rect 291498 280046 322038 280102
rect 322094 280046 322162 280102
rect 322218 280046 352758 280102
rect 352814 280046 352882 280102
rect 352938 280046 377874 280102
rect 377930 280046 377998 280102
rect 378054 280046 378122 280102
rect 378178 280046 378246 280102
rect 378302 280046 399878 280102
rect 399934 280046 400002 280102
rect 400058 280046 430598 280102
rect 430654 280046 430722 280102
rect 430778 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 470034 280102
rect 470090 280046 470158 280102
rect 470214 280046 470282 280102
rect 470338 280046 470406 280102
rect 470462 280046 500754 280102
rect 500810 280046 500878 280102
rect 500934 280046 501002 280102
rect 501058 280046 501126 280102
rect 501182 280046 531474 280102
rect 531530 280046 531598 280102
rect 531654 280046 531722 280102
rect 531778 280046 531846 280102
rect 531902 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 70674 279978
rect 70730 279922 70798 279978
rect 70854 279922 70922 279978
rect 70978 279922 71046 279978
rect 71102 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 229878 279978
rect 229934 279922 230002 279978
rect 230058 279922 260598 279978
rect 260654 279922 260722 279978
rect 260778 279922 291318 279978
rect 291374 279922 291442 279978
rect 291498 279922 322038 279978
rect 322094 279922 322162 279978
rect 322218 279922 352758 279978
rect 352814 279922 352882 279978
rect 352938 279922 377874 279978
rect 377930 279922 377998 279978
rect 378054 279922 378122 279978
rect 378178 279922 378246 279978
rect 378302 279922 399878 279978
rect 399934 279922 400002 279978
rect 400058 279922 430598 279978
rect 430654 279922 430722 279978
rect 430778 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 470034 279978
rect 470090 279922 470158 279978
rect 470214 279922 470282 279978
rect 470338 279922 470406 279978
rect 470462 279922 500754 279978
rect 500810 279922 500878 279978
rect 500934 279922 501002 279978
rect 501058 279922 501126 279978
rect 501182 279922 531474 279978
rect 531530 279922 531598 279978
rect 531654 279922 531722 279978
rect 531778 279922 531846 279978
rect 531902 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect 106636 279658 201812 279674
rect 106636 279602 106652 279658
rect 106708 279602 201740 279658
rect 201796 279602 201812 279658
rect 106636 279586 201812 279602
rect 108540 279478 202148 279494
rect 108540 279422 108556 279478
rect 108612 279422 202076 279478
rect 202132 279422 202148 279478
rect 108540 279406 202148 279422
rect 118620 278578 155444 278594
rect 118620 278522 118636 278578
rect 118692 278522 155372 278578
rect 155428 278522 155444 278578
rect 118620 278506 155444 278522
rect 109996 278398 174708 278414
rect 109996 278342 110012 278398
rect 110068 278342 174636 278398
rect 174692 278342 174708 278398
rect 109996 278326 174708 278342
rect 74156 278218 110980 278234
rect 74156 278162 74172 278218
rect 74228 278162 110908 278218
rect 110964 278162 110980 278218
rect 74156 278146 110980 278162
rect 120188 278218 187476 278234
rect 120188 278162 120204 278218
rect 120260 278162 187404 278218
rect 187460 278162 187476 278218
rect 120188 278146 187476 278162
rect 4940 278038 137076 278054
rect 4940 277982 4956 278038
rect 5012 277982 137004 278038
rect 137060 277982 137076 278038
rect 4940 277966 137076 277982
rect 7740 277318 63940 277334
rect 7740 277262 7756 277318
rect 7812 277262 63868 277318
rect 63924 277262 63940 277318
rect 7740 277246 63940 277262
rect 115036 277318 175380 277334
rect 115036 277262 115052 277318
rect 115108 277262 175308 277318
rect 175364 277262 175380 277318
rect 115036 277246 175380 277262
rect 45260 277138 63716 277154
rect 45260 277082 45276 277138
rect 45332 277082 63644 277138
rect 63700 277082 63716 277138
rect 45260 277066 63716 277082
rect 118732 277138 165972 277154
rect 118732 277082 118748 277138
rect 118804 277082 165900 277138
rect 165956 277082 165972 277138
rect 118732 277066 165972 277082
rect 209564 277138 213460 277154
rect 209564 277082 209580 277138
rect 209636 277082 213388 277138
rect 213444 277082 213460 277138
rect 209564 277066 213460 277082
rect 48620 276958 73124 276974
rect 48620 276902 48636 276958
rect 48692 276902 63532 276958
rect 63588 276902 73052 276958
rect 73108 276902 73124 276958
rect 48620 276886 73124 276902
rect 119852 276958 165300 276974
rect 119852 276902 119868 276958
rect 119924 276902 165228 276958
rect 165284 276902 165300 276958
rect 119852 276886 165300 276902
rect 64188 276778 70436 276794
rect 64188 276722 64204 276778
rect 64260 276722 70364 276778
rect 70420 276722 70436 276778
rect 64188 276706 70436 276722
rect 119628 276778 160036 276794
rect 119628 276722 119644 276778
rect 119700 276722 159964 276778
rect 160020 276722 160036 276778
rect 119628 276706 160036 276722
rect 189516 276778 212116 276794
rect 189516 276722 189532 276778
rect 189588 276722 212044 276778
rect 212100 276722 212116 276778
rect 189516 276706 212116 276722
rect 48732 276598 62260 276614
rect 48732 276542 48748 276598
rect 48804 276542 62188 276598
rect 62244 276542 62260 276598
rect 48732 276526 62260 276542
rect 119180 276598 158020 276614
rect 119180 276542 119196 276598
rect 119252 276542 157948 276598
rect 158004 276542 158020 276598
rect 119180 276526 158020 276542
rect 189516 276598 209652 276614
rect 189516 276542 189532 276598
rect 189588 276542 209580 276598
rect 209636 276542 209652 276598
rect 189516 276526 209652 276542
rect 209788 276598 212004 276614
rect 209788 276542 211932 276598
rect 211988 276542 212004 276598
rect 209788 276526 212004 276542
rect 209788 276434 209876 276526
rect 58028 276418 74804 276434
rect 58028 276362 58044 276418
rect 58100 276362 74732 276418
rect 74788 276362 74804 276418
rect 58028 276346 74804 276362
rect 120524 276418 151188 276434
rect 120524 276362 120540 276418
rect 120596 276362 151116 276418
rect 151172 276362 151188 276418
rect 120524 276346 151188 276362
rect 173836 276418 209876 276434
rect 173836 276362 173852 276418
rect 173908 276362 209876 276418
rect 173836 276346 209876 276362
rect 210684 276418 213572 276434
rect 210684 276362 210700 276418
rect 210756 276362 213500 276418
rect 213556 276362 213572 276418
rect 210684 276346 213572 276362
rect 63628 276238 69764 276254
rect 63628 276182 63644 276238
rect 63700 276182 69692 276238
rect 69748 276182 69764 276238
rect 63628 276166 69764 276182
rect 60380 276058 70436 276074
rect 60380 276002 60396 276058
rect 60452 276002 70364 276058
rect 70420 276002 70436 276058
rect 60380 275986 70436 276002
rect 7068 275518 63492 275534
rect 7068 275462 7084 275518
rect 7140 275462 63420 275518
rect 63476 275462 63492 275518
rect 7068 275446 63492 275462
rect 111900 274618 202260 274634
rect 111900 274562 111916 274618
rect 111972 274562 202188 274618
rect 202244 274562 202260 274618
rect 111900 274546 202260 274562
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 66954 274350
rect 67010 274294 67078 274350
rect 67134 274294 67202 274350
rect 67258 274294 67326 274350
rect 67382 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 214518 274350
rect 214574 274294 214642 274350
rect 214698 274294 245238 274350
rect 245294 274294 245362 274350
rect 245418 274294 275958 274350
rect 276014 274294 276082 274350
rect 276138 274294 306678 274350
rect 306734 274294 306802 274350
rect 306858 274294 337398 274350
rect 337454 274294 337522 274350
rect 337578 274294 368118 274350
rect 368174 274294 368242 274350
rect 368298 274294 374154 274350
rect 374210 274294 374278 274350
rect 374334 274294 374402 274350
rect 374458 274294 374526 274350
rect 374582 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 466314 274350
rect 466370 274294 466438 274350
rect 466494 274294 466562 274350
rect 466618 274294 466686 274350
rect 466742 274294 497034 274350
rect 497090 274294 497158 274350
rect 497214 274294 497282 274350
rect 497338 274294 497406 274350
rect 497462 274294 527754 274350
rect 527810 274294 527878 274350
rect 527934 274294 528002 274350
rect 528058 274294 528126 274350
rect 528182 274294 558474 274350
rect 558530 274294 558598 274350
rect 558654 274294 558722 274350
rect 558778 274294 558846 274350
rect 558902 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 66954 274226
rect 67010 274170 67078 274226
rect 67134 274170 67202 274226
rect 67258 274170 67326 274226
rect 67382 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 214518 274226
rect 214574 274170 214642 274226
rect 214698 274170 245238 274226
rect 245294 274170 245362 274226
rect 245418 274170 275958 274226
rect 276014 274170 276082 274226
rect 276138 274170 306678 274226
rect 306734 274170 306802 274226
rect 306858 274170 337398 274226
rect 337454 274170 337522 274226
rect 337578 274170 368118 274226
rect 368174 274170 368242 274226
rect 368298 274170 374154 274226
rect 374210 274170 374278 274226
rect 374334 274170 374402 274226
rect 374458 274170 374526 274226
rect 374582 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 466314 274226
rect 466370 274170 466438 274226
rect 466494 274170 466562 274226
rect 466618 274170 466686 274226
rect 466742 274170 497034 274226
rect 497090 274170 497158 274226
rect 497214 274170 497282 274226
rect 497338 274170 497406 274226
rect 497462 274170 527754 274226
rect 527810 274170 527878 274226
rect 527934 274170 528002 274226
rect 528058 274170 528126 274226
rect 528182 274170 558474 274226
rect 558530 274170 558598 274226
rect 558654 274170 558722 274226
rect 558778 274170 558846 274226
rect 558902 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 66954 274102
rect 67010 274046 67078 274102
rect 67134 274046 67202 274102
rect 67258 274046 67326 274102
rect 67382 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 214518 274102
rect 214574 274046 214642 274102
rect 214698 274046 245238 274102
rect 245294 274046 245362 274102
rect 245418 274046 275958 274102
rect 276014 274046 276082 274102
rect 276138 274046 306678 274102
rect 306734 274046 306802 274102
rect 306858 274046 337398 274102
rect 337454 274046 337522 274102
rect 337578 274046 368118 274102
rect 368174 274046 368242 274102
rect 368298 274046 374154 274102
rect 374210 274046 374278 274102
rect 374334 274046 374402 274102
rect 374458 274046 374526 274102
rect 374582 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 466314 274102
rect 466370 274046 466438 274102
rect 466494 274046 466562 274102
rect 466618 274046 466686 274102
rect 466742 274046 497034 274102
rect 497090 274046 497158 274102
rect 497214 274046 497282 274102
rect 497338 274046 497406 274102
rect 497462 274046 527754 274102
rect 527810 274046 527878 274102
rect 527934 274046 528002 274102
rect 528058 274046 528126 274102
rect 528182 274046 558474 274102
rect 558530 274046 558598 274102
rect 558654 274046 558722 274102
rect 558778 274046 558846 274102
rect 558902 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 66954 273978
rect 67010 273922 67078 273978
rect 67134 273922 67202 273978
rect 67258 273922 67326 273978
rect 67382 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 214518 273978
rect 214574 273922 214642 273978
rect 214698 273922 245238 273978
rect 245294 273922 245362 273978
rect 245418 273922 275958 273978
rect 276014 273922 276082 273978
rect 276138 273922 306678 273978
rect 306734 273922 306802 273978
rect 306858 273922 337398 273978
rect 337454 273922 337522 273978
rect 337578 273922 368118 273978
rect 368174 273922 368242 273978
rect 368298 273922 374154 273978
rect 374210 273922 374278 273978
rect 374334 273922 374402 273978
rect 374458 273922 374526 273978
rect 374582 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 466314 273978
rect 466370 273922 466438 273978
rect 466494 273922 466562 273978
rect 466618 273922 466686 273978
rect 466742 273922 497034 273978
rect 497090 273922 497158 273978
rect 497214 273922 497282 273978
rect 497338 273922 497406 273978
rect 497462 273922 527754 273978
rect 527810 273922 527878 273978
rect 527934 273922 528002 273978
rect 528058 273922 528126 273978
rect 528182 273922 558474 273978
rect 558530 273922 558598 273978
rect 558654 273922 558722 273978
rect 558778 273922 558846 273978
rect 558902 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect 2476 273718 186804 273734
rect 2476 273662 2492 273718
rect 2548 273662 186732 273718
rect 186788 273662 186804 273718
rect 2476 273646 186804 273662
rect 12 273538 176052 273554
rect 12 273482 28 273538
rect 84 273482 175980 273538
rect 176036 273482 176052 273538
rect 12 273466 176052 273482
rect 108316 273358 197108 273374
rect 108316 273302 108332 273358
rect 108388 273302 197036 273358
rect 197092 273302 197108 273358
rect 108316 273286 197108 273302
rect 4268 272098 188148 272114
rect 4268 272042 4284 272098
rect 4340 272042 188076 272098
rect 188132 272042 188148 272098
rect 4268 272026 188148 272042
rect 124 271918 184788 271934
rect 124 271862 140 271918
rect 196 271862 184716 271918
rect 184772 271862 184788 271918
rect 124 271846 184788 271862
rect 111676 271738 188820 271754
rect 111676 271682 111692 271738
rect 111748 271682 188748 271738
rect 188804 271682 188820 271738
rect 111676 271666 188820 271682
rect 120076 271558 177396 271574
rect 120076 271502 120092 271558
rect 120148 271502 177324 271558
rect 177380 271502 177396 271558
rect 120076 271486 177396 271502
rect 70348 271378 103588 271394
rect 70348 271322 70364 271378
rect 70420 271322 103516 271378
rect 103572 271322 103588 271378
rect 70348 271306 103588 271322
rect 370844 270658 385492 270674
rect 370844 270602 370860 270658
rect 370916 270602 385420 270658
rect 385476 270602 385492 270658
rect 370844 270586 385492 270602
rect 4380 270478 184900 270494
rect 4380 270422 4396 270478
rect 4452 270422 184828 270478
rect 184884 270422 184900 270478
rect 4380 270406 184900 270422
rect 4156 270298 183220 270314
rect 4156 270242 4172 270298
rect 4228 270242 183148 270298
rect 183204 270242 183220 270298
rect 4156 270226 183220 270242
rect 118844 270118 194644 270134
rect 118844 270062 118860 270118
rect 118916 270062 194572 270118
rect 194628 270062 194644 270118
rect 118844 270046 194644 270062
rect 111788 269938 176612 269954
rect 111788 269882 111804 269938
rect 111860 269882 176540 269938
rect 176596 269882 176612 269938
rect 111788 269866 176612 269882
rect 375436 268858 388068 268874
rect 375436 268802 375452 268858
rect 375508 268802 387996 268858
rect 388052 268802 388068 268858
rect 375436 268786 388068 268802
rect 109996 268498 189492 268514
rect 109996 268442 110012 268498
rect 110068 268442 189420 268498
rect 189476 268442 189492 268498
rect 109996 268426 189492 268442
rect 4268 268318 169332 268334
rect 4268 268262 4284 268318
rect 4340 268262 169260 268318
rect 169316 268262 169332 268318
rect 4268 268246 169332 268262
rect 10876 268138 180084 268154
rect 10876 268082 10892 268138
rect 10948 268082 180012 268138
rect 180068 268082 180084 268138
rect 10876 268066 180084 268082
rect 379916 268138 416404 268154
rect 379916 268082 379932 268138
rect 379988 268082 416332 268138
rect 416388 268082 416404 268138
rect 379916 268066 416404 268082
rect 12 267958 178180 267974
rect 12 267902 28 267958
rect 84 267902 178108 267958
rect 178164 267902 178180 267958
rect 12 267886 178180 267902
rect 379804 267958 424692 267974
rect 379804 267902 379820 267958
rect 379876 267902 424620 267958
rect 424676 267902 424692 267958
rect 379804 267886 424692 267902
rect 378796 267238 420436 267254
rect 378796 267182 378812 267238
rect 378868 267182 420364 267238
rect 420420 267182 420436 267238
rect 378796 267166 420436 267182
rect 108316 266878 190500 266894
rect 108316 266822 108332 266878
rect 108388 266822 190428 266878
rect 190484 266822 190500 266878
rect 108316 266806 190500 266822
rect 4156 266698 163844 266714
rect 4156 266642 4172 266698
rect 4228 266642 163772 266698
rect 163828 266642 163844 266698
rect 4156 266626 163844 266642
rect 124 266518 168212 266534
rect 124 266462 140 266518
rect 196 266462 168140 266518
rect 168196 266462 168212 266518
rect 124 266446 168212 266462
rect 7516 266338 179972 266354
rect 7516 266282 7532 266338
rect 7588 266282 179900 266338
rect 179956 266282 179972 266338
rect 7516 266266 179972 266282
rect 127580 265078 197892 265094
rect 127580 265022 127596 265078
rect 127652 265022 197820 265078
rect 197876 265022 197892 265078
rect 127580 265006 197892 265022
rect 103276 264898 179860 264914
rect 103276 264842 103292 264898
rect 103348 264842 179788 264898
rect 179844 264842 179860 264898
rect 103276 264826 179860 264842
rect 7628 264718 169780 264734
rect 7628 264662 7644 264718
rect 7700 264662 169708 264718
rect 169764 264662 169780 264718
rect 7628 264646 169780 264662
rect 10988 264538 181540 264554
rect 10988 264482 11004 264538
rect 11060 264482 181468 264538
rect 181524 264482 181540 264538
rect 10988 264466 181540 264482
rect 379468 264538 413380 264554
rect 379468 264482 379484 264538
rect 379540 264482 413308 264538
rect 413364 264482 413380 264538
rect 379468 264466 413380 264482
rect 113356 262918 184004 262934
rect 113356 262862 113372 262918
rect 113428 262862 183932 262918
rect 183988 262862 184004 262918
rect 113356 262846 184004 262862
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 70674 262350
rect 70730 262294 70798 262350
rect 70854 262294 70922 262350
rect 70978 262294 71046 262350
rect 71102 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 229878 262350
rect 229934 262294 230002 262350
rect 230058 262294 260598 262350
rect 260654 262294 260722 262350
rect 260778 262294 291318 262350
rect 291374 262294 291442 262350
rect 291498 262294 322038 262350
rect 322094 262294 322162 262350
rect 322218 262294 352758 262350
rect 352814 262294 352882 262350
rect 352938 262294 377874 262350
rect 377930 262294 377998 262350
rect 378054 262294 378122 262350
rect 378178 262294 378246 262350
rect 378302 262294 408594 262350
rect 408650 262294 408718 262350
rect 408774 262294 408842 262350
rect 408898 262294 408966 262350
rect 409022 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 470034 262350
rect 470090 262294 470158 262350
rect 470214 262294 470282 262350
rect 470338 262294 470406 262350
rect 470462 262294 500754 262350
rect 500810 262294 500878 262350
rect 500934 262294 501002 262350
rect 501058 262294 501126 262350
rect 501182 262294 531474 262350
rect 531530 262294 531598 262350
rect 531654 262294 531722 262350
rect 531778 262294 531846 262350
rect 531902 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 70674 262226
rect 70730 262170 70798 262226
rect 70854 262170 70922 262226
rect 70978 262170 71046 262226
rect 71102 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 229878 262226
rect 229934 262170 230002 262226
rect 230058 262170 260598 262226
rect 260654 262170 260722 262226
rect 260778 262170 291318 262226
rect 291374 262170 291442 262226
rect 291498 262170 322038 262226
rect 322094 262170 322162 262226
rect 322218 262170 352758 262226
rect 352814 262170 352882 262226
rect 352938 262170 377874 262226
rect 377930 262170 377998 262226
rect 378054 262170 378122 262226
rect 378178 262170 378246 262226
rect 378302 262170 408594 262226
rect 408650 262170 408718 262226
rect 408774 262170 408842 262226
rect 408898 262170 408966 262226
rect 409022 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 470034 262226
rect 470090 262170 470158 262226
rect 470214 262170 470282 262226
rect 470338 262170 470406 262226
rect 470462 262170 500754 262226
rect 500810 262170 500878 262226
rect 500934 262170 501002 262226
rect 501058 262170 501126 262226
rect 501182 262170 531474 262226
rect 531530 262170 531598 262226
rect 531654 262170 531722 262226
rect 531778 262170 531846 262226
rect 531902 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 70674 262102
rect 70730 262046 70798 262102
rect 70854 262046 70922 262102
rect 70978 262046 71046 262102
rect 71102 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 229878 262102
rect 229934 262046 230002 262102
rect 230058 262046 260598 262102
rect 260654 262046 260722 262102
rect 260778 262046 291318 262102
rect 291374 262046 291442 262102
rect 291498 262046 322038 262102
rect 322094 262046 322162 262102
rect 322218 262046 352758 262102
rect 352814 262046 352882 262102
rect 352938 262046 377874 262102
rect 377930 262046 377998 262102
rect 378054 262046 378122 262102
rect 378178 262046 378246 262102
rect 378302 262046 408594 262102
rect 408650 262046 408718 262102
rect 408774 262046 408842 262102
rect 408898 262046 408966 262102
rect 409022 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 470034 262102
rect 470090 262046 470158 262102
rect 470214 262046 470282 262102
rect 470338 262046 470406 262102
rect 470462 262046 500754 262102
rect 500810 262046 500878 262102
rect 500934 262046 501002 262102
rect 501058 262046 501126 262102
rect 501182 262046 531474 262102
rect 531530 262046 531598 262102
rect 531654 262046 531722 262102
rect 531778 262046 531846 262102
rect 531902 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 70674 261978
rect 70730 261922 70798 261978
rect 70854 261922 70922 261978
rect 70978 261922 71046 261978
rect 71102 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 229878 261978
rect 229934 261922 230002 261978
rect 230058 261922 260598 261978
rect 260654 261922 260722 261978
rect 260778 261922 291318 261978
rect 291374 261922 291442 261978
rect 291498 261922 322038 261978
rect 322094 261922 322162 261978
rect 322218 261922 352758 261978
rect 352814 261922 352882 261978
rect 352938 261922 377874 261978
rect 377930 261922 377998 261978
rect 378054 261922 378122 261978
rect 378178 261922 378246 261978
rect 378302 261922 408594 261978
rect 408650 261922 408718 261978
rect 408774 261922 408842 261978
rect 408898 261922 408966 261978
rect 409022 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 470034 261978
rect 470090 261922 470158 261978
rect 470214 261922 470282 261978
rect 470338 261922 470406 261978
rect 470462 261922 500754 261978
rect 500810 261922 500878 261978
rect 500934 261922 501002 261978
rect 501058 261922 501126 261978
rect 501182 261922 531474 261978
rect 531530 261922 531598 261978
rect 531654 261922 531722 261978
rect 531778 261922 531846 261978
rect 531902 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect 112684 261658 173924 261674
rect 112684 261602 112700 261658
rect 112756 261602 173852 261658
rect 173908 261602 173924 261658
rect 112684 261586 173924 261602
rect 377564 261658 387508 261674
rect 377564 261602 377580 261658
rect 377636 261602 387436 261658
rect 387492 261602 387508 261658
rect 377564 261586 387508 261602
rect 379580 261298 403636 261314
rect 379580 261242 379596 261298
rect 379652 261242 403564 261298
rect 403620 261242 403636 261298
rect 379580 261226 403636 261242
rect 61388 260398 187364 260414
rect 61388 260342 61404 260398
rect 61460 260342 186172 260398
rect 186228 260342 187292 260398
rect 187348 260342 187364 260398
rect 61388 260326 187364 260342
rect 377116 260398 383924 260414
rect 377116 260342 377132 260398
rect 377188 260342 383852 260398
rect 383908 260342 383924 260398
rect 377116 260326 383924 260342
rect 4940 257878 160596 257894
rect 4940 257822 4956 257878
rect 5012 257822 160524 257878
rect 160580 257822 160596 257878
rect 4940 257806 160596 257822
rect 210684 257878 211892 257894
rect 210684 257822 210700 257878
rect 210756 257822 211820 257878
rect 211876 257822 211892 257878
rect 210684 257806 211892 257822
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 13760 256350
rect 13816 256294 13884 256350
rect 13940 256294 14008 256350
rect 14064 256294 14132 256350
rect 14188 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 66954 256350
rect 67010 256294 67078 256350
rect 67134 256294 67202 256350
rect 67258 256294 67326 256350
rect 67382 256294 98442 256350
rect 98498 256294 98566 256350
rect 98622 256294 98690 256350
rect 98746 256294 98814 256350
rect 98870 256294 113760 256350
rect 113816 256294 113884 256350
rect 113940 256294 114008 256350
rect 114064 256294 114132 256350
rect 114188 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 198442 256350
rect 198498 256294 198566 256350
rect 198622 256294 198690 256350
rect 198746 256294 198814 256350
rect 198870 256294 214518 256350
rect 214574 256294 214642 256350
rect 214698 256294 245238 256350
rect 245294 256294 245362 256350
rect 245418 256294 275958 256350
rect 276014 256294 276082 256350
rect 276138 256294 306678 256350
rect 306734 256294 306802 256350
rect 306858 256294 337398 256350
rect 337454 256294 337522 256350
rect 337578 256294 368118 256350
rect 368174 256294 368242 256350
rect 368298 256294 374154 256350
rect 374210 256294 374278 256350
rect 374334 256294 374402 256350
rect 374458 256294 374526 256350
rect 374582 256294 384518 256350
rect 384574 256294 384642 256350
rect 384698 256294 415238 256350
rect 415294 256294 415362 256350
rect 415418 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 466314 256350
rect 466370 256294 466438 256350
rect 466494 256294 466562 256350
rect 466618 256294 466686 256350
rect 466742 256294 497034 256350
rect 497090 256294 497158 256350
rect 497214 256294 497282 256350
rect 497338 256294 497406 256350
rect 497462 256294 527754 256350
rect 527810 256294 527878 256350
rect 527934 256294 528002 256350
rect 528058 256294 528126 256350
rect 528182 256294 558474 256350
rect 558530 256294 558598 256350
rect 558654 256294 558722 256350
rect 558778 256294 558846 256350
rect 558902 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 13760 256226
rect 13816 256170 13884 256226
rect 13940 256170 14008 256226
rect 14064 256170 14132 256226
rect 14188 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 66954 256226
rect 67010 256170 67078 256226
rect 67134 256170 67202 256226
rect 67258 256170 67326 256226
rect 67382 256170 98442 256226
rect 98498 256170 98566 256226
rect 98622 256170 98690 256226
rect 98746 256170 98814 256226
rect 98870 256170 113760 256226
rect 113816 256170 113884 256226
rect 113940 256170 114008 256226
rect 114064 256170 114132 256226
rect 114188 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 198442 256226
rect 198498 256170 198566 256226
rect 198622 256170 198690 256226
rect 198746 256170 198814 256226
rect 198870 256170 214518 256226
rect 214574 256170 214642 256226
rect 214698 256170 245238 256226
rect 245294 256170 245362 256226
rect 245418 256170 275958 256226
rect 276014 256170 276082 256226
rect 276138 256170 306678 256226
rect 306734 256170 306802 256226
rect 306858 256170 337398 256226
rect 337454 256170 337522 256226
rect 337578 256170 368118 256226
rect 368174 256170 368242 256226
rect 368298 256170 374154 256226
rect 374210 256170 374278 256226
rect 374334 256170 374402 256226
rect 374458 256170 374526 256226
rect 374582 256170 384518 256226
rect 384574 256170 384642 256226
rect 384698 256170 415238 256226
rect 415294 256170 415362 256226
rect 415418 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 466314 256226
rect 466370 256170 466438 256226
rect 466494 256170 466562 256226
rect 466618 256170 466686 256226
rect 466742 256170 497034 256226
rect 497090 256170 497158 256226
rect 497214 256170 497282 256226
rect 497338 256170 497406 256226
rect 497462 256170 527754 256226
rect 527810 256170 527878 256226
rect 527934 256170 528002 256226
rect 528058 256170 528126 256226
rect 528182 256170 558474 256226
rect 558530 256170 558598 256226
rect 558654 256170 558722 256226
rect 558778 256170 558846 256226
rect 558902 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 13760 256102
rect 13816 256046 13884 256102
rect 13940 256046 14008 256102
rect 14064 256046 14132 256102
rect 14188 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 66954 256102
rect 67010 256046 67078 256102
rect 67134 256046 67202 256102
rect 67258 256046 67326 256102
rect 67382 256046 98442 256102
rect 98498 256046 98566 256102
rect 98622 256046 98690 256102
rect 98746 256046 98814 256102
rect 98870 256046 113760 256102
rect 113816 256046 113884 256102
rect 113940 256046 114008 256102
rect 114064 256046 114132 256102
rect 114188 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 198442 256102
rect 198498 256046 198566 256102
rect 198622 256046 198690 256102
rect 198746 256046 198814 256102
rect 198870 256046 214518 256102
rect 214574 256046 214642 256102
rect 214698 256046 245238 256102
rect 245294 256046 245362 256102
rect 245418 256046 275958 256102
rect 276014 256046 276082 256102
rect 276138 256046 306678 256102
rect 306734 256046 306802 256102
rect 306858 256046 337398 256102
rect 337454 256046 337522 256102
rect 337578 256046 368118 256102
rect 368174 256046 368242 256102
rect 368298 256046 374154 256102
rect 374210 256046 374278 256102
rect 374334 256046 374402 256102
rect 374458 256046 374526 256102
rect 374582 256046 384518 256102
rect 384574 256046 384642 256102
rect 384698 256046 415238 256102
rect 415294 256046 415362 256102
rect 415418 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 466314 256102
rect 466370 256046 466438 256102
rect 466494 256046 466562 256102
rect 466618 256046 466686 256102
rect 466742 256046 497034 256102
rect 497090 256046 497158 256102
rect 497214 256046 497282 256102
rect 497338 256046 497406 256102
rect 497462 256046 527754 256102
rect 527810 256046 527878 256102
rect 527934 256046 528002 256102
rect 528058 256046 528126 256102
rect 528182 256046 558474 256102
rect 558530 256046 558598 256102
rect 558654 256046 558722 256102
rect 558778 256046 558846 256102
rect 558902 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 13760 255978
rect 13816 255922 13884 255978
rect 13940 255922 14008 255978
rect 14064 255922 14132 255978
rect 14188 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 66954 255978
rect 67010 255922 67078 255978
rect 67134 255922 67202 255978
rect 67258 255922 67326 255978
rect 67382 255922 98442 255978
rect 98498 255922 98566 255978
rect 98622 255922 98690 255978
rect 98746 255922 98814 255978
rect 98870 255922 113760 255978
rect 113816 255922 113884 255978
rect 113940 255922 114008 255978
rect 114064 255922 114132 255978
rect 114188 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 198442 255978
rect 198498 255922 198566 255978
rect 198622 255922 198690 255978
rect 198746 255922 198814 255978
rect 198870 255922 214518 255978
rect 214574 255922 214642 255978
rect 214698 255922 245238 255978
rect 245294 255922 245362 255978
rect 245418 255922 275958 255978
rect 276014 255922 276082 255978
rect 276138 255922 306678 255978
rect 306734 255922 306802 255978
rect 306858 255922 337398 255978
rect 337454 255922 337522 255978
rect 337578 255922 368118 255978
rect 368174 255922 368242 255978
rect 368298 255922 374154 255978
rect 374210 255922 374278 255978
rect 374334 255922 374402 255978
rect 374458 255922 374526 255978
rect 374582 255922 384518 255978
rect 384574 255922 384642 255978
rect 384698 255922 415238 255978
rect 415294 255922 415362 255978
rect 415418 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 466314 255978
rect 466370 255922 466438 255978
rect 466494 255922 466562 255978
rect 466618 255922 466686 255978
rect 466742 255922 497034 255978
rect 497090 255922 497158 255978
rect 497214 255922 497282 255978
rect 497338 255922 497406 255978
rect 497462 255922 527754 255978
rect 527810 255922 527878 255978
rect 527934 255922 528002 255978
rect 528058 255922 528126 255978
rect 528182 255922 558474 255978
rect 558530 255922 558598 255978
rect 558654 255922 558722 255978
rect 558778 255922 558846 255978
rect 558902 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect 115036 255358 168100 255374
rect 115036 255302 115052 255358
rect 115108 255302 168028 255358
rect 168084 255302 168100 255358
rect 115036 255286 168100 255302
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 12960 244350
rect 13016 244294 13084 244350
rect 13140 244294 13208 244350
rect 13264 244294 13332 244350
rect 13388 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 97642 244350
rect 97698 244294 97766 244350
rect 97822 244294 97890 244350
rect 97946 244294 98014 244350
rect 98070 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 112960 244350
rect 113016 244294 113084 244350
rect 113140 244294 113208 244350
rect 113264 244294 113332 244350
rect 113388 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 197642 244350
rect 197698 244294 197766 244350
rect 197822 244294 197890 244350
rect 197946 244294 198014 244350
rect 198070 244294 229878 244350
rect 229934 244294 230002 244350
rect 230058 244294 260598 244350
rect 260654 244294 260722 244350
rect 260778 244294 291318 244350
rect 291374 244294 291442 244350
rect 291498 244294 322038 244350
rect 322094 244294 322162 244350
rect 322218 244294 352758 244350
rect 352814 244294 352882 244350
rect 352938 244294 377874 244350
rect 377930 244294 377998 244350
rect 378054 244294 378122 244350
rect 378178 244294 378246 244350
rect 378302 244294 399878 244350
rect 399934 244294 400002 244350
rect 400058 244294 430598 244350
rect 430654 244294 430722 244350
rect 430778 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 470034 244350
rect 470090 244294 470158 244350
rect 470214 244294 470282 244350
rect 470338 244294 470406 244350
rect 470462 244294 500754 244350
rect 500810 244294 500878 244350
rect 500934 244294 501002 244350
rect 501058 244294 501126 244350
rect 501182 244294 531474 244350
rect 531530 244294 531598 244350
rect 531654 244294 531722 244350
rect 531778 244294 531846 244350
rect 531902 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 12960 244226
rect 13016 244170 13084 244226
rect 13140 244170 13208 244226
rect 13264 244170 13332 244226
rect 13388 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 97642 244226
rect 97698 244170 97766 244226
rect 97822 244170 97890 244226
rect 97946 244170 98014 244226
rect 98070 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 112960 244226
rect 113016 244170 113084 244226
rect 113140 244170 113208 244226
rect 113264 244170 113332 244226
rect 113388 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 197642 244226
rect 197698 244170 197766 244226
rect 197822 244170 197890 244226
rect 197946 244170 198014 244226
rect 198070 244170 229878 244226
rect 229934 244170 230002 244226
rect 230058 244170 260598 244226
rect 260654 244170 260722 244226
rect 260778 244170 291318 244226
rect 291374 244170 291442 244226
rect 291498 244170 322038 244226
rect 322094 244170 322162 244226
rect 322218 244170 352758 244226
rect 352814 244170 352882 244226
rect 352938 244170 377874 244226
rect 377930 244170 377998 244226
rect 378054 244170 378122 244226
rect 378178 244170 378246 244226
rect 378302 244170 399878 244226
rect 399934 244170 400002 244226
rect 400058 244170 430598 244226
rect 430654 244170 430722 244226
rect 430778 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 470034 244226
rect 470090 244170 470158 244226
rect 470214 244170 470282 244226
rect 470338 244170 470406 244226
rect 470462 244170 500754 244226
rect 500810 244170 500878 244226
rect 500934 244170 501002 244226
rect 501058 244170 501126 244226
rect 501182 244170 531474 244226
rect 531530 244170 531598 244226
rect 531654 244170 531722 244226
rect 531778 244170 531846 244226
rect 531902 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 12960 244102
rect 13016 244046 13084 244102
rect 13140 244046 13208 244102
rect 13264 244046 13332 244102
rect 13388 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 97642 244102
rect 97698 244046 97766 244102
rect 97822 244046 97890 244102
rect 97946 244046 98014 244102
rect 98070 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 112960 244102
rect 113016 244046 113084 244102
rect 113140 244046 113208 244102
rect 113264 244046 113332 244102
rect 113388 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 197642 244102
rect 197698 244046 197766 244102
rect 197822 244046 197890 244102
rect 197946 244046 198014 244102
rect 198070 244046 229878 244102
rect 229934 244046 230002 244102
rect 230058 244046 260598 244102
rect 260654 244046 260722 244102
rect 260778 244046 291318 244102
rect 291374 244046 291442 244102
rect 291498 244046 322038 244102
rect 322094 244046 322162 244102
rect 322218 244046 352758 244102
rect 352814 244046 352882 244102
rect 352938 244046 377874 244102
rect 377930 244046 377998 244102
rect 378054 244046 378122 244102
rect 378178 244046 378246 244102
rect 378302 244046 399878 244102
rect 399934 244046 400002 244102
rect 400058 244046 430598 244102
rect 430654 244046 430722 244102
rect 430778 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 470034 244102
rect 470090 244046 470158 244102
rect 470214 244046 470282 244102
rect 470338 244046 470406 244102
rect 470462 244046 500754 244102
rect 500810 244046 500878 244102
rect 500934 244046 501002 244102
rect 501058 244046 501126 244102
rect 501182 244046 531474 244102
rect 531530 244046 531598 244102
rect 531654 244046 531722 244102
rect 531778 244046 531846 244102
rect 531902 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 12960 243978
rect 13016 243922 13084 243978
rect 13140 243922 13208 243978
rect 13264 243922 13332 243978
rect 13388 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 97642 243978
rect 97698 243922 97766 243978
rect 97822 243922 97890 243978
rect 97946 243922 98014 243978
rect 98070 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 112960 243978
rect 113016 243922 113084 243978
rect 113140 243922 113208 243978
rect 113264 243922 113332 243978
rect 113388 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 197642 243978
rect 197698 243922 197766 243978
rect 197822 243922 197890 243978
rect 197946 243922 198014 243978
rect 198070 243922 229878 243978
rect 229934 243922 230002 243978
rect 230058 243922 260598 243978
rect 260654 243922 260722 243978
rect 260778 243922 291318 243978
rect 291374 243922 291442 243978
rect 291498 243922 322038 243978
rect 322094 243922 322162 243978
rect 322218 243922 352758 243978
rect 352814 243922 352882 243978
rect 352938 243922 377874 243978
rect 377930 243922 377998 243978
rect 378054 243922 378122 243978
rect 378178 243922 378246 243978
rect 378302 243922 399878 243978
rect 399934 243922 400002 243978
rect 400058 243922 430598 243978
rect 430654 243922 430722 243978
rect 430778 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 470034 243978
rect 470090 243922 470158 243978
rect 470214 243922 470282 243978
rect 470338 243922 470406 243978
rect 470462 243922 500754 243978
rect 500810 243922 500878 243978
rect 500934 243922 501002 243978
rect 501058 243922 501126 243978
rect 501182 243922 531474 243978
rect 531530 243922 531598 243978
rect 531654 243922 531722 243978
rect 531778 243922 531846 243978
rect 531902 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect 430988 242758 440260 242774
rect 430988 242702 431004 242758
rect 431060 242702 436828 242758
rect 436884 242702 440188 242758
rect 440244 242702 440260 242758
rect 430988 242686 440260 242702
rect 380028 241858 381572 241874
rect 380028 241802 380044 241858
rect 380100 241802 381500 241858
rect 381556 241802 381572 241858
rect 380028 241786 381572 241802
rect 434236 240058 440036 240074
rect 434236 240002 434252 240058
rect 434308 240002 439964 240058
rect 440020 240002 440036 240058
rect 434236 239986 440036 240002
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 13760 238350
rect 13816 238294 13884 238350
rect 13940 238294 14008 238350
rect 14064 238294 14132 238350
rect 14188 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 98442 238350
rect 98498 238294 98566 238350
rect 98622 238294 98690 238350
rect 98746 238294 98814 238350
rect 98870 238294 113760 238350
rect 113816 238294 113884 238350
rect 113940 238294 114008 238350
rect 114064 238294 114132 238350
rect 114188 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 198442 238350
rect 198498 238294 198566 238350
rect 198622 238294 198690 238350
rect 198746 238294 198814 238350
rect 198870 238294 214518 238350
rect 214574 238294 214642 238350
rect 214698 238294 245238 238350
rect 245294 238294 245362 238350
rect 245418 238294 275958 238350
rect 276014 238294 276082 238350
rect 276138 238294 306678 238350
rect 306734 238294 306802 238350
rect 306858 238294 337398 238350
rect 337454 238294 337522 238350
rect 337578 238294 368118 238350
rect 368174 238294 368242 238350
rect 368298 238294 374154 238350
rect 374210 238294 374278 238350
rect 374334 238294 374402 238350
rect 374458 238294 374526 238350
rect 374582 238294 384518 238350
rect 384574 238294 384642 238350
rect 384698 238294 415238 238350
rect 415294 238294 415362 238350
rect 415418 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 466314 238350
rect 466370 238294 466438 238350
rect 466494 238294 466562 238350
rect 466618 238294 466686 238350
rect 466742 238294 497034 238350
rect 497090 238294 497158 238350
rect 497214 238294 497282 238350
rect 497338 238294 497406 238350
rect 497462 238294 527754 238350
rect 527810 238294 527878 238350
rect 527934 238294 528002 238350
rect 528058 238294 528126 238350
rect 528182 238294 558474 238350
rect 558530 238294 558598 238350
rect 558654 238294 558722 238350
rect 558778 238294 558846 238350
rect 558902 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 13760 238226
rect 13816 238170 13884 238226
rect 13940 238170 14008 238226
rect 14064 238170 14132 238226
rect 14188 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 98442 238226
rect 98498 238170 98566 238226
rect 98622 238170 98690 238226
rect 98746 238170 98814 238226
rect 98870 238170 113760 238226
rect 113816 238170 113884 238226
rect 113940 238170 114008 238226
rect 114064 238170 114132 238226
rect 114188 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 198442 238226
rect 198498 238170 198566 238226
rect 198622 238170 198690 238226
rect 198746 238170 198814 238226
rect 198870 238170 214518 238226
rect 214574 238170 214642 238226
rect 214698 238170 245238 238226
rect 245294 238170 245362 238226
rect 245418 238170 275958 238226
rect 276014 238170 276082 238226
rect 276138 238170 306678 238226
rect 306734 238170 306802 238226
rect 306858 238170 337398 238226
rect 337454 238170 337522 238226
rect 337578 238170 368118 238226
rect 368174 238170 368242 238226
rect 368298 238170 374154 238226
rect 374210 238170 374278 238226
rect 374334 238170 374402 238226
rect 374458 238170 374526 238226
rect 374582 238170 384518 238226
rect 384574 238170 384642 238226
rect 384698 238170 415238 238226
rect 415294 238170 415362 238226
rect 415418 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 466314 238226
rect 466370 238170 466438 238226
rect 466494 238170 466562 238226
rect 466618 238170 466686 238226
rect 466742 238170 497034 238226
rect 497090 238170 497158 238226
rect 497214 238170 497282 238226
rect 497338 238170 497406 238226
rect 497462 238170 527754 238226
rect 527810 238170 527878 238226
rect 527934 238170 528002 238226
rect 528058 238170 528126 238226
rect 528182 238170 558474 238226
rect 558530 238170 558598 238226
rect 558654 238170 558722 238226
rect 558778 238170 558846 238226
rect 558902 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 13760 238102
rect 13816 238046 13884 238102
rect 13940 238046 14008 238102
rect 14064 238046 14132 238102
rect 14188 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 98442 238102
rect 98498 238046 98566 238102
rect 98622 238046 98690 238102
rect 98746 238046 98814 238102
rect 98870 238046 113760 238102
rect 113816 238046 113884 238102
rect 113940 238046 114008 238102
rect 114064 238046 114132 238102
rect 114188 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 198442 238102
rect 198498 238046 198566 238102
rect 198622 238046 198690 238102
rect 198746 238046 198814 238102
rect 198870 238046 214518 238102
rect 214574 238046 214642 238102
rect 214698 238046 245238 238102
rect 245294 238046 245362 238102
rect 245418 238046 275958 238102
rect 276014 238046 276082 238102
rect 276138 238046 306678 238102
rect 306734 238046 306802 238102
rect 306858 238046 337398 238102
rect 337454 238046 337522 238102
rect 337578 238046 368118 238102
rect 368174 238046 368242 238102
rect 368298 238046 374154 238102
rect 374210 238046 374278 238102
rect 374334 238046 374402 238102
rect 374458 238046 374526 238102
rect 374582 238046 384518 238102
rect 384574 238046 384642 238102
rect 384698 238046 415238 238102
rect 415294 238046 415362 238102
rect 415418 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 466314 238102
rect 466370 238046 466438 238102
rect 466494 238046 466562 238102
rect 466618 238046 466686 238102
rect 466742 238046 497034 238102
rect 497090 238046 497158 238102
rect 497214 238046 497282 238102
rect 497338 238046 497406 238102
rect 497462 238046 527754 238102
rect 527810 238046 527878 238102
rect 527934 238046 528002 238102
rect 528058 238046 528126 238102
rect 528182 238046 558474 238102
rect 558530 238046 558598 238102
rect 558654 238046 558722 238102
rect 558778 238046 558846 238102
rect 558902 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 13760 237978
rect 13816 237922 13884 237978
rect 13940 237922 14008 237978
rect 14064 237922 14132 237978
rect 14188 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 98442 237978
rect 98498 237922 98566 237978
rect 98622 237922 98690 237978
rect 98746 237922 98814 237978
rect 98870 237922 113760 237978
rect 113816 237922 113884 237978
rect 113940 237922 114008 237978
rect 114064 237922 114132 237978
rect 114188 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 198442 237978
rect 198498 237922 198566 237978
rect 198622 237922 198690 237978
rect 198746 237922 198814 237978
rect 198870 237922 214518 237978
rect 214574 237922 214642 237978
rect 214698 237922 245238 237978
rect 245294 237922 245362 237978
rect 245418 237922 275958 237978
rect 276014 237922 276082 237978
rect 276138 237922 306678 237978
rect 306734 237922 306802 237978
rect 306858 237922 337398 237978
rect 337454 237922 337522 237978
rect 337578 237922 368118 237978
rect 368174 237922 368242 237978
rect 368298 237922 374154 237978
rect 374210 237922 374278 237978
rect 374334 237922 374402 237978
rect 374458 237922 374526 237978
rect 374582 237922 384518 237978
rect 384574 237922 384642 237978
rect 384698 237922 415238 237978
rect 415294 237922 415362 237978
rect 415418 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 466314 237978
rect 466370 237922 466438 237978
rect 466494 237922 466562 237978
rect 466618 237922 466686 237978
rect 466742 237922 497034 237978
rect 497090 237922 497158 237978
rect 497214 237922 497282 237978
rect 497338 237922 497406 237978
rect 497462 237922 527754 237978
rect 527810 237922 527878 237978
rect 527934 237922 528002 237978
rect 528058 237922 528126 237978
rect 528182 237922 558474 237978
rect 558530 237922 558598 237978
rect 558654 237922 558722 237978
rect 558778 237922 558846 237978
rect 558902 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect 210684 236098 211780 236114
rect 210684 236042 210700 236098
rect 210756 236042 211708 236098
rect 211764 236042 211780 236098
rect 210684 236026 211780 236042
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 12960 226350
rect 13016 226294 13084 226350
rect 13140 226294 13208 226350
rect 13264 226294 13332 226350
rect 13388 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 97642 226350
rect 97698 226294 97766 226350
rect 97822 226294 97890 226350
rect 97946 226294 98014 226350
rect 98070 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 112960 226350
rect 113016 226294 113084 226350
rect 113140 226294 113208 226350
rect 113264 226294 113332 226350
rect 113388 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 197642 226350
rect 197698 226294 197766 226350
rect 197822 226294 197890 226350
rect 197946 226294 198014 226350
rect 198070 226294 229878 226350
rect 229934 226294 230002 226350
rect 230058 226294 260598 226350
rect 260654 226294 260722 226350
rect 260778 226294 291318 226350
rect 291374 226294 291442 226350
rect 291498 226294 322038 226350
rect 322094 226294 322162 226350
rect 322218 226294 352758 226350
rect 352814 226294 352882 226350
rect 352938 226294 377874 226350
rect 377930 226294 377998 226350
rect 378054 226294 378122 226350
rect 378178 226294 378246 226350
rect 378302 226294 399878 226350
rect 399934 226294 400002 226350
rect 400058 226294 430598 226350
rect 430654 226294 430722 226350
rect 430778 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 470034 226350
rect 470090 226294 470158 226350
rect 470214 226294 470282 226350
rect 470338 226294 470406 226350
rect 470462 226294 500754 226350
rect 500810 226294 500878 226350
rect 500934 226294 501002 226350
rect 501058 226294 501126 226350
rect 501182 226294 531474 226350
rect 531530 226294 531598 226350
rect 531654 226294 531722 226350
rect 531778 226294 531846 226350
rect 531902 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 12960 226226
rect 13016 226170 13084 226226
rect 13140 226170 13208 226226
rect 13264 226170 13332 226226
rect 13388 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 97642 226226
rect 97698 226170 97766 226226
rect 97822 226170 97890 226226
rect 97946 226170 98014 226226
rect 98070 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 112960 226226
rect 113016 226170 113084 226226
rect 113140 226170 113208 226226
rect 113264 226170 113332 226226
rect 113388 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 197642 226226
rect 197698 226170 197766 226226
rect 197822 226170 197890 226226
rect 197946 226170 198014 226226
rect 198070 226170 229878 226226
rect 229934 226170 230002 226226
rect 230058 226170 260598 226226
rect 260654 226170 260722 226226
rect 260778 226170 291318 226226
rect 291374 226170 291442 226226
rect 291498 226170 322038 226226
rect 322094 226170 322162 226226
rect 322218 226170 352758 226226
rect 352814 226170 352882 226226
rect 352938 226170 377874 226226
rect 377930 226170 377998 226226
rect 378054 226170 378122 226226
rect 378178 226170 378246 226226
rect 378302 226170 399878 226226
rect 399934 226170 400002 226226
rect 400058 226170 430598 226226
rect 430654 226170 430722 226226
rect 430778 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 470034 226226
rect 470090 226170 470158 226226
rect 470214 226170 470282 226226
rect 470338 226170 470406 226226
rect 470462 226170 500754 226226
rect 500810 226170 500878 226226
rect 500934 226170 501002 226226
rect 501058 226170 501126 226226
rect 501182 226170 531474 226226
rect 531530 226170 531598 226226
rect 531654 226170 531722 226226
rect 531778 226170 531846 226226
rect 531902 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 12960 226102
rect 13016 226046 13084 226102
rect 13140 226046 13208 226102
rect 13264 226046 13332 226102
rect 13388 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 97642 226102
rect 97698 226046 97766 226102
rect 97822 226046 97890 226102
rect 97946 226046 98014 226102
rect 98070 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 112960 226102
rect 113016 226046 113084 226102
rect 113140 226046 113208 226102
rect 113264 226046 113332 226102
rect 113388 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 197642 226102
rect 197698 226046 197766 226102
rect 197822 226046 197890 226102
rect 197946 226046 198014 226102
rect 198070 226046 229878 226102
rect 229934 226046 230002 226102
rect 230058 226046 260598 226102
rect 260654 226046 260722 226102
rect 260778 226046 291318 226102
rect 291374 226046 291442 226102
rect 291498 226046 322038 226102
rect 322094 226046 322162 226102
rect 322218 226046 352758 226102
rect 352814 226046 352882 226102
rect 352938 226046 377874 226102
rect 377930 226046 377998 226102
rect 378054 226046 378122 226102
rect 378178 226046 378246 226102
rect 378302 226046 399878 226102
rect 399934 226046 400002 226102
rect 400058 226046 430598 226102
rect 430654 226046 430722 226102
rect 430778 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 470034 226102
rect 470090 226046 470158 226102
rect 470214 226046 470282 226102
rect 470338 226046 470406 226102
rect 470462 226046 500754 226102
rect 500810 226046 500878 226102
rect 500934 226046 501002 226102
rect 501058 226046 501126 226102
rect 501182 226046 531474 226102
rect 531530 226046 531598 226102
rect 531654 226046 531722 226102
rect 531778 226046 531846 226102
rect 531902 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 12960 225978
rect 13016 225922 13084 225978
rect 13140 225922 13208 225978
rect 13264 225922 13332 225978
rect 13388 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 97642 225978
rect 97698 225922 97766 225978
rect 97822 225922 97890 225978
rect 97946 225922 98014 225978
rect 98070 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 112960 225978
rect 113016 225922 113084 225978
rect 113140 225922 113208 225978
rect 113264 225922 113332 225978
rect 113388 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 197642 225978
rect 197698 225922 197766 225978
rect 197822 225922 197890 225978
rect 197946 225922 198014 225978
rect 198070 225922 229878 225978
rect 229934 225922 230002 225978
rect 230058 225922 260598 225978
rect 260654 225922 260722 225978
rect 260778 225922 291318 225978
rect 291374 225922 291442 225978
rect 291498 225922 322038 225978
rect 322094 225922 322162 225978
rect 322218 225922 352758 225978
rect 352814 225922 352882 225978
rect 352938 225922 377874 225978
rect 377930 225922 377998 225978
rect 378054 225922 378122 225978
rect 378178 225922 378246 225978
rect 378302 225922 399878 225978
rect 399934 225922 400002 225978
rect 400058 225922 430598 225978
rect 430654 225922 430722 225978
rect 430778 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 470034 225978
rect 470090 225922 470158 225978
rect 470214 225922 470282 225978
rect 470338 225922 470406 225978
rect 470462 225922 500754 225978
rect 500810 225922 500878 225978
rect 500934 225922 501002 225978
rect 501058 225922 501126 225978
rect 501182 225922 531474 225978
rect 531530 225922 531598 225978
rect 531654 225922 531722 225978
rect 531778 225922 531846 225978
rect 531902 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect 187388 225118 192404 225134
rect 187388 225062 187404 225118
rect 187460 225062 192332 225118
rect 192388 225062 192404 225118
rect 187388 225046 192404 225062
rect 192316 223498 205060 223514
rect 192316 223442 192332 223498
rect 192388 223442 204988 223498
rect 205044 223442 205060 223498
rect 192316 223426 205060 223442
rect 183916 222598 205060 222614
rect 183916 222542 183932 222598
rect 183988 222542 184716 222598
rect 184772 222542 204988 222598
rect 205044 222542 205060 222598
rect 183916 222526 205060 222542
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 13760 220350
rect 13816 220294 13884 220350
rect 13940 220294 14008 220350
rect 14064 220294 14132 220350
rect 14188 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 98442 220350
rect 98498 220294 98566 220350
rect 98622 220294 98690 220350
rect 98746 220294 98814 220350
rect 98870 220294 113760 220350
rect 113816 220294 113884 220350
rect 113940 220294 114008 220350
rect 114064 220294 114132 220350
rect 114188 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 198442 220350
rect 198498 220294 198566 220350
rect 198622 220294 198690 220350
rect 198746 220294 198814 220350
rect 198870 220294 214518 220350
rect 214574 220294 214642 220350
rect 214698 220294 245238 220350
rect 245294 220294 245362 220350
rect 245418 220294 275958 220350
rect 276014 220294 276082 220350
rect 276138 220294 306678 220350
rect 306734 220294 306802 220350
rect 306858 220294 337398 220350
rect 337454 220294 337522 220350
rect 337578 220294 368118 220350
rect 368174 220294 368242 220350
rect 368298 220294 374154 220350
rect 374210 220294 374278 220350
rect 374334 220294 374402 220350
rect 374458 220294 374526 220350
rect 374582 220294 384518 220350
rect 384574 220294 384642 220350
rect 384698 220294 415238 220350
rect 415294 220294 415362 220350
rect 415418 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 466314 220350
rect 466370 220294 466438 220350
rect 466494 220294 466562 220350
rect 466618 220294 466686 220350
rect 466742 220294 497034 220350
rect 497090 220294 497158 220350
rect 497214 220294 497282 220350
rect 497338 220294 497406 220350
rect 497462 220294 527754 220350
rect 527810 220294 527878 220350
rect 527934 220294 528002 220350
rect 528058 220294 528126 220350
rect 528182 220294 558474 220350
rect 558530 220294 558598 220350
rect 558654 220294 558722 220350
rect 558778 220294 558846 220350
rect 558902 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 13760 220226
rect 13816 220170 13884 220226
rect 13940 220170 14008 220226
rect 14064 220170 14132 220226
rect 14188 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 98442 220226
rect 98498 220170 98566 220226
rect 98622 220170 98690 220226
rect 98746 220170 98814 220226
rect 98870 220170 113760 220226
rect 113816 220170 113884 220226
rect 113940 220170 114008 220226
rect 114064 220170 114132 220226
rect 114188 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 198442 220226
rect 198498 220170 198566 220226
rect 198622 220170 198690 220226
rect 198746 220170 198814 220226
rect 198870 220170 214518 220226
rect 214574 220170 214642 220226
rect 214698 220170 245238 220226
rect 245294 220170 245362 220226
rect 245418 220170 275958 220226
rect 276014 220170 276082 220226
rect 276138 220170 306678 220226
rect 306734 220170 306802 220226
rect 306858 220170 337398 220226
rect 337454 220170 337522 220226
rect 337578 220170 368118 220226
rect 368174 220170 368242 220226
rect 368298 220170 374154 220226
rect 374210 220170 374278 220226
rect 374334 220170 374402 220226
rect 374458 220170 374526 220226
rect 374582 220170 384518 220226
rect 384574 220170 384642 220226
rect 384698 220170 415238 220226
rect 415294 220170 415362 220226
rect 415418 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 466314 220226
rect 466370 220170 466438 220226
rect 466494 220170 466562 220226
rect 466618 220170 466686 220226
rect 466742 220170 497034 220226
rect 497090 220170 497158 220226
rect 497214 220170 497282 220226
rect 497338 220170 497406 220226
rect 497462 220170 527754 220226
rect 527810 220170 527878 220226
rect 527934 220170 528002 220226
rect 528058 220170 528126 220226
rect 528182 220170 558474 220226
rect 558530 220170 558598 220226
rect 558654 220170 558722 220226
rect 558778 220170 558846 220226
rect 558902 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 13760 220102
rect 13816 220046 13884 220102
rect 13940 220046 14008 220102
rect 14064 220046 14132 220102
rect 14188 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 98442 220102
rect 98498 220046 98566 220102
rect 98622 220046 98690 220102
rect 98746 220046 98814 220102
rect 98870 220046 113760 220102
rect 113816 220046 113884 220102
rect 113940 220046 114008 220102
rect 114064 220046 114132 220102
rect 114188 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 198442 220102
rect 198498 220046 198566 220102
rect 198622 220046 198690 220102
rect 198746 220046 198814 220102
rect 198870 220046 214518 220102
rect 214574 220046 214642 220102
rect 214698 220046 245238 220102
rect 245294 220046 245362 220102
rect 245418 220046 275958 220102
rect 276014 220046 276082 220102
rect 276138 220046 306678 220102
rect 306734 220046 306802 220102
rect 306858 220046 337398 220102
rect 337454 220046 337522 220102
rect 337578 220046 368118 220102
rect 368174 220046 368242 220102
rect 368298 220046 374154 220102
rect 374210 220046 374278 220102
rect 374334 220046 374402 220102
rect 374458 220046 374526 220102
rect 374582 220046 384518 220102
rect 384574 220046 384642 220102
rect 384698 220046 415238 220102
rect 415294 220046 415362 220102
rect 415418 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 466314 220102
rect 466370 220046 466438 220102
rect 466494 220046 466562 220102
rect 466618 220046 466686 220102
rect 466742 220046 497034 220102
rect 497090 220046 497158 220102
rect 497214 220046 497282 220102
rect 497338 220046 497406 220102
rect 497462 220046 527754 220102
rect 527810 220046 527878 220102
rect 527934 220046 528002 220102
rect 528058 220046 528126 220102
rect 528182 220046 558474 220102
rect 558530 220046 558598 220102
rect 558654 220046 558722 220102
rect 558778 220046 558846 220102
rect 558902 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 13760 219978
rect 13816 219922 13884 219978
rect 13940 219922 14008 219978
rect 14064 219922 14132 219978
rect 14188 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 98442 219978
rect 98498 219922 98566 219978
rect 98622 219922 98690 219978
rect 98746 219922 98814 219978
rect 98870 219922 113760 219978
rect 113816 219922 113884 219978
rect 113940 219922 114008 219978
rect 114064 219922 114132 219978
rect 114188 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 198442 219978
rect 198498 219922 198566 219978
rect 198622 219922 198690 219978
rect 198746 219922 198814 219978
rect 198870 219922 214518 219978
rect 214574 219922 214642 219978
rect 214698 219922 245238 219978
rect 245294 219922 245362 219978
rect 245418 219922 275958 219978
rect 276014 219922 276082 219978
rect 276138 219922 306678 219978
rect 306734 219922 306802 219978
rect 306858 219922 337398 219978
rect 337454 219922 337522 219978
rect 337578 219922 368118 219978
rect 368174 219922 368242 219978
rect 368298 219922 374154 219978
rect 374210 219922 374278 219978
rect 374334 219922 374402 219978
rect 374458 219922 374526 219978
rect 374582 219922 384518 219978
rect 384574 219922 384642 219978
rect 384698 219922 415238 219978
rect 415294 219922 415362 219978
rect 415418 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 466314 219978
rect 466370 219922 466438 219978
rect 466494 219922 466562 219978
rect 466618 219922 466686 219978
rect 466742 219922 497034 219978
rect 497090 219922 497158 219978
rect 497214 219922 497282 219978
rect 497338 219922 497406 219978
rect 497462 219922 527754 219978
rect 527810 219922 527878 219978
rect 527934 219922 528002 219978
rect 528058 219922 528126 219978
rect 528182 219922 558474 219978
rect 558530 219922 558598 219978
rect 558654 219922 558722 219978
rect 558778 219922 558846 219978
rect 558902 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect 183020 219178 206740 219194
rect 183020 219122 183036 219178
rect 183092 219122 206668 219178
rect 206724 219122 206740 219178
rect 183020 219106 206740 219122
rect 373868 218458 381460 218474
rect 373868 218402 373884 218458
rect 373940 218402 381388 218458
rect 381444 218402 381460 218458
rect 373868 218386 381460 218402
rect 176412 218278 206740 218294
rect 176412 218222 176428 218278
rect 176484 218222 206668 218278
rect 206724 218222 206740 218278
rect 176412 218206 206740 218222
rect 379692 217738 383924 217754
rect 379692 217682 379708 217738
rect 379764 217682 383852 217738
rect 383908 217682 383924 217738
rect 379692 217666 383924 217682
rect 372860 217558 384148 217574
rect 372860 217502 372876 217558
rect 372932 217502 384076 217558
rect 384132 217502 384148 217558
rect 372860 217486 384148 217502
rect 384676 217378 445412 217394
rect 384676 217322 445340 217378
rect 445396 217322 445412 217378
rect 384676 217306 445412 217322
rect 384676 217214 384764 217306
rect 379468 217198 384764 217214
rect 379468 217142 379484 217198
rect 379540 217142 384764 217198
rect 379468 217126 384764 217142
rect 376108 217018 381796 217034
rect 376108 216962 376124 217018
rect 376180 216962 381724 217018
rect 381780 216962 381796 217018
rect 376108 216946 381796 216962
rect 380364 216838 381572 216854
rect 380364 216782 380380 216838
rect 380436 216782 381500 216838
rect 381556 216782 381572 216838
rect 380364 216766 381572 216782
rect 369388 216658 373844 216674
rect 369388 216602 369404 216658
rect 369460 216602 373772 216658
rect 373828 216602 373844 216658
rect 369388 216586 373844 216602
rect 379468 216658 443620 216674
rect 379468 216602 443548 216658
rect 443604 216602 443620 216658
rect 379468 216586 443620 216602
rect 379468 216478 379556 216586
rect 379468 216422 379484 216478
rect 379540 216422 379556 216478
rect 379468 216406 379556 216422
rect 380364 216478 445300 216494
rect 380364 216422 380380 216478
rect 380436 216422 445228 216478
rect 445284 216422 445300 216478
rect 380364 216406 445300 216422
rect 381372 215938 442164 215954
rect 381372 215882 381388 215938
rect 381444 215882 442092 215938
rect 442148 215882 442164 215938
rect 381372 215866 442164 215882
rect 379244 215578 382132 215594
rect 379244 215522 379260 215578
rect 379316 215522 382060 215578
rect 382116 215522 382132 215578
rect 379244 215506 382132 215522
rect 379468 215398 381908 215414
rect 379468 215342 379484 215398
rect 379540 215342 381836 215398
rect 381892 215342 381908 215398
rect 379468 215326 381908 215342
rect 380252 215218 381684 215234
rect 380252 215162 380268 215218
rect 380324 215162 381612 215218
rect 381668 215162 381684 215218
rect 380252 215146 381684 215162
rect 172996 215038 206740 215054
rect 172996 214982 206668 215038
rect 206724 214982 206740 215038
rect 172996 214966 206740 214982
rect 172996 214154 173084 214966
rect 373644 214318 395796 214334
rect 373644 214262 373660 214318
rect 373716 214262 395724 214318
rect 395780 214262 395796 214318
rect 373644 214246 395796 214262
rect 160508 214138 173084 214154
rect 160508 214082 160524 214138
rect 160580 214082 168028 214138
rect 168084 214082 173084 214138
rect 160508 214066 173084 214082
rect 378684 214138 442612 214154
rect 378684 214082 378700 214138
rect 378756 214082 442540 214138
rect 442596 214082 442612 214138
rect 378684 214066 442612 214082
rect 380252 213598 382020 213614
rect 380252 213542 380268 213598
rect 380324 213542 381948 213598
rect 382004 213542 382020 213598
rect 380252 213526 382020 213542
rect 373868 213418 418420 213434
rect 373868 213362 373884 213418
rect 373940 213362 418348 213418
rect 418404 213362 418420 213418
rect 373868 213346 418420 213362
rect 374988 213238 382580 213254
rect 374988 213182 375004 213238
rect 375060 213182 382508 213238
rect 382564 213182 382580 213238
rect 374988 213166 382580 213182
rect 173836 212518 206740 212534
rect 173836 212462 173852 212518
rect 173908 212462 206668 212518
rect 206724 212462 206740 212518
rect 173836 212446 206740 212462
rect 379692 212518 442724 212534
rect 379692 212462 379708 212518
rect 379764 212462 442652 212518
rect 442708 212462 442724 212518
rect 379692 212446 442724 212462
rect 375660 212158 386836 212174
rect 375660 212102 375676 212158
rect 375732 212102 386764 212158
rect 386820 212102 386836 212158
rect 375660 212086 386836 212102
rect 373868 211978 392324 211994
rect 373868 211922 373884 211978
rect 373940 211922 392252 211978
rect 392308 211922 392324 211978
rect 373868 211906 392324 211922
rect 380252 211798 383476 211814
rect 380252 211742 380268 211798
rect 380324 211742 383404 211798
rect 383460 211742 383476 211798
rect 380252 211726 383476 211742
rect 378908 211078 389524 211094
rect 378908 211022 378924 211078
rect 378980 211022 389452 211078
rect 389508 211022 389524 211078
rect 378908 211006 389524 211022
rect 372412 210898 386164 210914
rect 372412 210842 372428 210898
rect 372484 210842 386092 210898
rect 386148 210842 386164 210898
rect 372412 210826 386164 210842
rect 177196 209998 206740 210014
rect 177196 209942 177212 209998
rect 177268 209942 178892 209998
rect 178948 209942 206668 209998
rect 206724 209942 206740 209998
rect 177196 209926 206740 209942
rect 372748 209278 380340 209294
rect 372748 209222 372764 209278
rect 372820 209222 380268 209278
rect 380324 209222 380340 209278
rect 372748 209206 380340 209222
rect 370956 209098 381236 209114
rect 370956 209042 370972 209098
rect 371028 209042 381164 209098
rect 381220 209042 381236 209098
rect 370956 209026 381236 209042
rect -1916 208393 597980 208446
rect -1916 208350 399836 208393
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 12960 208350
rect 13016 208294 13084 208350
rect 13140 208294 13208 208350
rect 13264 208294 13332 208350
rect 13388 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 70674 208350
rect 70730 208294 70798 208350
rect 70854 208294 70922 208350
rect 70978 208294 71046 208350
rect 71102 208294 97642 208350
rect 97698 208294 97766 208350
rect 97822 208294 97890 208350
rect 97946 208294 98014 208350
rect 98070 208294 101394 208350
rect 101450 208294 101518 208350
rect 101574 208294 101642 208350
rect 101698 208294 101766 208350
rect 101822 208294 112960 208350
rect 113016 208294 113084 208350
rect 113140 208294 113208 208350
rect 113264 208294 113332 208350
rect 113388 208294 132114 208350
rect 132170 208294 132238 208350
rect 132294 208294 132362 208350
rect 132418 208294 132486 208350
rect 132542 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 193554 208350
rect 193610 208294 193678 208350
rect 193734 208294 193802 208350
rect 193858 208294 193926 208350
rect 193982 208294 197642 208350
rect 197698 208294 197766 208350
rect 197822 208294 197890 208350
rect 197946 208294 198014 208350
rect 198070 208294 229878 208350
rect 229934 208294 230002 208350
rect 230058 208294 260598 208350
rect 260654 208294 260722 208350
rect 260778 208294 291318 208350
rect 291374 208294 291442 208350
rect 291498 208294 322038 208350
rect 322094 208294 322162 208350
rect 322218 208294 352758 208350
rect 352814 208294 352882 208350
rect 352938 208294 377874 208350
rect 377930 208294 377998 208350
rect 378054 208294 378122 208350
rect 378178 208294 378246 208350
rect 378302 208337 399836 208350
rect 399892 208337 399940 208393
rect 399996 208337 400044 208393
rect 400100 208350 430556 208393
rect 400100 208337 408594 208350
rect 378302 208294 408594 208337
rect 408650 208294 408718 208350
rect 408774 208294 408842 208350
rect 408898 208294 408966 208350
rect 409022 208337 430556 208350
rect 430612 208337 430660 208393
rect 430716 208337 430764 208393
rect 430820 208350 597980 208393
rect 430820 208337 439314 208350
rect 409022 208294 439314 208337
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 470034 208350
rect 470090 208294 470158 208350
rect 470214 208294 470282 208350
rect 470338 208294 470406 208350
rect 470462 208294 500754 208350
rect 500810 208294 500878 208350
rect 500934 208294 501002 208350
rect 501058 208294 501126 208350
rect 501182 208294 531474 208350
rect 531530 208294 531598 208350
rect 531654 208294 531722 208350
rect 531778 208294 531846 208350
rect 531902 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208289 597980 208294
rect -1916 208233 399836 208289
rect 399892 208233 399940 208289
rect 399996 208233 400044 208289
rect 400100 208233 430556 208289
rect 430612 208233 430660 208289
rect 430716 208233 430764 208289
rect 430820 208233 597980 208289
rect -1916 208226 597980 208233
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 12960 208226
rect 13016 208170 13084 208226
rect 13140 208170 13208 208226
rect 13264 208170 13332 208226
rect 13388 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 70674 208226
rect 70730 208170 70798 208226
rect 70854 208170 70922 208226
rect 70978 208170 71046 208226
rect 71102 208170 97642 208226
rect 97698 208170 97766 208226
rect 97822 208170 97890 208226
rect 97946 208170 98014 208226
rect 98070 208170 101394 208226
rect 101450 208170 101518 208226
rect 101574 208170 101642 208226
rect 101698 208170 101766 208226
rect 101822 208170 112960 208226
rect 113016 208170 113084 208226
rect 113140 208170 113208 208226
rect 113264 208170 113332 208226
rect 113388 208170 132114 208226
rect 132170 208170 132238 208226
rect 132294 208170 132362 208226
rect 132418 208170 132486 208226
rect 132542 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 193554 208226
rect 193610 208170 193678 208226
rect 193734 208170 193802 208226
rect 193858 208170 193926 208226
rect 193982 208170 197642 208226
rect 197698 208170 197766 208226
rect 197822 208170 197890 208226
rect 197946 208170 198014 208226
rect 198070 208170 229878 208226
rect 229934 208170 230002 208226
rect 230058 208170 260598 208226
rect 260654 208170 260722 208226
rect 260778 208170 291318 208226
rect 291374 208170 291442 208226
rect 291498 208170 322038 208226
rect 322094 208170 322162 208226
rect 322218 208170 352758 208226
rect 352814 208170 352882 208226
rect 352938 208170 377874 208226
rect 377930 208170 377998 208226
rect 378054 208170 378122 208226
rect 378178 208170 378246 208226
rect 378302 208185 408594 208226
rect 378302 208170 399836 208185
rect -1916 208129 399836 208170
rect 399892 208129 399940 208185
rect 399996 208129 400044 208185
rect 400100 208170 408594 208185
rect 408650 208170 408718 208226
rect 408774 208170 408842 208226
rect 408898 208170 408966 208226
rect 409022 208185 439314 208226
rect 409022 208170 430556 208185
rect 400100 208129 430556 208170
rect 430612 208129 430660 208185
rect 430716 208129 430764 208185
rect 430820 208170 439314 208185
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 470034 208226
rect 470090 208170 470158 208226
rect 470214 208170 470282 208226
rect 470338 208170 470406 208226
rect 470462 208170 500754 208226
rect 500810 208170 500878 208226
rect 500934 208170 501002 208226
rect 501058 208170 501126 208226
rect 501182 208170 531474 208226
rect 531530 208170 531598 208226
rect 531654 208170 531722 208226
rect 531778 208170 531846 208226
rect 531902 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 430820 208129 597980 208170
rect -1916 208102 597980 208129
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 12960 208102
rect 13016 208046 13084 208102
rect 13140 208046 13208 208102
rect 13264 208046 13332 208102
rect 13388 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 70674 208102
rect 70730 208046 70798 208102
rect 70854 208046 70922 208102
rect 70978 208046 71046 208102
rect 71102 208046 97642 208102
rect 97698 208046 97766 208102
rect 97822 208046 97890 208102
rect 97946 208046 98014 208102
rect 98070 208046 101394 208102
rect 101450 208046 101518 208102
rect 101574 208046 101642 208102
rect 101698 208046 101766 208102
rect 101822 208046 112960 208102
rect 113016 208046 113084 208102
rect 113140 208046 113208 208102
rect 113264 208046 113332 208102
rect 113388 208046 132114 208102
rect 132170 208046 132238 208102
rect 132294 208046 132362 208102
rect 132418 208046 132486 208102
rect 132542 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 193554 208102
rect 193610 208046 193678 208102
rect 193734 208046 193802 208102
rect 193858 208046 193926 208102
rect 193982 208046 197642 208102
rect 197698 208046 197766 208102
rect 197822 208046 197890 208102
rect 197946 208046 198014 208102
rect 198070 208046 229878 208102
rect 229934 208046 230002 208102
rect 230058 208046 260598 208102
rect 260654 208046 260722 208102
rect 260778 208046 291318 208102
rect 291374 208046 291442 208102
rect 291498 208046 322038 208102
rect 322094 208046 322162 208102
rect 322218 208046 352758 208102
rect 352814 208046 352882 208102
rect 352938 208046 377874 208102
rect 377930 208046 377998 208102
rect 378054 208046 378122 208102
rect 378178 208046 378246 208102
rect 378302 208046 408594 208102
rect 408650 208046 408718 208102
rect 408774 208046 408842 208102
rect 408898 208046 408966 208102
rect 409022 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 470034 208102
rect 470090 208046 470158 208102
rect 470214 208046 470282 208102
rect 470338 208046 470406 208102
rect 470462 208046 500754 208102
rect 500810 208046 500878 208102
rect 500934 208046 501002 208102
rect 501058 208046 501126 208102
rect 501182 208046 531474 208102
rect 531530 208046 531598 208102
rect 531654 208046 531722 208102
rect 531778 208046 531846 208102
rect 531902 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 12960 207978
rect 13016 207922 13084 207978
rect 13140 207922 13208 207978
rect 13264 207922 13332 207978
rect 13388 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 70674 207978
rect 70730 207922 70798 207978
rect 70854 207922 70922 207978
rect 70978 207922 71046 207978
rect 71102 207922 97642 207978
rect 97698 207922 97766 207978
rect 97822 207922 97890 207978
rect 97946 207922 98014 207978
rect 98070 207922 101394 207978
rect 101450 207922 101518 207978
rect 101574 207922 101642 207978
rect 101698 207922 101766 207978
rect 101822 207922 112960 207978
rect 113016 207922 113084 207978
rect 113140 207922 113208 207978
rect 113264 207922 113332 207978
rect 113388 207922 132114 207978
rect 132170 207922 132238 207978
rect 132294 207922 132362 207978
rect 132418 207922 132486 207978
rect 132542 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 193554 207978
rect 193610 207922 193678 207978
rect 193734 207922 193802 207978
rect 193858 207922 193926 207978
rect 193982 207922 197642 207978
rect 197698 207922 197766 207978
rect 197822 207922 197890 207978
rect 197946 207922 198014 207978
rect 198070 207922 229878 207978
rect 229934 207922 230002 207978
rect 230058 207922 260598 207978
rect 260654 207922 260722 207978
rect 260778 207922 291318 207978
rect 291374 207922 291442 207978
rect 291498 207922 322038 207978
rect 322094 207922 322162 207978
rect 322218 207922 352758 207978
rect 352814 207922 352882 207978
rect 352938 207922 377874 207978
rect 377930 207922 377998 207978
rect 378054 207922 378122 207978
rect 378178 207922 378246 207978
rect 378302 207922 408594 207978
rect 408650 207922 408718 207978
rect 408774 207922 408842 207978
rect 408898 207922 408966 207978
rect 409022 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 470034 207978
rect 470090 207922 470158 207978
rect 470214 207922 470282 207978
rect 470338 207922 470406 207978
rect 470462 207922 500754 207978
rect 500810 207922 500878 207978
rect 500934 207922 501002 207978
rect 501058 207922 501126 207978
rect 501182 207922 531474 207978
rect 531530 207922 531598 207978
rect 531654 207922 531722 207978
rect 531778 207922 531846 207978
rect 531902 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect 4156 206578 111764 206594
rect 4156 206522 4172 206578
rect 4228 206522 111692 206578
rect 111748 206522 111764 206578
rect 4156 206506 111764 206522
rect 103612 205858 126044 205874
rect 103612 205802 103628 205858
rect 103684 205802 120092 205858
rect 120148 205802 126044 205858
rect 103612 205786 126044 205802
rect 125956 205154 126044 205786
rect 125956 205138 202484 205154
rect 125956 205082 202412 205138
rect 202468 205082 202484 205138
rect 125956 205066 202484 205082
rect 94876 204958 204948 204974
rect 94876 204902 94892 204958
rect 94948 204902 204876 204958
rect 204932 204902 204948 204958
rect 94876 204886 204948 204902
rect 402204 204058 432196 204074
rect 402204 204002 402220 204058
rect 402276 204002 432124 204058
rect 432180 204002 432196 204058
rect 402204 203986 432196 204002
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 13760 202350
rect 13816 202294 13884 202350
rect 13940 202294 14008 202350
rect 14064 202294 14132 202350
rect 14188 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 66954 202350
rect 67010 202294 67078 202350
rect 67134 202294 67202 202350
rect 67258 202294 67326 202350
rect 67382 202294 98442 202350
rect 98498 202294 98566 202350
rect 98622 202294 98690 202350
rect 98746 202294 98814 202350
rect 98870 202294 113760 202350
rect 113816 202294 113884 202350
rect 113940 202294 114008 202350
rect 114064 202294 114132 202350
rect 114188 202294 128394 202350
rect 128450 202294 128518 202350
rect 128574 202294 128642 202350
rect 128698 202294 128766 202350
rect 128822 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 189834 202350
rect 189890 202294 189958 202350
rect 190014 202294 190082 202350
rect 190138 202294 190206 202350
rect 190262 202294 198442 202350
rect 198498 202294 198566 202350
rect 198622 202294 198690 202350
rect 198746 202294 198814 202350
rect 198870 202294 214518 202350
rect 214574 202294 214642 202350
rect 214698 202294 245238 202350
rect 245294 202294 245362 202350
rect 245418 202294 275958 202350
rect 276014 202294 276082 202350
rect 276138 202294 306678 202350
rect 306734 202294 306802 202350
rect 306858 202294 337398 202350
rect 337454 202294 337522 202350
rect 337578 202294 368118 202350
rect 368174 202294 368242 202350
rect 368298 202294 374154 202350
rect 374210 202294 374278 202350
rect 374334 202294 374402 202350
rect 374458 202294 374526 202350
rect 374582 202294 404874 202350
rect 404930 202294 404998 202350
rect 405054 202294 405122 202350
rect 405178 202294 405246 202350
rect 405302 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 466314 202350
rect 466370 202294 466438 202350
rect 466494 202294 466562 202350
rect 466618 202294 466686 202350
rect 466742 202294 497034 202350
rect 497090 202294 497158 202350
rect 497214 202294 497282 202350
rect 497338 202294 497406 202350
rect 497462 202294 527754 202350
rect 527810 202294 527878 202350
rect 527934 202294 528002 202350
rect 528058 202294 528126 202350
rect 528182 202294 558474 202350
rect 558530 202294 558598 202350
rect 558654 202294 558722 202350
rect 558778 202294 558846 202350
rect 558902 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 13760 202226
rect 13816 202170 13884 202226
rect 13940 202170 14008 202226
rect 14064 202170 14132 202226
rect 14188 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 66954 202226
rect 67010 202170 67078 202226
rect 67134 202170 67202 202226
rect 67258 202170 67326 202226
rect 67382 202170 98442 202226
rect 98498 202170 98566 202226
rect 98622 202170 98690 202226
rect 98746 202170 98814 202226
rect 98870 202170 113760 202226
rect 113816 202170 113884 202226
rect 113940 202170 114008 202226
rect 114064 202170 114132 202226
rect 114188 202170 128394 202226
rect 128450 202170 128518 202226
rect 128574 202170 128642 202226
rect 128698 202170 128766 202226
rect 128822 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 189834 202226
rect 189890 202170 189958 202226
rect 190014 202170 190082 202226
rect 190138 202170 190206 202226
rect 190262 202170 198442 202226
rect 198498 202170 198566 202226
rect 198622 202170 198690 202226
rect 198746 202170 198814 202226
rect 198870 202170 214518 202226
rect 214574 202170 214642 202226
rect 214698 202170 245238 202226
rect 245294 202170 245362 202226
rect 245418 202170 275958 202226
rect 276014 202170 276082 202226
rect 276138 202170 306678 202226
rect 306734 202170 306802 202226
rect 306858 202170 337398 202226
rect 337454 202170 337522 202226
rect 337578 202170 368118 202226
rect 368174 202170 368242 202226
rect 368298 202170 374154 202226
rect 374210 202170 374278 202226
rect 374334 202170 374402 202226
rect 374458 202170 374526 202226
rect 374582 202170 404874 202226
rect 404930 202170 404998 202226
rect 405054 202170 405122 202226
rect 405178 202170 405246 202226
rect 405302 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 466314 202226
rect 466370 202170 466438 202226
rect 466494 202170 466562 202226
rect 466618 202170 466686 202226
rect 466742 202170 497034 202226
rect 497090 202170 497158 202226
rect 497214 202170 497282 202226
rect 497338 202170 497406 202226
rect 497462 202170 527754 202226
rect 527810 202170 527878 202226
rect 527934 202170 528002 202226
rect 528058 202170 528126 202226
rect 528182 202170 558474 202226
rect 558530 202170 558598 202226
rect 558654 202170 558722 202226
rect 558778 202170 558846 202226
rect 558902 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 13760 202102
rect 13816 202046 13884 202102
rect 13940 202046 14008 202102
rect 14064 202046 14132 202102
rect 14188 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 66954 202102
rect 67010 202046 67078 202102
rect 67134 202046 67202 202102
rect 67258 202046 67326 202102
rect 67382 202046 98442 202102
rect 98498 202046 98566 202102
rect 98622 202046 98690 202102
rect 98746 202046 98814 202102
rect 98870 202046 113760 202102
rect 113816 202046 113884 202102
rect 113940 202046 114008 202102
rect 114064 202046 114132 202102
rect 114188 202046 128394 202102
rect 128450 202046 128518 202102
rect 128574 202046 128642 202102
rect 128698 202046 128766 202102
rect 128822 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 189834 202102
rect 189890 202046 189958 202102
rect 190014 202046 190082 202102
rect 190138 202046 190206 202102
rect 190262 202046 198442 202102
rect 198498 202046 198566 202102
rect 198622 202046 198690 202102
rect 198746 202046 198814 202102
rect 198870 202046 214518 202102
rect 214574 202046 214642 202102
rect 214698 202046 245238 202102
rect 245294 202046 245362 202102
rect 245418 202046 275958 202102
rect 276014 202046 276082 202102
rect 276138 202046 306678 202102
rect 306734 202046 306802 202102
rect 306858 202046 337398 202102
rect 337454 202046 337522 202102
rect 337578 202046 368118 202102
rect 368174 202046 368242 202102
rect 368298 202046 374154 202102
rect 374210 202046 374278 202102
rect 374334 202046 374402 202102
rect 374458 202046 374526 202102
rect 374582 202046 404874 202102
rect 404930 202046 404998 202102
rect 405054 202046 405122 202102
rect 405178 202046 405246 202102
rect 405302 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 466314 202102
rect 466370 202046 466438 202102
rect 466494 202046 466562 202102
rect 466618 202046 466686 202102
rect 466742 202046 497034 202102
rect 497090 202046 497158 202102
rect 497214 202046 497282 202102
rect 497338 202046 497406 202102
rect 497462 202046 527754 202102
rect 527810 202046 527878 202102
rect 527934 202046 528002 202102
rect 528058 202046 528126 202102
rect 528182 202046 558474 202102
rect 558530 202046 558598 202102
rect 558654 202046 558722 202102
rect 558778 202046 558846 202102
rect 558902 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 13760 201978
rect 13816 201922 13884 201978
rect 13940 201922 14008 201978
rect 14064 201922 14132 201978
rect 14188 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 66954 201978
rect 67010 201922 67078 201978
rect 67134 201922 67202 201978
rect 67258 201922 67326 201978
rect 67382 201922 98442 201978
rect 98498 201922 98566 201978
rect 98622 201922 98690 201978
rect 98746 201922 98814 201978
rect 98870 201922 113760 201978
rect 113816 201922 113884 201978
rect 113940 201922 114008 201978
rect 114064 201922 114132 201978
rect 114188 201922 128394 201978
rect 128450 201922 128518 201978
rect 128574 201922 128642 201978
rect 128698 201922 128766 201978
rect 128822 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 189834 201978
rect 189890 201922 189958 201978
rect 190014 201922 190082 201978
rect 190138 201922 190206 201978
rect 190262 201922 198442 201978
rect 198498 201922 198566 201978
rect 198622 201922 198690 201978
rect 198746 201922 198814 201978
rect 198870 201922 214518 201978
rect 214574 201922 214642 201978
rect 214698 201922 245238 201978
rect 245294 201922 245362 201978
rect 245418 201922 275958 201978
rect 276014 201922 276082 201978
rect 276138 201922 306678 201978
rect 306734 201922 306802 201978
rect 306858 201922 337398 201978
rect 337454 201922 337522 201978
rect 337578 201922 368118 201978
rect 368174 201922 368242 201978
rect 368298 201922 374154 201978
rect 374210 201922 374278 201978
rect 374334 201922 374402 201978
rect 374458 201922 374526 201978
rect 374582 201922 404874 201978
rect 404930 201922 404998 201978
rect 405054 201922 405122 201978
rect 405178 201922 405246 201978
rect 405302 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 466314 201978
rect 466370 201922 466438 201978
rect 466494 201922 466562 201978
rect 466618 201922 466686 201978
rect 466742 201922 497034 201978
rect 497090 201922 497158 201978
rect 497214 201922 497282 201978
rect 497338 201922 497406 201978
rect 497462 201922 527754 201978
rect 527810 201922 527878 201978
rect 527934 201922 528002 201978
rect 528058 201922 528126 201978
rect 528182 201922 558474 201978
rect 558530 201922 558598 201978
rect 558654 201922 558722 201978
rect 558778 201922 558846 201978
rect 558902 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect 84796 201538 205060 201554
rect 84796 201482 84812 201538
rect 84868 201482 186284 201538
rect 186340 201482 204988 201538
rect 205044 201482 205060 201538
rect 84796 201466 205060 201482
rect 82220 199018 206740 199034
rect 82220 198962 82236 199018
rect 82292 198962 206668 199018
rect 206724 198962 206740 199018
rect 82220 198946 206740 198962
rect 389772 198118 430180 198134
rect 389772 198062 389788 198118
rect 389844 198062 430108 198118
rect 430164 198062 430180 198118
rect 389772 198046 430180 198062
rect 72140 195778 206964 195794
rect 72140 195722 72156 195778
rect 72212 195722 206892 195778
rect 206948 195722 206964 195778
rect 72140 195706 206964 195722
rect 369500 193978 426764 193994
rect 369500 193922 369516 193978
rect 369572 193922 426764 193978
rect 369500 193906 426764 193922
rect 426676 193274 426764 193906
rect 426676 193258 442052 193274
rect 426676 193202 441980 193258
rect 442036 193202 442052 193258
rect 426676 193186 442052 193202
rect 39660 193078 205284 193094
rect 39660 193022 39676 193078
rect 39732 193022 205212 193078
rect 205268 193022 205284 193078
rect 39660 193006 205284 193022
rect 28460 191458 205060 191474
rect 28460 191402 28476 191458
rect 28532 191402 186396 191458
rect 186452 191402 204988 191458
rect 205044 191402 205060 191458
rect 28460 191386 205060 191402
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 12960 190350
rect 13016 190294 13084 190350
rect 13140 190294 13208 190350
rect 13264 190294 13332 190350
rect 13388 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 70674 190350
rect 70730 190294 70798 190350
rect 70854 190294 70922 190350
rect 70978 190294 71046 190350
rect 71102 190294 97642 190350
rect 97698 190294 97766 190350
rect 97822 190294 97890 190350
rect 97946 190294 98014 190350
rect 98070 190294 101394 190350
rect 101450 190294 101518 190350
rect 101574 190294 101642 190350
rect 101698 190294 101766 190350
rect 101822 190294 112960 190350
rect 113016 190294 113084 190350
rect 113140 190294 113208 190350
rect 113264 190294 113332 190350
rect 113388 190294 132114 190350
rect 132170 190294 132238 190350
rect 132294 190294 132362 190350
rect 132418 190294 132486 190350
rect 132542 190294 162834 190350
rect 162890 190294 162958 190350
rect 163014 190294 163082 190350
rect 163138 190294 163206 190350
rect 163262 190294 193554 190350
rect 193610 190294 193678 190350
rect 193734 190294 193802 190350
rect 193858 190294 193926 190350
rect 193982 190294 197642 190350
rect 197698 190294 197766 190350
rect 197822 190294 197890 190350
rect 197946 190294 198014 190350
rect 198070 190294 229878 190350
rect 229934 190294 230002 190350
rect 230058 190294 260598 190350
rect 260654 190294 260722 190350
rect 260778 190294 291318 190350
rect 291374 190294 291442 190350
rect 291498 190294 322038 190350
rect 322094 190294 322162 190350
rect 322218 190294 352758 190350
rect 352814 190294 352882 190350
rect 352938 190294 377874 190350
rect 377930 190294 377998 190350
rect 378054 190294 378122 190350
rect 378178 190294 378246 190350
rect 378302 190294 399878 190350
rect 399934 190294 400002 190350
rect 400058 190294 408594 190350
rect 408650 190294 408718 190350
rect 408774 190294 408842 190350
rect 408898 190294 408966 190350
rect 409022 190294 430598 190350
rect 430654 190294 430722 190350
rect 430778 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 470034 190350
rect 470090 190294 470158 190350
rect 470214 190294 470282 190350
rect 470338 190294 470406 190350
rect 470462 190294 500754 190350
rect 500810 190294 500878 190350
rect 500934 190294 501002 190350
rect 501058 190294 501126 190350
rect 501182 190294 531474 190350
rect 531530 190294 531598 190350
rect 531654 190294 531722 190350
rect 531778 190294 531846 190350
rect 531902 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 12960 190226
rect 13016 190170 13084 190226
rect 13140 190170 13208 190226
rect 13264 190170 13332 190226
rect 13388 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 70674 190226
rect 70730 190170 70798 190226
rect 70854 190170 70922 190226
rect 70978 190170 71046 190226
rect 71102 190170 97642 190226
rect 97698 190170 97766 190226
rect 97822 190170 97890 190226
rect 97946 190170 98014 190226
rect 98070 190170 101394 190226
rect 101450 190170 101518 190226
rect 101574 190170 101642 190226
rect 101698 190170 101766 190226
rect 101822 190170 112960 190226
rect 113016 190170 113084 190226
rect 113140 190170 113208 190226
rect 113264 190170 113332 190226
rect 113388 190170 132114 190226
rect 132170 190170 132238 190226
rect 132294 190170 132362 190226
rect 132418 190170 132486 190226
rect 132542 190170 162834 190226
rect 162890 190170 162958 190226
rect 163014 190170 163082 190226
rect 163138 190170 163206 190226
rect 163262 190170 193554 190226
rect 193610 190170 193678 190226
rect 193734 190170 193802 190226
rect 193858 190170 193926 190226
rect 193982 190170 197642 190226
rect 197698 190170 197766 190226
rect 197822 190170 197890 190226
rect 197946 190170 198014 190226
rect 198070 190170 229878 190226
rect 229934 190170 230002 190226
rect 230058 190170 260598 190226
rect 260654 190170 260722 190226
rect 260778 190170 291318 190226
rect 291374 190170 291442 190226
rect 291498 190170 322038 190226
rect 322094 190170 322162 190226
rect 322218 190170 352758 190226
rect 352814 190170 352882 190226
rect 352938 190170 377874 190226
rect 377930 190170 377998 190226
rect 378054 190170 378122 190226
rect 378178 190170 378246 190226
rect 378302 190170 399878 190226
rect 399934 190170 400002 190226
rect 400058 190170 408594 190226
rect 408650 190170 408718 190226
rect 408774 190170 408842 190226
rect 408898 190170 408966 190226
rect 409022 190170 430598 190226
rect 430654 190170 430722 190226
rect 430778 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 470034 190226
rect 470090 190170 470158 190226
rect 470214 190170 470282 190226
rect 470338 190170 470406 190226
rect 470462 190170 500754 190226
rect 500810 190170 500878 190226
rect 500934 190170 501002 190226
rect 501058 190170 501126 190226
rect 501182 190170 531474 190226
rect 531530 190170 531598 190226
rect 531654 190170 531722 190226
rect 531778 190170 531846 190226
rect 531902 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 12960 190102
rect 13016 190046 13084 190102
rect 13140 190046 13208 190102
rect 13264 190046 13332 190102
rect 13388 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 70674 190102
rect 70730 190046 70798 190102
rect 70854 190046 70922 190102
rect 70978 190046 71046 190102
rect 71102 190046 97642 190102
rect 97698 190046 97766 190102
rect 97822 190046 97890 190102
rect 97946 190046 98014 190102
rect 98070 190046 101394 190102
rect 101450 190046 101518 190102
rect 101574 190046 101642 190102
rect 101698 190046 101766 190102
rect 101822 190046 112960 190102
rect 113016 190046 113084 190102
rect 113140 190046 113208 190102
rect 113264 190046 113332 190102
rect 113388 190046 132114 190102
rect 132170 190046 132238 190102
rect 132294 190046 132362 190102
rect 132418 190046 132486 190102
rect 132542 190046 162834 190102
rect 162890 190046 162958 190102
rect 163014 190046 163082 190102
rect 163138 190046 163206 190102
rect 163262 190046 193554 190102
rect 193610 190046 193678 190102
rect 193734 190046 193802 190102
rect 193858 190046 193926 190102
rect 193982 190046 197642 190102
rect 197698 190046 197766 190102
rect 197822 190046 197890 190102
rect 197946 190046 198014 190102
rect 198070 190046 229878 190102
rect 229934 190046 230002 190102
rect 230058 190046 260598 190102
rect 260654 190046 260722 190102
rect 260778 190046 291318 190102
rect 291374 190046 291442 190102
rect 291498 190046 322038 190102
rect 322094 190046 322162 190102
rect 322218 190046 352758 190102
rect 352814 190046 352882 190102
rect 352938 190046 377874 190102
rect 377930 190046 377998 190102
rect 378054 190046 378122 190102
rect 378178 190046 378246 190102
rect 378302 190046 399878 190102
rect 399934 190046 400002 190102
rect 400058 190046 408594 190102
rect 408650 190046 408718 190102
rect 408774 190046 408842 190102
rect 408898 190046 408966 190102
rect 409022 190046 430598 190102
rect 430654 190046 430722 190102
rect 430778 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 470034 190102
rect 470090 190046 470158 190102
rect 470214 190046 470282 190102
rect 470338 190046 470406 190102
rect 470462 190046 500754 190102
rect 500810 190046 500878 190102
rect 500934 190046 501002 190102
rect 501058 190046 501126 190102
rect 501182 190046 531474 190102
rect 531530 190046 531598 190102
rect 531654 190046 531722 190102
rect 531778 190046 531846 190102
rect 531902 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 12960 189978
rect 13016 189922 13084 189978
rect 13140 189922 13208 189978
rect 13264 189922 13332 189978
rect 13388 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 70674 189978
rect 70730 189922 70798 189978
rect 70854 189922 70922 189978
rect 70978 189922 71046 189978
rect 71102 189922 97642 189978
rect 97698 189922 97766 189978
rect 97822 189922 97890 189978
rect 97946 189922 98014 189978
rect 98070 189922 101394 189978
rect 101450 189922 101518 189978
rect 101574 189922 101642 189978
rect 101698 189922 101766 189978
rect 101822 189922 112960 189978
rect 113016 189922 113084 189978
rect 113140 189922 113208 189978
rect 113264 189922 113332 189978
rect 113388 189922 132114 189978
rect 132170 189922 132238 189978
rect 132294 189922 132362 189978
rect 132418 189922 132486 189978
rect 132542 189922 162834 189978
rect 162890 189922 162958 189978
rect 163014 189922 163082 189978
rect 163138 189922 163206 189978
rect 163262 189922 193554 189978
rect 193610 189922 193678 189978
rect 193734 189922 193802 189978
rect 193858 189922 193926 189978
rect 193982 189922 197642 189978
rect 197698 189922 197766 189978
rect 197822 189922 197890 189978
rect 197946 189922 198014 189978
rect 198070 189922 229878 189978
rect 229934 189922 230002 189978
rect 230058 189922 260598 189978
rect 260654 189922 260722 189978
rect 260778 189922 291318 189978
rect 291374 189922 291442 189978
rect 291498 189922 322038 189978
rect 322094 189922 322162 189978
rect 322218 189922 352758 189978
rect 352814 189922 352882 189978
rect 352938 189922 377874 189978
rect 377930 189922 377998 189978
rect 378054 189922 378122 189978
rect 378178 189922 378246 189978
rect 378302 189922 399878 189978
rect 399934 189922 400002 189978
rect 400058 189922 408594 189978
rect 408650 189922 408718 189978
rect 408774 189922 408842 189978
rect 408898 189922 408966 189978
rect 409022 189922 430598 189978
rect 430654 189922 430722 189978
rect 430778 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 470034 189978
rect 470090 189922 470158 189978
rect 470214 189922 470282 189978
rect 470338 189922 470406 189978
rect 470462 189922 500754 189978
rect 500810 189922 500878 189978
rect 500934 189922 501002 189978
rect 501058 189922 501126 189978
rect 501182 189922 531474 189978
rect 531530 189922 531598 189978
rect 531654 189922 531722 189978
rect 531778 189922 531846 189978
rect 531902 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect 375212 188038 431076 188054
rect 375212 187982 375228 188038
rect 375284 187982 431004 188038
rect 431060 187982 431076 188038
rect 375212 187966 431076 187982
rect 373420 187858 384148 187874
rect 373420 187802 373436 187858
rect 373492 187802 384076 187858
rect 384132 187802 384148 187858
rect 373420 187786 384148 187802
rect 26780 187318 203492 187334
rect 26780 187262 26796 187318
rect 26852 187262 203420 187318
rect 203476 187262 203492 187318
rect 26780 187246 203492 187262
rect 21740 185698 205060 185714
rect 21740 185642 21756 185698
rect 21812 185642 204988 185698
rect 205044 185642 205060 185698
rect 21740 185626 205060 185642
rect 373868 184978 443732 184994
rect 373868 184922 373884 184978
rect 373940 184922 443660 184978
rect 443716 184922 443732 184978
rect 373868 184906 443732 184922
rect -1916 184386 597980 184446
rect -1916 184350 404874 184386
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 13760 184350
rect 13816 184294 13884 184350
rect 13940 184294 14008 184350
rect 14064 184294 14132 184350
rect 14188 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 66954 184350
rect 67010 184294 67078 184350
rect 67134 184294 67202 184350
rect 67258 184294 67326 184350
rect 67382 184294 98442 184350
rect 98498 184294 98566 184350
rect 98622 184294 98690 184350
rect 98746 184294 98814 184350
rect 98870 184294 113760 184350
rect 113816 184294 113884 184350
rect 113940 184294 114008 184350
rect 114064 184294 114132 184350
rect 114188 184294 128394 184350
rect 128450 184294 128518 184350
rect 128574 184294 128642 184350
rect 128698 184294 128766 184350
rect 128822 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 189834 184350
rect 189890 184294 189958 184350
rect 190014 184294 190082 184350
rect 190138 184294 190206 184350
rect 190262 184294 198442 184350
rect 198498 184294 198566 184350
rect 198622 184294 198690 184350
rect 198746 184294 198814 184350
rect 198870 184294 214518 184350
rect 214574 184294 214642 184350
rect 214698 184294 245238 184350
rect 245294 184294 245362 184350
rect 245418 184294 275958 184350
rect 276014 184294 276082 184350
rect 276138 184294 306678 184350
rect 306734 184294 306802 184350
rect 306858 184294 337398 184350
rect 337454 184294 337522 184350
rect 337578 184294 368118 184350
rect 368174 184294 368242 184350
rect 368298 184294 374154 184350
rect 374210 184294 374278 184350
rect 374334 184294 374402 184350
rect 374458 184294 374526 184350
rect 374582 184294 384518 184350
rect 384574 184294 384642 184350
rect 384698 184330 404874 184350
rect 404930 184330 404998 184386
rect 405054 184330 405122 184386
rect 405178 184330 405246 184386
rect 405302 184350 597980 184386
rect 405302 184330 415238 184350
rect 384698 184294 415238 184330
rect 415294 184294 415362 184350
rect 415418 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 466314 184350
rect 466370 184294 466438 184350
rect 466494 184294 466562 184350
rect 466618 184294 466686 184350
rect 466742 184294 497034 184350
rect 497090 184294 497158 184350
rect 497214 184294 497282 184350
rect 497338 184294 497406 184350
rect 497462 184294 527754 184350
rect 527810 184294 527878 184350
rect 527934 184294 528002 184350
rect 528058 184294 528126 184350
rect 528182 184294 558474 184350
rect 558530 184294 558598 184350
rect 558654 184294 558722 184350
rect 558778 184294 558846 184350
rect 558902 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184262 597980 184294
rect -1916 184226 404874 184262
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 13760 184226
rect 13816 184170 13884 184226
rect 13940 184170 14008 184226
rect 14064 184170 14132 184226
rect 14188 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 66954 184226
rect 67010 184170 67078 184226
rect 67134 184170 67202 184226
rect 67258 184170 67326 184226
rect 67382 184170 98442 184226
rect 98498 184170 98566 184226
rect 98622 184170 98690 184226
rect 98746 184170 98814 184226
rect 98870 184170 113760 184226
rect 113816 184170 113884 184226
rect 113940 184170 114008 184226
rect 114064 184170 114132 184226
rect 114188 184170 128394 184226
rect 128450 184170 128518 184226
rect 128574 184170 128642 184226
rect 128698 184170 128766 184226
rect 128822 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 189834 184226
rect 189890 184170 189958 184226
rect 190014 184170 190082 184226
rect 190138 184170 190206 184226
rect 190262 184170 198442 184226
rect 198498 184170 198566 184226
rect 198622 184170 198690 184226
rect 198746 184170 198814 184226
rect 198870 184170 214518 184226
rect 214574 184170 214642 184226
rect 214698 184170 245238 184226
rect 245294 184170 245362 184226
rect 245418 184170 275958 184226
rect 276014 184170 276082 184226
rect 276138 184170 306678 184226
rect 306734 184170 306802 184226
rect 306858 184170 337398 184226
rect 337454 184170 337522 184226
rect 337578 184170 368118 184226
rect 368174 184170 368242 184226
rect 368298 184170 374154 184226
rect 374210 184170 374278 184226
rect 374334 184170 374402 184226
rect 374458 184170 374526 184226
rect 374582 184170 384518 184226
rect 384574 184170 384642 184226
rect 384698 184206 404874 184226
rect 404930 184206 404998 184262
rect 405054 184206 405122 184262
rect 405178 184206 405246 184262
rect 405302 184226 597980 184262
rect 405302 184206 415238 184226
rect 384698 184170 415238 184206
rect 415294 184170 415362 184226
rect 415418 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 466314 184226
rect 466370 184170 466438 184226
rect 466494 184170 466562 184226
rect 466618 184170 466686 184226
rect 466742 184170 497034 184226
rect 497090 184170 497158 184226
rect 497214 184170 497282 184226
rect 497338 184170 497406 184226
rect 497462 184170 527754 184226
rect 527810 184170 527878 184226
rect 527934 184170 528002 184226
rect 528058 184170 528126 184226
rect 528182 184170 558474 184226
rect 558530 184170 558598 184226
rect 558654 184170 558722 184226
rect 558778 184170 558846 184226
rect 558902 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184138 597980 184170
rect -1916 184102 404874 184138
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 13760 184102
rect 13816 184046 13884 184102
rect 13940 184046 14008 184102
rect 14064 184046 14132 184102
rect 14188 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 66954 184102
rect 67010 184046 67078 184102
rect 67134 184046 67202 184102
rect 67258 184046 67326 184102
rect 67382 184046 98442 184102
rect 98498 184046 98566 184102
rect 98622 184046 98690 184102
rect 98746 184046 98814 184102
rect 98870 184046 113760 184102
rect 113816 184046 113884 184102
rect 113940 184046 114008 184102
rect 114064 184046 114132 184102
rect 114188 184046 128394 184102
rect 128450 184046 128518 184102
rect 128574 184046 128642 184102
rect 128698 184046 128766 184102
rect 128822 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 189834 184102
rect 189890 184046 189958 184102
rect 190014 184046 190082 184102
rect 190138 184046 190206 184102
rect 190262 184046 198442 184102
rect 198498 184046 198566 184102
rect 198622 184046 198690 184102
rect 198746 184046 198814 184102
rect 198870 184046 214518 184102
rect 214574 184046 214642 184102
rect 214698 184046 245238 184102
rect 245294 184046 245362 184102
rect 245418 184046 275958 184102
rect 276014 184046 276082 184102
rect 276138 184046 306678 184102
rect 306734 184046 306802 184102
rect 306858 184046 337398 184102
rect 337454 184046 337522 184102
rect 337578 184046 368118 184102
rect 368174 184046 368242 184102
rect 368298 184046 374154 184102
rect 374210 184046 374278 184102
rect 374334 184046 374402 184102
rect 374458 184046 374526 184102
rect 374582 184046 384518 184102
rect 384574 184046 384642 184102
rect 384698 184082 404874 184102
rect 404930 184082 404998 184138
rect 405054 184082 405122 184138
rect 405178 184082 405246 184138
rect 405302 184102 597980 184138
rect 405302 184082 415238 184102
rect 384698 184046 415238 184082
rect 415294 184046 415362 184102
rect 415418 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 466314 184102
rect 466370 184046 466438 184102
rect 466494 184046 466562 184102
rect 466618 184046 466686 184102
rect 466742 184046 497034 184102
rect 497090 184046 497158 184102
rect 497214 184046 497282 184102
rect 497338 184046 497406 184102
rect 497462 184046 527754 184102
rect 527810 184046 527878 184102
rect 527934 184046 528002 184102
rect 528058 184046 528126 184102
rect 528182 184046 558474 184102
rect 558530 184046 558598 184102
rect 558654 184046 558722 184102
rect 558778 184046 558846 184102
rect 558902 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 13760 183978
rect 13816 183922 13884 183978
rect 13940 183922 14008 183978
rect 14064 183922 14132 183978
rect 14188 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 66954 183978
rect 67010 183922 67078 183978
rect 67134 183922 67202 183978
rect 67258 183922 67326 183978
rect 67382 183922 98442 183978
rect 98498 183922 98566 183978
rect 98622 183922 98690 183978
rect 98746 183922 98814 183978
rect 98870 183922 113760 183978
rect 113816 183922 113884 183978
rect 113940 183922 114008 183978
rect 114064 183922 114132 183978
rect 114188 183922 128394 183978
rect 128450 183922 128518 183978
rect 128574 183922 128642 183978
rect 128698 183922 128766 183978
rect 128822 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 189834 183978
rect 189890 183922 189958 183978
rect 190014 183922 190082 183978
rect 190138 183922 190206 183978
rect 190262 183922 198442 183978
rect 198498 183922 198566 183978
rect 198622 183922 198690 183978
rect 198746 183922 198814 183978
rect 198870 183922 214518 183978
rect 214574 183922 214642 183978
rect 214698 183922 245238 183978
rect 245294 183922 245362 183978
rect 245418 183922 275958 183978
rect 276014 183922 276082 183978
rect 276138 183922 306678 183978
rect 306734 183922 306802 183978
rect 306858 183922 337398 183978
rect 337454 183922 337522 183978
rect 337578 183922 368118 183978
rect 368174 183922 368242 183978
rect 368298 183922 374154 183978
rect 374210 183922 374278 183978
rect 374334 183922 374402 183978
rect 374458 183922 374526 183978
rect 374582 183922 384518 183978
rect 384574 183922 384642 183978
rect 384698 183922 415238 183978
rect 415294 183922 415362 183978
rect 415418 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 466314 183978
rect 466370 183922 466438 183978
rect 466494 183922 466562 183978
rect 466618 183922 466686 183978
rect 466742 183922 497034 183978
rect 497090 183922 497158 183978
rect 497214 183922 497282 183978
rect 497338 183922 497406 183978
rect 497462 183922 527754 183978
rect 527810 183922 527878 183978
rect 527934 183922 528002 183978
rect 528058 183922 528126 183978
rect 528182 183922 558474 183978
rect 558530 183922 558598 183978
rect 558654 183922 558722 183978
rect 558778 183922 558846 183978
rect 558902 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect 379356 182278 395684 182294
rect 379356 182222 379372 182278
rect 379428 182222 395612 182278
rect 395668 182222 395684 182278
rect 379356 182206 395684 182222
rect 104956 181558 203492 181574
rect 104956 181502 104972 181558
rect 105028 181502 118636 181558
rect 118692 181502 203420 181558
rect 203476 181502 203492 181558
rect 104956 181486 203492 181502
rect 100028 178858 126044 178874
rect 100028 178802 100044 178858
rect 100100 178802 126044 178858
rect 100028 178786 126044 178802
rect 125956 178154 126044 178786
rect 125956 178138 205060 178154
rect 125956 178082 126812 178138
rect 126868 178082 204988 178138
rect 205044 178082 205060 178138
rect 125956 178066 205060 178082
rect 103500 177238 126044 177254
rect 103500 177182 103516 177238
rect 103572 177182 126044 177238
rect 103500 177166 126044 177182
rect 125956 176534 126044 177166
rect 125956 176518 206740 176534
rect 125956 176462 129052 176518
rect 129108 176462 206668 176518
rect 206724 176462 206740 176518
rect 125956 176446 206740 176462
rect 99916 173818 126044 173834
rect 99916 173762 99932 173818
rect 99988 173762 126044 173818
rect 99916 173746 126044 173762
rect 125956 173114 126044 173746
rect 125956 173098 206964 173114
rect 125956 173042 138572 173098
rect 138628 173042 206892 173098
rect 206948 173042 206964 173098
rect 125956 173026 206964 173042
rect 187276 172738 205060 172754
rect 187276 172682 187292 172738
rect 187348 172682 204988 172738
rect 205044 172682 205060 172738
rect 187276 172666 205060 172682
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 12960 172350
rect 13016 172294 13084 172350
rect 13140 172294 13208 172350
rect 13264 172294 13332 172350
rect 13388 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 70674 172350
rect 70730 172294 70798 172350
rect 70854 172294 70922 172350
rect 70978 172294 71046 172350
rect 71102 172294 97642 172350
rect 97698 172294 97766 172350
rect 97822 172294 97890 172350
rect 97946 172294 98014 172350
rect 98070 172294 101394 172350
rect 101450 172294 101518 172350
rect 101574 172294 101642 172350
rect 101698 172294 101766 172350
rect 101822 172294 112960 172350
rect 113016 172294 113084 172350
rect 113140 172294 113208 172350
rect 113264 172294 113332 172350
rect 113388 172294 132114 172350
rect 132170 172294 132238 172350
rect 132294 172294 132362 172350
rect 132418 172294 132486 172350
rect 132542 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 193554 172350
rect 193610 172294 193678 172350
rect 193734 172294 193802 172350
rect 193858 172294 193926 172350
rect 193982 172294 197642 172350
rect 197698 172294 197766 172350
rect 197822 172294 197890 172350
rect 197946 172294 198014 172350
rect 198070 172294 229878 172350
rect 229934 172294 230002 172350
rect 230058 172294 260598 172350
rect 260654 172294 260722 172350
rect 260778 172294 291318 172350
rect 291374 172294 291442 172350
rect 291498 172294 322038 172350
rect 322094 172294 322162 172350
rect 322218 172294 352758 172350
rect 352814 172294 352882 172350
rect 352938 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 399878 172350
rect 399934 172294 400002 172350
rect 400058 172294 430598 172350
rect 430654 172294 430722 172350
rect 430778 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 12960 172226
rect 13016 172170 13084 172226
rect 13140 172170 13208 172226
rect 13264 172170 13332 172226
rect 13388 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 70674 172226
rect 70730 172170 70798 172226
rect 70854 172170 70922 172226
rect 70978 172170 71046 172226
rect 71102 172170 97642 172226
rect 97698 172170 97766 172226
rect 97822 172170 97890 172226
rect 97946 172170 98014 172226
rect 98070 172170 101394 172226
rect 101450 172170 101518 172226
rect 101574 172170 101642 172226
rect 101698 172170 101766 172226
rect 101822 172170 112960 172226
rect 113016 172170 113084 172226
rect 113140 172170 113208 172226
rect 113264 172170 113332 172226
rect 113388 172170 132114 172226
rect 132170 172170 132238 172226
rect 132294 172170 132362 172226
rect 132418 172170 132486 172226
rect 132542 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 193554 172226
rect 193610 172170 193678 172226
rect 193734 172170 193802 172226
rect 193858 172170 193926 172226
rect 193982 172170 197642 172226
rect 197698 172170 197766 172226
rect 197822 172170 197890 172226
rect 197946 172170 198014 172226
rect 198070 172170 229878 172226
rect 229934 172170 230002 172226
rect 230058 172170 260598 172226
rect 260654 172170 260722 172226
rect 260778 172170 291318 172226
rect 291374 172170 291442 172226
rect 291498 172170 322038 172226
rect 322094 172170 322162 172226
rect 322218 172170 352758 172226
rect 352814 172170 352882 172226
rect 352938 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 399878 172226
rect 399934 172170 400002 172226
rect 400058 172170 430598 172226
rect 430654 172170 430722 172226
rect 430778 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 12960 172102
rect 13016 172046 13084 172102
rect 13140 172046 13208 172102
rect 13264 172046 13332 172102
rect 13388 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 70674 172102
rect 70730 172046 70798 172102
rect 70854 172046 70922 172102
rect 70978 172046 71046 172102
rect 71102 172046 97642 172102
rect 97698 172046 97766 172102
rect 97822 172046 97890 172102
rect 97946 172046 98014 172102
rect 98070 172046 101394 172102
rect 101450 172046 101518 172102
rect 101574 172046 101642 172102
rect 101698 172046 101766 172102
rect 101822 172046 112960 172102
rect 113016 172046 113084 172102
rect 113140 172046 113208 172102
rect 113264 172046 113332 172102
rect 113388 172046 132114 172102
rect 132170 172046 132238 172102
rect 132294 172046 132362 172102
rect 132418 172046 132486 172102
rect 132542 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 193554 172102
rect 193610 172046 193678 172102
rect 193734 172046 193802 172102
rect 193858 172046 193926 172102
rect 193982 172046 197642 172102
rect 197698 172046 197766 172102
rect 197822 172046 197890 172102
rect 197946 172046 198014 172102
rect 198070 172046 229878 172102
rect 229934 172046 230002 172102
rect 230058 172046 260598 172102
rect 260654 172046 260722 172102
rect 260778 172046 291318 172102
rect 291374 172046 291442 172102
rect 291498 172046 322038 172102
rect 322094 172046 322162 172102
rect 322218 172046 352758 172102
rect 352814 172046 352882 172102
rect 352938 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 399878 172102
rect 399934 172046 400002 172102
rect 400058 172046 430598 172102
rect 430654 172046 430722 172102
rect 430778 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 12960 171978
rect 13016 171922 13084 171978
rect 13140 171922 13208 171978
rect 13264 171922 13332 171978
rect 13388 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 70674 171978
rect 70730 171922 70798 171978
rect 70854 171922 70922 171978
rect 70978 171922 71046 171978
rect 71102 171922 97642 171978
rect 97698 171922 97766 171978
rect 97822 171922 97890 171978
rect 97946 171922 98014 171978
rect 98070 171922 101394 171978
rect 101450 171922 101518 171978
rect 101574 171922 101642 171978
rect 101698 171922 101766 171978
rect 101822 171922 112960 171978
rect 113016 171922 113084 171978
rect 113140 171922 113208 171978
rect 113264 171922 113332 171978
rect 113388 171922 132114 171978
rect 132170 171922 132238 171978
rect 132294 171922 132362 171978
rect 132418 171922 132486 171978
rect 132542 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 193554 171978
rect 193610 171922 193678 171978
rect 193734 171922 193802 171978
rect 193858 171922 193926 171978
rect 193982 171922 197642 171978
rect 197698 171922 197766 171978
rect 197822 171922 197890 171978
rect 197946 171922 198014 171978
rect 198070 171922 229878 171978
rect 229934 171922 230002 171978
rect 230058 171922 260598 171978
rect 260654 171922 260722 171978
rect 260778 171922 291318 171978
rect 291374 171922 291442 171978
rect 291498 171922 322038 171978
rect 322094 171922 322162 171978
rect 322218 171922 352758 171978
rect 352814 171922 352882 171978
rect 352938 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 399878 171978
rect 399934 171922 400002 171978
rect 400058 171922 430598 171978
rect 430654 171922 430722 171978
rect 430778 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect 189068 168778 201588 168794
rect 189068 168722 189084 168778
rect 189140 168722 201516 168778
rect 201572 168722 201588 168778
rect 189068 168706 201588 168722
rect 380364 166618 381796 166634
rect 380364 166562 380380 166618
rect 380436 166562 381724 166618
rect 381780 166562 381796 166618
rect 380364 166546 381796 166562
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 66954 166350
rect 67010 166294 67078 166350
rect 67134 166294 67202 166350
rect 67258 166294 67326 166350
rect 67382 166294 97674 166350
rect 97730 166294 97798 166350
rect 97854 166294 97922 166350
rect 97978 166294 98046 166350
rect 98102 166294 128394 166350
rect 128450 166294 128518 166350
rect 128574 166294 128642 166350
rect 128698 166294 128766 166350
rect 128822 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 189834 166350
rect 189890 166294 189958 166350
rect 190014 166294 190082 166350
rect 190138 166294 190206 166350
rect 190262 166294 214518 166350
rect 214574 166294 214642 166350
rect 214698 166294 245238 166350
rect 245294 166294 245362 166350
rect 245418 166294 275958 166350
rect 276014 166294 276082 166350
rect 276138 166294 306678 166350
rect 306734 166294 306802 166350
rect 306858 166294 337398 166350
rect 337454 166294 337522 166350
rect 337578 166294 368118 166350
rect 368174 166294 368242 166350
rect 368298 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 384518 166350
rect 384574 166294 384642 166350
rect 384698 166294 415238 166350
rect 415294 166294 415362 166350
rect 415418 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 466314 166350
rect 466370 166294 466438 166350
rect 466494 166294 466562 166350
rect 466618 166294 466686 166350
rect 466742 166294 497034 166350
rect 497090 166294 497158 166350
rect 497214 166294 497282 166350
rect 497338 166294 497406 166350
rect 497462 166294 527754 166350
rect 527810 166294 527878 166350
rect 527934 166294 528002 166350
rect 528058 166294 528126 166350
rect 528182 166294 558474 166350
rect 558530 166294 558598 166350
rect 558654 166294 558722 166350
rect 558778 166294 558846 166350
rect 558902 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 66954 166226
rect 67010 166170 67078 166226
rect 67134 166170 67202 166226
rect 67258 166170 67326 166226
rect 67382 166170 97674 166226
rect 97730 166170 97798 166226
rect 97854 166170 97922 166226
rect 97978 166170 98046 166226
rect 98102 166170 128394 166226
rect 128450 166170 128518 166226
rect 128574 166170 128642 166226
rect 128698 166170 128766 166226
rect 128822 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 189834 166226
rect 189890 166170 189958 166226
rect 190014 166170 190082 166226
rect 190138 166170 190206 166226
rect 190262 166170 214518 166226
rect 214574 166170 214642 166226
rect 214698 166170 245238 166226
rect 245294 166170 245362 166226
rect 245418 166170 275958 166226
rect 276014 166170 276082 166226
rect 276138 166170 306678 166226
rect 306734 166170 306802 166226
rect 306858 166170 337398 166226
rect 337454 166170 337522 166226
rect 337578 166170 368118 166226
rect 368174 166170 368242 166226
rect 368298 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 384518 166226
rect 384574 166170 384642 166226
rect 384698 166170 415238 166226
rect 415294 166170 415362 166226
rect 415418 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 466314 166226
rect 466370 166170 466438 166226
rect 466494 166170 466562 166226
rect 466618 166170 466686 166226
rect 466742 166170 497034 166226
rect 497090 166170 497158 166226
rect 497214 166170 497282 166226
rect 497338 166170 497406 166226
rect 497462 166170 527754 166226
rect 527810 166170 527878 166226
rect 527934 166170 528002 166226
rect 528058 166170 528126 166226
rect 528182 166170 558474 166226
rect 558530 166170 558598 166226
rect 558654 166170 558722 166226
rect 558778 166170 558846 166226
rect 558902 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 66954 166102
rect 67010 166046 67078 166102
rect 67134 166046 67202 166102
rect 67258 166046 67326 166102
rect 67382 166046 97674 166102
rect 97730 166046 97798 166102
rect 97854 166046 97922 166102
rect 97978 166046 98046 166102
rect 98102 166046 128394 166102
rect 128450 166046 128518 166102
rect 128574 166046 128642 166102
rect 128698 166046 128766 166102
rect 128822 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 189834 166102
rect 189890 166046 189958 166102
rect 190014 166046 190082 166102
rect 190138 166046 190206 166102
rect 190262 166046 214518 166102
rect 214574 166046 214642 166102
rect 214698 166046 245238 166102
rect 245294 166046 245362 166102
rect 245418 166046 275958 166102
rect 276014 166046 276082 166102
rect 276138 166046 306678 166102
rect 306734 166046 306802 166102
rect 306858 166046 337398 166102
rect 337454 166046 337522 166102
rect 337578 166046 368118 166102
rect 368174 166046 368242 166102
rect 368298 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 384518 166102
rect 384574 166046 384642 166102
rect 384698 166046 415238 166102
rect 415294 166046 415362 166102
rect 415418 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 466314 166102
rect 466370 166046 466438 166102
rect 466494 166046 466562 166102
rect 466618 166046 466686 166102
rect 466742 166046 497034 166102
rect 497090 166046 497158 166102
rect 497214 166046 497282 166102
rect 497338 166046 497406 166102
rect 497462 166046 527754 166102
rect 527810 166046 527878 166102
rect 527934 166046 528002 166102
rect 528058 166046 528126 166102
rect 528182 166046 558474 166102
rect 558530 166046 558598 166102
rect 558654 166046 558722 166102
rect 558778 166046 558846 166102
rect 558902 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 66954 165978
rect 67010 165922 67078 165978
rect 67134 165922 67202 165978
rect 67258 165922 67326 165978
rect 67382 165922 97674 165978
rect 97730 165922 97798 165978
rect 97854 165922 97922 165978
rect 97978 165922 98046 165978
rect 98102 165922 128394 165978
rect 128450 165922 128518 165978
rect 128574 165922 128642 165978
rect 128698 165922 128766 165978
rect 128822 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 189834 165978
rect 189890 165922 189958 165978
rect 190014 165922 190082 165978
rect 190138 165922 190206 165978
rect 190262 165922 214518 165978
rect 214574 165922 214642 165978
rect 214698 165922 245238 165978
rect 245294 165922 245362 165978
rect 245418 165922 275958 165978
rect 276014 165922 276082 165978
rect 276138 165922 306678 165978
rect 306734 165922 306802 165978
rect 306858 165922 337398 165978
rect 337454 165922 337522 165978
rect 337578 165922 368118 165978
rect 368174 165922 368242 165978
rect 368298 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 384518 165978
rect 384574 165922 384642 165978
rect 384698 165922 415238 165978
rect 415294 165922 415362 165978
rect 415418 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 466314 165978
rect 466370 165922 466438 165978
rect 466494 165922 466562 165978
rect 466618 165922 466686 165978
rect 466742 165922 497034 165978
rect 497090 165922 497158 165978
rect 497214 165922 497282 165978
rect 497338 165922 497406 165978
rect 497462 165922 527754 165978
rect 527810 165922 527878 165978
rect 527934 165922 528002 165978
rect 528058 165922 528126 165978
rect 528182 165922 558474 165978
rect 558530 165922 558598 165978
rect 558654 165922 558722 165978
rect 558778 165922 558846 165978
rect 558902 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect 20844 162838 111988 162854
rect 20844 162782 20860 162838
rect 20916 162782 111916 162838
rect 111972 162782 111988 162838
rect 20844 162766 111988 162782
rect 126236 162838 206852 162854
rect 126236 162782 126252 162838
rect 126308 162782 206780 162838
rect 206836 162782 206852 162838
rect 126236 162766 206852 162782
rect 27116 162658 103476 162674
rect 27116 162602 27132 162658
rect 27188 162602 103404 162658
rect 103460 162602 103476 162658
rect 27116 162586 103476 162602
rect 377340 156358 381684 156374
rect 377340 156302 377356 156358
rect 377412 156302 381612 156358
rect 381668 156302 381684 156358
rect 377340 156286 381684 156302
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 70674 154350
rect 70730 154294 70798 154350
rect 70854 154294 70922 154350
rect 70978 154294 71046 154350
rect 71102 154294 101394 154350
rect 101450 154294 101518 154350
rect 101574 154294 101642 154350
rect 101698 154294 101766 154350
rect 101822 154294 132114 154350
rect 132170 154294 132238 154350
rect 132294 154294 132362 154350
rect 132418 154294 132486 154350
rect 132542 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 193554 154350
rect 193610 154294 193678 154350
rect 193734 154294 193802 154350
rect 193858 154294 193926 154350
rect 193982 154294 229878 154350
rect 229934 154294 230002 154350
rect 230058 154294 260598 154350
rect 260654 154294 260722 154350
rect 260778 154294 291318 154350
rect 291374 154294 291442 154350
rect 291498 154294 322038 154350
rect 322094 154294 322162 154350
rect 322218 154294 352758 154350
rect 352814 154294 352882 154350
rect 352938 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 399878 154350
rect 399934 154294 400002 154350
rect 400058 154294 430598 154350
rect 430654 154294 430722 154350
rect 430778 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 70674 154226
rect 70730 154170 70798 154226
rect 70854 154170 70922 154226
rect 70978 154170 71046 154226
rect 71102 154170 101394 154226
rect 101450 154170 101518 154226
rect 101574 154170 101642 154226
rect 101698 154170 101766 154226
rect 101822 154170 132114 154226
rect 132170 154170 132238 154226
rect 132294 154170 132362 154226
rect 132418 154170 132486 154226
rect 132542 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 193554 154226
rect 193610 154170 193678 154226
rect 193734 154170 193802 154226
rect 193858 154170 193926 154226
rect 193982 154170 229878 154226
rect 229934 154170 230002 154226
rect 230058 154170 260598 154226
rect 260654 154170 260722 154226
rect 260778 154170 291318 154226
rect 291374 154170 291442 154226
rect 291498 154170 322038 154226
rect 322094 154170 322162 154226
rect 322218 154170 352758 154226
rect 352814 154170 352882 154226
rect 352938 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 399878 154226
rect 399934 154170 400002 154226
rect 400058 154170 430598 154226
rect 430654 154170 430722 154226
rect 430778 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 70674 154102
rect 70730 154046 70798 154102
rect 70854 154046 70922 154102
rect 70978 154046 71046 154102
rect 71102 154046 101394 154102
rect 101450 154046 101518 154102
rect 101574 154046 101642 154102
rect 101698 154046 101766 154102
rect 101822 154046 132114 154102
rect 132170 154046 132238 154102
rect 132294 154046 132362 154102
rect 132418 154046 132486 154102
rect 132542 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 193554 154102
rect 193610 154046 193678 154102
rect 193734 154046 193802 154102
rect 193858 154046 193926 154102
rect 193982 154046 229878 154102
rect 229934 154046 230002 154102
rect 230058 154046 260598 154102
rect 260654 154046 260722 154102
rect 260778 154046 291318 154102
rect 291374 154046 291442 154102
rect 291498 154046 322038 154102
rect 322094 154046 322162 154102
rect 322218 154046 352758 154102
rect 352814 154046 352882 154102
rect 352938 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 399878 154102
rect 399934 154046 400002 154102
rect 400058 154046 430598 154102
rect 430654 154046 430722 154102
rect 430778 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 70674 153978
rect 70730 153922 70798 153978
rect 70854 153922 70922 153978
rect 70978 153922 71046 153978
rect 71102 153922 101394 153978
rect 101450 153922 101518 153978
rect 101574 153922 101642 153978
rect 101698 153922 101766 153978
rect 101822 153922 132114 153978
rect 132170 153922 132238 153978
rect 132294 153922 132362 153978
rect 132418 153922 132486 153978
rect 132542 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 193554 153978
rect 193610 153922 193678 153978
rect 193734 153922 193802 153978
rect 193858 153922 193926 153978
rect 193982 153922 229878 153978
rect 229934 153922 230002 153978
rect 230058 153922 260598 153978
rect 260654 153922 260722 153978
rect 260778 153922 291318 153978
rect 291374 153922 291442 153978
rect 291498 153922 322038 153978
rect 322094 153922 322162 153978
rect 322218 153922 352758 153978
rect 352814 153922 352882 153978
rect 352938 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 399878 153978
rect 399934 153922 400002 153978
rect 400058 153922 430598 153978
rect 430654 153922 430722 153978
rect 430778 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect 379580 151138 382580 151154
rect 379580 151082 379596 151138
rect 379652 151082 382508 151138
rect 382564 151082 382580 151138
rect 379580 151066 382580 151082
rect 380588 149878 381572 149894
rect 380588 149822 380604 149878
rect 380660 149822 381500 149878
rect 381556 149822 381572 149878
rect 380588 149806 381572 149822
rect 72028 149518 110196 149534
rect 72028 149462 72044 149518
rect 72100 149462 110124 149518
rect 110180 149462 110196 149518
rect 72028 149446 110196 149462
rect 112460 149518 118820 149534
rect 112460 149462 112476 149518
rect 112532 149462 118748 149518
rect 118804 149462 118820 149518
rect 112460 149446 118820 149462
rect 81436 149338 110420 149354
rect 81436 149282 81452 149338
rect 81508 149282 110348 149338
rect 110404 149282 110420 149338
rect 81436 149266 110420 149282
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 66954 148350
rect 67010 148294 67078 148350
rect 67134 148294 67202 148350
rect 67258 148294 67326 148350
rect 67382 148294 97674 148350
rect 97730 148294 97798 148350
rect 97854 148294 97922 148350
rect 97978 148294 98046 148350
rect 98102 148294 128394 148350
rect 128450 148294 128518 148350
rect 128574 148294 128642 148350
rect 128698 148294 128766 148350
rect 128822 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 189834 148350
rect 189890 148294 189958 148350
rect 190014 148294 190082 148350
rect 190138 148294 190206 148350
rect 190262 148294 214518 148350
rect 214574 148294 214642 148350
rect 214698 148294 245238 148350
rect 245294 148294 245362 148350
rect 245418 148294 275958 148350
rect 276014 148294 276082 148350
rect 276138 148294 306678 148350
rect 306734 148294 306802 148350
rect 306858 148294 337398 148350
rect 337454 148294 337522 148350
rect 337578 148294 368118 148350
rect 368174 148294 368242 148350
rect 368298 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 384518 148350
rect 384574 148294 384642 148350
rect 384698 148294 415238 148350
rect 415294 148294 415362 148350
rect 415418 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 466314 148350
rect 466370 148294 466438 148350
rect 466494 148294 466562 148350
rect 466618 148294 466686 148350
rect 466742 148294 497034 148350
rect 497090 148294 497158 148350
rect 497214 148294 497282 148350
rect 497338 148294 497406 148350
rect 497462 148294 527754 148350
rect 527810 148294 527878 148350
rect 527934 148294 528002 148350
rect 528058 148294 528126 148350
rect 528182 148294 558474 148350
rect 558530 148294 558598 148350
rect 558654 148294 558722 148350
rect 558778 148294 558846 148350
rect 558902 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 66954 148226
rect 67010 148170 67078 148226
rect 67134 148170 67202 148226
rect 67258 148170 67326 148226
rect 67382 148170 97674 148226
rect 97730 148170 97798 148226
rect 97854 148170 97922 148226
rect 97978 148170 98046 148226
rect 98102 148170 128394 148226
rect 128450 148170 128518 148226
rect 128574 148170 128642 148226
rect 128698 148170 128766 148226
rect 128822 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 189834 148226
rect 189890 148170 189958 148226
rect 190014 148170 190082 148226
rect 190138 148170 190206 148226
rect 190262 148170 214518 148226
rect 214574 148170 214642 148226
rect 214698 148170 245238 148226
rect 245294 148170 245362 148226
rect 245418 148170 275958 148226
rect 276014 148170 276082 148226
rect 276138 148170 306678 148226
rect 306734 148170 306802 148226
rect 306858 148170 337398 148226
rect 337454 148170 337522 148226
rect 337578 148170 368118 148226
rect 368174 148170 368242 148226
rect 368298 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 384518 148226
rect 384574 148170 384642 148226
rect 384698 148170 415238 148226
rect 415294 148170 415362 148226
rect 415418 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 466314 148226
rect 466370 148170 466438 148226
rect 466494 148170 466562 148226
rect 466618 148170 466686 148226
rect 466742 148170 497034 148226
rect 497090 148170 497158 148226
rect 497214 148170 497282 148226
rect 497338 148170 497406 148226
rect 497462 148170 527754 148226
rect 527810 148170 527878 148226
rect 527934 148170 528002 148226
rect 528058 148170 528126 148226
rect 528182 148170 558474 148226
rect 558530 148170 558598 148226
rect 558654 148170 558722 148226
rect 558778 148170 558846 148226
rect 558902 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 66954 148102
rect 67010 148046 67078 148102
rect 67134 148046 67202 148102
rect 67258 148046 67326 148102
rect 67382 148046 97674 148102
rect 97730 148046 97798 148102
rect 97854 148046 97922 148102
rect 97978 148046 98046 148102
rect 98102 148046 128394 148102
rect 128450 148046 128518 148102
rect 128574 148046 128642 148102
rect 128698 148046 128766 148102
rect 128822 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 189834 148102
rect 189890 148046 189958 148102
rect 190014 148046 190082 148102
rect 190138 148046 190206 148102
rect 190262 148046 214518 148102
rect 214574 148046 214642 148102
rect 214698 148046 245238 148102
rect 245294 148046 245362 148102
rect 245418 148046 275958 148102
rect 276014 148046 276082 148102
rect 276138 148046 306678 148102
rect 306734 148046 306802 148102
rect 306858 148046 337398 148102
rect 337454 148046 337522 148102
rect 337578 148046 368118 148102
rect 368174 148046 368242 148102
rect 368298 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 384518 148102
rect 384574 148046 384642 148102
rect 384698 148046 415238 148102
rect 415294 148046 415362 148102
rect 415418 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 466314 148102
rect 466370 148046 466438 148102
rect 466494 148046 466562 148102
rect 466618 148046 466686 148102
rect 466742 148046 497034 148102
rect 497090 148046 497158 148102
rect 497214 148046 497282 148102
rect 497338 148046 497406 148102
rect 497462 148046 527754 148102
rect 527810 148046 527878 148102
rect 527934 148046 528002 148102
rect 528058 148046 528126 148102
rect 528182 148046 558474 148102
rect 558530 148046 558598 148102
rect 558654 148046 558722 148102
rect 558778 148046 558846 148102
rect 558902 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 66954 147978
rect 67010 147922 67078 147978
rect 67134 147922 67202 147978
rect 67258 147922 67326 147978
rect 67382 147922 97674 147978
rect 97730 147922 97798 147978
rect 97854 147922 97922 147978
rect 97978 147922 98046 147978
rect 98102 147922 128394 147978
rect 128450 147922 128518 147978
rect 128574 147922 128642 147978
rect 128698 147922 128766 147978
rect 128822 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 189834 147978
rect 189890 147922 189958 147978
rect 190014 147922 190082 147978
rect 190138 147922 190206 147978
rect 190262 147922 214518 147978
rect 214574 147922 214642 147978
rect 214698 147922 245238 147978
rect 245294 147922 245362 147978
rect 245418 147922 275958 147978
rect 276014 147922 276082 147978
rect 276138 147922 306678 147978
rect 306734 147922 306802 147978
rect 306858 147922 337398 147978
rect 337454 147922 337522 147978
rect 337578 147922 368118 147978
rect 368174 147922 368242 147978
rect 368298 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 384518 147978
rect 384574 147922 384642 147978
rect 384698 147922 415238 147978
rect 415294 147922 415362 147978
rect 415418 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 466314 147978
rect 466370 147922 466438 147978
rect 466494 147922 466562 147978
rect 466618 147922 466686 147978
rect 466742 147922 497034 147978
rect 497090 147922 497158 147978
rect 497214 147922 497282 147978
rect 497338 147922 497406 147978
rect 497462 147922 527754 147978
rect 527810 147922 527878 147978
rect 527934 147922 528002 147978
rect 528058 147922 528126 147978
rect 528182 147922 558474 147978
rect 558530 147922 558598 147978
rect 558654 147922 558722 147978
rect 558778 147922 558846 147978
rect 558902 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect 380588 145018 382356 145034
rect 380588 144962 380604 145018
rect 380660 144962 382284 145018
rect 382340 144962 382356 145018
rect 380588 144946 382356 144962
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 11930 136350
rect 11986 136294 12054 136350
rect 12110 136294 12178 136350
rect 12234 136294 12302 136350
rect 12358 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 70674 136350
rect 70730 136294 70798 136350
rect 70854 136294 70922 136350
rect 70978 136294 71046 136350
rect 71102 136294 96612 136350
rect 96668 136294 96736 136350
rect 96792 136294 96860 136350
rect 96916 136294 96984 136350
rect 97040 136294 101394 136350
rect 101450 136294 101518 136350
rect 101574 136294 101642 136350
rect 101698 136294 101766 136350
rect 101822 136294 111930 136350
rect 111986 136294 112054 136350
rect 112110 136294 112178 136350
rect 112234 136294 112302 136350
rect 112358 136294 132114 136350
rect 132170 136294 132238 136350
rect 132294 136294 132362 136350
rect 132418 136294 132486 136350
rect 132542 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 193554 136350
rect 193610 136294 193678 136350
rect 193734 136294 193802 136350
rect 193858 136294 193926 136350
rect 193982 136294 196612 136350
rect 196668 136294 196736 136350
rect 196792 136294 196860 136350
rect 196916 136294 196984 136350
rect 197040 136294 229878 136350
rect 229934 136294 230002 136350
rect 230058 136294 260598 136350
rect 260654 136294 260722 136350
rect 260778 136294 291318 136350
rect 291374 136294 291442 136350
rect 291498 136294 322038 136350
rect 322094 136294 322162 136350
rect 322218 136294 352758 136350
rect 352814 136294 352882 136350
rect 352938 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 470034 136350
rect 470090 136294 470158 136350
rect 470214 136294 470282 136350
rect 470338 136294 470406 136350
rect 470462 136294 500754 136350
rect 500810 136294 500878 136350
rect 500934 136294 501002 136350
rect 501058 136294 501126 136350
rect 501182 136294 531474 136350
rect 531530 136294 531598 136350
rect 531654 136294 531722 136350
rect 531778 136294 531846 136350
rect 531902 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 11930 136226
rect 11986 136170 12054 136226
rect 12110 136170 12178 136226
rect 12234 136170 12302 136226
rect 12358 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 70674 136226
rect 70730 136170 70798 136226
rect 70854 136170 70922 136226
rect 70978 136170 71046 136226
rect 71102 136170 96612 136226
rect 96668 136170 96736 136226
rect 96792 136170 96860 136226
rect 96916 136170 96984 136226
rect 97040 136170 101394 136226
rect 101450 136170 101518 136226
rect 101574 136170 101642 136226
rect 101698 136170 101766 136226
rect 101822 136170 111930 136226
rect 111986 136170 112054 136226
rect 112110 136170 112178 136226
rect 112234 136170 112302 136226
rect 112358 136170 132114 136226
rect 132170 136170 132238 136226
rect 132294 136170 132362 136226
rect 132418 136170 132486 136226
rect 132542 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 193554 136226
rect 193610 136170 193678 136226
rect 193734 136170 193802 136226
rect 193858 136170 193926 136226
rect 193982 136170 196612 136226
rect 196668 136170 196736 136226
rect 196792 136170 196860 136226
rect 196916 136170 196984 136226
rect 197040 136170 229878 136226
rect 229934 136170 230002 136226
rect 230058 136170 260598 136226
rect 260654 136170 260722 136226
rect 260778 136170 291318 136226
rect 291374 136170 291442 136226
rect 291498 136170 322038 136226
rect 322094 136170 322162 136226
rect 322218 136170 352758 136226
rect 352814 136170 352882 136226
rect 352938 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 470034 136226
rect 470090 136170 470158 136226
rect 470214 136170 470282 136226
rect 470338 136170 470406 136226
rect 470462 136170 500754 136226
rect 500810 136170 500878 136226
rect 500934 136170 501002 136226
rect 501058 136170 501126 136226
rect 501182 136170 531474 136226
rect 531530 136170 531598 136226
rect 531654 136170 531722 136226
rect 531778 136170 531846 136226
rect 531902 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 11930 136102
rect 11986 136046 12054 136102
rect 12110 136046 12178 136102
rect 12234 136046 12302 136102
rect 12358 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 70674 136102
rect 70730 136046 70798 136102
rect 70854 136046 70922 136102
rect 70978 136046 71046 136102
rect 71102 136046 96612 136102
rect 96668 136046 96736 136102
rect 96792 136046 96860 136102
rect 96916 136046 96984 136102
rect 97040 136046 101394 136102
rect 101450 136046 101518 136102
rect 101574 136046 101642 136102
rect 101698 136046 101766 136102
rect 101822 136046 111930 136102
rect 111986 136046 112054 136102
rect 112110 136046 112178 136102
rect 112234 136046 112302 136102
rect 112358 136046 132114 136102
rect 132170 136046 132238 136102
rect 132294 136046 132362 136102
rect 132418 136046 132486 136102
rect 132542 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 193554 136102
rect 193610 136046 193678 136102
rect 193734 136046 193802 136102
rect 193858 136046 193926 136102
rect 193982 136046 196612 136102
rect 196668 136046 196736 136102
rect 196792 136046 196860 136102
rect 196916 136046 196984 136102
rect 197040 136046 229878 136102
rect 229934 136046 230002 136102
rect 230058 136046 260598 136102
rect 260654 136046 260722 136102
rect 260778 136046 291318 136102
rect 291374 136046 291442 136102
rect 291498 136046 322038 136102
rect 322094 136046 322162 136102
rect 322218 136046 352758 136102
rect 352814 136046 352882 136102
rect 352938 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 470034 136102
rect 470090 136046 470158 136102
rect 470214 136046 470282 136102
rect 470338 136046 470406 136102
rect 470462 136046 500754 136102
rect 500810 136046 500878 136102
rect 500934 136046 501002 136102
rect 501058 136046 501126 136102
rect 501182 136046 531474 136102
rect 531530 136046 531598 136102
rect 531654 136046 531722 136102
rect 531778 136046 531846 136102
rect 531902 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 11930 135978
rect 11986 135922 12054 135978
rect 12110 135922 12178 135978
rect 12234 135922 12302 135978
rect 12358 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 70674 135978
rect 70730 135922 70798 135978
rect 70854 135922 70922 135978
rect 70978 135922 71046 135978
rect 71102 135922 96612 135978
rect 96668 135922 96736 135978
rect 96792 135922 96860 135978
rect 96916 135922 96984 135978
rect 97040 135922 101394 135978
rect 101450 135922 101518 135978
rect 101574 135922 101642 135978
rect 101698 135922 101766 135978
rect 101822 135922 111930 135978
rect 111986 135922 112054 135978
rect 112110 135922 112178 135978
rect 112234 135922 112302 135978
rect 112358 135922 132114 135978
rect 132170 135922 132238 135978
rect 132294 135922 132362 135978
rect 132418 135922 132486 135978
rect 132542 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 193554 135978
rect 193610 135922 193678 135978
rect 193734 135922 193802 135978
rect 193858 135922 193926 135978
rect 193982 135922 196612 135978
rect 196668 135922 196736 135978
rect 196792 135922 196860 135978
rect 196916 135922 196984 135978
rect 197040 135922 229878 135978
rect 229934 135922 230002 135978
rect 230058 135922 260598 135978
rect 260654 135922 260722 135978
rect 260778 135922 291318 135978
rect 291374 135922 291442 135978
rect 291498 135922 322038 135978
rect 322094 135922 322162 135978
rect 322218 135922 352758 135978
rect 352814 135922 352882 135978
rect 352938 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 470034 135978
rect 470090 135922 470158 135978
rect 470214 135922 470282 135978
rect 470338 135922 470406 135978
rect 470462 135922 500754 135978
rect 500810 135922 500878 135978
rect 500934 135922 501002 135978
rect 501058 135922 501126 135978
rect 501182 135922 531474 135978
rect 531530 135922 531598 135978
rect 531654 135922 531722 135978
rect 531778 135922 531846 135978
rect 531902 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect 376892 133678 441940 133694
rect 376892 133622 376908 133678
rect 376964 133622 441868 133678
rect 441924 133622 441940 133678
rect 376892 133606 441940 133622
rect 375324 133498 442052 133514
rect 375324 133442 375340 133498
rect 375396 133442 441980 133498
rect 442036 133442 442052 133498
rect 375324 133426 442052 133442
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 11130 130350
rect 11186 130294 11254 130350
rect 11310 130294 11378 130350
rect 11434 130294 11502 130350
rect 11558 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 66954 130350
rect 67010 130294 67078 130350
rect 67134 130294 67202 130350
rect 67258 130294 67326 130350
rect 67382 130294 95812 130350
rect 95868 130294 95936 130350
rect 95992 130294 96060 130350
rect 96116 130294 96184 130350
rect 96240 130294 97674 130350
rect 97730 130294 97798 130350
rect 97854 130294 97922 130350
rect 97978 130294 98046 130350
rect 98102 130294 111130 130350
rect 111186 130294 111254 130350
rect 111310 130294 111378 130350
rect 111434 130294 111502 130350
rect 111558 130294 128394 130350
rect 128450 130294 128518 130350
rect 128574 130294 128642 130350
rect 128698 130294 128766 130350
rect 128822 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 189834 130350
rect 189890 130294 189958 130350
rect 190014 130294 190082 130350
rect 190138 130294 190206 130350
rect 190262 130294 195812 130350
rect 195868 130294 195936 130350
rect 195992 130294 196060 130350
rect 196116 130294 196184 130350
rect 196240 130294 214518 130350
rect 214574 130294 214642 130350
rect 214698 130294 245238 130350
rect 245294 130294 245362 130350
rect 245418 130294 275958 130350
rect 276014 130294 276082 130350
rect 276138 130294 306678 130350
rect 306734 130294 306802 130350
rect 306858 130294 337398 130350
rect 337454 130294 337522 130350
rect 337578 130294 368118 130350
rect 368174 130294 368242 130350
rect 368298 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 466314 130350
rect 466370 130294 466438 130350
rect 466494 130294 466562 130350
rect 466618 130294 466686 130350
rect 466742 130294 497034 130350
rect 497090 130294 497158 130350
rect 497214 130294 497282 130350
rect 497338 130294 497406 130350
rect 497462 130294 527754 130350
rect 527810 130294 527878 130350
rect 527934 130294 528002 130350
rect 528058 130294 528126 130350
rect 528182 130294 558474 130350
rect 558530 130294 558598 130350
rect 558654 130294 558722 130350
rect 558778 130294 558846 130350
rect 558902 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 11130 130226
rect 11186 130170 11254 130226
rect 11310 130170 11378 130226
rect 11434 130170 11502 130226
rect 11558 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 66954 130226
rect 67010 130170 67078 130226
rect 67134 130170 67202 130226
rect 67258 130170 67326 130226
rect 67382 130170 95812 130226
rect 95868 130170 95936 130226
rect 95992 130170 96060 130226
rect 96116 130170 96184 130226
rect 96240 130170 97674 130226
rect 97730 130170 97798 130226
rect 97854 130170 97922 130226
rect 97978 130170 98046 130226
rect 98102 130170 111130 130226
rect 111186 130170 111254 130226
rect 111310 130170 111378 130226
rect 111434 130170 111502 130226
rect 111558 130170 128394 130226
rect 128450 130170 128518 130226
rect 128574 130170 128642 130226
rect 128698 130170 128766 130226
rect 128822 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 189834 130226
rect 189890 130170 189958 130226
rect 190014 130170 190082 130226
rect 190138 130170 190206 130226
rect 190262 130170 195812 130226
rect 195868 130170 195936 130226
rect 195992 130170 196060 130226
rect 196116 130170 196184 130226
rect 196240 130170 214518 130226
rect 214574 130170 214642 130226
rect 214698 130170 245238 130226
rect 245294 130170 245362 130226
rect 245418 130170 275958 130226
rect 276014 130170 276082 130226
rect 276138 130170 306678 130226
rect 306734 130170 306802 130226
rect 306858 130170 337398 130226
rect 337454 130170 337522 130226
rect 337578 130170 368118 130226
rect 368174 130170 368242 130226
rect 368298 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 466314 130226
rect 466370 130170 466438 130226
rect 466494 130170 466562 130226
rect 466618 130170 466686 130226
rect 466742 130170 497034 130226
rect 497090 130170 497158 130226
rect 497214 130170 497282 130226
rect 497338 130170 497406 130226
rect 497462 130170 527754 130226
rect 527810 130170 527878 130226
rect 527934 130170 528002 130226
rect 528058 130170 528126 130226
rect 528182 130170 558474 130226
rect 558530 130170 558598 130226
rect 558654 130170 558722 130226
rect 558778 130170 558846 130226
rect 558902 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 11130 130102
rect 11186 130046 11254 130102
rect 11310 130046 11378 130102
rect 11434 130046 11502 130102
rect 11558 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 66954 130102
rect 67010 130046 67078 130102
rect 67134 130046 67202 130102
rect 67258 130046 67326 130102
rect 67382 130046 95812 130102
rect 95868 130046 95936 130102
rect 95992 130046 96060 130102
rect 96116 130046 96184 130102
rect 96240 130046 97674 130102
rect 97730 130046 97798 130102
rect 97854 130046 97922 130102
rect 97978 130046 98046 130102
rect 98102 130046 111130 130102
rect 111186 130046 111254 130102
rect 111310 130046 111378 130102
rect 111434 130046 111502 130102
rect 111558 130046 128394 130102
rect 128450 130046 128518 130102
rect 128574 130046 128642 130102
rect 128698 130046 128766 130102
rect 128822 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 189834 130102
rect 189890 130046 189958 130102
rect 190014 130046 190082 130102
rect 190138 130046 190206 130102
rect 190262 130046 195812 130102
rect 195868 130046 195936 130102
rect 195992 130046 196060 130102
rect 196116 130046 196184 130102
rect 196240 130046 214518 130102
rect 214574 130046 214642 130102
rect 214698 130046 245238 130102
rect 245294 130046 245362 130102
rect 245418 130046 275958 130102
rect 276014 130046 276082 130102
rect 276138 130046 306678 130102
rect 306734 130046 306802 130102
rect 306858 130046 337398 130102
rect 337454 130046 337522 130102
rect 337578 130046 368118 130102
rect 368174 130046 368242 130102
rect 368298 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 466314 130102
rect 466370 130046 466438 130102
rect 466494 130046 466562 130102
rect 466618 130046 466686 130102
rect 466742 130046 497034 130102
rect 497090 130046 497158 130102
rect 497214 130046 497282 130102
rect 497338 130046 497406 130102
rect 497462 130046 527754 130102
rect 527810 130046 527878 130102
rect 527934 130046 528002 130102
rect 528058 130046 528126 130102
rect 528182 130046 558474 130102
rect 558530 130046 558598 130102
rect 558654 130046 558722 130102
rect 558778 130046 558846 130102
rect 558902 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 11130 129978
rect 11186 129922 11254 129978
rect 11310 129922 11378 129978
rect 11434 129922 11502 129978
rect 11558 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 66954 129978
rect 67010 129922 67078 129978
rect 67134 129922 67202 129978
rect 67258 129922 67326 129978
rect 67382 129922 95812 129978
rect 95868 129922 95936 129978
rect 95992 129922 96060 129978
rect 96116 129922 96184 129978
rect 96240 129922 97674 129978
rect 97730 129922 97798 129978
rect 97854 129922 97922 129978
rect 97978 129922 98046 129978
rect 98102 129922 111130 129978
rect 111186 129922 111254 129978
rect 111310 129922 111378 129978
rect 111434 129922 111502 129978
rect 111558 129922 128394 129978
rect 128450 129922 128518 129978
rect 128574 129922 128642 129978
rect 128698 129922 128766 129978
rect 128822 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 189834 129978
rect 189890 129922 189958 129978
rect 190014 129922 190082 129978
rect 190138 129922 190206 129978
rect 190262 129922 195812 129978
rect 195868 129922 195936 129978
rect 195992 129922 196060 129978
rect 196116 129922 196184 129978
rect 196240 129922 214518 129978
rect 214574 129922 214642 129978
rect 214698 129922 245238 129978
rect 245294 129922 245362 129978
rect 245418 129922 275958 129978
rect 276014 129922 276082 129978
rect 276138 129922 306678 129978
rect 306734 129922 306802 129978
rect 306858 129922 337398 129978
rect 337454 129922 337522 129978
rect 337578 129922 368118 129978
rect 368174 129922 368242 129978
rect 368298 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 466314 129978
rect 466370 129922 466438 129978
rect 466494 129922 466562 129978
rect 466618 129922 466686 129978
rect 466742 129922 497034 129978
rect 497090 129922 497158 129978
rect 497214 129922 497282 129978
rect 497338 129922 497406 129978
rect 497462 129922 527754 129978
rect 527810 129922 527878 129978
rect 527934 129922 528002 129978
rect 528058 129922 528126 129978
rect 528182 129922 558474 129978
rect 558530 129922 558598 129978
rect 558654 129922 558722 129978
rect 558778 129922 558846 129978
rect 558902 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect 373868 120898 440708 120914
rect 373868 120842 373884 120898
rect 373940 120842 440636 120898
rect 440692 120842 440708 120898
rect 373868 120826 440708 120842
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 11930 118350
rect 11986 118294 12054 118350
rect 12110 118294 12178 118350
rect 12234 118294 12302 118350
rect 12358 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 70674 118350
rect 70730 118294 70798 118350
rect 70854 118294 70922 118350
rect 70978 118294 71046 118350
rect 71102 118294 96612 118350
rect 96668 118294 96736 118350
rect 96792 118294 96860 118350
rect 96916 118294 96984 118350
rect 97040 118294 101394 118350
rect 101450 118294 101518 118350
rect 101574 118294 101642 118350
rect 101698 118294 101766 118350
rect 101822 118294 111930 118350
rect 111986 118294 112054 118350
rect 112110 118294 112178 118350
rect 112234 118294 112302 118350
rect 112358 118294 132114 118350
rect 132170 118294 132238 118350
rect 132294 118294 132362 118350
rect 132418 118294 132486 118350
rect 132542 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 193554 118350
rect 193610 118294 193678 118350
rect 193734 118294 193802 118350
rect 193858 118294 193926 118350
rect 193982 118294 196612 118350
rect 196668 118294 196736 118350
rect 196792 118294 196860 118350
rect 196916 118294 196984 118350
rect 197040 118294 229878 118350
rect 229934 118294 230002 118350
rect 230058 118294 260598 118350
rect 260654 118294 260722 118350
rect 260778 118294 291318 118350
rect 291374 118294 291442 118350
rect 291498 118294 322038 118350
rect 322094 118294 322162 118350
rect 322218 118294 352758 118350
rect 352814 118294 352882 118350
rect 352938 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 399878 118350
rect 399934 118294 400002 118350
rect 400058 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 430598 118350
rect 430654 118294 430722 118350
rect 430778 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 470034 118350
rect 470090 118294 470158 118350
rect 470214 118294 470282 118350
rect 470338 118294 470406 118350
rect 470462 118294 500754 118350
rect 500810 118294 500878 118350
rect 500934 118294 501002 118350
rect 501058 118294 501126 118350
rect 501182 118294 531474 118350
rect 531530 118294 531598 118350
rect 531654 118294 531722 118350
rect 531778 118294 531846 118350
rect 531902 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 11930 118226
rect 11986 118170 12054 118226
rect 12110 118170 12178 118226
rect 12234 118170 12302 118226
rect 12358 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 70674 118226
rect 70730 118170 70798 118226
rect 70854 118170 70922 118226
rect 70978 118170 71046 118226
rect 71102 118170 96612 118226
rect 96668 118170 96736 118226
rect 96792 118170 96860 118226
rect 96916 118170 96984 118226
rect 97040 118170 101394 118226
rect 101450 118170 101518 118226
rect 101574 118170 101642 118226
rect 101698 118170 101766 118226
rect 101822 118170 111930 118226
rect 111986 118170 112054 118226
rect 112110 118170 112178 118226
rect 112234 118170 112302 118226
rect 112358 118170 132114 118226
rect 132170 118170 132238 118226
rect 132294 118170 132362 118226
rect 132418 118170 132486 118226
rect 132542 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 193554 118226
rect 193610 118170 193678 118226
rect 193734 118170 193802 118226
rect 193858 118170 193926 118226
rect 193982 118170 196612 118226
rect 196668 118170 196736 118226
rect 196792 118170 196860 118226
rect 196916 118170 196984 118226
rect 197040 118170 229878 118226
rect 229934 118170 230002 118226
rect 230058 118170 260598 118226
rect 260654 118170 260722 118226
rect 260778 118170 291318 118226
rect 291374 118170 291442 118226
rect 291498 118170 322038 118226
rect 322094 118170 322162 118226
rect 322218 118170 352758 118226
rect 352814 118170 352882 118226
rect 352938 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 399878 118226
rect 399934 118170 400002 118226
rect 400058 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 430598 118226
rect 430654 118170 430722 118226
rect 430778 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 470034 118226
rect 470090 118170 470158 118226
rect 470214 118170 470282 118226
rect 470338 118170 470406 118226
rect 470462 118170 500754 118226
rect 500810 118170 500878 118226
rect 500934 118170 501002 118226
rect 501058 118170 501126 118226
rect 501182 118170 531474 118226
rect 531530 118170 531598 118226
rect 531654 118170 531722 118226
rect 531778 118170 531846 118226
rect 531902 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 11930 118102
rect 11986 118046 12054 118102
rect 12110 118046 12178 118102
rect 12234 118046 12302 118102
rect 12358 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 70674 118102
rect 70730 118046 70798 118102
rect 70854 118046 70922 118102
rect 70978 118046 71046 118102
rect 71102 118046 96612 118102
rect 96668 118046 96736 118102
rect 96792 118046 96860 118102
rect 96916 118046 96984 118102
rect 97040 118046 101394 118102
rect 101450 118046 101518 118102
rect 101574 118046 101642 118102
rect 101698 118046 101766 118102
rect 101822 118046 111930 118102
rect 111986 118046 112054 118102
rect 112110 118046 112178 118102
rect 112234 118046 112302 118102
rect 112358 118046 132114 118102
rect 132170 118046 132238 118102
rect 132294 118046 132362 118102
rect 132418 118046 132486 118102
rect 132542 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 193554 118102
rect 193610 118046 193678 118102
rect 193734 118046 193802 118102
rect 193858 118046 193926 118102
rect 193982 118046 196612 118102
rect 196668 118046 196736 118102
rect 196792 118046 196860 118102
rect 196916 118046 196984 118102
rect 197040 118046 229878 118102
rect 229934 118046 230002 118102
rect 230058 118046 260598 118102
rect 260654 118046 260722 118102
rect 260778 118046 291318 118102
rect 291374 118046 291442 118102
rect 291498 118046 322038 118102
rect 322094 118046 322162 118102
rect 322218 118046 352758 118102
rect 352814 118046 352882 118102
rect 352938 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 399878 118102
rect 399934 118046 400002 118102
rect 400058 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 430598 118102
rect 430654 118046 430722 118102
rect 430778 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 470034 118102
rect 470090 118046 470158 118102
rect 470214 118046 470282 118102
rect 470338 118046 470406 118102
rect 470462 118046 500754 118102
rect 500810 118046 500878 118102
rect 500934 118046 501002 118102
rect 501058 118046 501126 118102
rect 501182 118046 531474 118102
rect 531530 118046 531598 118102
rect 531654 118046 531722 118102
rect 531778 118046 531846 118102
rect 531902 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 11930 117978
rect 11986 117922 12054 117978
rect 12110 117922 12178 117978
rect 12234 117922 12302 117978
rect 12358 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 70674 117978
rect 70730 117922 70798 117978
rect 70854 117922 70922 117978
rect 70978 117922 71046 117978
rect 71102 117922 96612 117978
rect 96668 117922 96736 117978
rect 96792 117922 96860 117978
rect 96916 117922 96984 117978
rect 97040 117922 101394 117978
rect 101450 117922 101518 117978
rect 101574 117922 101642 117978
rect 101698 117922 101766 117978
rect 101822 117922 111930 117978
rect 111986 117922 112054 117978
rect 112110 117922 112178 117978
rect 112234 117922 112302 117978
rect 112358 117922 132114 117978
rect 132170 117922 132238 117978
rect 132294 117922 132362 117978
rect 132418 117922 132486 117978
rect 132542 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 193554 117978
rect 193610 117922 193678 117978
rect 193734 117922 193802 117978
rect 193858 117922 193926 117978
rect 193982 117922 196612 117978
rect 196668 117922 196736 117978
rect 196792 117922 196860 117978
rect 196916 117922 196984 117978
rect 197040 117922 229878 117978
rect 229934 117922 230002 117978
rect 230058 117922 260598 117978
rect 260654 117922 260722 117978
rect 260778 117922 291318 117978
rect 291374 117922 291442 117978
rect 291498 117922 322038 117978
rect 322094 117922 322162 117978
rect 322218 117922 352758 117978
rect 352814 117922 352882 117978
rect 352938 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 399878 117978
rect 399934 117922 400002 117978
rect 400058 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 430598 117978
rect 430654 117922 430722 117978
rect 430778 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 470034 117978
rect 470090 117922 470158 117978
rect 470214 117922 470282 117978
rect 470338 117922 470406 117978
rect 470462 117922 500754 117978
rect 500810 117922 500878 117978
rect 500934 117922 501002 117978
rect 501058 117922 501126 117978
rect 501182 117922 531474 117978
rect 531530 117922 531598 117978
rect 531654 117922 531722 117978
rect 531778 117922 531846 117978
rect 531902 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect 380140 117478 442164 117494
rect 380140 117422 380156 117478
rect 380212 117422 442092 117478
rect 442148 117422 442164 117478
rect 380140 117406 442164 117422
rect 396380 116038 398260 116054
rect 396380 115982 396396 116038
rect 396452 115982 398188 116038
rect 398244 115982 398260 116038
rect 396380 115966 398260 115982
rect 379580 115858 440596 115874
rect 379580 115802 379596 115858
rect 379652 115802 440524 115858
rect 440580 115802 440596 115858
rect 379580 115786 440596 115802
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 11130 112350
rect 11186 112294 11254 112350
rect 11310 112294 11378 112350
rect 11434 112294 11502 112350
rect 11558 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 66954 112350
rect 67010 112294 67078 112350
rect 67134 112294 67202 112350
rect 67258 112294 67326 112350
rect 67382 112294 95812 112350
rect 95868 112294 95936 112350
rect 95992 112294 96060 112350
rect 96116 112294 96184 112350
rect 96240 112294 97674 112350
rect 97730 112294 97798 112350
rect 97854 112294 97922 112350
rect 97978 112294 98046 112350
rect 98102 112294 111130 112350
rect 111186 112294 111254 112350
rect 111310 112294 111378 112350
rect 111434 112294 111502 112350
rect 111558 112294 128394 112350
rect 128450 112294 128518 112350
rect 128574 112294 128642 112350
rect 128698 112294 128766 112350
rect 128822 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 189834 112350
rect 189890 112294 189958 112350
rect 190014 112294 190082 112350
rect 190138 112294 190206 112350
rect 190262 112294 195812 112350
rect 195868 112294 195936 112350
rect 195992 112294 196060 112350
rect 196116 112294 196184 112350
rect 196240 112294 214518 112350
rect 214574 112294 214642 112350
rect 214698 112294 245238 112350
rect 245294 112294 245362 112350
rect 245418 112294 275958 112350
rect 276014 112294 276082 112350
rect 276138 112294 306678 112350
rect 306734 112294 306802 112350
rect 306858 112294 337398 112350
rect 337454 112294 337522 112350
rect 337578 112294 368118 112350
rect 368174 112294 368242 112350
rect 368298 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 384518 112350
rect 384574 112294 384642 112350
rect 384698 112294 415238 112350
rect 415294 112294 415362 112350
rect 415418 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 466314 112350
rect 466370 112294 466438 112350
rect 466494 112294 466562 112350
rect 466618 112294 466686 112350
rect 466742 112294 497034 112350
rect 497090 112294 497158 112350
rect 497214 112294 497282 112350
rect 497338 112294 497406 112350
rect 497462 112294 527754 112350
rect 527810 112294 527878 112350
rect 527934 112294 528002 112350
rect 528058 112294 528126 112350
rect 528182 112294 558474 112350
rect 558530 112294 558598 112350
rect 558654 112294 558722 112350
rect 558778 112294 558846 112350
rect 558902 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 11130 112226
rect 11186 112170 11254 112226
rect 11310 112170 11378 112226
rect 11434 112170 11502 112226
rect 11558 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 66954 112226
rect 67010 112170 67078 112226
rect 67134 112170 67202 112226
rect 67258 112170 67326 112226
rect 67382 112170 95812 112226
rect 95868 112170 95936 112226
rect 95992 112170 96060 112226
rect 96116 112170 96184 112226
rect 96240 112170 97674 112226
rect 97730 112170 97798 112226
rect 97854 112170 97922 112226
rect 97978 112170 98046 112226
rect 98102 112170 111130 112226
rect 111186 112170 111254 112226
rect 111310 112170 111378 112226
rect 111434 112170 111502 112226
rect 111558 112170 128394 112226
rect 128450 112170 128518 112226
rect 128574 112170 128642 112226
rect 128698 112170 128766 112226
rect 128822 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 189834 112226
rect 189890 112170 189958 112226
rect 190014 112170 190082 112226
rect 190138 112170 190206 112226
rect 190262 112170 195812 112226
rect 195868 112170 195936 112226
rect 195992 112170 196060 112226
rect 196116 112170 196184 112226
rect 196240 112170 214518 112226
rect 214574 112170 214642 112226
rect 214698 112170 245238 112226
rect 245294 112170 245362 112226
rect 245418 112170 275958 112226
rect 276014 112170 276082 112226
rect 276138 112170 306678 112226
rect 306734 112170 306802 112226
rect 306858 112170 337398 112226
rect 337454 112170 337522 112226
rect 337578 112170 368118 112226
rect 368174 112170 368242 112226
rect 368298 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 384518 112226
rect 384574 112170 384642 112226
rect 384698 112170 415238 112226
rect 415294 112170 415362 112226
rect 415418 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 466314 112226
rect 466370 112170 466438 112226
rect 466494 112170 466562 112226
rect 466618 112170 466686 112226
rect 466742 112170 497034 112226
rect 497090 112170 497158 112226
rect 497214 112170 497282 112226
rect 497338 112170 497406 112226
rect 497462 112170 527754 112226
rect 527810 112170 527878 112226
rect 527934 112170 528002 112226
rect 528058 112170 528126 112226
rect 528182 112170 558474 112226
rect 558530 112170 558598 112226
rect 558654 112170 558722 112226
rect 558778 112170 558846 112226
rect 558902 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 11130 112102
rect 11186 112046 11254 112102
rect 11310 112046 11378 112102
rect 11434 112046 11502 112102
rect 11558 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 66954 112102
rect 67010 112046 67078 112102
rect 67134 112046 67202 112102
rect 67258 112046 67326 112102
rect 67382 112046 95812 112102
rect 95868 112046 95936 112102
rect 95992 112046 96060 112102
rect 96116 112046 96184 112102
rect 96240 112046 97674 112102
rect 97730 112046 97798 112102
rect 97854 112046 97922 112102
rect 97978 112046 98046 112102
rect 98102 112046 111130 112102
rect 111186 112046 111254 112102
rect 111310 112046 111378 112102
rect 111434 112046 111502 112102
rect 111558 112046 128394 112102
rect 128450 112046 128518 112102
rect 128574 112046 128642 112102
rect 128698 112046 128766 112102
rect 128822 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 189834 112102
rect 189890 112046 189958 112102
rect 190014 112046 190082 112102
rect 190138 112046 190206 112102
rect 190262 112046 195812 112102
rect 195868 112046 195936 112102
rect 195992 112046 196060 112102
rect 196116 112046 196184 112102
rect 196240 112046 214518 112102
rect 214574 112046 214642 112102
rect 214698 112046 245238 112102
rect 245294 112046 245362 112102
rect 245418 112046 275958 112102
rect 276014 112046 276082 112102
rect 276138 112046 306678 112102
rect 306734 112046 306802 112102
rect 306858 112046 337398 112102
rect 337454 112046 337522 112102
rect 337578 112046 368118 112102
rect 368174 112046 368242 112102
rect 368298 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 384518 112102
rect 384574 112046 384642 112102
rect 384698 112046 415238 112102
rect 415294 112046 415362 112102
rect 415418 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 466314 112102
rect 466370 112046 466438 112102
rect 466494 112046 466562 112102
rect 466618 112046 466686 112102
rect 466742 112046 497034 112102
rect 497090 112046 497158 112102
rect 497214 112046 497282 112102
rect 497338 112046 497406 112102
rect 497462 112046 527754 112102
rect 527810 112046 527878 112102
rect 527934 112046 528002 112102
rect 528058 112046 528126 112102
rect 528182 112046 558474 112102
rect 558530 112046 558598 112102
rect 558654 112046 558722 112102
rect 558778 112046 558846 112102
rect 558902 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 11130 111978
rect 11186 111922 11254 111978
rect 11310 111922 11378 111978
rect 11434 111922 11502 111978
rect 11558 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 66954 111978
rect 67010 111922 67078 111978
rect 67134 111922 67202 111978
rect 67258 111922 67326 111978
rect 67382 111922 95812 111978
rect 95868 111922 95936 111978
rect 95992 111922 96060 111978
rect 96116 111922 96184 111978
rect 96240 111922 97674 111978
rect 97730 111922 97798 111978
rect 97854 111922 97922 111978
rect 97978 111922 98046 111978
rect 98102 111922 111130 111978
rect 111186 111922 111254 111978
rect 111310 111922 111378 111978
rect 111434 111922 111502 111978
rect 111558 111922 128394 111978
rect 128450 111922 128518 111978
rect 128574 111922 128642 111978
rect 128698 111922 128766 111978
rect 128822 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 189834 111978
rect 189890 111922 189958 111978
rect 190014 111922 190082 111978
rect 190138 111922 190206 111978
rect 190262 111922 195812 111978
rect 195868 111922 195936 111978
rect 195992 111922 196060 111978
rect 196116 111922 196184 111978
rect 196240 111922 214518 111978
rect 214574 111922 214642 111978
rect 214698 111922 245238 111978
rect 245294 111922 245362 111978
rect 245418 111922 275958 111978
rect 276014 111922 276082 111978
rect 276138 111922 306678 111978
rect 306734 111922 306802 111978
rect 306858 111922 337398 111978
rect 337454 111922 337522 111978
rect 337578 111922 368118 111978
rect 368174 111922 368242 111978
rect 368298 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 384518 111978
rect 384574 111922 384642 111978
rect 384698 111922 415238 111978
rect 415294 111922 415362 111978
rect 415418 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 466314 111978
rect 466370 111922 466438 111978
rect 466494 111922 466562 111978
rect 466618 111922 466686 111978
rect 466742 111922 497034 111978
rect 497090 111922 497158 111978
rect 497214 111922 497282 111978
rect 497338 111922 497406 111978
rect 497462 111922 527754 111978
rect 527810 111922 527878 111978
rect 527934 111922 528002 111978
rect 528058 111922 528126 111978
rect 528182 111922 558474 111978
rect 558530 111922 558598 111978
rect 558654 111922 558722 111978
rect 558778 111922 558846 111978
rect 558902 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect 376108 105778 392436 105794
rect 376108 105722 376124 105778
rect 376180 105722 392364 105778
rect 392420 105722 392436 105778
rect 376108 105706 392436 105722
rect 377564 101638 384764 101654
rect 377564 101582 377580 101638
rect 377636 101582 384764 101638
rect 377564 101566 384764 101582
rect 384676 100934 384764 101566
rect 384676 100918 392548 100934
rect 384676 100862 391468 100918
rect 391524 100862 392476 100918
rect 392532 100862 392548 100918
rect 384676 100846 392548 100862
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 11930 100350
rect 11986 100294 12054 100350
rect 12110 100294 12178 100350
rect 12234 100294 12302 100350
rect 12358 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 70674 100350
rect 70730 100294 70798 100350
rect 70854 100294 70922 100350
rect 70978 100294 71046 100350
rect 71102 100294 96612 100350
rect 96668 100294 96736 100350
rect 96792 100294 96860 100350
rect 96916 100294 96984 100350
rect 97040 100294 101394 100350
rect 101450 100294 101518 100350
rect 101574 100294 101642 100350
rect 101698 100294 101766 100350
rect 101822 100294 111930 100350
rect 111986 100294 112054 100350
rect 112110 100294 112178 100350
rect 112234 100294 112302 100350
rect 112358 100294 132114 100350
rect 132170 100294 132238 100350
rect 132294 100294 132362 100350
rect 132418 100294 132486 100350
rect 132542 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 193554 100350
rect 193610 100294 193678 100350
rect 193734 100294 193802 100350
rect 193858 100294 193926 100350
rect 193982 100294 196612 100350
rect 196668 100294 196736 100350
rect 196792 100294 196860 100350
rect 196916 100294 196984 100350
rect 197040 100294 229878 100350
rect 229934 100294 230002 100350
rect 230058 100294 260598 100350
rect 260654 100294 260722 100350
rect 260778 100294 291318 100350
rect 291374 100294 291442 100350
rect 291498 100294 322038 100350
rect 322094 100294 322162 100350
rect 322218 100294 352758 100350
rect 352814 100294 352882 100350
rect 352938 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 399878 100350
rect 399934 100294 400002 100350
rect 400058 100294 430598 100350
rect 430654 100294 430722 100350
rect 430778 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 470034 100350
rect 470090 100294 470158 100350
rect 470214 100294 470282 100350
rect 470338 100294 470406 100350
rect 470462 100294 500754 100350
rect 500810 100294 500878 100350
rect 500934 100294 501002 100350
rect 501058 100294 501126 100350
rect 501182 100294 531474 100350
rect 531530 100294 531598 100350
rect 531654 100294 531722 100350
rect 531778 100294 531846 100350
rect 531902 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 11930 100226
rect 11986 100170 12054 100226
rect 12110 100170 12178 100226
rect 12234 100170 12302 100226
rect 12358 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 70674 100226
rect 70730 100170 70798 100226
rect 70854 100170 70922 100226
rect 70978 100170 71046 100226
rect 71102 100170 96612 100226
rect 96668 100170 96736 100226
rect 96792 100170 96860 100226
rect 96916 100170 96984 100226
rect 97040 100170 101394 100226
rect 101450 100170 101518 100226
rect 101574 100170 101642 100226
rect 101698 100170 101766 100226
rect 101822 100170 111930 100226
rect 111986 100170 112054 100226
rect 112110 100170 112178 100226
rect 112234 100170 112302 100226
rect 112358 100170 132114 100226
rect 132170 100170 132238 100226
rect 132294 100170 132362 100226
rect 132418 100170 132486 100226
rect 132542 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 193554 100226
rect 193610 100170 193678 100226
rect 193734 100170 193802 100226
rect 193858 100170 193926 100226
rect 193982 100170 196612 100226
rect 196668 100170 196736 100226
rect 196792 100170 196860 100226
rect 196916 100170 196984 100226
rect 197040 100170 229878 100226
rect 229934 100170 230002 100226
rect 230058 100170 260598 100226
rect 260654 100170 260722 100226
rect 260778 100170 291318 100226
rect 291374 100170 291442 100226
rect 291498 100170 322038 100226
rect 322094 100170 322162 100226
rect 322218 100170 352758 100226
rect 352814 100170 352882 100226
rect 352938 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 399878 100226
rect 399934 100170 400002 100226
rect 400058 100170 430598 100226
rect 430654 100170 430722 100226
rect 430778 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 470034 100226
rect 470090 100170 470158 100226
rect 470214 100170 470282 100226
rect 470338 100170 470406 100226
rect 470462 100170 500754 100226
rect 500810 100170 500878 100226
rect 500934 100170 501002 100226
rect 501058 100170 501126 100226
rect 501182 100170 531474 100226
rect 531530 100170 531598 100226
rect 531654 100170 531722 100226
rect 531778 100170 531846 100226
rect 531902 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 11930 100102
rect 11986 100046 12054 100102
rect 12110 100046 12178 100102
rect 12234 100046 12302 100102
rect 12358 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 70674 100102
rect 70730 100046 70798 100102
rect 70854 100046 70922 100102
rect 70978 100046 71046 100102
rect 71102 100046 96612 100102
rect 96668 100046 96736 100102
rect 96792 100046 96860 100102
rect 96916 100046 96984 100102
rect 97040 100046 101394 100102
rect 101450 100046 101518 100102
rect 101574 100046 101642 100102
rect 101698 100046 101766 100102
rect 101822 100046 111930 100102
rect 111986 100046 112054 100102
rect 112110 100046 112178 100102
rect 112234 100046 112302 100102
rect 112358 100046 132114 100102
rect 132170 100046 132238 100102
rect 132294 100046 132362 100102
rect 132418 100046 132486 100102
rect 132542 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 193554 100102
rect 193610 100046 193678 100102
rect 193734 100046 193802 100102
rect 193858 100046 193926 100102
rect 193982 100046 196612 100102
rect 196668 100046 196736 100102
rect 196792 100046 196860 100102
rect 196916 100046 196984 100102
rect 197040 100046 229878 100102
rect 229934 100046 230002 100102
rect 230058 100046 260598 100102
rect 260654 100046 260722 100102
rect 260778 100046 291318 100102
rect 291374 100046 291442 100102
rect 291498 100046 322038 100102
rect 322094 100046 322162 100102
rect 322218 100046 352758 100102
rect 352814 100046 352882 100102
rect 352938 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 399878 100102
rect 399934 100046 400002 100102
rect 400058 100046 430598 100102
rect 430654 100046 430722 100102
rect 430778 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 470034 100102
rect 470090 100046 470158 100102
rect 470214 100046 470282 100102
rect 470338 100046 470406 100102
rect 470462 100046 500754 100102
rect 500810 100046 500878 100102
rect 500934 100046 501002 100102
rect 501058 100046 501126 100102
rect 501182 100046 531474 100102
rect 531530 100046 531598 100102
rect 531654 100046 531722 100102
rect 531778 100046 531846 100102
rect 531902 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 11930 99978
rect 11986 99922 12054 99978
rect 12110 99922 12178 99978
rect 12234 99922 12302 99978
rect 12358 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 70674 99978
rect 70730 99922 70798 99978
rect 70854 99922 70922 99978
rect 70978 99922 71046 99978
rect 71102 99922 96612 99978
rect 96668 99922 96736 99978
rect 96792 99922 96860 99978
rect 96916 99922 96984 99978
rect 97040 99922 101394 99978
rect 101450 99922 101518 99978
rect 101574 99922 101642 99978
rect 101698 99922 101766 99978
rect 101822 99922 111930 99978
rect 111986 99922 112054 99978
rect 112110 99922 112178 99978
rect 112234 99922 112302 99978
rect 112358 99922 132114 99978
rect 132170 99922 132238 99978
rect 132294 99922 132362 99978
rect 132418 99922 132486 99978
rect 132542 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99922 193554 99978
rect 193610 99922 193678 99978
rect 193734 99922 193802 99978
rect 193858 99922 193926 99978
rect 193982 99922 196612 99978
rect 196668 99922 196736 99978
rect 196792 99922 196860 99978
rect 196916 99922 196984 99978
rect 197040 99922 229878 99978
rect 229934 99922 230002 99978
rect 230058 99922 260598 99978
rect 260654 99922 260722 99978
rect 260778 99922 291318 99978
rect 291374 99922 291442 99978
rect 291498 99922 322038 99978
rect 322094 99922 322162 99978
rect 322218 99922 352758 99978
rect 352814 99922 352882 99978
rect 352938 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 399878 99978
rect 399934 99922 400002 99978
rect 400058 99922 430598 99978
rect 430654 99922 430722 99978
rect 430778 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 470034 99978
rect 470090 99922 470158 99978
rect 470214 99922 470282 99978
rect 470338 99922 470406 99978
rect 470462 99922 500754 99978
rect 500810 99922 500878 99978
rect 500934 99922 501002 99978
rect 501058 99922 501126 99978
rect 501182 99922 531474 99978
rect 531530 99922 531598 99978
rect 531654 99922 531722 99978
rect 531778 99922 531846 99978
rect 531902 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 11130 94350
rect 11186 94294 11254 94350
rect 11310 94294 11378 94350
rect 11434 94294 11502 94350
rect 11558 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 66954 94350
rect 67010 94294 67078 94350
rect 67134 94294 67202 94350
rect 67258 94294 67326 94350
rect 67382 94294 95812 94350
rect 95868 94294 95936 94350
rect 95992 94294 96060 94350
rect 96116 94294 96184 94350
rect 96240 94294 97674 94350
rect 97730 94294 97798 94350
rect 97854 94294 97922 94350
rect 97978 94294 98046 94350
rect 98102 94294 111130 94350
rect 111186 94294 111254 94350
rect 111310 94294 111378 94350
rect 111434 94294 111502 94350
rect 111558 94294 128394 94350
rect 128450 94294 128518 94350
rect 128574 94294 128642 94350
rect 128698 94294 128766 94350
rect 128822 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 195812 94350
rect 195868 94294 195936 94350
rect 195992 94294 196060 94350
rect 196116 94294 196184 94350
rect 196240 94294 214518 94350
rect 214574 94294 214642 94350
rect 214698 94294 245238 94350
rect 245294 94294 245362 94350
rect 245418 94294 275958 94350
rect 276014 94294 276082 94350
rect 276138 94294 306678 94350
rect 306734 94294 306802 94350
rect 306858 94294 337398 94350
rect 337454 94294 337522 94350
rect 337578 94294 368118 94350
rect 368174 94294 368242 94350
rect 368298 94294 374154 94350
rect 374210 94294 374278 94350
rect 374334 94294 374402 94350
rect 374458 94294 374526 94350
rect 374582 94294 384518 94350
rect 384574 94294 384642 94350
rect 384698 94294 415238 94350
rect 415294 94294 415362 94350
rect 415418 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 466314 94350
rect 466370 94294 466438 94350
rect 466494 94294 466562 94350
rect 466618 94294 466686 94350
rect 466742 94294 497034 94350
rect 497090 94294 497158 94350
rect 497214 94294 497282 94350
rect 497338 94294 497406 94350
rect 497462 94294 527754 94350
rect 527810 94294 527878 94350
rect 527934 94294 528002 94350
rect 528058 94294 528126 94350
rect 528182 94294 558474 94350
rect 558530 94294 558598 94350
rect 558654 94294 558722 94350
rect 558778 94294 558846 94350
rect 558902 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 11130 94226
rect 11186 94170 11254 94226
rect 11310 94170 11378 94226
rect 11434 94170 11502 94226
rect 11558 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 66954 94226
rect 67010 94170 67078 94226
rect 67134 94170 67202 94226
rect 67258 94170 67326 94226
rect 67382 94170 95812 94226
rect 95868 94170 95936 94226
rect 95992 94170 96060 94226
rect 96116 94170 96184 94226
rect 96240 94170 97674 94226
rect 97730 94170 97798 94226
rect 97854 94170 97922 94226
rect 97978 94170 98046 94226
rect 98102 94170 111130 94226
rect 111186 94170 111254 94226
rect 111310 94170 111378 94226
rect 111434 94170 111502 94226
rect 111558 94170 128394 94226
rect 128450 94170 128518 94226
rect 128574 94170 128642 94226
rect 128698 94170 128766 94226
rect 128822 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 195812 94226
rect 195868 94170 195936 94226
rect 195992 94170 196060 94226
rect 196116 94170 196184 94226
rect 196240 94170 214518 94226
rect 214574 94170 214642 94226
rect 214698 94170 245238 94226
rect 245294 94170 245362 94226
rect 245418 94170 275958 94226
rect 276014 94170 276082 94226
rect 276138 94170 306678 94226
rect 306734 94170 306802 94226
rect 306858 94170 337398 94226
rect 337454 94170 337522 94226
rect 337578 94170 368118 94226
rect 368174 94170 368242 94226
rect 368298 94170 374154 94226
rect 374210 94170 374278 94226
rect 374334 94170 374402 94226
rect 374458 94170 374526 94226
rect 374582 94170 384518 94226
rect 384574 94170 384642 94226
rect 384698 94170 415238 94226
rect 415294 94170 415362 94226
rect 415418 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 466314 94226
rect 466370 94170 466438 94226
rect 466494 94170 466562 94226
rect 466618 94170 466686 94226
rect 466742 94170 497034 94226
rect 497090 94170 497158 94226
rect 497214 94170 497282 94226
rect 497338 94170 497406 94226
rect 497462 94170 527754 94226
rect 527810 94170 527878 94226
rect 527934 94170 528002 94226
rect 528058 94170 528126 94226
rect 528182 94170 558474 94226
rect 558530 94170 558598 94226
rect 558654 94170 558722 94226
rect 558778 94170 558846 94226
rect 558902 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 11130 94102
rect 11186 94046 11254 94102
rect 11310 94046 11378 94102
rect 11434 94046 11502 94102
rect 11558 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 66954 94102
rect 67010 94046 67078 94102
rect 67134 94046 67202 94102
rect 67258 94046 67326 94102
rect 67382 94046 95812 94102
rect 95868 94046 95936 94102
rect 95992 94046 96060 94102
rect 96116 94046 96184 94102
rect 96240 94046 97674 94102
rect 97730 94046 97798 94102
rect 97854 94046 97922 94102
rect 97978 94046 98046 94102
rect 98102 94046 111130 94102
rect 111186 94046 111254 94102
rect 111310 94046 111378 94102
rect 111434 94046 111502 94102
rect 111558 94046 128394 94102
rect 128450 94046 128518 94102
rect 128574 94046 128642 94102
rect 128698 94046 128766 94102
rect 128822 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 195812 94102
rect 195868 94046 195936 94102
rect 195992 94046 196060 94102
rect 196116 94046 196184 94102
rect 196240 94046 214518 94102
rect 214574 94046 214642 94102
rect 214698 94046 245238 94102
rect 245294 94046 245362 94102
rect 245418 94046 275958 94102
rect 276014 94046 276082 94102
rect 276138 94046 306678 94102
rect 306734 94046 306802 94102
rect 306858 94046 337398 94102
rect 337454 94046 337522 94102
rect 337578 94046 368118 94102
rect 368174 94046 368242 94102
rect 368298 94046 374154 94102
rect 374210 94046 374278 94102
rect 374334 94046 374402 94102
rect 374458 94046 374526 94102
rect 374582 94046 384518 94102
rect 384574 94046 384642 94102
rect 384698 94046 415238 94102
rect 415294 94046 415362 94102
rect 415418 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 466314 94102
rect 466370 94046 466438 94102
rect 466494 94046 466562 94102
rect 466618 94046 466686 94102
rect 466742 94046 497034 94102
rect 497090 94046 497158 94102
rect 497214 94046 497282 94102
rect 497338 94046 497406 94102
rect 497462 94046 527754 94102
rect 527810 94046 527878 94102
rect 527934 94046 528002 94102
rect 528058 94046 528126 94102
rect 528182 94046 558474 94102
rect 558530 94046 558598 94102
rect 558654 94046 558722 94102
rect 558778 94046 558846 94102
rect 558902 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 11130 93978
rect 11186 93922 11254 93978
rect 11310 93922 11378 93978
rect 11434 93922 11502 93978
rect 11558 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 66954 93978
rect 67010 93922 67078 93978
rect 67134 93922 67202 93978
rect 67258 93922 67326 93978
rect 67382 93922 95812 93978
rect 95868 93922 95936 93978
rect 95992 93922 96060 93978
rect 96116 93922 96184 93978
rect 96240 93922 97674 93978
rect 97730 93922 97798 93978
rect 97854 93922 97922 93978
rect 97978 93922 98046 93978
rect 98102 93922 111130 93978
rect 111186 93922 111254 93978
rect 111310 93922 111378 93978
rect 111434 93922 111502 93978
rect 111558 93922 128394 93978
rect 128450 93922 128518 93978
rect 128574 93922 128642 93978
rect 128698 93922 128766 93978
rect 128822 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 195812 93978
rect 195868 93922 195936 93978
rect 195992 93922 196060 93978
rect 196116 93922 196184 93978
rect 196240 93922 214518 93978
rect 214574 93922 214642 93978
rect 214698 93922 245238 93978
rect 245294 93922 245362 93978
rect 245418 93922 275958 93978
rect 276014 93922 276082 93978
rect 276138 93922 306678 93978
rect 306734 93922 306802 93978
rect 306858 93922 337398 93978
rect 337454 93922 337522 93978
rect 337578 93922 368118 93978
rect 368174 93922 368242 93978
rect 368298 93922 374154 93978
rect 374210 93922 374278 93978
rect 374334 93922 374402 93978
rect 374458 93922 374526 93978
rect 374582 93922 384518 93978
rect 384574 93922 384642 93978
rect 384698 93922 415238 93978
rect 415294 93922 415362 93978
rect 415418 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 466314 93978
rect 466370 93922 466438 93978
rect 466494 93922 466562 93978
rect 466618 93922 466686 93978
rect 466742 93922 497034 93978
rect 497090 93922 497158 93978
rect 497214 93922 497282 93978
rect 497338 93922 497406 93978
rect 497462 93922 527754 93978
rect 527810 93922 527878 93978
rect 527934 93922 528002 93978
rect 528058 93922 528126 93978
rect 528182 93922 558474 93978
rect 558530 93922 558598 93978
rect 558654 93922 558722 93978
rect 558778 93922 558846 93978
rect 558902 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect 376108 91558 394228 91574
rect 376108 91502 376124 91558
rect 376180 91502 394156 91558
rect 394212 91502 394228 91558
rect 376108 91486 394228 91502
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 11930 82350
rect 11986 82294 12054 82350
rect 12110 82294 12178 82350
rect 12234 82294 12302 82350
rect 12358 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 70674 82350
rect 70730 82294 70798 82350
rect 70854 82294 70922 82350
rect 70978 82294 71046 82350
rect 71102 82294 96612 82350
rect 96668 82294 96736 82350
rect 96792 82294 96860 82350
rect 96916 82294 96984 82350
rect 97040 82294 101394 82350
rect 101450 82294 101518 82350
rect 101574 82294 101642 82350
rect 101698 82294 101766 82350
rect 101822 82294 111930 82350
rect 111986 82294 112054 82350
rect 112110 82294 112178 82350
rect 112234 82294 112302 82350
rect 112358 82294 132114 82350
rect 132170 82294 132238 82350
rect 132294 82294 132362 82350
rect 132418 82294 132486 82350
rect 132542 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 193554 82350
rect 193610 82294 193678 82350
rect 193734 82294 193802 82350
rect 193858 82294 193926 82350
rect 193982 82294 196612 82350
rect 196668 82294 196736 82350
rect 196792 82294 196860 82350
rect 196916 82294 196984 82350
rect 197040 82294 229878 82350
rect 229934 82294 230002 82350
rect 230058 82294 260598 82350
rect 260654 82294 260722 82350
rect 260778 82294 291318 82350
rect 291374 82294 291442 82350
rect 291498 82294 322038 82350
rect 322094 82294 322162 82350
rect 322218 82294 352758 82350
rect 352814 82294 352882 82350
rect 352938 82294 377874 82350
rect 377930 82294 377998 82350
rect 378054 82294 378122 82350
rect 378178 82294 378246 82350
rect 378302 82294 399878 82350
rect 399934 82294 400002 82350
rect 400058 82294 430598 82350
rect 430654 82294 430722 82350
rect 430778 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 470034 82350
rect 470090 82294 470158 82350
rect 470214 82294 470282 82350
rect 470338 82294 470406 82350
rect 470462 82294 479878 82350
rect 479934 82294 480002 82350
rect 480058 82294 500754 82350
rect 500810 82294 500878 82350
rect 500934 82294 501002 82350
rect 501058 82294 501126 82350
rect 501182 82294 531474 82350
rect 531530 82294 531598 82350
rect 531654 82294 531722 82350
rect 531778 82294 531846 82350
rect 531902 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 11930 82226
rect 11986 82170 12054 82226
rect 12110 82170 12178 82226
rect 12234 82170 12302 82226
rect 12358 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 70674 82226
rect 70730 82170 70798 82226
rect 70854 82170 70922 82226
rect 70978 82170 71046 82226
rect 71102 82170 96612 82226
rect 96668 82170 96736 82226
rect 96792 82170 96860 82226
rect 96916 82170 96984 82226
rect 97040 82170 101394 82226
rect 101450 82170 101518 82226
rect 101574 82170 101642 82226
rect 101698 82170 101766 82226
rect 101822 82170 111930 82226
rect 111986 82170 112054 82226
rect 112110 82170 112178 82226
rect 112234 82170 112302 82226
rect 112358 82170 132114 82226
rect 132170 82170 132238 82226
rect 132294 82170 132362 82226
rect 132418 82170 132486 82226
rect 132542 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 193554 82226
rect 193610 82170 193678 82226
rect 193734 82170 193802 82226
rect 193858 82170 193926 82226
rect 193982 82170 196612 82226
rect 196668 82170 196736 82226
rect 196792 82170 196860 82226
rect 196916 82170 196984 82226
rect 197040 82170 229878 82226
rect 229934 82170 230002 82226
rect 230058 82170 260598 82226
rect 260654 82170 260722 82226
rect 260778 82170 291318 82226
rect 291374 82170 291442 82226
rect 291498 82170 322038 82226
rect 322094 82170 322162 82226
rect 322218 82170 352758 82226
rect 352814 82170 352882 82226
rect 352938 82170 377874 82226
rect 377930 82170 377998 82226
rect 378054 82170 378122 82226
rect 378178 82170 378246 82226
rect 378302 82170 399878 82226
rect 399934 82170 400002 82226
rect 400058 82170 430598 82226
rect 430654 82170 430722 82226
rect 430778 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 470034 82226
rect 470090 82170 470158 82226
rect 470214 82170 470282 82226
rect 470338 82170 470406 82226
rect 470462 82170 479878 82226
rect 479934 82170 480002 82226
rect 480058 82170 500754 82226
rect 500810 82170 500878 82226
rect 500934 82170 501002 82226
rect 501058 82170 501126 82226
rect 501182 82170 531474 82226
rect 531530 82170 531598 82226
rect 531654 82170 531722 82226
rect 531778 82170 531846 82226
rect 531902 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 11930 82102
rect 11986 82046 12054 82102
rect 12110 82046 12178 82102
rect 12234 82046 12302 82102
rect 12358 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 70674 82102
rect 70730 82046 70798 82102
rect 70854 82046 70922 82102
rect 70978 82046 71046 82102
rect 71102 82046 96612 82102
rect 96668 82046 96736 82102
rect 96792 82046 96860 82102
rect 96916 82046 96984 82102
rect 97040 82046 101394 82102
rect 101450 82046 101518 82102
rect 101574 82046 101642 82102
rect 101698 82046 101766 82102
rect 101822 82046 111930 82102
rect 111986 82046 112054 82102
rect 112110 82046 112178 82102
rect 112234 82046 112302 82102
rect 112358 82046 132114 82102
rect 132170 82046 132238 82102
rect 132294 82046 132362 82102
rect 132418 82046 132486 82102
rect 132542 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 193554 82102
rect 193610 82046 193678 82102
rect 193734 82046 193802 82102
rect 193858 82046 193926 82102
rect 193982 82046 196612 82102
rect 196668 82046 196736 82102
rect 196792 82046 196860 82102
rect 196916 82046 196984 82102
rect 197040 82046 229878 82102
rect 229934 82046 230002 82102
rect 230058 82046 260598 82102
rect 260654 82046 260722 82102
rect 260778 82046 291318 82102
rect 291374 82046 291442 82102
rect 291498 82046 322038 82102
rect 322094 82046 322162 82102
rect 322218 82046 352758 82102
rect 352814 82046 352882 82102
rect 352938 82046 377874 82102
rect 377930 82046 377998 82102
rect 378054 82046 378122 82102
rect 378178 82046 378246 82102
rect 378302 82046 399878 82102
rect 399934 82046 400002 82102
rect 400058 82046 430598 82102
rect 430654 82046 430722 82102
rect 430778 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 470034 82102
rect 470090 82046 470158 82102
rect 470214 82046 470282 82102
rect 470338 82046 470406 82102
rect 470462 82046 479878 82102
rect 479934 82046 480002 82102
rect 480058 82046 500754 82102
rect 500810 82046 500878 82102
rect 500934 82046 501002 82102
rect 501058 82046 501126 82102
rect 501182 82046 531474 82102
rect 531530 82046 531598 82102
rect 531654 82046 531722 82102
rect 531778 82046 531846 82102
rect 531902 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 11930 81978
rect 11986 81922 12054 81978
rect 12110 81922 12178 81978
rect 12234 81922 12302 81978
rect 12358 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 70674 81978
rect 70730 81922 70798 81978
rect 70854 81922 70922 81978
rect 70978 81922 71046 81978
rect 71102 81922 96612 81978
rect 96668 81922 96736 81978
rect 96792 81922 96860 81978
rect 96916 81922 96984 81978
rect 97040 81922 101394 81978
rect 101450 81922 101518 81978
rect 101574 81922 101642 81978
rect 101698 81922 101766 81978
rect 101822 81922 111930 81978
rect 111986 81922 112054 81978
rect 112110 81922 112178 81978
rect 112234 81922 112302 81978
rect 112358 81922 132114 81978
rect 132170 81922 132238 81978
rect 132294 81922 132362 81978
rect 132418 81922 132486 81978
rect 132542 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 193554 81978
rect 193610 81922 193678 81978
rect 193734 81922 193802 81978
rect 193858 81922 193926 81978
rect 193982 81922 196612 81978
rect 196668 81922 196736 81978
rect 196792 81922 196860 81978
rect 196916 81922 196984 81978
rect 197040 81922 229878 81978
rect 229934 81922 230002 81978
rect 230058 81922 260598 81978
rect 260654 81922 260722 81978
rect 260778 81922 291318 81978
rect 291374 81922 291442 81978
rect 291498 81922 322038 81978
rect 322094 81922 322162 81978
rect 322218 81922 352758 81978
rect 352814 81922 352882 81978
rect 352938 81922 377874 81978
rect 377930 81922 377998 81978
rect 378054 81922 378122 81978
rect 378178 81922 378246 81978
rect 378302 81922 399878 81978
rect 399934 81922 400002 81978
rect 400058 81922 430598 81978
rect 430654 81922 430722 81978
rect 430778 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 470034 81978
rect 470090 81922 470158 81978
rect 470214 81922 470282 81978
rect 470338 81922 470406 81978
rect 470462 81922 479878 81978
rect 479934 81922 480002 81978
rect 480058 81922 500754 81978
rect 500810 81922 500878 81978
rect 500934 81922 501002 81978
rect 501058 81922 501126 81978
rect 501182 81922 531474 81978
rect 531530 81922 531598 81978
rect 531654 81922 531722 81978
rect 531778 81922 531846 81978
rect 531902 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect 378796 81658 386612 81674
rect 378796 81602 378812 81658
rect 378868 81602 386540 81658
rect 386596 81602 386612 81658
rect 378796 81586 386612 81602
rect 378796 80758 386500 80774
rect 378796 80702 378812 80758
rect 378868 80702 386428 80758
rect 386484 80702 386500 80758
rect 378796 80686 386500 80702
rect 378796 80578 389972 80594
rect 378796 80522 378812 80578
rect 378868 80522 385644 80578
rect 385700 80522 389900 80578
rect 389956 80522 389972 80578
rect 378796 80506 389972 80522
rect 378796 78418 385044 78434
rect 378796 78362 378812 78418
rect 378868 78362 384972 78418
rect 385028 78362 385044 78418
rect 378796 78346 385044 78362
rect 378796 78058 390084 78074
rect 378796 78002 378812 78058
rect 378868 78002 385644 78058
rect 385700 78002 390012 78058
rect 390068 78002 390084 78058
rect 378796 77986 390084 78002
rect 379580 76618 383140 76634
rect 379580 76562 379596 76618
rect 379652 76562 383068 76618
rect 383124 76562 383140 76618
rect 379580 76546 383140 76562
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 11130 76350
rect 11186 76294 11254 76350
rect 11310 76294 11378 76350
rect 11434 76294 11502 76350
rect 11558 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 66954 76350
rect 67010 76294 67078 76350
rect 67134 76294 67202 76350
rect 67258 76294 67326 76350
rect 67382 76294 95812 76350
rect 95868 76294 95936 76350
rect 95992 76294 96060 76350
rect 96116 76294 96184 76350
rect 96240 76294 97674 76350
rect 97730 76294 97798 76350
rect 97854 76294 97922 76350
rect 97978 76294 98046 76350
rect 98102 76294 111130 76350
rect 111186 76294 111254 76350
rect 111310 76294 111378 76350
rect 111434 76294 111502 76350
rect 111558 76294 128394 76350
rect 128450 76294 128518 76350
rect 128574 76294 128642 76350
rect 128698 76294 128766 76350
rect 128822 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 195812 76350
rect 195868 76294 195936 76350
rect 195992 76294 196060 76350
rect 196116 76294 196184 76350
rect 196240 76294 214518 76350
rect 214574 76294 214642 76350
rect 214698 76294 245238 76350
rect 245294 76294 245362 76350
rect 245418 76294 275958 76350
rect 276014 76294 276082 76350
rect 276138 76294 306678 76350
rect 306734 76294 306802 76350
rect 306858 76294 337398 76350
rect 337454 76294 337522 76350
rect 337578 76294 368118 76350
rect 368174 76294 368242 76350
rect 368298 76294 374154 76350
rect 374210 76294 374278 76350
rect 374334 76294 374402 76350
rect 374458 76294 374526 76350
rect 374582 76294 384518 76350
rect 384574 76294 384642 76350
rect 384698 76294 415238 76350
rect 415294 76294 415362 76350
rect 415418 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 464518 76350
rect 464574 76294 464642 76350
rect 464698 76294 466314 76350
rect 466370 76294 466438 76350
rect 466494 76294 466562 76350
rect 466618 76294 466686 76350
rect 466742 76294 495238 76350
rect 495294 76294 495362 76350
rect 495418 76294 497034 76350
rect 497090 76294 497158 76350
rect 497214 76294 497282 76350
rect 497338 76294 497406 76350
rect 497462 76294 527754 76350
rect 527810 76294 527878 76350
rect 527934 76294 528002 76350
rect 528058 76294 528126 76350
rect 528182 76294 558474 76350
rect 558530 76294 558598 76350
rect 558654 76294 558722 76350
rect 558778 76294 558846 76350
rect 558902 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 11130 76226
rect 11186 76170 11254 76226
rect 11310 76170 11378 76226
rect 11434 76170 11502 76226
rect 11558 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 66954 76226
rect 67010 76170 67078 76226
rect 67134 76170 67202 76226
rect 67258 76170 67326 76226
rect 67382 76170 95812 76226
rect 95868 76170 95936 76226
rect 95992 76170 96060 76226
rect 96116 76170 96184 76226
rect 96240 76170 97674 76226
rect 97730 76170 97798 76226
rect 97854 76170 97922 76226
rect 97978 76170 98046 76226
rect 98102 76170 111130 76226
rect 111186 76170 111254 76226
rect 111310 76170 111378 76226
rect 111434 76170 111502 76226
rect 111558 76170 128394 76226
rect 128450 76170 128518 76226
rect 128574 76170 128642 76226
rect 128698 76170 128766 76226
rect 128822 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 195812 76226
rect 195868 76170 195936 76226
rect 195992 76170 196060 76226
rect 196116 76170 196184 76226
rect 196240 76170 214518 76226
rect 214574 76170 214642 76226
rect 214698 76170 245238 76226
rect 245294 76170 245362 76226
rect 245418 76170 275958 76226
rect 276014 76170 276082 76226
rect 276138 76170 306678 76226
rect 306734 76170 306802 76226
rect 306858 76170 337398 76226
rect 337454 76170 337522 76226
rect 337578 76170 368118 76226
rect 368174 76170 368242 76226
rect 368298 76170 374154 76226
rect 374210 76170 374278 76226
rect 374334 76170 374402 76226
rect 374458 76170 374526 76226
rect 374582 76170 384518 76226
rect 384574 76170 384642 76226
rect 384698 76170 415238 76226
rect 415294 76170 415362 76226
rect 415418 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 464518 76226
rect 464574 76170 464642 76226
rect 464698 76170 466314 76226
rect 466370 76170 466438 76226
rect 466494 76170 466562 76226
rect 466618 76170 466686 76226
rect 466742 76170 495238 76226
rect 495294 76170 495362 76226
rect 495418 76170 497034 76226
rect 497090 76170 497158 76226
rect 497214 76170 497282 76226
rect 497338 76170 497406 76226
rect 497462 76170 527754 76226
rect 527810 76170 527878 76226
rect 527934 76170 528002 76226
rect 528058 76170 528126 76226
rect 528182 76170 558474 76226
rect 558530 76170 558598 76226
rect 558654 76170 558722 76226
rect 558778 76170 558846 76226
rect 558902 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 11130 76102
rect 11186 76046 11254 76102
rect 11310 76046 11378 76102
rect 11434 76046 11502 76102
rect 11558 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 66954 76102
rect 67010 76046 67078 76102
rect 67134 76046 67202 76102
rect 67258 76046 67326 76102
rect 67382 76046 95812 76102
rect 95868 76046 95936 76102
rect 95992 76046 96060 76102
rect 96116 76046 96184 76102
rect 96240 76046 97674 76102
rect 97730 76046 97798 76102
rect 97854 76046 97922 76102
rect 97978 76046 98046 76102
rect 98102 76046 111130 76102
rect 111186 76046 111254 76102
rect 111310 76046 111378 76102
rect 111434 76046 111502 76102
rect 111558 76046 128394 76102
rect 128450 76046 128518 76102
rect 128574 76046 128642 76102
rect 128698 76046 128766 76102
rect 128822 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 195812 76102
rect 195868 76046 195936 76102
rect 195992 76046 196060 76102
rect 196116 76046 196184 76102
rect 196240 76046 214518 76102
rect 214574 76046 214642 76102
rect 214698 76046 245238 76102
rect 245294 76046 245362 76102
rect 245418 76046 275958 76102
rect 276014 76046 276082 76102
rect 276138 76046 306678 76102
rect 306734 76046 306802 76102
rect 306858 76046 337398 76102
rect 337454 76046 337522 76102
rect 337578 76046 368118 76102
rect 368174 76046 368242 76102
rect 368298 76046 374154 76102
rect 374210 76046 374278 76102
rect 374334 76046 374402 76102
rect 374458 76046 374526 76102
rect 374582 76046 384518 76102
rect 384574 76046 384642 76102
rect 384698 76046 415238 76102
rect 415294 76046 415362 76102
rect 415418 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 464518 76102
rect 464574 76046 464642 76102
rect 464698 76046 466314 76102
rect 466370 76046 466438 76102
rect 466494 76046 466562 76102
rect 466618 76046 466686 76102
rect 466742 76046 495238 76102
rect 495294 76046 495362 76102
rect 495418 76046 497034 76102
rect 497090 76046 497158 76102
rect 497214 76046 497282 76102
rect 497338 76046 497406 76102
rect 497462 76046 527754 76102
rect 527810 76046 527878 76102
rect 527934 76046 528002 76102
rect 528058 76046 528126 76102
rect 528182 76046 558474 76102
rect 558530 76046 558598 76102
rect 558654 76046 558722 76102
rect 558778 76046 558846 76102
rect 558902 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 11130 75978
rect 11186 75922 11254 75978
rect 11310 75922 11378 75978
rect 11434 75922 11502 75978
rect 11558 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 66954 75978
rect 67010 75922 67078 75978
rect 67134 75922 67202 75978
rect 67258 75922 67326 75978
rect 67382 75922 95812 75978
rect 95868 75922 95936 75978
rect 95992 75922 96060 75978
rect 96116 75922 96184 75978
rect 96240 75922 97674 75978
rect 97730 75922 97798 75978
rect 97854 75922 97922 75978
rect 97978 75922 98046 75978
rect 98102 75922 111130 75978
rect 111186 75922 111254 75978
rect 111310 75922 111378 75978
rect 111434 75922 111502 75978
rect 111558 75922 128394 75978
rect 128450 75922 128518 75978
rect 128574 75922 128642 75978
rect 128698 75922 128766 75978
rect 128822 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 195812 75978
rect 195868 75922 195936 75978
rect 195992 75922 196060 75978
rect 196116 75922 196184 75978
rect 196240 75922 214518 75978
rect 214574 75922 214642 75978
rect 214698 75922 245238 75978
rect 245294 75922 245362 75978
rect 245418 75922 275958 75978
rect 276014 75922 276082 75978
rect 276138 75922 306678 75978
rect 306734 75922 306802 75978
rect 306858 75922 337398 75978
rect 337454 75922 337522 75978
rect 337578 75922 368118 75978
rect 368174 75922 368242 75978
rect 368298 75922 374154 75978
rect 374210 75922 374278 75978
rect 374334 75922 374402 75978
rect 374458 75922 374526 75978
rect 374582 75922 384518 75978
rect 384574 75922 384642 75978
rect 384698 75922 415238 75978
rect 415294 75922 415362 75978
rect 415418 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 464518 75978
rect 464574 75922 464642 75978
rect 464698 75922 466314 75978
rect 466370 75922 466438 75978
rect 466494 75922 466562 75978
rect 466618 75922 466686 75978
rect 466742 75922 495238 75978
rect 495294 75922 495362 75978
rect 495418 75922 497034 75978
rect 497090 75922 497158 75978
rect 497214 75922 497282 75978
rect 497338 75922 497406 75978
rect 497462 75922 527754 75978
rect 527810 75922 527878 75978
rect 527934 75922 528002 75978
rect 528058 75922 528126 75978
rect 528182 75922 558474 75978
rect 558530 75922 558598 75978
rect 558654 75922 558722 75978
rect 558778 75922 558846 75978
rect 558902 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect 378572 74278 381572 74294
rect 378572 74222 378588 74278
rect 378644 74222 381500 74278
rect 381556 74222 381572 74278
rect 378572 74206 381572 74222
rect 379580 74098 393220 74114
rect 379580 74042 379596 74098
rect 379652 74042 383852 74098
rect 383908 74042 393148 74098
rect 393204 74042 393220 74098
rect 379580 74026 393220 74042
rect 378796 72838 381908 72854
rect 378796 72782 378812 72838
rect 378868 72782 381836 72838
rect 381892 72782 381908 72838
rect 378796 72766 381908 72782
rect 379916 72118 381460 72134
rect 379916 72062 379932 72118
rect 379988 72062 381388 72118
rect 381444 72062 381460 72118
rect 379916 72046 381460 72062
rect 377564 71398 388404 71414
rect 377564 71342 377580 71398
rect 377636 71342 381388 71398
rect 381444 71342 388332 71398
rect 388388 71342 388404 71398
rect 377564 71326 388404 71342
rect 377564 64918 388404 64934
rect 377564 64862 377580 64918
rect 377636 64862 388332 64918
rect 388388 64862 388404 64918
rect 377564 64846 388404 64862
rect 377564 64738 388180 64754
rect 377564 64682 377580 64738
rect 377636 64682 388108 64738
rect 388164 64682 388180 64738
rect 377564 64666 388180 64682
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 11930 64350
rect 11986 64294 12054 64350
rect 12110 64294 12178 64350
rect 12234 64294 12302 64350
rect 12358 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 70674 64350
rect 70730 64294 70798 64350
rect 70854 64294 70922 64350
rect 70978 64294 71046 64350
rect 71102 64294 96612 64350
rect 96668 64294 96736 64350
rect 96792 64294 96860 64350
rect 96916 64294 96984 64350
rect 97040 64294 101394 64350
rect 101450 64294 101518 64350
rect 101574 64294 101642 64350
rect 101698 64294 101766 64350
rect 101822 64294 111930 64350
rect 111986 64294 112054 64350
rect 112110 64294 112178 64350
rect 112234 64294 112302 64350
rect 112358 64294 132114 64350
rect 132170 64294 132238 64350
rect 132294 64294 132362 64350
rect 132418 64294 132486 64350
rect 132542 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 193554 64350
rect 193610 64294 193678 64350
rect 193734 64294 193802 64350
rect 193858 64294 193926 64350
rect 193982 64294 196612 64350
rect 196668 64294 196736 64350
rect 196792 64294 196860 64350
rect 196916 64294 196984 64350
rect 197040 64294 229878 64350
rect 229934 64294 230002 64350
rect 230058 64294 260598 64350
rect 260654 64294 260722 64350
rect 260778 64294 291318 64350
rect 291374 64294 291442 64350
rect 291498 64294 322038 64350
rect 322094 64294 322162 64350
rect 322218 64294 352758 64350
rect 352814 64294 352882 64350
rect 352938 64294 377874 64350
rect 377930 64294 377998 64350
rect 378054 64294 378122 64350
rect 378178 64294 378246 64350
rect 378302 64294 399878 64350
rect 399934 64294 400002 64350
rect 400058 64294 430598 64350
rect 430654 64294 430722 64350
rect 430778 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 470034 64350
rect 470090 64294 470158 64350
rect 470214 64294 470282 64350
rect 470338 64294 470406 64350
rect 470462 64294 479878 64350
rect 479934 64294 480002 64350
rect 480058 64294 500754 64350
rect 500810 64294 500878 64350
rect 500934 64294 501002 64350
rect 501058 64294 501126 64350
rect 501182 64294 531474 64350
rect 531530 64294 531598 64350
rect 531654 64294 531722 64350
rect 531778 64294 531846 64350
rect 531902 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 11930 64226
rect 11986 64170 12054 64226
rect 12110 64170 12178 64226
rect 12234 64170 12302 64226
rect 12358 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 70674 64226
rect 70730 64170 70798 64226
rect 70854 64170 70922 64226
rect 70978 64170 71046 64226
rect 71102 64170 96612 64226
rect 96668 64170 96736 64226
rect 96792 64170 96860 64226
rect 96916 64170 96984 64226
rect 97040 64170 101394 64226
rect 101450 64170 101518 64226
rect 101574 64170 101642 64226
rect 101698 64170 101766 64226
rect 101822 64170 111930 64226
rect 111986 64170 112054 64226
rect 112110 64170 112178 64226
rect 112234 64170 112302 64226
rect 112358 64170 132114 64226
rect 132170 64170 132238 64226
rect 132294 64170 132362 64226
rect 132418 64170 132486 64226
rect 132542 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 193554 64226
rect 193610 64170 193678 64226
rect 193734 64170 193802 64226
rect 193858 64170 193926 64226
rect 193982 64170 196612 64226
rect 196668 64170 196736 64226
rect 196792 64170 196860 64226
rect 196916 64170 196984 64226
rect 197040 64170 229878 64226
rect 229934 64170 230002 64226
rect 230058 64170 260598 64226
rect 260654 64170 260722 64226
rect 260778 64170 291318 64226
rect 291374 64170 291442 64226
rect 291498 64170 322038 64226
rect 322094 64170 322162 64226
rect 322218 64170 352758 64226
rect 352814 64170 352882 64226
rect 352938 64170 377874 64226
rect 377930 64170 377998 64226
rect 378054 64170 378122 64226
rect 378178 64170 378246 64226
rect 378302 64170 399878 64226
rect 399934 64170 400002 64226
rect 400058 64170 430598 64226
rect 430654 64170 430722 64226
rect 430778 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 470034 64226
rect 470090 64170 470158 64226
rect 470214 64170 470282 64226
rect 470338 64170 470406 64226
rect 470462 64170 479878 64226
rect 479934 64170 480002 64226
rect 480058 64170 500754 64226
rect 500810 64170 500878 64226
rect 500934 64170 501002 64226
rect 501058 64170 501126 64226
rect 501182 64170 531474 64226
rect 531530 64170 531598 64226
rect 531654 64170 531722 64226
rect 531778 64170 531846 64226
rect 531902 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 11930 64102
rect 11986 64046 12054 64102
rect 12110 64046 12178 64102
rect 12234 64046 12302 64102
rect 12358 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 70674 64102
rect 70730 64046 70798 64102
rect 70854 64046 70922 64102
rect 70978 64046 71046 64102
rect 71102 64046 96612 64102
rect 96668 64046 96736 64102
rect 96792 64046 96860 64102
rect 96916 64046 96984 64102
rect 97040 64046 101394 64102
rect 101450 64046 101518 64102
rect 101574 64046 101642 64102
rect 101698 64046 101766 64102
rect 101822 64046 111930 64102
rect 111986 64046 112054 64102
rect 112110 64046 112178 64102
rect 112234 64046 112302 64102
rect 112358 64046 132114 64102
rect 132170 64046 132238 64102
rect 132294 64046 132362 64102
rect 132418 64046 132486 64102
rect 132542 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 193554 64102
rect 193610 64046 193678 64102
rect 193734 64046 193802 64102
rect 193858 64046 193926 64102
rect 193982 64046 196612 64102
rect 196668 64046 196736 64102
rect 196792 64046 196860 64102
rect 196916 64046 196984 64102
rect 197040 64046 229878 64102
rect 229934 64046 230002 64102
rect 230058 64046 260598 64102
rect 260654 64046 260722 64102
rect 260778 64046 291318 64102
rect 291374 64046 291442 64102
rect 291498 64046 322038 64102
rect 322094 64046 322162 64102
rect 322218 64046 352758 64102
rect 352814 64046 352882 64102
rect 352938 64046 377874 64102
rect 377930 64046 377998 64102
rect 378054 64046 378122 64102
rect 378178 64046 378246 64102
rect 378302 64046 399878 64102
rect 399934 64046 400002 64102
rect 400058 64046 430598 64102
rect 430654 64046 430722 64102
rect 430778 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 470034 64102
rect 470090 64046 470158 64102
rect 470214 64046 470282 64102
rect 470338 64046 470406 64102
rect 470462 64046 479878 64102
rect 479934 64046 480002 64102
rect 480058 64046 500754 64102
rect 500810 64046 500878 64102
rect 500934 64046 501002 64102
rect 501058 64046 501126 64102
rect 501182 64046 531474 64102
rect 531530 64046 531598 64102
rect 531654 64046 531722 64102
rect 531778 64046 531846 64102
rect 531902 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 11930 63978
rect 11986 63922 12054 63978
rect 12110 63922 12178 63978
rect 12234 63922 12302 63978
rect 12358 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 70674 63978
rect 70730 63922 70798 63978
rect 70854 63922 70922 63978
rect 70978 63922 71046 63978
rect 71102 63922 96612 63978
rect 96668 63922 96736 63978
rect 96792 63922 96860 63978
rect 96916 63922 96984 63978
rect 97040 63922 101394 63978
rect 101450 63922 101518 63978
rect 101574 63922 101642 63978
rect 101698 63922 101766 63978
rect 101822 63922 111930 63978
rect 111986 63922 112054 63978
rect 112110 63922 112178 63978
rect 112234 63922 112302 63978
rect 112358 63922 132114 63978
rect 132170 63922 132238 63978
rect 132294 63922 132362 63978
rect 132418 63922 132486 63978
rect 132542 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 193554 63978
rect 193610 63922 193678 63978
rect 193734 63922 193802 63978
rect 193858 63922 193926 63978
rect 193982 63922 196612 63978
rect 196668 63922 196736 63978
rect 196792 63922 196860 63978
rect 196916 63922 196984 63978
rect 197040 63922 229878 63978
rect 229934 63922 230002 63978
rect 230058 63922 260598 63978
rect 260654 63922 260722 63978
rect 260778 63922 291318 63978
rect 291374 63922 291442 63978
rect 291498 63922 322038 63978
rect 322094 63922 322162 63978
rect 322218 63922 352758 63978
rect 352814 63922 352882 63978
rect 352938 63922 377874 63978
rect 377930 63922 377998 63978
rect 378054 63922 378122 63978
rect 378178 63922 378246 63978
rect 378302 63922 399878 63978
rect 399934 63922 400002 63978
rect 400058 63922 430598 63978
rect 430654 63922 430722 63978
rect 430778 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 470034 63978
rect 470090 63922 470158 63978
rect 470214 63922 470282 63978
rect 470338 63922 470406 63978
rect 470462 63922 479878 63978
rect 479934 63922 480002 63978
rect 480058 63922 500754 63978
rect 500810 63922 500878 63978
rect 500934 63922 501002 63978
rect 501058 63922 501126 63978
rect 501182 63922 531474 63978
rect 531530 63922 531598 63978
rect 531654 63922 531722 63978
rect 531778 63922 531846 63978
rect 531902 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect 377564 62938 389860 62954
rect 377564 62882 377580 62938
rect 377636 62882 389788 62938
rect 389844 62882 389860 62938
rect 377564 62866 389860 62882
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 11130 58350
rect 11186 58294 11254 58350
rect 11310 58294 11378 58350
rect 11434 58294 11502 58350
rect 11558 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 66954 58350
rect 67010 58294 67078 58350
rect 67134 58294 67202 58350
rect 67258 58294 67326 58350
rect 67382 58294 95812 58350
rect 95868 58294 95936 58350
rect 95992 58294 96060 58350
rect 96116 58294 96184 58350
rect 96240 58294 97674 58350
rect 97730 58294 97798 58350
rect 97854 58294 97922 58350
rect 97978 58294 98046 58350
rect 98102 58294 111130 58350
rect 111186 58294 111254 58350
rect 111310 58294 111378 58350
rect 111434 58294 111502 58350
rect 111558 58294 128394 58350
rect 128450 58294 128518 58350
rect 128574 58294 128642 58350
rect 128698 58294 128766 58350
rect 128822 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 189834 58350
rect 189890 58294 189958 58350
rect 190014 58294 190082 58350
rect 190138 58294 190206 58350
rect 190262 58294 195812 58350
rect 195868 58294 195936 58350
rect 195992 58294 196060 58350
rect 196116 58294 196184 58350
rect 196240 58294 214518 58350
rect 214574 58294 214642 58350
rect 214698 58294 245238 58350
rect 245294 58294 245362 58350
rect 245418 58294 275958 58350
rect 276014 58294 276082 58350
rect 276138 58294 306678 58350
rect 306734 58294 306802 58350
rect 306858 58294 337398 58350
rect 337454 58294 337522 58350
rect 337578 58294 368118 58350
rect 368174 58294 368242 58350
rect 368298 58294 374154 58350
rect 374210 58294 374278 58350
rect 374334 58294 374402 58350
rect 374458 58294 374526 58350
rect 374582 58294 384518 58350
rect 384574 58294 384642 58350
rect 384698 58294 415238 58350
rect 415294 58294 415362 58350
rect 415418 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 464518 58350
rect 464574 58294 464642 58350
rect 464698 58294 466314 58350
rect 466370 58294 466438 58350
rect 466494 58294 466562 58350
rect 466618 58294 466686 58350
rect 466742 58294 495238 58350
rect 495294 58294 495362 58350
rect 495418 58294 497034 58350
rect 497090 58294 497158 58350
rect 497214 58294 497282 58350
rect 497338 58294 497406 58350
rect 497462 58294 527754 58350
rect 527810 58294 527878 58350
rect 527934 58294 528002 58350
rect 528058 58294 528126 58350
rect 528182 58294 558474 58350
rect 558530 58294 558598 58350
rect 558654 58294 558722 58350
rect 558778 58294 558846 58350
rect 558902 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 11130 58226
rect 11186 58170 11254 58226
rect 11310 58170 11378 58226
rect 11434 58170 11502 58226
rect 11558 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 66954 58226
rect 67010 58170 67078 58226
rect 67134 58170 67202 58226
rect 67258 58170 67326 58226
rect 67382 58170 95812 58226
rect 95868 58170 95936 58226
rect 95992 58170 96060 58226
rect 96116 58170 96184 58226
rect 96240 58170 97674 58226
rect 97730 58170 97798 58226
rect 97854 58170 97922 58226
rect 97978 58170 98046 58226
rect 98102 58170 111130 58226
rect 111186 58170 111254 58226
rect 111310 58170 111378 58226
rect 111434 58170 111502 58226
rect 111558 58170 128394 58226
rect 128450 58170 128518 58226
rect 128574 58170 128642 58226
rect 128698 58170 128766 58226
rect 128822 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 189834 58226
rect 189890 58170 189958 58226
rect 190014 58170 190082 58226
rect 190138 58170 190206 58226
rect 190262 58170 195812 58226
rect 195868 58170 195936 58226
rect 195992 58170 196060 58226
rect 196116 58170 196184 58226
rect 196240 58170 214518 58226
rect 214574 58170 214642 58226
rect 214698 58170 245238 58226
rect 245294 58170 245362 58226
rect 245418 58170 275958 58226
rect 276014 58170 276082 58226
rect 276138 58170 306678 58226
rect 306734 58170 306802 58226
rect 306858 58170 337398 58226
rect 337454 58170 337522 58226
rect 337578 58170 368118 58226
rect 368174 58170 368242 58226
rect 368298 58170 374154 58226
rect 374210 58170 374278 58226
rect 374334 58170 374402 58226
rect 374458 58170 374526 58226
rect 374582 58170 384518 58226
rect 384574 58170 384642 58226
rect 384698 58170 415238 58226
rect 415294 58170 415362 58226
rect 415418 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 464518 58226
rect 464574 58170 464642 58226
rect 464698 58170 466314 58226
rect 466370 58170 466438 58226
rect 466494 58170 466562 58226
rect 466618 58170 466686 58226
rect 466742 58170 495238 58226
rect 495294 58170 495362 58226
rect 495418 58170 497034 58226
rect 497090 58170 497158 58226
rect 497214 58170 497282 58226
rect 497338 58170 497406 58226
rect 497462 58170 527754 58226
rect 527810 58170 527878 58226
rect 527934 58170 528002 58226
rect 528058 58170 528126 58226
rect 528182 58170 558474 58226
rect 558530 58170 558598 58226
rect 558654 58170 558722 58226
rect 558778 58170 558846 58226
rect 558902 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 11130 58102
rect 11186 58046 11254 58102
rect 11310 58046 11378 58102
rect 11434 58046 11502 58102
rect 11558 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 66954 58102
rect 67010 58046 67078 58102
rect 67134 58046 67202 58102
rect 67258 58046 67326 58102
rect 67382 58046 95812 58102
rect 95868 58046 95936 58102
rect 95992 58046 96060 58102
rect 96116 58046 96184 58102
rect 96240 58046 97674 58102
rect 97730 58046 97798 58102
rect 97854 58046 97922 58102
rect 97978 58046 98046 58102
rect 98102 58046 111130 58102
rect 111186 58046 111254 58102
rect 111310 58046 111378 58102
rect 111434 58046 111502 58102
rect 111558 58046 128394 58102
rect 128450 58046 128518 58102
rect 128574 58046 128642 58102
rect 128698 58046 128766 58102
rect 128822 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 189834 58102
rect 189890 58046 189958 58102
rect 190014 58046 190082 58102
rect 190138 58046 190206 58102
rect 190262 58046 195812 58102
rect 195868 58046 195936 58102
rect 195992 58046 196060 58102
rect 196116 58046 196184 58102
rect 196240 58046 214518 58102
rect 214574 58046 214642 58102
rect 214698 58046 245238 58102
rect 245294 58046 245362 58102
rect 245418 58046 275958 58102
rect 276014 58046 276082 58102
rect 276138 58046 306678 58102
rect 306734 58046 306802 58102
rect 306858 58046 337398 58102
rect 337454 58046 337522 58102
rect 337578 58046 368118 58102
rect 368174 58046 368242 58102
rect 368298 58046 374154 58102
rect 374210 58046 374278 58102
rect 374334 58046 374402 58102
rect 374458 58046 374526 58102
rect 374582 58046 384518 58102
rect 384574 58046 384642 58102
rect 384698 58046 415238 58102
rect 415294 58046 415362 58102
rect 415418 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 464518 58102
rect 464574 58046 464642 58102
rect 464698 58046 466314 58102
rect 466370 58046 466438 58102
rect 466494 58046 466562 58102
rect 466618 58046 466686 58102
rect 466742 58046 495238 58102
rect 495294 58046 495362 58102
rect 495418 58046 497034 58102
rect 497090 58046 497158 58102
rect 497214 58046 497282 58102
rect 497338 58046 497406 58102
rect 497462 58046 527754 58102
rect 527810 58046 527878 58102
rect 527934 58046 528002 58102
rect 528058 58046 528126 58102
rect 528182 58046 558474 58102
rect 558530 58046 558598 58102
rect 558654 58046 558722 58102
rect 558778 58046 558846 58102
rect 558902 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 11130 57978
rect 11186 57922 11254 57978
rect 11310 57922 11378 57978
rect 11434 57922 11502 57978
rect 11558 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 66954 57978
rect 67010 57922 67078 57978
rect 67134 57922 67202 57978
rect 67258 57922 67326 57978
rect 67382 57922 95812 57978
rect 95868 57922 95936 57978
rect 95992 57922 96060 57978
rect 96116 57922 96184 57978
rect 96240 57922 97674 57978
rect 97730 57922 97798 57978
rect 97854 57922 97922 57978
rect 97978 57922 98046 57978
rect 98102 57922 111130 57978
rect 111186 57922 111254 57978
rect 111310 57922 111378 57978
rect 111434 57922 111502 57978
rect 111558 57922 128394 57978
rect 128450 57922 128518 57978
rect 128574 57922 128642 57978
rect 128698 57922 128766 57978
rect 128822 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 189834 57978
rect 189890 57922 189958 57978
rect 190014 57922 190082 57978
rect 190138 57922 190206 57978
rect 190262 57922 195812 57978
rect 195868 57922 195936 57978
rect 195992 57922 196060 57978
rect 196116 57922 196184 57978
rect 196240 57922 214518 57978
rect 214574 57922 214642 57978
rect 214698 57922 245238 57978
rect 245294 57922 245362 57978
rect 245418 57922 275958 57978
rect 276014 57922 276082 57978
rect 276138 57922 306678 57978
rect 306734 57922 306802 57978
rect 306858 57922 337398 57978
rect 337454 57922 337522 57978
rect 337578 57922 368118 57978
rect 368174 57922 368242 57978
rect 368298 57922 374154 57978
rect 374210 57922 374278 57978
rect 374334 57922 374402 57978
rect 374458 57922 374526 57978
rect 374582 57922 384518 57978
rect 384574 57922 384642 57978
rect 384698 57922 415238 57978
rect 415294 57922 415362 57978
rect 415418 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 464518 57978
rect 464574 57922 464642 57978
rect 464698 57922 466314 57978
rect 466370 57922 466438 57978
rect 466494 57922 466562 57978
rect 466618 57922 466686 57978
rect 466742 57922 495238 57978
rect 495294 57922 495362 57978
rect 495418 57922 497034 57978
rect 497090 57922 497158 57978
rect 497214 57922 497282 57978
rect 497338 57922 497406 57978
rect 497462 57922 527754 57978
rect 527810 57922 527878 57978
rect 527934 57922 528002 57978
rect 528058 57922 528126 57978
rect 528182 57922 558474 57978
rect 558530 57922 558598 57978
rect 558654 57922 558722 57978
rect 558778 57922 558846 57978
rect 558902 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect 209900 56998 370484 57014
rect 209900 56942 209916 56998
rect 209972 56942 370412 56998
rect 370468 56942 370484 56998
rect 209900 56926 370484 56942
rect 376220 52138 394900 52154
rect 376220 52082 376236 52138
rect 376292 52082 394828 52138
rect 394884 52082 394900 52138
rect 376220 52066 394900 52082
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46198 439314 46226
rect 378302 46170 408594 46198
rect -1916 46142 408594 46170
rect 408650 46142 408718 46198
rect 408774 46142 408842 46198
rect 408898 46142 408966 46198
rect 409022 46170 439314 46198
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 409022 46142 597980 46170
rect -1916 46102 597980 46142
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46074 439314 46102
rect 378302 46046 408594 46074
rect -1916 46018 408594 46046
rect 408650 46018 408718 46074
rect 408774 46018 408842 46074
rect 408898 46018 408966 46074
rect 409022 46046 439314 46074
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 409022 46018 597980 46046
rect -1916 45978 597980 46018
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45950 439314 45978
rect 378302 45922 408594 45950
rect -1916 45894 408594 45922
rect 408650 45894 408718 45950
rect 408774 45894 408842 45950
rect 408898 45894 408966 45950
rect 409022 45922 439314 45950
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 409022 45894 597980 45922
rect -1916 45826 597980 45894
rect 379692 43678 419764 43694
rect 379692 43622 379708 43678
rect 379764 43622 419692 43678
rect 419748 43622 419764 43678
rect 379692 43606 419764 43622
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 150558 28350
rect 150614 28294 150682 28350
rect 150738 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 279862 28350
rect 279918 28294 279986 28350
rect 280042 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 409166 28350
rect 409222 28294 409290 28350
rect 409346 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 538470 28350
rect 538526 28294 538594 28350
rect 538650 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 150558 28226
rect 150614 28170 150682 28226
rect 150738 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 279862 28226
rect 279918 28170 279986 28226
rect 280042 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 409166 28226
rect 409222 28170 409290 28226
rect 409346 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 538470 28226
rect 538526 28170 538594 28226
rect 538650 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 150558 28102
rect 150614 28046 150682 28102
rect 150738 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 279862 28102
rect 279918 28046 279986 28102
rect 280042 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 409166 28102
rect 409222 28046 409290 28102
rect 409346 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 538470 28102
rect 538526 28046 538594 28102
rect 538650 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 150558 27978
rect 150614 27922 150682 27978
rect 150738 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 279862 27978
rect 279918 27922 279986 27978
rect 280042 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 409166 27978
rect 409222 27922 409290 27978
rect 409346 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 538470 27978
rect 538526 27922 538594 27978
rect 538650 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 85906 22350
rect 85962 22294 86030 22350
rect 86086 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 215210 22350
rect 215266 22294 215334 22350
rect 215390 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 344514 22350
rect 344570 22294 344638 22350
rect 344694 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 473818 22350
rect 473874 22294 473942 22350
rect 473998 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 85906 22226
rect 85962 22170 86030 22226
rect 86086 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 215210 22226
rect 215266 22170 215334 22226
rect 215390 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 344514 22226
rect 344570 22170 344638 22226
rect 344694 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 473818 22226
rect 473874 22170 473942 22226
rect 473998 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 85906 22102
rect 85962 22046 86030 22102
rect 86086 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 215210 22102
rect 215266 22046 215334 22102
rect 215390 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 344514 22102
rect 344570 22046 344638 22102
rect 344694 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 473818 22102
rect 473874 22046 473942 22102
rect 473998 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 85906 21978
rect 85962 21922 86030 21978
rect 86086 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 215210 21978
rect 215266 21922 215334 21978
rect 215390 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 344514 21978
rect 344570 21922 344638 21978
rect 344694 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 473818 21978
rect 473874 21922 473942 21978
rect 473998 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 150558 10350
rect 150614 10294 150682 10350
rect 150738 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 279862 10350
rect 279918 10294 279986 10350
rect 280042 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 409166 10350
rect 409222 10294 409290 10350
rect 409346 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 538470 10350
rect 538526 10294 538594 10350
rect 538650 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 150558 10226
rect 150614 10170 150682 10226
rect 150738 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 279862 10226
rect 279918 10170 279986 10226
rect 280042 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 409166 10226
rect 409222 10170 409290 10226
rect 409346 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 538470 10226
rect 538526 10170 538594 10226
rect 538650 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 150558 10102
rect 150614 10046 150682 10102
rect 150738 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 279862 10102
rect 279918 10046 279986 10102
rect 280042 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 409166 10102
rect 409222 10046 409290 10102
rect 409346 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 538470 10102
rect 538526 10046 538594 10102
rect 538650 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 150558 9978
rect 150614 9922 150682 9978
rect 150738 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 279862 9978
rect 279918 9922 279986 9978
rect 280042 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 409166 9978
rect 409222 9922 409290 9978
rect 409346 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 538470 9978
rect 538526 9922 538594 9978
rect 538650 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect 475452 5338 529300 5354
rect 475452 5282 475468 5338
rect 475524 5282 529228 5338
rect 529284 5282 529300 5338
rect 475452 5266 529300 5282
rect 442972 5158 495028 5174
rect 442972 5102 442988 5158
rect 443044 5102 494956 5158
rect 495012 5102 495028 5158
rect 442972 5086 495028 5102
rect 498972 5158 557860 5174
rect 498972 5102 498988 5158
rect 499044 5102 557788 5158
rect 557844 5102 557860 5158
rect 498972 5086 557860 5102
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect 447676 3358 499060 3374
rect 447676 3302 447692 3358
rect 447748 3302 498988 3358
rect 499044 3302 499060 3358
rect 447676 3286 499060 3302
rect 501660 3358 565476 3374
rect 501660 3302 501676 3358
rect 501732 3302 565404 3358
rect 565460 3302 565476 3358
rect 501660 3286 565476 3302
rect 499420 3178 563572 3194
rect 499420 3122 499436 3178
rect 499492 3122 563500 3178
rect 563556 3122 563572 3178
rect 499420 3106 563572 3122
rect 457084 478 512164 494
rect 457084 422 457100 478
rect 457156 422 512092 478
rect 512148 422 512164 478
rect 457084 406 512164 422
rect 510732 298 571300 314
rect 510732 242 510748 298
rect 510804 242 571228 298
rect 571284 242 571300 298
rect 510732 226 571300 242
rect 504124 118 569284 134
rect 504124 62 504140 118
rect 504196 62 569212 118
rect 569268 62 569284 118
rect 504124 46 569284 62
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use cpu  cpu_inst_0
timestamp 0
transform 1 0 210000 0 1 45000
box 0 2688 160000 280000
use ctrl  ctrl_inst_0
timestamp 0
transform 1 0 460000 0 1 45000
box 0 0 50000 46316
use pcpi_approx_mul  pcpi_approx_mul_inst_0
timestamp 0
transform 1 0 380000 0 1 275000
box 0 0 60000 50000
use pcpi_div  pcpi_div_inst_0
timestamp 0
transform 1 0 380000 0 1 135000
box 0 0 60000 60000
use pcpi_exact_mul  pcpi_exact_mul_inst_0
timestamp 0
transform 1 0 380000 0 1 205000
box 0 0 60000 60000
use pcpi_mul  pcpi_mul_inst_0
timestamp 0
transform 1 0 380000 0 1 45000
box 0 0 60000 76892
use simple_interconnect  simple_interconnect_inst_0
timestamp 0
transform -1 0 200000 0 -1 360000
box 0 0 80000 80000
use simpleuart  simpleuart
timestamp 0
transform 1 0 60000 0 1 280000
box 0 0 50000 50000
use spimemio  spimemio
timestamp 0
transform 1 0 5000 0 1 280000
box 0 0 50000 50000
use gf180_ram_512x8x1  sram512x8_0
timestamp 0
transform 1 0 10000 0 1 45000
box 1000 1000 87372 100000
use gf180_ram_512x8x1  sram512x8_1
timestamp 0
transform 1 0 110000 0 1 45000
box 1000 1000 87372 100000
use gf180_ram_512x8x1  sram512x8_2
timestamp 0
transform -1 0 100000 0 -1 265000
box 1000 1000 87372 100000
use gf180_ram_512x8x1  sram512x8_3
timestamp 0
transform -1 0 200000 0 -1 265000
box 1000 1000 87372 100000
use user_proj_example  user_proj_example_inst_0
timestamp 0
transform 1 0 20000 0 1 5000
box 1258 0 520000 27888
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5418 -1644 6038 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 -1644 36758 281266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 326670 36758 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 -1644 67478 286194 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 330590 67478 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 -1644 98198 166456 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 330590 98198 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 -1644 128918 281298 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 358958 128918 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 -1644 159638 281298 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 358958 159638 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 -1644 190358 281298 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 358958 190358 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 -1644 221078 56794 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 321718 221078 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 -1644 251798 56794 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 321718 251798 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 -1644 282518 56794 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 321718 282518 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 -1644 313238 56794 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 321718 313238 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 -1644 343958 56794 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 321718 343958 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 -1644 374678 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 -1644 405398 46266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 184022 405398 215898 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 311926 405398 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 -1644 436118 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 -1644 466838 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 -1644 497558 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 -1644 528278 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 -1644 558998 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 589098 -1644 589718 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 -1644 9758 280964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 328428 9758 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 -1644 40478 280964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 328428 40478 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 -1644 71198 286194 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 330590 71198 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 -1644 101918 286194 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 330590 101918 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 -1644 132638 281298 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 358958 132638 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 -1644 163358 281298 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 358958 163358 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 -1644 194078 281298 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 358958 194078 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 -1644 224798 56794 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 321718 224798 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 -1644 255518 56794 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 321718 255518 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 -1644 286238 56794 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 321718 286238 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 -1644 316958 56794 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 321718 316958 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 -1644 347678 56794 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 321718 347678 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 -1644 378398 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 33828 409118 46266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 116310 409118 136602 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 184022 409118 215898 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 261638 409118 275930 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 311926 409118 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 -1644 439838 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 -1644 470558 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 -1644 501278 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 -1644 531998 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 -1644 562718 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 592818 -1644 593438 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 528154 22322 528154 22322 0 vdd
rlabel via4 538622 28322 538622 28322 0 vss
rlabel metal3 567784 7112 567784 7112 0 io_in[0]
rlabel metal3 4144 280504 4144 280504 0 io_in[10]
rlabel metal2 20552 278978 20552 278978 0 io_in[11]
rlabel metal3 56350 304920 56350 304920 0 io_in[12]
rlabel metal3 54936 304486 54936 304486 0 io_in[13]
rlabel metal3 593138 562184 593138 562184 0 io_in[14]
rlabel metal2 584696 592914 584696 592914 0 io_in[15]
rlabel metal2 518504 593138 518504 593138 0 io_in[16]
rlabel metal2 93688 351022 93688 351022 0 io_in[17]
rlabel metal2 217224 334278 217224 334278 0 io_in[18]
rlabel metal3 275184 330120 275184 330120 0 io_in[19]
rlabel metal3 593138 46760 593138 46760 0 io_in[1]
rlabel metal3 248696 589624 248696 589624 0 io_in[20]
rlabel metal2 187544 484722 187544 484722 0 io_in[21]
rlabel metal2 121576 593194 121576 593194 0 io_in[22]
rlabel metal2 55160 553602 55160 553602 0 io_in[23]
rlabel metal5 199024 305730 199024 305730 0 io_in[24]
rlabel metal3 54390 544824 54390 544824 0 io_in[25]
rlabel metal3 56910 502488 56910 502488 0 io_in[26]
rlabel metal2 196168 276066 196168 276066 0 io_in[27]
rlabel metal2 195496 276850 195496 276850 0 io_in[28]
rlabel metal2 194824 276682 194824 276682 0 io_in[29]
rlabel metal3 548422 13832 548422 13832 0 io_in[2]
rlabel metal3 2366 333144 2366 333144 0 io_in[30]
rlabel metal5 6216 290790 6216 290790 0 io_in[31]
rlabel metal3 2702 248584 2702 248584 0 io_in[32]
rlabel metal3 2310 206360 2310 206360 0 io_in[33]
rlabel metal3 190960 275576 190960 275576 0 io_in[34]
rlabel metal3 3990 121688 3990 121688 0 io_in[35]
rlabel metal3 2310 79352 2310 79352 0 io_in[36]
rlabel metal4 189448 272023 189448 272023 0 io_in[37]
rlabel metal4 572040 71624 572040 71624 0 io_in[3]
rlabel metal3 542150 20552 542150 20552 0 io_in[4]
rlabel metal3 550102 23912 550102 23912 0 io_in[5]
rlabel metal3 542094 27272 542094 27272 0 io_in[6]
rlabel metal4 565320 157640 565320 157640 0 io_in[7]
rlabel metal1 44520 163128 44520 163128 0 io_in[8]
rlabel metal3 593082 363944 593082 363944 0 io_in[9]
rlabel metal3 545118 9352 545118 9352 0 io_oeb[0]
rlabel metal3 326802 430136 326802 430136 0 io_oeb[10]
rlabel metal3 3290 284760 3290 284760 0 io_oeb[11]
rlabel metal4 45416 280672 45416 280672 0 io_oeb[12]
rlabel metal3 49112 280616 49112 280616 0 io_oeb[13]
rlabel metal3 54824 288246 54824 288246 0 io_oeb[14]
rlabel metal2 540568 487242 540568 487242 0 io_oeb[15]
rlabel metal2 101080 278586 101080 278586 0 io_oeb[16]
rlabel metal2 408296 592242 408296 592242 0 io_oeb[17]
rlabel metal2 270088 333438 270088 333438 0 io_oeb[18]
rlabel metal2 283304 327614 283304 327614 0 io_oeb[19]
rlabel metal3 542542 12712 542542 12712 0 io_oeb[1]
rlabel metal2 209608 478002 209608 478002 0 io_oeb[20]
rlabel metal2 143416 488082 143416 488082 0 io_oeb[21]
rlabel metal2 77448 593250 77448 593250 0 io_oeb[22]
rlabel metal2 11256 593194 11256 593194 0 io_oeb[23]
rlabel metal2 176610 280056 176610 280056 0 io_oeb[24]
rlabel metal3 280 516488 280 516488 0 io_oeb[25]
rlabel metal4 115080 277721 115080 277721 0 io_oeb[26]
rlabel metal3 55230 431928 55230 431928 0 io_oeb[27]
rlabel metal3 56126 389592 56126 389592 0 io_oeb[28]
rlabel metal3 59654 347256 59654 347256 0 io_oeb[29]
rlabel metal3 543382 16072 543382 16072 0 io_oeb[2]
rlabel metal3 280 304808 280 304808 0 io_oeb[30]
rlabel metal3 3598 262808 3598 262808 0 io_oeb[31]
rlabel metal3 4102 220472 4102 220472 0 io_oeb[32]
rlabel metal3 4046 178024 4046 178024 0 io_oeb[33]
rlabel metal2 169834 280056 169834 280056 0 io_oeb[34]
rlabel metal3 2366 93464 2366 93464 0 io_oeb[35]
rlabel metal3 336 51240 336 51240 0 io_oeb[36]
rlabel metal3 2366 8792 2366 8792 0 io_oeb[37]
rlabel metal3 541870 19432 541870 19432 0 io_oeb[3]
rlabel metal3 544222 22792 544222 22792 0 io_oeb[4]
rlabel metal3 541758 26152 541758 26152 0 io_oeb[5]
rlabel metal3 545062 29512 545062 29512 0 io_oeb[6]
rlabel metal3 541702 32872 541702 32872 0 io_oeb[7]
rlabel metal2 540120 197176 540120 197176 0 io_oeb[8]
rlabel metal3 511574 70616 511574 70616 0 io_oeb[9]
rlabel metal3 544222 8232 544222 8232 0 io_out[0]
rlabel metal3 49392 280392 49392 280392 0 io_out[10]
rlabel metal2 42728 279146 42728 279146 0 io_out[11]
rlabel metal4 49560 388192 49560 388192 0 io_out[12]
rlabel metal4 25928 281064 25928 281064 0 io_out[13]
rlabel metal2 31304 279314 31304 279314 0 io_out[14]
rlabel metal2 562632 593082 562632 593082 0 io_out[15]
rlabel metal3 495600 590184 495600 590184 0 io_out[16]
rlabel metal2 430248 490602 430248 490602 0 io_out[17]
rlabel metal2 364056 593194 364056 593194 0 io_out[18]
rlabel metal2 336168 340998 336168 340998 0 io_out[19]
rlabel metal3 541982 11592 541982 11592 0 io_out[1]
rlabel metal3 290528 336840 290528 336840 0 io_out[20]
rlabel metal2 165704 593250 165704 593250 0 io_out[21]
rlabel metal2 99512 593306 99512 593306 0 io_out[22]
rlabel metal2 188104 277970 188104 277970 0 io_out[23]
rlabel metal4 187432 278339 187432 278339 0 io_out[24]
rlabel metal3 1470 530712 1470 530712 0 io_out[25]
rlabel metal3 2310 488376 2310 488376 0 io_out[26]
rlabel metal3 2422 446040 2422 446040 0 io_out[27]
rlabel metal3 336 403592 336 403592 0 io_out[28]
rlabel metal3 59542 361368 59542 361368 0 io_out[29]
rlabel metal4 590184 98952 590184 98952 0 io_out[2]
rlabel metal3 2366 319032 2366 319032 0 io_out[30]
rlabel metal3 4214 276696 4214 276696 0 io_out[31]
rlabel metal3 5726 234584 5726 234584 0 io_out[32]
rlabel metal3 5670 192248 5670 192248 0 io_out[33]
rlabel metal5 141568 264870 141568 264870 0 io_out[34]
rlabel metal3 3990 107464 3990 107464 0 io_out[35]
rlabel metal3 2310 65240 2310 65240 0 io_out[36]
rlabel metal3 280 23016 280 23016 0 io_out[37]
rlabel metal3 541926 18312 541926 18312 0 io_out[3]
rlabel metal3 546742 21672 546742 21672 0 io_out[4]
rlabel metal3 541814 25032 541814 25032 0 io_out[5]
rlabel metal3 547582 28392 547582 28392 0 io_out[6]
rlabel metal4 563640 164136 563640 164136 0 io_out[7]
rlabel metal3 529648 45080 529648 45080 0 io_out[8]
rlabel metal3 553602 377160 553602 377160 0 io_out[9]
rlabel metal2 213192 1974 213192 1974 0 la_data_in[0]
rlabel metal2 257992 3850 257992 3850 0 la_data_in[10]
rlabel metal2 262696 3962 262696 3962 0 la_data_in[11]
rlabel metal2 281736 1414 281736 1414 0 la_data_in[12]
rlabel metal2 287448 1806 287448 1806 0 la_data_in[13]
rlabel metal2 276808 4018 276808 4018 0 la_data_in[14]
rlabel metal2 281512 4522 281512 4522 0 la_data_in[15]
rlabel metal2 286216 3850 286216 3850 0 la_data_in[16]
rlabel metal2 310296 2366 310296 2366 0 la_data_in[17]
rlabel metal2 295624 4746 295624 4746 0 la_data_in[18]
rlabel metal2 300328 4130 300328 4130 0 la_data_in[19]
rlabel metal2 218904 1918 218904 1918 0 la_data_in[1]
rlabel metal2 305032 4970 305032 4970 0 la_data_in[20]
rlabel metal2 309736 3962 309736 3962 0 la_data_in[21]
rlabel metal2 314440 4522 314440 4522 0 la_data_in[22]
rlabel metal2 319144 4634 319144 4634 0 la_data_in[23]
rlabel metal2 350280 1862 350280 1862 0 la_data_in[24]
rlabel metal2 328552 4858 328552 4858 0 la_data_in[25]
rlabel metal2 361704 2758 361704 2758 0 la_data_in[26]
rlabel metal2 337960 4970 337960 4970 0 la_data_in[27]
rlabel metal2 373016 336 373016 336 0 la_data_in[28]
rlabel metal2 378840 574 378840 574 0 la_data_in[29]
rlabel metal2 224616 1918 224616 1918 0 la_data_in[2]
rlabel metal2 352072 2954 352072 2954 0 la_data_in[30]
rlabel metal2 356776 2786 356776 2786 0 la_data_in[31]
rlabel metal2 364504 1232 364504 1232 0 la_data_in[32]
rlabel metal2 401688 518 401688 518 0 la_data_in[33]
rlabel metal2 407288 392 407288 392 0 la_data_in[34]
rlabel metal2 376264 2632 376264 2632 0 la_data_in[35]
rlabel metal2 380072 2576 380072 2576 0 la_data_in[36]
rlabel metal2 424536 966 424536 966 0 la_data_in[37]
rlabel metal2 430248 2310 430248 2310 0 la_data_in[38]
rlabel metal2 394408 3346 394408 3346 0 la_data_in[39]
rlabel metal2 230328 1470 230328 1470 0 la_data_in[3]
rlabel metal2 399112 2898 399112 2898 0 la_data_in[40]
rlabel metal2 403816 2954 403816 2954 0 la_data_in[41]
rlabel metal2 453096 518 453096 518 0 la_data_in[42]
rlabel metal3 420000 1064 420000 1064 0 la_data_in[43]
rlabel metal2 417928 2786 417928 2786 0 la_data_in[44]
rlabel metal2 423304 3248 423304 3248 0 la_data_in[45]
rlabel metal2 427336 2730 427336 2730 0 la_data_in[46]
rlabel metal2 433048 2688 433048 2688 0 la_data_in[47]
rlabel metal4 436856 1008 436856 1008 0 la_data_in[48]
rlabel metal2 493080 1918 493080 1918 0 la_data_in[49]
rlabel metal2 236040 1638 236040 1638 0 la_data_in[4]
rlabel metal2 446152 2898 446152 2898 0 la_data_in[50]
rlabel metal2 450856 2954 450856 2954 0 la_data_in[51]
rlabel metal2 455560 3178 455560 3178 0 la_data_in[52]
rlabel metal2 515928 1918 515928 1918 0 la_data_in[53]
rlabel metal2 521640 518 521640 518 0 la_data_in[54]
rlabel metal2 469672 2786 469672 2786 0 la_data_in[55]
rlabel metal2 533064 2870 533064 2870 0 la_data_in[56]
rlabel metal2 538776 518 538776 518 0 la_data_in[57]
rlabel metal2 544376 392 544376 392 0 la_data_in[58]
rlabel metal2 488488 2618 488488 2618 0 la_data_in[59]
rlabel metal2 241752 1526 241752 1526 0 la_data_in[5]
rlabel metal2 555912 2814 555912 2814 0 la_data_in[60]
rlabel metal2 497896 3346 497896 3346 0 la_data_in[61]
rlabel metal2 567224 280 567224 280 0 la_data_in[62]
rlabel metal2 573048 2758 573048 2758 0 la_data_in[63]
rlabel metal2 239176 4746 239176 4746 0 la_data_in[6]
rlabel metal2 253176 2030 253176 2030 0 la_data_in[7]
rlabel metal2 258888 1582 258888 1582 0 la_data_in[8]
rlabel metal2 264600 1862 264600 1862 0 la_data_in[9]
rlabel metal2 215096 1918 215096 1918 0 la_data_out[0]
rlabel metal2 259560 4018 259560 4018 0 la_data_out[10]
rlabel metal2 264264 3906 264264 3906 0 la_data_out[11]
rlabel metal2 283640 1862 283640 1862 0 la_data_out[12]
rlabel metal2 289352 1750 289352 1750 0 la_data_out[13]
rlabel metal2 278376 3962 278376 3962 0 la_data_out[14]
rlabel metal2 283080 4914 283080 4914 0 la_data_out[15]
rlabel metal2 287784 4578 287784 4578 0 la_data_out[16]
rlabel metal2 312200 1470 312200 1470 0 la_data_out[17]
rlabel metal2 297192 4802 297192 4802 0 la_data_out[18]
rlabel metal2 301896 4914 301896 4914 0 la_data_out[19]
rlabel metal2 217224 4298 217224 4298 0 la_data_out[1]
rlabel metal2 306600 4018 306600 4018 0 la_data_out[20]
rlabel metal2 311304 3906 311304 3906 0 la_data_out[21]
rlabel metal2 316680 5040 316680 5040 0 la_data_out[22]
rlabel metal2 320712 4690 320712 4690 0 la_data_out[23]
rlabel metal2 352184 1806 352184 1806 0 la_data_out[24]
rlabel metal2 330120 4074 330120 4074 0 la_data_out[25]
rlabel metal2 334824 4018 334824 4018 0 la_data_out[26]
rlabel metal2 339528 3962 339528 3962 0 la_data_out[27]
rlabel metal2 375032 1470 375032 1470 0 la_data_out[28]
rlabel metal2 380744 1582 380744 1582 0 la_data_out[29]
rlabel metal2 226520 1974 226520 1974 0 la_data_out[2]
rlabel metal2 386680 2814 386680 2814 0 la_data_out[30]
rlabel metal2 358344 3738 358344 3738 0 la_data_out[31]
rlabel metal2 397880 1526 397880 1526 0 la_data_out[32]
rlabel metal2 403200 5096 403200 5096 0 la_data_out[33]
rlabel metal2 381416 3472 381416 3472 0 la_data_out[34]
rlabel metal2 377160 3794 377160 3794 0 la_data_out[35]
rlabel metal2 382214 5320 382214 5320 0 la_data_out[36]
rlabel metal2 426440 1750 426440 1750 0 la_data_out[37]
rlabel metal2 391272 3626 391272 3626 0 la_data_out[38]
rlabel metal2 396214 5544 396214 5544 0 la_data_out[39]
rlabel metal2 232232 1526 232232 1526 0 la_data_out[3]
rlabel metal2 401030 5432 401030 5432 0 la_data_out[40]
rlabel metal2 405384 4018 405384 4018 0 la_data_out[41]
rlabel metal3 449288 3304 449288 3304 0 la_data_out[42]
rlabel metal2 414792 3906 414792 3906 0 la_data_out[43]
rlabel metal2 419846 5320 419846 5320 0 la_data_out[44]
rlabel metal2 424200 3850 424200 3850 0 la_data_out[45]
rlabel metal2 429254 5208 429254 5208 0 la_data_out[46]
rlabel metal3 443240 5040 443240 5040 0 la_data_out[47]
rlabel metal2 438312 3794 438312 3794 0 la_data_out[48]
rlabel metal4 494984 4273 494984 4273 0 la_data_out[49]
rlabel metal2 237944 1582 237944 1582 0 la_data_out[4]
rlabel via4 447720 3317 447720 3317 0 la_data_out[50]
rlabel metal2 452424 4130 452424 4130 0 la_data_out[51]
rlabel metal4 457128 1709 457128 1709 0 la_data_out[52]
rlabel metal2 517832 1246 517832 1246 0 la_data_out[53]
rlabel metal2 523544 2982 523544 2982 0 la_data_out[54]
rlabel metal4 475496 4307 475496 4307 0 la_data_out[55]
rlabel metal2 475944 3850 475944 3850 0 la_data_out[56]
rlabel metal2 540680 574 540680 574 0 la_data_out[57]
rlabel metal2 546392 1750 546392 1750 0 la_data_out[58]
rlabel metal2 490056 4018 490056 4018 0 la_data_out[59]
rlabel metal2 236040 4242 236040 4242 0 la_data_out[5]
rlabel via4 499016 5113 499016 5113 0 la_data_out[60]
rlabel metal4 499464 3227 499464 3227 0 la_data_out[61]
rlabel metal4 569240 353 569240 353 0 la_data_out[62]
rlabel metal2 508872 3906 508872 3906 0 la_data_out[63]
rlabel metal2 240744 4802 240744 4802 0 la_data_out[6]
rlabel metal2 255080 2086 255080 2086 0 la_data_out[7]
rlabel metal2 260792 1470 260792 1470 0 la_data_out[8]
rlabel metal2 266504 1806 266504 1806 0 la_data_out[9]
rlabel metal2 217000 1974 217000 1974 0 la_oenb[0]
rlabel metal2 261128 3794 261128 3794 0 la_oenb[10]
rlabel metal2 265832 3682 265832 3682 0 la_oenb[11]
rlabel metal2 285656 1526 285656 1526 0 la_oenb[12]
rlabel metal2 275240 3794 275240 3794 0 la_oenb[13]
rlabel metal2 279944 3906 279944 3906 0 la_oenb[14]
rlabel metal2 284648 4970 284648 4970 0 la_oenb[15]
rlabel metal2 289352 4634 289352 4634 0 la_oenb[16]
rlabel metal2 294728 5040 294728 5040 0 la_oenb[17]
rlabel metal2 298760 4858 298760 4858 0 la_oenb[18]
rlabel metal2 303464 4074 303464 4074 0 la_oenb[19]
rlabel metal2 218792 4354 218792 4354 0 la_oenb[1]
rlabel metal2 308168 3850 308168 3850 0 la_oenb[20]
rlabel metal2 312872 3794 312872 3794 0 la_oenb[21]
rlabel metal2 317576 4578 317576 4578 0 la_oenb[22]
rlabel metal2 322280 4746 322280 4746 0 la_oenb[23]
rlabel metal2 326984 4802 326984 4802 0 la_oenb[24]
rlabel metal2 331688 3850 331688 3850 0 la_oenb[25]
rlabel metal2 336392 4914 336392 4914 0 la_oenb[26]
rlabel metal2 341768 5040 341768 5040 0 la_oenb[27]
rlabel metal2 359576 2912 359576 2912 0 la_oenb[28]
rlabel metal2 351064 4480 351064 4480 0 la_oenb[29]
rlabel metal2 228536 2030 228536 2030 0 la_oenb[2]
rlabel metal2 355208 4130 355208 4130 0 la_oenb[30]
rlabel metal2 359912 4186 359912 4186 0 la_oenb[31]
rlabel metal2 399896 2198 399896 2198 0 la_oenb[32]
rlabel metal2 405496 1358 405496 1358 0 la_oenb[33]
rlabel metal2 377944 3416 377944 3416 0 la_oenb[34]
rlabel metal2 378728 4018 378728 4018 0 la_oenb[35]
rlabel metal2 383432 4186 383432 4186 0 la_oenb[36]
rlabel metal2 428568 2086 428568 2086 0 la_oenb[37]
rlabel metal2 393064 5040 393064 5040 0 la_oenb[38]
rlabel metal2 397544 3570 397544 3570 0 la_oenb[39]
rlabel metal2 234136 1414 234136 1414 0 la_oenb[3]
rlabel metal2 402248 3962 402248 3962 0 la_oenb[40]
rlabel metal2 407624 4368 407624 4368 0 la_oenb[41]
rlabel metal2 412328 4536 412328 4536 0 la_oenb[42]
rlabel metal2 450296 2912 450296 2912 0 la_oenb[43]
rlabel metal2 421064 3682 421064 3682 0 la_oenb[44]
rlabel metal2 425768 4970 425768 4970 0 la_oenb[45]
rlabel metal2 430472 3514 430472 3514 0 la_oenb[46]
rlabel metal2 435848 4424 435848 4424 0 la_oenb[47]
rlabel metal2 491176 2030 491176 2030 0 la_oenb[48]
rlabel metal2 444584 4690 444584 4690 0 la_oenb[49]
rlabel metal2 239848 1470 239848 1470 0 la_oenb[4]
rlabel metal2 449288 3458 449288 3458 0 la_oenb[50]
rlabel metal2 454664 5040 454664 5040 0 la_oenb[51]
rlabel metal2 514136 2086 514136 2086 0 la_oenb[52]
rlabel metal2 519736 2422 519736 2422 0 la_oenb[53]
rlabel metal2 468104 4802 468104 4802 0 la_oenb[54]
rlabel metal2 472808 3738 472808 3738 0 la_oenb[55]
rlabel metal2 477512 4858 477512 4858 0 la_oenb[56]
rlabel metal2 542640 1736 542640 1736 0 la_oenb[57]
rlabel metal2 548296 2590 548296 2590 0 la_oenb[58]
rlabel metal2 491624 3962 491624 3962 0 la_oenb[59]
rlabel metal2 237608 4298 237608 4298 0 la_oenb[5]
rlabel metal2 496328 4970 496328 4970 0 la_oenb[60]
rlabel via4 501704 3317 501704 3317 0 la_oenb[61]
rlabel metal4 571256 443 571256 443 0 la_oenb[62]
rlabel metal2 510440 3850 510440 3850 0 la_oenb[63]
rlabel metal2 242312 4858 242312 4858 0 la_oenb[6]
rlabel metal2 257096 1918 257096 1918 0 la_oenb[7]
rlabel metal2 262696 1414 262696 1414 0 la_oenb[8]
rlabel metal2 256424 4074 256424 4074 0 la_oenb[9]
rlabel metal3 3906 305592 3906 305592 0 mem_addr\[0\]
rlabel metal2 44184 164010 44184 164010 0 mem_addr\[10\]
rlabel metal4 166152 359113 166152 359113 0 mem_addr\[11\]
rlabel metal3 4186 315672 4186 315672 0 mem_addr\[12\]
rlabel metal3 4130 312312 4130 312312 0 mem_addr\[13\]
rlabel metal3 4074 310968 4074 310968 0 mem_addr\[14\]
rlabel metal4 5096 325095 5096 325095 0 mem_addr\[15\]
rlabel metal3 5544 319942 5544 319942 0 mem_addr\[16\]
rlabel metal3 3850 312984 3850 312984 0 mem_addr\[17\]
rlabel metal2 161448 360542 161448 360542 0 mem_addr\[18\]
rlabel metal3 3962 304920 3962 304920 0 mem_addr\[19\]
rlabel metal3 5656 303814 5656 303814 0 mem_addr\[1\]
rlabel metal3 5320 308518 5320 308518 0 mem_addr\[20\]
rlabel metal3 4858 313656 4858 313656 0 mem_addr\[21\]
rlabel metal3 4914 311640 4914 311640 0 mem_addr\[22\]
rlabel metal3 3906 310296 3906 310296 0 mem_addr\[23\]
rlabel metal2 157654 359912 157654 359912 0 mem_addr\[24\]
rlabel metal3 209650 123032 209650 123032 0 mem_addr\[25\]
rlabel metal2 156142 359912 156142 359912 0 mem_addr\[26\]
rlabel metal3 209762 128408 209762 128408 0 mem_addr\[27\]
rlabel metal2 154728 361718 154728 361718 0 mem_addr\[28\]
rlabel metal3 209874 133784 209874 133784 0 mem_addr\[29\]
rlabel metal3 3290 308952 3290 308952 0 mem_addr\[2\]
rlabel metal3 154560 362152 154560 362152 0 mem_addr\[30\]
rlabel metal3 207130 139160 207130 139160 0 mem_addr\[31\]
rlabel metal3 4018 306264 4018 306264 0 mem_addr\[3\]
rlabel metal3 4186 307608 4186 307608 0 mem_addr\[4\]
rlabel metal2 166600 163170 166600 163170 0 mem_addr\[5\]
rlabel metal2 43918 144872 43918 144872 0 mem_addr\[6\]
rlabel metal2 44366 144872 44366 144872 0 mem_addr\[7\]
rlabel metal2 44814 144872 44814 144872 0 mem_addr\[8\]
rlabel metal2 44506 165032 44506 165032 0 mem_addr\[9\]
rlabel metal3 208810 50456 208810 50456 0 mem_instr
rlabel metal2 147336 363286 147336 363286 0 mem_rdata\[0\]
rlabel metal3 210000 266056 210000 266056 0 mem_rdata\[10\]
rlabel metal2 139944 363230 139944 363230 0 mem_rdata\[11\]
rlabel metal2 139272 365694 139272 365694 0 mem_rdata\[12\]
rlabel metal2 138600 363510 138600 363510 0 mem_rdata\[13\]
rlabel metal2 137928 362390 137928 362390 0 mem_rdata\[14\]
rlabel metal3 208138 278936 208138 278936 0 mem_rdata\[15\]
rlabel metal3 207186 281624 207186 281624 0 mem_rdata\[16\]
rlabel metal3 210056 284662 210056 284662 0 mem_rdata\[17\]
rlabel metal3 209706 287000 209706 287000 0 mem_rdata\[18\]
rlabel metal2 134568 360094 134568 360094 0 mem_rdata\[19\]
rlabel metal2 146664 363342 146664 363342 0 mem_rdata\[1\]
rlabel metal2 133896 365750 133896 365750 0 mem_rdata\[20\]
rlabel metal3 208194 295064 208194 295064 0 mem_rdata\[21\]
rlabel metal2 132552 362502 132552 362502 0 mem_rdata\[22\]
rlabel metal2 132118 359912 132118 359912 0 mem_rdata\[23\]
rlabel metal3 205394 303128 205394 303128 0 mem_rdata\[24\]
rlabel metal3 208306 305816 208306 305816 0 mem_rdata\[25\]
rlabel metal2 129864 360038 129864 360038 0 mem_rdata\[26\]
rlabel metal3 208810 311192 208810 311192 0 mem_rdata\[27\]
rlabel metal3 205618 313880 205618 313880 0 mem_rdata\[28\]
rlabel metal2 143640 362600 143640 362600 0 mem_rdata\[29\]
rlabel metal2 145992 361606 145992 361606 0 mem_rdata\[2\]
rlabel metal3 210280 319606 210280 319606 0 mem_rdata\[30\]
rlabel metal3 210168 322238 210168 322238 0 mem_rdata\[31\]
rlabel metal2 145320 361550 145320 361550 0 mem_rdata\[3\]
rlabel metal2 144648 364238 144648 364238 0 mem_rdata\[4\]
rlabel metal2 143976 364854 143976 364854 0 mem_rdata\[5\]
rlabel metal2 143304 361942 143304 361942 0 mem_rdata\[6\]
rlabel metal4 210728 257641 210728 257641 0 mem_rdata\[7\]
rlabel metal2 141960 365134 141960 365134 0 mem_rdata\[8\]
rlabel metal2 141288 360206 141288 360206 0 mem_rdata\[9\]
rlabel metal3 208754 53144 208754 53144 0 mem_ready
rlabel metal4 212296 344025 212296 344025 0 mem_valid
rlabel metal2 72856 331702 72856 331702 0 mem_wdata\[0\]
rlabel metal4 48776 276857 48776 276857 0 mem_wdata\[10\]
rlabel metal2 50120 278586 50120 278586 0 mem_wdata\[11\]
rlabel metal4 186984 358247 186984 358247 0 mem_wdata\[12\]
rlabel metal4 7112 276317 7112 276317 0 mem_wdata\[13\]
rlabel metal2 71750 280056 71750 280056 0 mem_wdata\[14\]
rlabel metal2 117880 146398 117880 146398 0 mem_wdata\[15\]
rlabel metal2 20566 165704 20566 165704 0 mem_wdata\[16\]
rlabel metal3 26768 165704 26768 165704 0 mem_wdata\[17\]
rlabel metal3 28280 165704 28280 165704 0 mem_wdata\[18\]
rlabel metal2 39270 165704 39270 165704 0 mem_wdata\[19\]
rlabel metal2 27272 279930 27272 279930 0 mem_wdata\[1\]
rlabel metal2 71638 165704 71638 165704 0 mem_wdata\[20\]
rlabel metal3 210056 198702 210056 198702 0 mem_wdata\[21\]
rlabel metal3 190680 280392 190680 280392 0 mem_wdata\[22\]
rlabel metal2 92120 164794 92120 164794 0 mem_wdata\[23\]
rlabel metal2 120274 165592 120274 165592 0 mem_wdata\[24\]
rlabel metal3 109704 279048 109704 279048 0 mem_wdata\[25\]
rlabel metal5 209832 276480 209832 276480 0 mem_wdata\[26\]
rlabel metal2 138824 164794 138824 164794 0 mem_wdata\[27\]
rlabel metal2 171528 164794 171528 164794 0 mem_wdata\[28\]
rlabel metal2 5768 278418 5768 278418 0 mem_wdata\[29\]
rlabel metal2 70392 333424 70392 333424 0 mem_wdata\[2\]
rlabel metal2 24584 278362 24584 278362 0 mem_wdata\[30\]
rlabel metal2 28966 280056 28966 280056 0 mem_wdata\[31\]
rlabel metal2 70504 332920 70504 332920 0 mem_wdata\[3\]
rlabel metal2 72184 331422 72184 331422 0 mem_wdata\[4\]
rlabel metal2 27790 144872 27790 144872 0 mem_wdata\[5\]
rlabel metal2 26446 144872 26446 144872 0 mem_wdata\[6\]
rlabel via4 190792 359563 190792 359563 0 mem_wdata\[7\]
rlabel metal4 189560 359147 189560 359147 0 mem_wdata\[8\]
rlabel metal4 189560 165256 189560 165256 0 mem_wdata\[9\]
rlabel metal2 150024 364350 150024 364350 0 mem_wstrb\[0\]
rlabel metal2 149352 365974 149352 365974 0 mem_wstrb\[1\]
rlabel metal2 148680 360878 148680 360878 0 mem_wstrb\[2\]
rlabel metal4 210728 235999 210728 235999 0 mem_wstrb\[3\]
rlabel metal4 374808 278320 374808 278320 0 pcpi_approx_mul_rd\[0\]
rlabel metal4 375704 283976 375704 283976 0 pcpi_approx_mul_rd\[10\]
rlabel metal3 371014 292376 371014 292376 0 pcpi_approx_mul_rd\[11\]
rlabel metal4 375480 285152 375480 285152 0 pcpi_approx_mul_rd\[12\]
rlabel metal4 373800 285768 373800 285768 0 pcpi_approx_mul_rd\[13\]
rlabel metal4 373800 303343 373800 303343 0 pcpi_approx_mul_rd\[14\]
rlabel metal3 371070 296856 371070 296856 0 pcpi_approx_mul_rd\[15\]
rlabel metal2 375816 285712 375816 285712 0 pcpi_approx_mul_rd\[16\]
rlabel metal3 380072 300314 380072 300314 0 pcpi_approx_mul_rd\[17\]
rlabel metal4 376488 301056 376488 301056 0 pcpi_approx_mul_rd\[18\]
rlabel metal3 380072 301294 380072 301294 0 pcpi_approx_mul_rd\[19\]
rlabel metal4 374920 278264 374920 278264 0 pcpi_approx_mul_rd\[1\]
rlabel metal3 378658 299880 378658 299880 0 pcpi_approx_mul_rd\[20\]
rlabel metal2 375592 288456 375592 288456 0 pcpi_approx_mul_rd\[21\]
rlabel metal2 375592 315392 375592 315392 0 pcpi_approx_mul_rd\[22\]
rlabel metal2 375816 316064 375816 316064 0 pcpi_approx_mul_rd\[23\]
rlabel metal3 376866 299208 376866 299208 0 pcpi_approx_mul_rd\[24\]
rlabel metal3 376978 298536 376978 298536 0 pcpi_approx_mul_rd\[25\]
rlabel metal4 375480 316008 375480 316008 0 pcpi_approx_mul_rd\[26\]
rlabel metal2 375704 317352 375704 317352 0 pcpi_approx_mul_rd\[27\]
rlabel metal4 378840 317184 378840 317184 0 pcpi_approx_mul_rd\[28\]
rlabel metal4 373800 313348 373800 313348 0 pcpi_approx_mul_rd\[29\]
rlabel metal4 373464 278712 373464 278712 0 pcpi_approx_mul_rd\[2\]
rlabel metal4 379064 318360 379064 318360 0 pcpi_approx_mul_rd\[30\]
rlabel metal4 373800 318696 373800 318696 0 pcpi_approx_mul_rd\[31\]
rlabel metal4 375592 279328 375592 279328 0 pcpi_approx_mul_rd\[3\]
rlabel metal4 373352 280784 373352 280784 0 pcpi_approx_mul_rd\[4\]
rlabel metal3 370958 285656 370958 285656 0 pcpi_approx_mul_rd\[5\]
rlabel metal3 371126 286776 371126 286776 0 pcpi_approx_mul_rd\[6\]
rlabel metal4 373912 280784 373912 280784 0 pcpi_approx_mul_rd\[7\]
rlabel metal3 371182 289016 371182 289016 0 pcpi_approx_mul_rd\[8\]
rlabel metal4 373688 282800 373688 282800 0 pcpi_approx_mul_rd\[9\]
rlabel metal4 377608 320376 377608 320376 0 pcpi_approx_mul_ready
rlabel metal2 375480 293552 375480 293552 0 pcpi_approx_mul_wait
rlabel metal4 373912 321384 373912 321384 0 pcpi_approx_mul_wr
rlabel metal2 384440 202776 384440 202776 0 pcpi_div_rd\[0\]
rlabel metal4 373912 213683 373912 213683 0 pcpi_div_rd\[10\]
rlabel metal3 370062 215096 370062 215096 0 pcpi_div_rd\[11\]
rlabel metal4 373128 208544 373128 208544 0 pcpi_div_rd\[12\]
rlabel metal3 374822 217336 374822 217336 0 pcpi_div_rd\[13\]
rlabel via4 373912 218443 373912 218443 0 pcpi_div_rd\[14\]
rlabel metal4 378728 216843 378728 216843 0 pcpi_div_rd\[15\]
rlabel metal4 369544 207323 369544 207323 0 pcpi_div_rd\[16\]
rlabel metal4 373744 195390 373744 195390 0 pcpi_div_rd\[17\]
rlabel metal3 441406 169960 441406 169960 0 pcpi_div_rd\[18\]
rlabel metal3 373800 202440 373800 202440 0 pcpi_div_rd\[19\]
rlabel metal2 375928 202440 375928 202440 0 pcpi_div_rd\[1\]
rlabel metal4 375256 215768 375256 215768 0 pcpi_div_rd\[20\]
rlabel metal3 370062 226296 370062 226296 0 pcpi_div_rd\[21\]
rlabel metal3 441070 172648 441070 172648 0 pcpi_div_rd\[22\]
rlabel metal3 370790 228536 370790 228536 0 pcpi_div_rd\[23\]
rlabel metal2 373464 208600 373464 208600 0 pcpi_div_rd\[24\]
rlabel metal3 370118 230776 370118 230776 0 pcpi_div_rd\[25\]
rlabel metal3 370902 231896 370902 231896 0 pcpi_div_rd\[26\]
rlabel metal4 373688 223653 373688 223653 0 pcpi_div_rd\[27\]
rlabel metal4 407624 205408 407624 205408 0 pcpi_div_rd\[28\]
rlabel metal2 375256 217336 375256 217336 0 pcpi_div_rd\[29\]
rlabel metal3 375256 205072 375256 205072 0 pcpi_div_rd\[2\]
rlabel metal3 377594 169960 377594 169960 0 pcpi_div_rd\[30\]
rlabel metal2 375872 204120 375872 204120 0 pcpi_div_rd\[31\]
rlabel metal4 403368 205632 403368 205632 0 pcpi_div_rd\[3\]
rlabel metal2 403592 196406 403592 196406 0 pcpi_div_rd\[4\]
rlabel metal2 375144 203112 375144 203112 0 pcpi_div_rd\[5\]
rlabel metal2 375480 203560 375480 203560 0 pcpi_div_rd\[6\]
rlabel metal4 373688 203280 373688 203280 0 pcpi_div_rd\[7\]
rlabel metal4 373912 203784 373912 203784 0 pcpi_div_rd\[8\]
rlabel metal4 373912 212403 373912 212403 0 pcpi_div_rd\[9\]
rlabel metal3 370006 239736 370006 239736 0 pcpi_div_ready
rlabel metal3 377818 174664 377818 174664 0 pcpi_div_wait
rlabel metal3 378770 178696 378770 178696 0 pcpi_div_wr
rlabel metal4 373464 241703 373464 241703 0 pcpi_exact_mul_rd\[0\]
rlabel metal4 376488 249704 376488 249704 0 pcpi_exact_mul_rd\[10\]
rlabel metal2 376152 259336 376152 259336 0 pcpi_exact_mul_rd\[11\]
rlabel metal3 378602 229880 378602 229880 0 pcpi_exact_mul_rd\[12\]
rlabel metal2 375368 260512 375368 260512 0 pcpi_exact_mul_rd\[13\]
rlabel metal2 375816 230440 375816 230440 0 pcpi_exact_mul_rd\[14\]
rlabel metal2 406952 204778 406952 204778 0 pcpi_exact_mul_rd\[15\]
rlabel metal3 376082 219800 376082 219800 0 pcpi_exact_mul_rd\[16\]
rlabel metal2 375592 232400 375592 232400 0 pcpi_exact_mul_rd\[17\]
rlabel metal4 373912 263088 373912 263088 0 pcpi_exact_mul_rd\[18\]
rlabel metal3 370174 262136 370174 262136 0 pcpi_exact_mul_rd\[19\]
rlabel metal4 373912 238000 373912 238000 0 pcpi_exact_mul_rd\[1\]
rlabel metal3 441448 235144 441448 235144 0 pcpi_exact_mul_rd\[20\]
rlabel metal3 371070 264376 371070 264376 0 pcpi_exact_mul_rd\[21\]
rlabel metal3 370006 265496 370006 265496 0 pcpi_exact_mul_rd\[22\]
rlabel metal2 375704 236320 375704 236320 0 pcpi_exact_mul_rd\[23\]
rlabel metal2 374696 267288 374696 267288 0 pcpi_exact_mul_rd\[24\]
rlabel metal3 440174 240632 440174 240632 0 pcpi_exact_mul_rd\[25\]
rlabel metal3 392798 269976 392798 269976 0 pcpi_exact_mul_rd\[26\]
rlabel metal2 381416 270480 381416 270480 0 pcpi_exact_mul_rd\[27\]
rlabel metal4 404040 268632 404040 268632 0 pcpi_exact_mul_rd\[28\]
rlabel metal4 373352 269864 373352 269864 0 pcpi_exact_mul_rd\[29\]
rlabel metal4 376264 239512 376264 239512 0 pcpi_exact_mul_rd\[2\]
rlabel metal4 375256 269528 375256 269528 0 pcpi_exact_mul_rd\[30\]
rlabel metal4 375144 271040 375144 271040 0 pcpi_exact_mul_rd\[31\]
rlabel metal4 373800 242370 373800 242370 0 pcpi_exact_mul_rd\[3\]
rlabel metal2 375256 256424 375256 256424 0 pcpi_exact_mul_rd\[4\]
rlabel metal4 376488 245560 376488 245560 0 pcpi_exact_mul_rd\[5\]
rlabel metal2 375480 256424 375480 256424 0 pcpi_exact_mul_rd\[6\]
rlabel metal2 407624 265174 407624 265174 0 pcpi_exact_mul_rd\[7\]
rlabel metal4 373016 245896 373016 245896 0 pcpi_exact_mul_rd\[8\]
rlabel metal4 373352 244776 373352 244776 0 pcpi_exact_mul_rd\[9\]
rlabel metal4 373576 271712 373576 271712 0 pcpi_exact_mul_ready
rlabel metal4 399560 206136 399560 206136 0 pcpi_exact_mul_wait
rlabel metal4 375032 276024 375032 276024 0 pcpi_exact_mul_wr
rlabel metal4 376320 75690 376320 75690 0 pcpi_insn\[0\]
rlabel metal5 380688 72090 380688 72090 0 pcpi_insn\[10\]
rlabel metal2 380688 67200 380688 67200 0 pcpi_insn\[11\]
rlabel metal3 378154 171976 378154 171976 0 pcpi_insn\[12\]
rlabel metal3 378042 91448 378042 91448 0 pcpi_insn\[13\]
rlabel metal3 376376 90832 376376 90832 0 pcpi_insn\[14\]
rlabel metal4 377608 71553 377608 71553 0 pcpi_insn\[15\]
rlabel via4 378840 72833 378840 72833 0 pcpi_insn\[16\]
rlabel metal4 378616 74169 378616 74169 0 pcpi_insn\[17\]
rlabel metal4 379624 74583 379624 74583 0 pcpi_insn\[18\]
rlabel metal4 379624 76403 379624 76403 0 pcpi_insn\[19\]
rlabel metal3 374752 233464 374752 233464 0 pcpi_insn\[1\]
rlabel metal4 378840 77683 378840 77683 0 pcpi_insn\[20\]
rlabel metal4 378840 78423 378840 78423 0 pcpi_insn\[21\]
rlabel metal4 378840 80063 378840 80063 0 pcpi_insn\[22\]
rlabel metal4 378840 80769 378840 80769 0 pcpi_insn\[23\]
rlabel metal4 378840 81723 378840 81723 0 pcpi_insn\[24\]
rlabel metal3 380072 96698 380072 96698 0 pcpi_insn\[25\]
rlabel metal4 373688 236320 373688 236320 0 pcpi_insn\[26\]
rlabel metal4 373016 94164 373016 94164 0 pcpi_insn\[27\]
rlabel metal3 376922 98168 376922 98168 0 pcpi_insn\[28\]
rlabel metal3 380072 88522 380072 88522 0 pcpi_insn\[29\]
rlabel via4 380408 216445 380408 216445 0 pcpi_insn\[2\]
rlabel metal3 378042 94808 378042 94808 0 pcpi_insn\[30\]
rlabel metal3 376586 97496 376586 97496 0 pcpi_insn\[31\]
rlabel metal3 377090 217112 377090 217112 0 pcpi_insn\[3\]
rlabel metal3 375480 72184 375480 72184 0 pcpi_insn\[4\]
rlabel metal2 373128 72968 373128 72968 0 pcpi_insn\[5\]
rlabel metal3 378098 225176 378098 225176 0 pcpi_insn\[6\]
rlabel metal4 377608 62843 377608 62843 0 pcpi_insn\[7\]
rlabel metal3 376432 217896 376432 217896 0 pcpi_insn\[8\]
rlabel metal3 377440 237720 377440 237720 0 pcpi_insn\[9\]
rlabel metal3 376026 93464 376026 93464 0 pcpi_mul_rd\[0\]
rlabel metal4 443800 112504 443800 112504 0 pcpi_mul_rd\[10\]
rlabel metal4 373352 141960 373352 141960 0 pcpi_mul_rd\[11\]
rlabel metal3 440902 76664 440902 76664 0 pcpi_mul_rd\[12\]
rlabel metal2 374024 186480 374024 186480 0 pcpi_mul_rd\[13\]
rlabel metal3 371854 179256 371854 179256 0 pcpi_mul_rd\[14\]
rlabel metal4 373688 178360 373688 178360 0 pcpi_mul_rd\[15\]
rlabel metal2 374136 186592 374136 186592 0 pcpi_mul_rd\[16\]
rlabel metal2 373128 191128 373128 191128 0 pcpi_mul_rd\[17\]
rlabel metal4 373688 187768 373688 187768 0 pcpi_mul_rd\[18\]
rlabel metal2 374472 189952 374472 189952 0 pcpi_mul_rd\[19\]
rlabel metal3 376138 92792 376138 92792 0 pcpi_mul_rd\[1\]
rlabel metal4 373912 185463 373912 185463 0 pcpi_mul_rd\[20\]
rlabel metal3 370622 187096 370622 187096 0 pcpi_mul_rd\[21\]
rlabel metal4 373912 191464 373912 191464 0 pcpi_mul_rd\[22\]
rlabel metal4 373800 192136 373800 192136 0 pcpi_mul_rd\[23\]
rlabel metal2 373240 193536 373240 193536 0 pcpi_mul_rd\[24\]
rlabel metal4 445368 139832 445368 139832 0 pcpi_mul_rd\[25\]
rlabel metal4 446936 139384 446936 139384 0 pcpi_mul_rd\[26\]
rlabel metal4 448616 139608 448616 139608 0 pcpi_mul_rd\[27\]
rlabel metal2 373128 195832 373128 195832 0 pcpi_mul_rd\[28\]
rlabel metal3 370678 196056 370678 196056 0 pcpi_mul_rd\[29\]
rlabel metal3 377930 92120 377930 92120 0 pcpi_mul_rd\[2\]
rlabel metal4 450296 141960 450296 141960 0 pcpi_mul_rd\[30\]
rlabel metal3 377762 81368 377762 81368 0 pcpi_mul_rd\[31\]
rlabel metal3 377874 88088 377874 88088 0 pcpi_mul_rd\[3\]
rlabel metal3 377818 76664 377818 76664 0 pcpi_mul_rd\[4\]
rlabel metal3 375074 78680 375074 78680 0 pcpi_mul_rd\[5\]
rlabel metal2 406280 44898 406280 44898 0 pcpi_mul_rd\[6\]
rlabel metal2 406952 44730 406952 44730 0 pcpi_mul_rd\[7\]
rlabel metal3 372638 172536 372638 172536 0 pcpi_mul_rd\[8\]
rlabel metal3 370902 173656 370902 173656 0 pcpi_mul_rd\[9\]
rlabel metal4 445256 140280 445256 140280 0 pcpi_mul_ready
rlabel metal3 376082 83384 376082 83384 0 pcpi_mul_wait
rlabel metal3 440174 79352 440174 79352 0 pcpi_mul_wr
rlabel metal4 376152 91153 376152 91153 0 pcpi_rs1\[0\]
rlabel metal4 377608 101793 377608 101793 0 pcpi_rs1\[10\]
rlabel metal3 378994 283752 378994 283752 0 pcpi_rs1\[11\]
rlabel metal3 379610 287784 379610 287784 0 pcpi_rs1\[12\]
rlabel metal3 379666 288456 379666 288456 0 pcpi_rs1\[13\]
rlabel metal3 377986 63224 377986 63224 0 pcpi_rs1\[14\]
rlabel metal3 377314 64568 377314 64568 0 pcpi_rs1\[15\]
rlabel metal3 376978 67256 376978 67256 0 pcpi_rs1\[16\]
rlabel metal5 380968 215190 380968 215190 0 pcpi_rs1\[17\]
rlabel metal3 377874 68600 377874 68600 0 pcpi_rs1\[18\]
rlabel metal3 377986 69272 377986 69272 0 pcpi_rs1\[19\]
rlabel metal2 379400 87472 379400 87472 0 pcpi_rs1\[1\]
rlabel metal3 380072 218582 380072 218582 0 pcpi_rs1\[20\]
rlabel metal3 377090 71288 377090 71288 0 pcpi_rs1\[21\]
rlabel metal3 380072 215166 380072 215166 0 pcpi_rs1\[22\]
rlabel metal3 377888 124488 377888 124488 0 pcpi_rs1\[23\]
rlabel metal4 380184 96488 380184 96488 0 pcpi_rs1\[24\]
rlabel metal3 379778 77336 379778 77336 0 pcpi_rs1\[25\]
rlabel metal4 373912 120383 373912 120383 0 pcpi_rs1\[26\]
rlabel metal3 424256 327656 424256 327656 0 pcpi_rs1\[27\]
rlabel metal3 378896 121016 378896 121016 0 pcpi_rs1\[28\]
rlabel metal3 377930 82712 377930 82712 0 pcpi_rs1\[29\]
rlabel metal3 380296 237454 380296 237454 0 pcpi_rs1\[2\]
rlabel metal3 373576 124376 373576 124376 0 pcpi_rs1\[30\]
rlabel metal3 420784 268744 420784 268744 0 pcpi_rs1\[31\]
rlabel metal2 377944 131264 377944 131264 0 pcpi_rs1\[3\]
rlabel metal2 379512 70728 379512 70728 0 pcpi_rs1\[4\]
rlabel metal3 376712 235144 376712 235144 0 pcpi_rs1\[5\]
rlabel metal3 384328 132160 384328 132160 0 pcpi_rs1\[6\]
rlabel metal3 380072 255766 380072 255766 0 pcpi_rs1\[7\]
rlabel metal3 378280 99176 378280 99176 0 pcpi_rs1\[8\]
rlabel metal3 379008 100856 379008 100856 0 pcpi_rs1\[9\]
rlabel metal3 378882 73976 378882 73976 0 pcpi_rs2\[0\]
rlabel metal3 378616 139384 378616 139384 0 pcpi_rs2\[10\]
rlabel metal5 378784 187830 378784 187830 0 pcpi_rs2\[11\]
rlabel metal3 378056 141064 378056 141064 0 pcpi_rs2\[12\]
rlabel metal3 378658 285096 378658 285096 0 pcpi_rs2\[13\]
rlabel metal3 373968 215096 373968 215096 0 pcpi_rs2\[14\]
rlabel metal3 379722 151144 379722 151144 0 pcpi_rs2\[15\]
rlabel metal4 380632 145043 380632 145043 0 pcpi_rs2\[16\]
rlabel metal3 377650 147112 377650 147112 0 pcpi_rs2\[17\]
rlabel metal3 380184 146314 380184 146314 0 pcpi_rs2\[18\]
rlabel metal3 378714 310632 378714 310632 0 pcpi_rs2\[19\]
rlabel metal3 378938 73304 378938 73304 0 pcpi_rs2\[1\]
rlabel metal5 380968 216810 380968 216810 0 pcpi_rs2\[20\]
rlabel metal3 379666 149128 379666 149128 0 pcpi_rs2\[21\]
rlabel metal3 379834 148456 379834 148456 0 pcpi_rs2\[22\]
rlabel metal3 378602 145768 378602 145768 0 pcpi_rs2\[23\]
rlabel metal4 406952 263816 406952 263816 0 pcpi_rs2\[24\]
rlabel metal3 380632 150766 380632 150766 0 pcpi_rs2\[25\]
rlabel metal4 379064 146552 379064 146552 0 pcpi_rs2\[26\]
rlabel metal4 408072 132160 408072 132160 0 pcpi_rs2\[27\]
rlabel metal3 423976 327768 423976 327768 0 pcpi_rs2\[28\]
rlabel metal3 378770 154504 378770 154504 0 pcpi_rs2\[29\]
rlabel metal3 378602 71960 378602 71960 0 pcpi_rs2\[2\]
rlabel metal4 375256 187273 375256 187273 0 pcpi_rs2\[30\]
rlabel metal2 426006 324408 426006 324408 0 pcpi_rs2\[31\]
rlabel metal3 378994 70616 378994 70616 0 pcpi_rs2\[3\]
rlabel metal3 377272 131040 377272 131040 0 pcpi_rs2\[4\]
rlabel metal3 378560 246680 378560 246680 0 pcpi_rs2\[5\]
rlabel metal4 403592 46872 403592 46872 0 pcpi_rs2\[6\]
rlabel metal4 403592 262767 403592 262767 0 pcpi_rs2\[7\]
rlabel metal3 378938 290472 378938 290472 0 pcpi_rs2\[8\]
rlabel metal3 378490 289800 378490 289800 0 pcpi_rs2\[9\]
rlabel metal4 377552 96570 377552 96570 0 pcpi_valid
rlabel metal2 56910 144872 56910 144872 0 ram_gwenb\[0\]
rlabel metal2 156856 152670 156856 152670 0 ram_gwenb\[1\]
rlabel metal2 53438 165032 53438 165032 0 ram_gwenb\[2\]
rlabel metal3 176064 278152 176064 278152 0 ram_gwenb\[3\]
rlabel metal2 88648 146734 88648 146734 0 ram_rdata\[0\]
rlabel metal2 181496 152726 181496 152726 0 ram_rdata\[10\]
rlabel metal2 172088 151886 172088 151886 0 ram_rdata\[11\]
rlabel metal3 169232 279720 169232 279720 0 ram_rdata\[12\]
rlabel metal2 128184 148582 128184 148582 0 ram_rdata\[13\]
rlabel metal2 125944 146734 125944 146734 0 ram_rdata\[14\]
rlabel metal2 118776 146510 118776 146510 0 ram_rdata\[15\]
rlabel metal2 21336 163786 21336 163786 0 ram_rdata\[16\]
rlabel metal2 26264 163842 26264 163842 0 ram_rdata\[17\]
rlabel metal2 28504 163058 28504 163058 0 ram_rdata\[18\]
rlabel metal4 172200 217224 172200 217224 0 ram_rdata\[19\]
rlabel metal2 83720 148526 83720 148526 0 ram_rdata\[1\]
rlabel metal2 72408 164458 72408 164458 0 ram_rdata\[20\]
rlabel metal2 81816 163674 81816 163674 0 ram_rdata\[21\]
rlabel metal3 201614 333032 201614 333032 0 ram_rdata\[22\]
rlabel metal2 91224 163954 91224 163954 0 ram_rdata\[23\]
rlabel metal2 121758 165592 121758 165592 0 ram_rdata\[24\]
rlabel metal4 126280 162857 126280 162857 0 ram_rdata\[25\]
rlabel metal4 210504 246400 210504 246400 0 ram_rdata\[26\]
rlabel metal2 137928 163506 137928 163506 0 ram_rdata\[27\]
rlabel metal2 172424 163786 172424 163786 0 ram_rdata\[28\]
rlabel metal2 181832 164458 181832 164458 0 ram_rdata\[29\]
rlabel metal2 81480 146398 81480 146398 0 ram_rdata\[2\]
rlabel metal2 184072 164794 184072 164794 0 ram_rdata\[30\]
rlabel metal2 191240 163954 191240 163954 0 ram_rdata\[31\]
rlabel metal3 200998 354312 200998 354312 0 ram_rdata\[3\]
rlabel metal4 54712 261016 54712 261016 0 ram_rdata\[4\]
rlabel metal2 28168 146790 28168 146790 0 ram_rdata\[5\]
rlabel metal2 25928 146846 25928 146846 0 ram_rdata\[6\]
rlabel metal4 2968 257647 2968 257647 0 ram_rdata\[7\]
rlabel metal2 188664 146734 188664 146734 0 ram_rdata\[8\]
rlabel metal3 183736 165424 183736 165424 0 ram_rdata\[9\]
rlabel metal2 89166 144872 89166 144872 0 ram_wenb\[0\]
rlabel metal3 202566 306152 202566 306152 0 ram_wenb\[10\]
rlabel metal2 171640 147630 171640 147630 0 ram_wenb\[11\]
rlabel metal3 169624 268408 169624 268408 0 ram_wenb\[12\]
rlabel metal2 208824 230888 208824 230888 0 ram_wenb\[13\]
rlabel metal2 126840 147798 126840 147798 0 ram_wenb\[14\]
rlabel metal2 118328 146454 118328 146454 0 ram_wenb\[15\]
rlabel metal4 20888 162857 20888 162857 0 ram_wenb\[16\]
rlabel metal4 27160 162767 27160 162767 0 ram_wenb\[17\]
rlabel metal2 27734 165032 27734 165032 0 ram_wenb\[18\]
rlabel metal2 38360 164514 38360 164514 0 ram_wenb\[19\]
rlabel metal2 82894 144872 82894 144872 0 ram_wenb\[1\]
rlabel metal2 71960 163730 71960 163730 0 ram_wenb\[20\]
rlabel metal2 82712 163842 82712 163842 0 ram_wenb\[21\]
rlabel metal2 83160 163786 83160 163786 0 ram_wenb\[22\]
rlabel metal2 91672 163898 91672 163898 0 ram_wenb\[23\]
rlabel metal2 120904 164570 120904 164570 0 ram_wenb\[24\]
rlabel metal2 127176 164402 127176 164402 0 ram_wenb\[25\]
rlabel metal5 162736 265050 162736 265050 0 ram_wenb\[26\]
rlabel metal2 138376 163898 138376 163898 0 ram_wenb\[27\]
rlabel metal2 171976 163730 171976 163730 0 ram_wenb\[28\]
rlabel metal2 182728 163618 182728 163618 0 ram_wenb\[29\]
rlabel metal2 82376 146398 82376 146398 0 ram_wenb\[2\]
rlabel metal2 183176 163898 183176 163898 0 ram_wenb\[30\]
rlabel metal2 191688 164738 191688 164738 0 ram_wenb\[31\]
rlabel metal3 201222 313992 201222 313992 0 ram_wenb\[3\]
rlabel metal2 38094 144872 38094 144872 0 ram_wenb\[4\]
rlabel metal2 27342 144872 27342 144872 0 ram_wenb\[5\]
rlabel metal2 26824 147686 26824 147686 0 ram_wenb\[6\]
rlabel metal2 18382 144872 18382 144872 0 ram_wenb\[7\]
rlabel metal2 189112 146902 189112 146902 0 ram_wenb\[8\]
rlabel metal3 200102 307272 200102 307272 0 ram_wenb\[9\]
rlabel metal2 45192 146398 45192 146398 0 reset
rlabel metal3 375424 52696 375424 52696 0 resetn
rlabel metal2 93016 330694 93016 330694 0 simpleuart_dat_re
rlabel metal3 117866 318920 117866 318920 0 simpleuart_dat_we
rlabel metal2 78232 344582 78232 344582 0 simpleuart_div_we\[0\]
rlabel metal3 66976 280728 66976 280728 0 simpleuart_div_we\[1\]
rlabel metal3 117642 357000 117642 357000 0 simpleuart_div_we\[2\]
rlabel metal3 118762 355880 118762 355880 0 simpleuart_div_we\[3\]
rlabel metal4 115864 315504 115864 315504 0 simpleuart_reg_dat_do\[0\]
rlabel metal3 117586 305480 117586 305480 0 simpleuart_reg_dat_do\[10\]
rlabel metal3 117922 304360 117922 304360 0 simpleuart_reg_dat_do\[11\]
rlabel metal3 119490 303240 119490 303240 0 simpleuart_reg_dat_do\[12\]
rlabel metal2 105112 330470 105112 330470 0 simpleuart_reg_dat_do\[13\]
rlabel metal2 100408 330582 100408 330582 0 simpleuart_reg_dat_do\[14\]
rlabel metal3 120120 299950 120120 299950 0 simpleuart_reg_dat_do\[15\]
rlabel metal3 118762 298760 118762 298760 0 simpleuart_reg_dat_do\[16\]
rlabel metal3 116074 297640 116074 297640 0 simpleuart_reg_dat_do\[17\]
rlabel metal2 102424 332430 102424 332430 0 simpleuart_reg_dat_do\[18\]
rlabel metal4 115864 297976 115864 297976 0 simpleuart_reg_dat_do\[19\]
rlabel metal4 117208 316960 117208 316960 0 simpleuart_reg_dat_do\[1\]
rlabel metal2 104440 330190 104440 330190 0 simpleuart_reg_dat_do\[20\]
rlabel metal3 116858 293160 116858 293160 0 simpleuart_reg_dat_do\[21\]
rlabel metal3 118650 292040 118650 292040 0 simpleuart_reg_dat_do\[22\]
rlabel metal3 117026 290920 117026 290920 0 simpleuart_reg_dat_do\[23\]
rlabel metal3 117418 289800 117418 289800 0 simpleuart_reg_dat_do\[24\]
rlabel metal3 117194 288680 117194 288680 0 simpleuart_reg_dat_do\[25\]
rlabel metal2 101080 332150 101080 332150 0 simpleuart_reg_dat_do\[26\]
rlabel metal2 101752 331366 101752 331366 0 simpleuart_reg_dat_do\[27\]
rlabel metal3 118650 285320 118650 285320 0 simpleuart_reg_dat_do\[28\]
rlabel metal3 117810 284200 117810 284200 0 simpleuart_reg_dat_do\[29\]
rlabel metal4 117320 317408 117320 317408 0 simpleuart_reg_dat_do\[2\]
rlabel metal3 118818 283080 118818 283080 0 simpleuart_reg_dat_do\[30\]
rlabel metal3 115584 282296 115584 282296 0 simpleuart_reg_dat_do\[31\]
rlabel metal3 118370 313320 118370 313320 0 simpleuart_reg_dat_do\[3\]
rlabel metal3 116634 312200 116634 312200 0 simpleuart_reg_dat_do\[4\]
rlabel metal3 116746 311080 116746 311080 0 simpleuart_reg_dat_do\[5\]
rlabel metal3 118034 309960 118034 309960 0 simpleuart_reg_dat_do\[6\]
rlabel metal2 95032 330974 95032 330974 0 simpleuart_reg_dat_do\[7\]
rlabel metal3 118370 307720 118370 307720 0 simpleuart_reg_dat_do\[8\]
rlabel metal3 118706 306600 118706 306600 0 simpleuart_reg_dat_do\[9\]
rlabel metal3 118482 280840 118482 280840 0 simpleuart_reg_dat_wait
rlabel metal3 89194 354760 89194 354760 0 simpleuart_reg_div_do\[0\]
rlabel metal3 57792 309176 57792 309176 0 simpleuart_reg_div_do\[10\]
rlabel metal3 58114 297528 58114 297528 0 simpleuart_reg_div_do\[11\]
rlabel metal2 70840 279930 70840 279930 0 simpleuart_reg_div_do\[12\]
rlabel metal2 72184 277298 72184 277298 0 simpleuart_reg_div_do\[13\]
rlabel metal3 118594 339080 118594 339080 0 simpleuart_reg_div_do\[14\]
rlabel metal3 118706 337960 118706 337960 0 simpleuart_reg_div_do\[15\]
rlabel metal3 118426 336840 118426 336840 0 simpleuart_reg_div_do\[16\]
rlabel metal3 116858 335720 116858 335720 0 simpleuart_reg_div_do\[17\]
rlabel metal3 117698 334600 117698 334600 0 simpleuart_reg_div_do\[18\]
rlabel metal3 118538 333480 118538 333480 0 simpleuart_reg_div_do\[19\]
rlabel metal3 89362 353640 89362 353640 0 simpleuart_reg_div_do\[1\]
rlabel metal2 119896 286244 119896 286244 0 simpleuart_reg_div_do\[20\]
rlabel metal2 93016 278082 93016 278082 0 simpleuart_reg_div_do\[21\]
rlabel metal2 94360 278474 94360 278474 0 simpleuart_reg_div_do\[22\]
rlabel metal2 97720 278418 97720 278418 0 simpleuart_reg_div_do\[23\]
rlabel metal3 111342 286104 111342 286104 0 simpleuart_reg_div_do\[24\]
rlabel metal3 112014 289464 112014 289464 0 simpleuart_reg_div_do\[25\]
rlabel metal3 111286 291480 111286 291480 0 simpleuart_reg_div_do\[26\]
rlabel metal3 112742 296184 112742 296184 0 simpleuart_reg_div_do\[27\]
rlabel metal3 111622 300216 111622 300216 0 simpleuart_reg_div_do\[28\]
rlabel metal3 112798 302904 112798 302904 0 simpleuart_reg_div_do\[29\]
rlabel metal3 118650 352520 118650 352520 0 simpleuart_reg_div_do\[2\]
rlabel metal3 112406 306264 112406 306264 0 simpleuart_reg_div_do\[30\]
rlabel metal3 117754 320040 117754 320040 0 simpleuart_reg_div_do\[31\]
rlabel metal4 91560 341600 91560 341600 0 simpleuart_reg_div_do\[3\]
rlabel metal3 118370 350280 118370 350280 0 simpleuart_reg_div_do\[4\]
rlabel metal2 76216 339542 76216 339542 0 simpleuart_reg_div_do\[5\]
rlabel metal3 58912 330792 58912 330792 0 simpleuart_reg_div_do\[6\]
rlabel metal3 58450 313656 58450 313656 0 simpleuart_reg_div_do\[7\]
rlabel metal3 58338 304248 58338 304248 0 simpleuart_reg_div_do\[8\]
rlabel metal3 60816 334376 60816 334376 0 simpleuart_reg_div_do\[9\]
rlabel metal2 28616 332374 28616 332374 0 spimem_rdata\[0\]
rlabel metal2 43400 330806 43400 330806 0 spimem_rdata\[10\]
rlabel metal2 44744 331534 44744 331534 0 spimem_rdata\[11\]
rlabel metal3 55678 319704 55678 319704 0 spimem_rdata\[12\]
rlabel metal3 57246 319032 57246 319032 0 spimem_rdata\[13\]
rlabel metal2 40040 331366 40040 331366 0 spimem_rdata\[14\]
rlabel metal4 51240 302568 51240 302568 0 spimem_rdata\[15\]
rlabel metal4 51464 302456 51464 302456 0 spimem_rdata\[16\]
rlabel metal2 41384 331478 41384 331478 0 spimem_rdata\[17\]
rlabel metal3 54936 321370 54936 321370 0 spimem_rdata\[18\]
rlabel metal1 52472 329336 52472 329336 0 spimem_rdata\[19\]
rlabel metal2 31304 330750 31304 330750 0 spimem_rdata\[1\]
rlabel metal3 54936 320250 54936 320250 0 spimem_rdata\[20\]
rlabel metal3 57694 315000 57694 315000 0 spimem_rdata\[21\]
rlabel metal2 35336 332206 35336 332206 0 spimem_rdata\[22\]
rlabel metal4 53032 301448 53032 301448 0 spimem_rdata\[23\]
rlabel metal3 118776 336112 118776 336112 0 spimem_rdata\[24\]
rlabel metal2 149128 278530 149128 278530 0 spimem_rdata\[25\]
rlabel metal3 54936 313530 54936 313530 0 spimem_rdata\[26\]
rlabel metal2 147784 274106 147784 274106 0 spimem_rdata\[27\]
rlabel metal2 147112 273378 147112 273378 0 spimem_rdata\[28\]
rlabel metal4 146440 281327 146440 281327 0 spimem_rdata\[29\]
rlabel metal3 54488 309386 54488 309386 0 spimem_rdata\[2\]
rlabel metal2 145768 278474 145768 278474 0 spimem_rdata\[30\]
rlabel metal2 145096 279314 145096 279314 0 spimem_rdata\[31\]
rlabel metal2 163912 275730 163912 275730 0 spimem_rdata\[3\]
rlabel metal2 163478 280504 163478 280504 0 spimem_rdata\[4\]
rlabel metal2 147896 275128 147896 275128 0 spimem_rdata\[5\]
rlabel metal2 161896 272650 161896 272650 0 spimem_rdata\[6\]
rlabel metal3 56686 308280 56686 308280 0 spimem_rdata\[7\]
rlabel metal2 30870 329896 30870 329896 0 spimem_rdata\[8\]
rlabel metal3 120568 279496 120568 279496 0 spimem_rdata\[9\]
rlabel metal3 4914 309624 4914 309624 0 spimem_ready
rlabel metal3 4858 306936 4858 306936 0 spimem_valid
rlabel metal3 56406 305592 56406 305592 0 spimemio_cfgreg_do\[0\]
rlabel metal4 68824 285169 68824 285169 0 spimemio_cfgreg_do\[10\]
rlabel metal3 56798 289464 56798 289464 0 spimemio_cfgreg_do\[11\]
rlabel metal4 5208 283431 5208 283431 0 spimemio_cfgreg_do\[12\]
rlabel metal3 5768 282506 5768 282506 0 spimemio_cfgreg_do\[13\]
rlabel metal2 119224 280672 119224 280672 0 spimemio_cfgreg_do\[14\]
rlabel metal3 5544 283962 5544 283962 0 spimemio_cfgreg_do\[15\]
rlabel metal2 16520 275954 16520 275954 0 spimemio_cfgreg_do\[16\]
rlabel metal3 75096 264824 75096 264824 0 spimemio_cfgreg_do\[17\]
rlabel metal2 18536 273938 18536 273938 0 spimemio_cfgreg_do\[18\]
rlabel metal2 21224 276402 21224 276402 0 spimemio_cfgreg_do\[19\]
rlabel metal4 141064 281867 141064 281867 0 spimemio_cfgreg_do\[1\]
rlabel metal3 4074 297528 4074 297528 0 spimemio_cfgreg_do\[20\]
rlabel metal2 14504 275114 14504 275114 0 spimemio_cfgreg_do\[21\]
rlabel metal2 22568 276346 22568 276346 0 spimemio_cfgreg_do\[22\]
rlabel metal3 56854 284760 56854 284760 0 spimemio_cfgreg_do\[23\]
rlabel metal2 125314 280056 125314 280056 0 spimemio_cfgreg_do\[24\]
rlabel metal2 124642 280056 124642 280056 0 spimemio_cfgreg_do\[25\]
rlabel metal2 123970 280056 123970 280056 0 spimemio_cfgreg_do\[26\]
rlabel metal2 123298 280056 123298 280056 0 spimemio_cfgreg_do\[27\]
rlabel metal2 122920 278026 122920 278026 0 spimemio_cfgreg_do\[28\]
rlabel metal2 122066 280056 122066 280056 0 spimemio_cfgreg_do\[29\]
rlabel metal3 54824 302106 54824 302106 0 spimemio_cfgreg_do\[2\]
rlabel metal4 5320 282603 5320 282603 0 spimemio_cfgreg_do\[30\]
rlabel metal2 120904 278418 120904 278418 0 spimemio_cfgreg_do\[31\]
rlabel metal4 139720 281777 139720 281777 0 spimemio_cfgreg_do\[3\]
rlabel metal2 139048 274218 139048 274218 0 spimemio_cfgreg_do\[4\]
rlabel metal2 138376 272594 138376 272594 0 spimemio_cfgreg_do\[5\]
rlabel metal4 127512 280280 127512 280280 0 spimemio_cfgreg_do\[6\]
rlabel metal3 5040 324632 5040 324632 0 spimemio_cfgreg_do\[7\]
rlabel metal2 46088 273434 46088 273434 0 spimemio_cfgreg_do\[8\]
rlabel metal2 46760 277466 46760 277466 0 spimemio_cfgreg_do\[9\]
rlabel metal2 144424 275898 144424 275898 0 spimemio_cfgreg_we\[0\]
rlabel metal2 49448 274162 49448 274162 0 spimemio_cfgreg_we\[1\]
rlabel metal2 143080 277746 143080 277746 0 spimemio_cfgreg_we\[2\]
rlabel metal2 27944 276010 27944 276010 0 spimemio_cfgreg_we\[3\]
rlabel metal2 512456 4368 512456 4368 0 user_irq[0]
rlabel metal2 513576 3794 513576 3794 0 user_irq[1]
rlabel metal2 515704 5040 515704 5040 0 user_irq[2]
rlabel metal2 44744 2562 44744 2562 0 wb_clk_i
rlabel metal2 46312 2618 46312 2618 0 wb_rst_i
rlabel metal2 15400 2758 15400 2758 0 wbs_ack_o
rlabel metal2 23128 392 23128 392 0 wbs_adr_i[0]
rlabel metal2 87752 1470 87752 1470 0 wbs_adr_i[10]
rlabel metal2 93464 1582 93464 1582 0 wbs_adr_i[11]
rlabel metal2 99064 2534 99064 2534 0 wbs_adr_i[12]
rlabel metal2 121576 4690 121576 4690 0 wbs_adr_i[13]
rlabel metal2 110600 2646 110600 2646 0 wbs_adr_i[14]
rlabel metal2 116312 1526 116312 1526 0 wbs_adr_i[15]
rlabel metal2 122024 1638 122024 1638 0 wbs_adr_i[16]
rlabel metal2 140392 4970 140392 4970 0 wbs_adr_i[17]
rlabel metal2 145096 3794 145096 3794 0 wbs_adr_i[18]
rlabel metal2 139160 2702 139160 2702 0 wbs_adr_i[19]
rlabel metal2 30632 2646 30632 2646 0 wbs_adr_i[1]
rlabel metal2 144872 2534 144872 2534 0 wbs_adr_i[20]
rlabel metal2 150584 2086 150584 2086 0 wbs_adr_i[21]
rlabel metal2 163912 4242 163912 4242 0 wbs_adr_i[22]
rlabel metal2 162008 2142 162008 2142 0 wbs_adr_i[23]
rlabel metal2 167720 1974 167720 1974 0 wbs_adr_i[24]
rlabel metal2 173432 1526 173432 1526 0 wbs_adr_i[25]
rlabel metal2 179144 1526 179144 1526 0 wbs_adr_i[26]
rlabel metal2 187432 3794 187432 3794 0 wbs_adr_i[27]
rlabel metal2 190568 462 190568 462 0 wbs_adr_i[28]
rlabel metal2 196280 1470 196280 1470 0 wbs_adr_i[29]
rlabel metal2 38248 1302 38248 1302 0 wbs_adr_i[2]
rlabel metal2 201768 2758 201768 2758 0 wbs_adr_i[30]
rlabel metal2 207480 462 207480 462 0 wbs_adr_i[31]
rlabel metal2 45864 2478 45864 2478 0 wbs_adr_i[3]
rlabel metal2 53480 2310 53480 2310 0 wbs_adr_i[4]
rlabel metal2 59192 1526 59192 1526 0 wbs_adr_i[5]
rlabel metal2 64904 2646 64904 2646 0 wbs_adr_i[6]
rlabel metal2 70504 2590 70504 2590 0 wbs_adr_i[7]
rlabel metal2 76328 2422 76328 2422 0 wbs_adr_i[8]
rlabel metal2 82040 2310 82040 2310 0 wbs_adr_i[9]
rlabel metal2 49448 3794 49448 3794 0 wbs_cyc_i
rlabel metal2 24920 1582 24920 1582 0 wbs_dat_i[0]
rlabel metal2 89656 2646 89656 2646 0 wbs_dat_i[10]
rlabel metal2 95368 2590 95368 2590 0 wbs_dat_i[11]
rlabel metal2 101080 2478 101080 2478 0 wbs_dat_i[12]
rlabel metal2 122696 5040 122696 5040 0 wbs_dat_i[13]
rlabel metal2 112504 2254 112504 2254 0 wbs_dat_i[14]
rlabel metal2 118216 1582 118216 1582 0 wbs_dat_i[15]
rlabel metal2 123928 2702 123928 2702 0 wbs_dat_i[16]
rlabel metal2 141960 4802 141960 4802 0 wbs_dat_i[17]
rlabel metal2 146664 3850 146664 3850 0 wbs_dat_i[18]
rlabel metal2 141064 2646 141064 2646 0 wbs_dat_i[19]
rlabel metal2 32536 1694 32536 1694 0 wbs_dat_i[1]
rlabel metal2 146776 2478 146776 2478 0 wbs_dat_i[20]
rlabel metal2 152488 2030 152488 2030 0 wbs_dat_i[21]
rlabel metal2 165480 4858 165480 4858 0 wbs_dat_i[22]
rlabel metal2 163912 462 163912 462 0 wbs_dat_i[23]
rlabel metal2 169624 1918 169624 1918 0 wbs_dat_i[24]
rlabel metal2 175336 1582 175336 1582 0 wbs_dat_i[25]
rlabel metal2 181048 1470 181048 1470 0 wbs_dat_i[26]
rlabel metal2 186760 1974 186760 1974 0 wbs_dat_i[27]
rlabel metal2 192472 462 192472 462 0 wbs_dat_i[28]
rlabel metal2 198184 2758 198184 2758 0 wbs_dat_i[29]
rlabel metal2 68264 4914 68264 4914 0 wbs_dat_i[2]
rlabel metal2 203672 2758 203672 2758 0 wbs_dat_i[30]
rlabel metal2 208376 2744 208376 2744 0 wbs_dat_i[31]
rlabel metal2 47768 2422 47768 2422 0 wbs_dat_i[3]
rlabel metal2 55384 1470 55384 1470 0 wbs_dat_i[4]
rlabel metal2 73080 4480 73080 4480 0 wbs_dat_i[5]
rlabel metal2 66808 1638 66808 1638 0 wbs_dat_i[6]
rlabel metal2 72520 2534 72520 2534 0 wbs_dat_i[7]
rlabel metal2 78232 2366 78232 2366 0 wbs_dat_i[8]
rlabel metal2 83944 2254 83944 2254 0 wbs_dat_i[9]
rlabel metal2 26824 1638 26824 1638 0 wbs_dat_o[0]
rlabel metal2 91560 1526 91560 1526 0 wbs_dat_o[10]
rlabel metal2 97272 1638 97272 1638 0 wbs_dat_o[11]
rlabel metal2 120008 4746 120008 4746 0 wbs_dat_o[12]
rlabel metal2 124712 4634 124712 4634 0 wbs_dat_o[13]
rlabel metal2 114408 1470 114408 1470 0 wbs_dat_o[14]
rlabel metal2 120120 2590 120120 2590 0 wbs_dat_o[15]
rlabel metal2 125832 2534 125832 2534 0 wbs_dat_o[16]
rlabel metal2 143528 4746 143528 4746 0 wbs_dat_o[17]
rlabel metal2 148232 3906 148232 3906 0 wbs_dat_o[18]
rlabel metal2 142968 2590 142968 2590 0 wbs_dat_o[19]
rlabel metal2 34440 1750 34440 1750 0 wbs_dat_o[1]
rlabel metal2 148680 2422 148680 2422 0 wbs_dat_o[20]
rlabel metal2 162344 4298 162344 4298 0 wbs_dat_o[21]
rlabel metal2 166376 5040 166376 5040 0 wbs_dat_o[22]
rlabel metal2 165816 2030 165816 2030 0 wbs_dat_o[23]
rlabel metal2 171528 1470 171528 1470 0 wbs_dat_o[24]
rlabel metal2 177240 1414 177240 1414 0 wbs_dat_o[25]
rlabel metal2 185864 3850 185864 3850 0 wbs_dat_o[26]
rlabel metal2 188664 1918 188664 1918 0 wbs_dat_o[27]
rlabel metal2 194376 462 194376 462 0 wbs_dat_o[28]
rlabel metal2 199976 2744 199976 2744 0 wbs_dat_o[29]
rlabel metal2 69832 3738 69832 3738 0 wbs_dat_o[2]
rlabel metal2 205576 462 205576 462 0 wbs_dat_o[30]
rlabel metal2 211288 1918 211288 1918 0 wbs_dat_o[31]
rlabel metal2 49672 1358 49672 1358 0 wbs_dat_o[3]
rlabel metal2 57288 1246 57288 1246 0 wbs_dat_o[4]
rlabel metal2 63000 1582 63000 1582 0 wbs_dat_o[5]
rlabel metal2 68712 2702 68712 2702 0 wbs_dat_o[6]
rlabel metal2 74424 2478 74424 2478 0 wbs_dat_o[7]
rlabel metal2 101192 4018 101192 4018 0 wbs_dat_o[8]
rlabel metal2 85848 2702 85848 2702 0 wbs_dat_o[9]
rlabel metal2 28728 2702 28728 2702 0 wbs_sel_i[0]
rlabel metal2 36344 1806 36344 1806 0 wbs_sel_i[1]
rlabel metal2 43960 2534 43960 2534 0 wbs_sel_i[2]
rlabel metal2 51576 2366 51576 2366 0 wbs_sel_i[3]
rlabel metal2 51016 3850 51016 3850 0 wbs_stb_i
rlabel metal2 21112 1918 21112 1918 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>

magic
tech gf180mcuD
magscale 1 5
timestamp 1702237551
<< obsm1 >>
rect 672 687 39312 38625
<< metal2 >>
rect 224 39600 280 40000
rect 560 39600 616 40000
rect 896 39600 952 40000
rect 1232 39600 1288 40000
rect 1568 39600 1624 40000
rect 1904 39600 1960 40000
rect 2240 39600 2296 40000
rect 2576 39600 2632 40000
rect 2912 39600 2968 40000
rect 3248 39600 3304 40000
rect 3584 39600 3640 40000
rect 3920 39600 3976 40000
rect 4256 39600 4312 40000
rect 4592 39600 4648 40000
rect 4928 39600 4984 40000
rect 5264 39600 5320 40000
rect 5600 39600 5656 40000
rect 5936 39600 5992 40000
rect 6272 39600 6328 40000
rect 6608 39600 6664 40000
rect 6944 39600 7000 40000
rect 7280 39600 7336 40000
rect 7616 39600 7672 40000
rect 7952 39600 8008 40000
rect 8288 39600 8344 40000
rect 8624 39600 8680 40000
rect 8960 39600 9016 40000
rect 9296 39600 9352 40000
rect 9632 39600 9688 40000
rect 9968 39600 10024 40000
rect 10304 39600 10360 40000
rect 10640 39600 10696 40000
rect 10976 39600 11032 40000
rect 11312 39600 11368 40000
rect 11648 39600 11704 40000
rect 11984 39600 12040 40000
rect 12320 39600 12376 40000
rect 12656 39600 12712 40000
rect 12992 39600 13048 40000
rect 13328 39600 13384 40000
rect 13664 39600 13720 40000
rect 14000 39600 14056 40000
rect 14336 39600 14392 40000
rect 14672 39600 14728 40000
rect 15008 39600 15064 40000
rect 15344 39600 15400 40000
rect 15680 39600 15736 40000
rect 16016 39600 16072 40000
rect 16352 39600 16408 40000
rect 16688 39600 16744 40000
rect 17024 39600 17080 40000
rect 17360 39600 17416 40000
rect 17696 39600 17752 40000
rect 18032 39600 18088 40000
rect 18368 39600 18424 40000
rect 18704 39600 18760 40000
rect 19040 39600 19096 40000
rect 19376 39600 19432 40000
rect 19712 39600 19768 40000
rect 20048 39600 20104 40000
rect 20384 39600 20440 40000
rect 20720 39600 20776 40000
rect 21056 39600 21112 40000
rect 21392 39600 21448 40000
rect 21728 39600 21784 40000
rect 22064 39600 22120 40000
rect 22400 39600 22456 40000
rect 22736 39600 22792 40000
rect 23072 39600 23128 40000
rect 23408 39600 23464 40000
rect 23744 39600 23800 40000
rect 24080 39600 24136 40000
rect 24416 39600 24472 40000
rect 24752 39600 24808 40000
rect 25088 39600 25144 40000
rect 25424 39600 25480 40000
rect 25760 39600 25816 40000
rect 26096 39600 26152 40000
rect 26432 39600 26488 40000
rect 26768 39600 26824 40000
rect 27104 39600 27160 40000
rect 27440 39600 27496 40000
rect 27776 39600 27832 40000
rect 28112 39600 28168 40000
rect 28448 39600 28504 40000
rect 28784 39600 28840 40000
rect 29120 39600 29176 40000
rect 29456 39600 29512 40000
rect 29792 39600 29848 40000
rect 30128 39600 30184 40000
rect 30464 39600 30520 40000
rect 30800 39600 30856 40000
rect 31136 39600 31192 40000
rect 31472 39600 31528 40000
rect 31808 39600 31864 40000
rect 32144 39600 32200 40000
rect 32480 39600 32536 40000
rect 32816 39600 32872 40000
rect 33152 39600 33208 40000
rect 33488 39600 33544 40000
rect 33824 39600 33880 40000
rect 34160 39600 34216 40000
rect 34496 39600 34552 40000
rect 34832 39600 34888 40000
rect 35168 39600 35224 40000
rect 35504 39600 35560 40000
rect 35840 39600 35896 40000
rect 36176 39600 36232 40000
rect 36512 39600 36568 40000
rect 36848 39600 36904 40000
rect 37184 39600 37240 40000
rect 37520 39600 37576 40000
rect 37856 39600 37912 40000
rect 38192 39600 38248 40000
rect 38528 39600 38584 40000
rect 38864 39600 38920 40000
rect 39200 39600 39256 40000
rect 39536 39600 39592 40000
rect 2464 0 2520 400
rect 2800 0 2856 400
rect 3136 0 3192 400
rect 3472 0 3528 400
rect 3808 0 3864 400
rect 4144 0 4200 400
rect 4480 0 4536 400
rect 4816 0 4872 400
rect 5152 0 5208 400
rect 5488 0 5544 400
rect 5824 0 5880 400
rect 6160 0 6216 400
rect 6496 0 6552 400
rect 6832 0 6888 400
rect 7168 0 7224 400
rect 7504 0 7560 400
rect 7840 0 7896 400
rect 8176 0 8232 400
rect 8512 0 8568 400
rect 8848 0 8904 400
rect 9184 0 9240 400
rect 9520 0 9576 400
rect 9856 0 9912 400
rect 10192 0 10248 400
rect 10528 0 10584 400
rect 10864 0 10920 400
rect 11200 0 11256 400
rect 11536 0 11592 400
rect 11872 0 11928 400
rect 12208 0 12264 400
rect 12544 0 12600 400
rect 12880 0 12936 400
rect 13216 0 13272 400
rect 13552 0 13608 400
rect 13888 0 13944 400
rect 14224 0 14280 400
rect 14560 0 14616 400
rect 14896 0 14952 400
rect 15232 0 15288 400
rect 15568 0 15624 400
rect 15904 0 15960 400
rect 16240 0 16296 400
rect 16576 0 16632 400
rect 16912 0 16968 400
rect 17248 0 17304 400
rect 17584 0 17640 400
rect 17920 0 17976 400
rect 18256 0 18312 400
rect 18592 0 18648 400
rect 18928 0 18984 400
rect 19264 0 19320 400
rect 19600 0 19656 400
rect 19936 0 19992 400
rect 20272 0 20328 400
rect 20608 0 20664 400
rect 20944 0 21000 400
rect 21280 0 21336 400
rect 21616 0 21672 400
rect 21952 0 22008 400
rect 22288 0 22344 400
rect 22624 0 22680 400
rect 22960 0 23016 400
rect 23296 0 23352 400
rect 23632 0 23688 400
rect 23968 0 24024 400
rect 24304 0 24360 400
rect 24640 0 24696 400
rect 24976 0 25032 400
rect 25312 0 25368 400
rect 25648 0 25704 400
rect 25984 0 26040 400
rect 26320 0 26376 400
rect 26656 0 26712 400
rect 26992 0 27048 400
rect 27328 0 27384 400
rect 27664 0 27720 400
rect 28000 0 28056 400
rect 28336 0 28392 400
rect 28672 0 28728 400
rect 29008 0 29064 400
rect 29344 0 29400 400
rect 29680 0 29736 400
rect 30016 0 30072 400
rect 30352 0 30408 400
rect 30688 0 30744 400
rect 31024 0 31080 400
rect 31360 0 31416 400
rect 31696 0 31752 400
rect 32032 0 32088 400
rect 32368 0 32424 400
rect 32704 0 32760 400
rect 33040 0 33096 400
rect 33376 0 33432 400
rect 33712 0 33768 400
rect 34048 0 34104 400
rect 34384 0 34440 400
rect 34720 0 34776 400
rect 35056 0 35112 400
rect 35392 0 35448 400
rect 35728 0 35784 400
rect 36064 0 36120 400
rect 36400 0 36456 400
rect 36736 0 36792 400
rect 37072 0 37128 400
rect 37408 0 37464 400
<< obsm2 >>
rect 854 39570 866 39600
rect 982 39570 1202 39600
rect 1318 39570 1538 39600
rect 1654 39570 1874 39600
rect 1990 39570 2210 39600
rect 2326 39570 2546 39600
rect 2662 39570 2882 39600
rect 2998 39570 3218 39600
rect 3334 39570 3554 39600
rect 3670 39570 3890 39600
rect 4006 39570 4226 39600
rect 4342 39570 4562 39600
rect 4678 39570 4898 39600
rect 5014 39570 5234 39600
rect 5350 39570 5570 39600
rect 5686 39570 5906 39600
rect 6022 39570 6242 39600
rect 6358 39570 6578 39600
rect 6694 39570 6914 39600
rect 7030 39570 7250 39600
rect 7366 39570 7586 39600
rect 7702 39570 7922 39600
rect 8038 39570 8258 39600
rect 8374 39570 8594 39600
rect 8710 39570 8930 39600
rect 9046 39570 9266 39600
rect 9382 39570 9602 39600
rect 9718 39570 9938 39600
rect 10054 39570 10274 39600
rect 10390 39570 10610 39600
rect 10726 39570 10946 39600
rect 11062 39570 11282 39600
rect 11398 39570 11618 39600
rect 11734 39570 11954 39600
rect 12070 39570 12290 39600
rect 12406 39570 12626 39600
rect 12742 39570 12962 39600
rect 13078 39570 13298 39600
rect 13414 39570 13634 39600
rect 13750 39570 13970 39600
rect 14086 39570 14306 39600
rect 14422 39570 14642 39600
rect 14758 39570 14978 39600
rect 15094 39570 15314 39600
rect 15430 39570 15650 39600
rect 15766 39570 15986 39600
rect 16102 39570 16322 39600
rect 16438 39570 16658 39600
rect 16774 39570 16994 39600
rect 17110 39570 17330 39600
rect 17446 39570 17666 39600
rect 17782 39570 18002 39600
rect 18118 39570 18338 39600
rect 18454 39570 18674 39600
rect 18790 39570 19010 39600
rect 19126 39570 19346 39600
rect 19462 39570 19682 39600
rect 19798 39570 20018 39600
rect 20134 39570 20354 39600
rect 20470 39570 20690 39600
rect 20806 39570 21026 39600
rect 21142 39570 21362 39600
rect 21478 39570 21698 39600
rect 21814 39570 22034 39600
rect 22150 39570 22370 39600
rect 22486 39570 22706 39600
rect 22822 39570 23042 39600
rect 23158 39570 23378 39600
rect 23494 39570 23714 39600
rect 23830 39570 24050 39600
rect 24166 39570 24386 39600
rect 24502 39570 24722 39600
rect 24838 39570 25058 39600
rect 25174 39570 25394 39600
rect 25510 39570 25730 39600
rect 25846 39570 26066 39600
rect 26182 39570 26402 39600
rect 26518 39570 26738 39600
rect 26854 39570 27074 39600
rect 27190 39570 27410 39600
rect 27526 39570 27746 39600
rect 27862 39570 28082 39600
rect 28198 39570 28418 39600
rect 28534 39570 28754 39600
rect 28870 39570 29090 39600
rect 29206 39570 29426 39600
rect 29542 39570 29762 39600
rect 29878 39570 30098 39600
rect 30214 39570 30434 39600
rect 30550 39570 30770 39600
rect 30886 39570 31106 39600
rect 31222 39570 31442 39600
rect 31558 39570 31778 39600
rect 31894 39570 32114 39600
rect 32230 39570 32450 39600
rect 32566 39570 32786 39600
rect 32902 39570 33122 39600
rect 33238 39570 33458 39600
rect 33574 39570 33794 39600
rect 33910 39570 34130 39600
rect 34246 39570 34466 39600
rect 34582 39570 34802 39600
rect 34918 39570 35138 39600
rect 35254 39570 35474 39600
rect 35590 39570 35810 39600
rect 35926 39570 36146 39600
rect 36262 39570 36482 39600
rect 36598 39570 36818 39600
rect 36934 39570 37154 39600
rect 37270 39570 37490 39600
rect 37606 39570 37826 39600
rect 37942 39570 38162 39600
rect 38278 39570 38498 39600
rect 38614 39570 38834 39600
rect 38950 39570 39170 39600
rect 39286 39570 39506 39600
rect 854 430 39578 39570
rect 854 350 2434 430
rect 2550 350 2770 430
rect 2886 350 3106 430
rect 3222 350 3442 430
rect 3558 350 3778 430
rect 3894 350 4114 430
rect 4230 350 4450 430
rect 4566 350 4786 430
rect 4902 350 5122 430
rect 5238 350 5458 430
rect 5574 350 5794 430
rect 5910 350 6130 430
rect 6246 350 6466 430
rect 6582 350 6802 430
rect 6918 350 7138 430
rect 7254 350 7474 430
rect 7590 350 7810 430
rect 7926 350 8146 430
rect 8262 350 8482 430
rect 8598 350 8818 430
rect 8934 350 9154 430
rect 9270 350 9490 430
rect 9606 350 9826 430
rect 9942 350 10162 430
rect 10278 350 10498 430
rect 10614 350 10834 430
rect 10950 350 11170 430
rect 11286 350 11506 430
rect 11622 350 11842 430
rect 11958 350 12178 430
rect 12294 350 12514 430
rect 12630 350 12850 430
rect 12966 350 13186 430
rect 13302 350 13522 430
rect 13638 350 13858 430
rect 13974 350 14194 430
rect 14310 350 14530 430
rect 14646 350 14866 430
rect 14982 350 15202 430
rect 15318 350 15538 430
rect 15654 350 15874 430
rect 15990 350 16210 430
rect 16326 350 16546 430
rect 16662 350 16882 430
rect 16998 350 17218 430
rect 17334 350 17554 430
rect 17670 350 17890 430
rect 18006 350 18226 430
rect 18342 350 18562 430
rect 18678 350 18898 430
rect 19014 350 19234 430
rect 19350 350 19570 430
rect 19686 350 19906 430
rect 20022 350 20242 430
rect 20358 350 20578 430
rect 20694 350 20914 430
rect 21030 350 21250 430
rect 21366 350 21586 430
rect 21702 350 21922 430
rect 22038 350 22258 430
rect 22374 350 22594 430
rect 22710 350 22930 430
rect 23046 350 23266 430
rect 23382 350 23602 430
rect 23718 350 23938 430
rect 24054 350 24274 430
rect 24390 350 24610 430
rect 24726 350 24946 430
rect 25062 350 25282 430
rect 25398 350 25618 430
rect 25734 350 25954 430
rect 26070 350 26290 430
rect 26406 350 26626 430
rect 26742 350 26962 430
rect 27078 350 27298 430
rect 27414 350 27634 430
rect 27750 350 27970 430
rect 28086 350 28306 430
rect 28422 350 28642 430
rect 28758 350 28978 430
rect 29094 350 29314 430
rect 29430 350 29650 430
rect 29766 350 29986 430
rect 30102 350 30322 430
rect 30438 350 30658 430
rect 30774 350 30994 430
rect 31110 350 31330 430
rect 31446 350 31666 430
rect 31782 350 32002 430
rect 32118 350 32338 430
rect 32454 350 32674 430
rect 32790 350 33010 430
rect 33126 350 33346 430
rect 33462 350 33682 430
rect 33798 350 34018 430
rect 34134 350 34354 430
rect 34470 350 34690 430
rect 34806 350 35026 430
rect 35142 350 35362 430
rect 35478 350 35698 430
rect 35814 350 36034 430
rect 36150 350 36370 430
rect 36486 350 36706 430
rect 36822 350 37042 430
rect 37158 350 37378 430
rect 37494 350 39578 430
<< metal3 >>
rect 39600 39536 40000 39592
rect 39600 38976 40000 39032
rect 0 38640 400 38696
rect 39600 38416 40000 38472
rect 0 38080 400 38136
rect 39600 37856 40000 37912
rect 0 37520 400 37576
rect 39600 37296 40000 37352
rect 0 36960 400 37016
rect 39600 36736 40000 36792
rect 0 36400 400 36456
rect 39600 36176 40000 36232
rect 0 35840 400 35896
rect 39600 35616 40000 35672
rect 0 35280 400 35336
rect 39600 35056 40000 35112
rect 0 34720 400 34776
rect 39600 34496 40000 34552
rect 0 34160 400 34216
rect 39600 33936 40000 33992
rect 0 33600 400 33656
rect 39600 33376 40000 33432
rect 0 33040 400 33096
rect 39600 32816 40000 32872
rect 0 32480 400 32536
rect 39600 32256 40000 32312
rect 0 31920 400 31976
rect 39600 31696 40000 31752
rect 0 31360 400 31416
rect 39600 31136 40000 31192
rect 0 30800 400 30856
rect 39600 30576 40000 30632
rect 0 30240 400 30296
rect 39600 30016 40000 30072
rect 0 29680 400 29736
rect 39600 29456 40000 29512
rect 0 29120 400 29176
rect 39600 28896 40000 28952
rect 0 28560 400 28616
rect 39600 28336 40000 28392
rect 0 28000 400 28056
rect 39600 27776 40000 27832
rect 0 27440 400 27496
rect 39600 27216 40000 27272
rect 0 26880 400 26936
rect 39600 26656 40000 26712
rect 0 26320 400 26376
rect 39600 26096 40000 26152
rect 0 25760 400 25816
rect 39600 25536 40000 25592
rect 0 25200 400 25256
rect 39600 24976 40000 25032
rect 0 24640 400 24696
rect 39600 24416 40000 24472
rect 0 24080 400 24136
rect 39600 23856 40000 23912
rect 0 23520 400 23576
rect 39600 23296 40000 23352
rect 0 22960 400 23016
rect 39600 22736 40000 22792
rect 0 22400 400 22456
rect 39600 22176 40000 22232
rect 0 21840 400 21896
rect 39600 21616 40000 21672
rect 0 21280 400 21336
rect 39600 21056 40000 21112
rect 0 20720 400 20776
rect 39600 20496 40000 20552
rect 0 20160 400 20216
rect 39600 19936 40000 19992
rect 0 19600 400 19656
rect 39600 19376 40000 19432
rect 0 19040 400 19096
rect 39600 18816 40000 18872
rect 0 18480 400 18536
rect 39600 18256 40000 18312
rect 0 17920 400 17976
rect 39600 17696 40000 17752
rect 0 17360 400 17416
rect 39600 17136 40000 17192
rect 0 16800 400 16856
rect 39600 16576 40000 16632
rect 0 16240 400 16296
rect 39600 16016 40000 16072
rect 0 15680 400 15736
rect 39600 15456 40000 15512
rect 0 15120 400 15176
rect 39600 14896 40000 14952
rect 0 14560 400 14616
rect 39600 14336 40000 14392
rect 0 14000 400 14056
rect 39600 13776 40000 13832
rect 0 13440 400 13496
rect 39600 13216 40000 13272
rect 0 12880 400 12936
rect 39600 12656 40000 12712
rect 0 12320 400 12376
rect 39600 12096 40000 12152
rect 0 11760 400 11816
rect 39600 11536 40000 11592
rect 0 11200 400 11256
rect 39600 10976 40000 11032
rect 0 10640 400 10696
rect 39600 10416 40000 10472
rect 0 10080 400 10136
rect 39600 9856 40000 9912
rect 0 9520 400 9576
rect 39600 9296 40000 9352
rect 0 8960 400 9016
rect 39600 8736 40000 8792
rect 0 8400 400 8456
rect 39600 8176 40000 8232
rect 0 7840 400 7896
rect 39600 7616 40000 7672
rect 0 7280 400 7336
rect 39600 7056 40000 7112
rect 0 6720 400 6776
rect 39600 6496 40000 6552
rect 0 6160 400 6216
rect 39600 5936 40000 5992
rect 0 5600 400 5656
rect 39600 5376 40000 5432
rect 0 5040 400 5096
rect 39600 4816 40000 4872
rect 0 4480 400 4536
rect 39600 4256 40000 4312
rect 0 3920 400 3976
rect 39600 3696 40000 3752
rect 0 3360 400 3416
rect 39600 3136 40000 3192
rect 0 2800 400 2856
rect 39600 2576 40000 2632
rect 0 2240 400 2296
rect 39600 2016 40000 2072
rect 0 1680 400 1736
rect 39600 1456 40000 1512
rect 0 1120 400 1176
rect 39600 896 40000 952
rect 39600 336 40000 392
<< obsm3 >>
rect 400 39506 39570 39578
rect 400 39062 39600 39506
rect 400 38946 39570 39062
rect 400 38726 39600 38946
rect 430 38610 39600 38726
rect 400 38502 39600 38610
rect 400 38386 39570 38502
rect 400 38166 39600 38386
rect 430 38050 39600 38166
rect 400 37942 39600 38050
rect 400 37826 39570 37942
rect 400 37606 39600 37826
rect 430 37490 39600 37606
rect 400 37382 39600 37490
rect 400 37266 39570 37382
rect 400 37046 39600 37266
rect 430 36930 39600 37046
rect 400 36822 39600 36930
rect 400 36706 39570 36822
rect 400 36486 39600 36706
rect 430 36370 39600 36486
rect 400 36262 39600 36370
rect 400 36146 39570 36262
rect 400 35926 39600 36146
rect 430 35810 39600 35926
rect 400 35702 39600 35810
rect 400 35586 39570 35702
rect 400 35366 39600 35586
rect 430 35250 39600 35366
rect 400 35142 39600 35250
rect 400 35026 39570 35142
rect 400 34806 39600 35026
rect 430 34690 39600 34806
rect 400 34582 39600 34690
rect 400 34466 39570 34582
rect 400 34246 39600 34466
rect 430 34130 39600 34246
rect 400 34022 39600 34130
rect 400 33906 39570 34022
rect 400 33686 39600 33906
rect 430 33570 39600 33686
rect 400 33462 39600 33570
rect 400 33346 39570 33462
rect 400 33126 39600 33346
rect 430 33010 39600 33126
rect 400 32902 39600 33010
rect 400 32786 39570 32902
rect 400 32566 39600 32786
rect 430 32450 39600 32566
rect 400 32342 39600 32450
rect 400 32226 39570 32342
rect 400 32006 39600 32226
rect 430 31890 39600 32006
rect 400 31782 39600 31890
rect 400 31666 39570 31782
rect 400 31446 39600 31666
rect 430 31330 39600 31446
rect 400 31222 39600 31330
rect 400 31106 39570 31222
rect 400 30886 39600 31106
rect 430 30770 39600 30886
rect 400 30662 39600 30770
rect 400 30546 39570 30662
rect 400 30326 39600 30546
rect 430 30210 39600 30326
rect 400 30102 39600 30210
rect 400 29986 39570 30102
rect 400 29766 39600 29986
rect 430 29650 39600 29766
rect 400 29542 39600 29650
rect 400 29426 39570 29542
rect 400 29206 39600 29426
rect 430 29090 39600 29206
rect 400 28982 39600 29090
rect 400 28866 39570 28982
rect 400 28646 39600 28866
rect 430 28530 39600 28646
rect 400 28422 39600 28530
rect 400 28306 39570 28422
rect 400 28086 39600 28306
rect 430 27970 39600 28086
rect 400 27862 39600 27970
rect 400 27746 39570 27862
rect 400 27526 39600 27746
rect 430 27410 39600 27526
rect 400 27302 39600 27410
rect 400 27186 39570 27302
rect 400 26966 39600 27186
rect 430 26850 39600 26966
rect 400 26742 39600 26850
rect 400 26626 39570 26742
rect 400 26406 39600 26626
rect 430 26290 39600 26406
rect 400 26182 39600 26290
rect 400 26066 39570 26182
rect 400 25846 39600 26066
rect 430 25730 39600 25846
rect 400 25622 39600 25730
rect 400 25506 39570 25622
rect 400 25286 39600 25506
rect 430 25170 39600 25286
rect 400 25062 39600 25170
rect 400 24946 39570 25062
rect 400 24726 39600 24946
rect 430 24610 39600 24726
rect 400 24502 39600 24610
rect 400 24386 39570 24502
rect 400 24166 39600 24386
rect 430 24050 39600 24166
rect 400 23942 39600 24050
rect 400 23826 39570 23942
rect 400 23606 39600 23826
rect 430 23490 39600 23606
rect 400 23382 39600 23490
rect 400 23266 39570 23382
rect 400 23046 39600 23266
rect 430 22930 39600 23046
rect 400 22822 39600 22930
rect 400 22706 39570 22822
rect 400 22486 39600 22706
rect 430 22370 39600 22486
rect 400 22262 39600 22370
rect 400 22146 39570 22262
rect 400 21926 39600 22146
rect 430 21810 39600 21926
rect 400 21702 39600 21810
rect 400 21586 39570 21702
rect 400 21366 39600 21586
rect 430 21250 39600 21366
rect 400 21142 39600 21250
rect 400 21026 39570 21142
rect 400 20806 39600 21026
rect 430 20690 39600 20806
rect 400 20582 39600 20690
rect 400 20466 39570 20582
rect 400 20246 39600 20466
rect 430 20130 39600 20246
rect 400 20022 39600 20130
rect 400 19906 39570 20022
rect 400 19686 39600 19906
rect 430 19570 39600 19686
rect 400 19462 39600 19570
rect 400 19346 39570 19462
rect 400 19126 39600 19346
rect 430 19010 39600 19126
rect 400 18902 39600 19010
rect 400 18786 39570 18902
rect 400 18566 39600 18786
rect 430 18450 39600 18566
rect 400 18342 39600 18450
rect 400 18226 39570 18342
rect 400 18006 39600 18226
rect 430 17890 39600 18006
rect 400 17782 39600 17890
rect 400 17666 39570 17782
rect 400 17446 39600 17666
rect 430 17330 39600 17446
rect 400 17222 39600 17330
rect 400 17106 39570 17222
rect 400 16886 39600 17106
rect 430 16770 39600 16886
rect 400 16662 39600 16770
rect 400 16546 39570 16662
rect 400 16326 39600 16546
rect 430 16210 39600 16326
rect 400 16102 39600 16210
rect 400 15986 39570 16102
rect 400 15766 39600 15986
rect 430 15650 39600 15766
rect 400 15542 39600 15650
rect 400 15426 39570 15542
rect 400 15206 39600 15426
rect 430 15090 39600 15206
rect 400 14982 39600 15090
rect 400 14866 39570 14982
rect 400 14646 39600 14866
rect 430 14530 39600 14646
rect 400 14422 39600 14530
rect 400 14306 39570 14422
rect 400 14086 39600 14306
rect 430 13970 39600 14086
rect 400 13862 39600 13970
rect 400 13746 39570 13862
rect 400 13526 39600 13746
rect 430 13410 39600 13526
rect 400 13302 39600 13410
rect 400 13186 39570 13302
rect 400 12966 39600 13186
rect 430 12850 39600 12966
rect 400 12742 39600 12850
rect 400 12626 39570 12742
rect 400 12406 39600 12626
rect 430 12290 39600 12406
rect 400 12182 39600 12290
rect 400 12066 39570 12182
rect 400 11846 39600 12066
rect 430 11730 39600 11846
rect 400 11622 39600 11730
rect 400 11506 39570 11622
rect 400 11286 39600 11506
rect 430 11170 39600 11286
rect 400 11062 39600 11170
rect 400 10946 39570 11062
rect 400 10726 39600 10946
rect 430 10610 39600 10726
rect 400 10502 39600 10610
rect 400 10386 39570 10502
rect 400 10166 39600 10386
rect 430 10050 39600 10166
rect 400 9942 39600 10050
rect 400 9826 39570 9942
rect 400 9606 39600 9826
rect 430 9490 39600 9606
rect 400 9382 39600 9490
rect 400 9266 39570 9382
rect 400 9046 39600 9266
rect 430 8930 39600 9046
rect 400 8822 39600 8930
rect 400 8706 39570 8822
rect 400 8486 39600 8706
rect 430 8370 39600 8486
rect 400 8262 39600 8370
rect 400 8146 39570 8262
rect 400 7926 39600 8146
rect 430 7810 39600 7926
rect 400 7702 39600 7810
rect 400 7586 39570 7702
rect 400 7366 39600 7586
rect 430 7250 39600 7366
rect 400 7142 39600 7250
rect 400 7026 39570 7142
rect 400 6806 39600 7026
rect 430 6690 39600 6806
rect 400 6582 39600 6690
rect 400 6466 39570 6582
rect 400 6246 39600 6466
rect 430 6130 39600 6246
rect 400 6022 39600 6130
rect 400 5906 39570 6022
rect 400 5686 39600 5906
rect 430 5570 39600 5686
rect 400 5462 39600 5570
rect 400 5346 39570 5462
rect 400 5126 39600 5346
rect 430 5010 39600 5126
rect 400 4902 39600 5010
rect 400 4786 39570 4902
rect 400 4566 39600 4786
rect 430 4450 39600 4566
rect 400 4342 39600 4450
rect 400 4226 39570 4342
rect 400 4006 39600 4226
rect 430 3890 39600 4006
rect 400 3782 39600 3890
rect 400 3666 39570 3782
rect 400 3446 39600 3666
rect 430 3330 39600 3446
rect 400 3222 39600 3330
rect 400 3106 39570 3222
rect 400 2886 39600 3106
rect 430 2770 39600 2886
rect 400 2662 39600 2770
rect 400 2546 39570 2662
rect 400 2326 39600 2546
rect 430 2210 39600 2326
rect 400 2102 39600 2210
rect 400 1986 39570 2102
rect 400 1766 39600 1986
rect 430 1650 39600 1766
rect 400 1542 39600 1650
rect 400 1426 39570 1542
rect 400 1206 39600 1426
rect 430 1090 39600 1206
rect 400 982 39600 1090
rect 400 866 39570 982
rect 400 422 39600 866
rect 400 350 39570 422
<< metal4 >>
rect 2224 1538 2384 38446
rect 9904 1538 10064 38446
rect 17584 1538 17744 38446
rect 25264 1538 25424 38446
rect 32944 1538 33104 38446
<< obsm4 >>
rect 3598 1577 9874 38295
rect 10094 1577 17554 38295
rect 17774 1577 25234 38295
rect 25454 1577 32914 38295
rect 33134 1577 38962 38295
<< labels >>
rlabel metal2 s 37072 0 37128 400 6 clk
port 1 nsew signal input
rlabel metal2 s 224 39600 280 40000 6 gpio_in[0]
port 2 nsew signal input
rlabel metal2 s 3584 39600 3640 40000 6 gpio_in[10]
port 3 nsew signal input
rlabel metal2 s 3920 39600 3976 40000 6 gpio_in[11]
port 4 nsew signal input
rlabel metal2 s 4256 39600 4312 40000 6 gpio_in[12]
port 5 nsew signal input
rlabel metal2 s 4592 39600 4648 40000 6 gpio_in[13]
port 6 nsew signal input
rlabel metal2 s 4928 39600 4984 40000 6 gpio_in[14]
port 7 nsew signal input
rlabel metal2 s 5264 39600 5320 40000 6 gpio_in[15]
port 8 nsew signal input
rlabel metal2 s 560 39600 616 40000 6 gpio_in[1]
port 9 nsew signal input
rlabel metal2 s 896 39600 952 40000 6 gpio_in[2]
port 10 nsew signal input
rlabel metal2 s 1232 39600 1288 40000 6 gpio_in[3]
port 11 nsew signal input
rlabel metal2 s 1568 39600 1624 40000 6 gpio_in[4]
port 12 nsew signal input
rlabel metal2 s 1904 39600 1960 40000 6 gpio_in[5]
port 13 nsew signal input
rlabel metal2 s 2240 39600 2296 40000 6 gpio_in[6]
port 14 nsew signal input
rlabel metal2 s 2576 39600 2632 40000 6 gpio_in[7]
port 15 nsew signal input
rlabel metal2 s 2912 39600 2968 40000 6 gpio_in[8]
port 16 nsew signal input
rlabel metal2 s 3248 39600 3304 40000 6 gpio_in[9]
port 17 nsew signal input
rlabel metal2 s 10976 39600 11032 40000 6 gpio_oeb[0]
port 18 nsew signal output
rlabel metal2 s 14336 39600 14392 40000 6 gpio_oeb[10]
port 19 nsew signal output
rlabel metal2 s 14672 39600 14728 40000 6 gpio_oeb[11]
port 20 nsew signal output
rlabel metal2 s 15008 39600 15064 40000 6 gpio_oeb[12]
port 21 nsew signal output
rlabel metal2 s 15344 39600 15400 40000 6 gpio_oeb[13]
port 22 nsew signal output
rlabel metal2 s 15680 39600 15736 40000 6 gpio_oeb[14]
port 23 nsew signal output
rlabel metal2 s 16016 39600 16072 40000 6 gpio_oeb[15]
port 24 nsew signal output
rlabel metal2 s 11312 39600 11368 40000 6 gpio_oeb[1]
port 25 nsew signal output
rlabel metal2 s 11648 39600 11704 40000 6 gpio_oeb[2]
port 26 nsew signal output
rlabel metal2 s 11984 39600 12040 40000 6 gpio_oeb[3]
port 27 nsew signal output
rlabel metal2 s 12320 39600 12376 40000 6 gpio_oeb[4]
port 28 nsew signal output
rlabel metal2 s 12656 39600 12712 40000 6 gpio_oeb[5]
port 29 nsew signal output
rlabel metal2 s 12992 39600 13048 40000 6 gpio_oeb[6]
port 30 nsew signal output
rlabel metal2 s 13328 39600 13384 40000 6 gpio_oeb[7]
port 31 nsew signal output
rlabel metal2 s 13664 39600 13720 40000 6 gpio_oeb[8]
port 32 nsew signal output
rlabel metal2 s 14000 39600 14056 40000 6 gpio_oeb[9]
port 33 nsew signal output
rlabel metal2 s 5600 39600 5656 40000 6 gpio_out[0]
port 34 nsew signal output
rlabel metal2 s 8960 39600 9016 40000 6 gpio_out[10]
port 35 nsew signal output
rlabel metal2 s 9296 39600 9352 40000 6 gpio_out[11]
port 36 nsew signal output
rlabel metal2 s 9632 39600 9688 40000 6 gpio_out[12]
port 37 nsew signal output
rlabel metal2 s 9968 39600 10024 40000 6 gpio_out[13]
port 38 nsew signal output
rlabel metal2 s 10304 39600 10360 40000 6 gpio_out[14]
port 39 nsew signal output
rlabel metal2 s 10640 39600 10696 40000 6 gpio_out[15]
port 40 nsew signal output
rlabel metal2 s 5936 39600 5992 40000 6 gpio_out[1]
port 41 nsew signal output
rlabel metal2 s 6272 39600 6328 40000 6 gpio_out[2]
port 42 nsew signal output
rlabel metal2 s 6608 39600 6664 40000 6 gpio_out[3]
port 43 nsew signal output
rlabel metal2 s 6944 39600 7000 40000 6 gpio_out[4]
port 44 nsew signal output
rlabel metal2 s 7280 39600 7336 40000 6 gpio_out[5]
port 45 nsew signal output
rlabel metal2 s 7616 39600 7672 40000 6 gpio_out[6]
port 46 nsew signal output
rlabel metal2 s 7952 39600 8008 40000 6 gpio_out[7]
port 47 nsew signal output
rlabel metal2 s 8288 39600 8344 40000 6 gpio_out[8]
port 48 nsew signal output
rlabel metal2 s 8624 39600 8680 40000 6 gpio_out[9]
port 49 nsew signal output
rlabel metal2 s 13216 0 13272 400 6 mem_addr[0]
port 50 nsew signal input
rlabel metal2 s 16576 0 16632 400 6 mem_addr[10]
port 51 nsew signal input
rlabel metal2 s 16912 0 16968 400 6 mem_addr[11]
port 52 nsew signal input
rlabel metal2 s 17248 0 17304 400 6 mem_addr[12]
port 53 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 mem_addr[13]
port 54 nsew signal input
rlabel metal2 s 17920 0 17976 400 6 mem_addr[14]
port 55 nsew signal input
rlabel metal2 s 18256 0 18312 400 6 mem_addr[15]
port 56 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 mem_addr[16]
port 57 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 mem_addr[17]
port 58 nsew signal input
rlabel metal2 s 19264 0 19320 400 6 mem_addr[18]
port 59 nsew signal input
rlabel metal2 s 19600 0 19656 400 6 mem_addr[19]
port 60 nsew signal input
rlabel metal2 s 13552 0 13608 400 6 mem_addr[1]
port 61 nsew signal input
rlabel metal2 s 19936 0 19992 400 6 mem_addr[20]
port 62 nsew signal input
rlabel metal2 s 20272 0 20328 400 6 mem_addr[21]
port 63 nsew signal input
rlabel metal2 s 20608 0 20664 400 6 mem_addr[22]
port 64 nsew signal input
rlabel metal2 s 20944 0 21000 400 6 mem_addr[23]
port 65 nsew signal input
rlabel metal2 s 21280 0 21336 400 6 mem_addr[24]
port 66 nsew signal input
rlabel metal2 s 21616 0 21672 400 6 mem_addr[25]
port 67 nsew signal input
rlabel metal2 s 21952 0 22008 400 6 mem_addr[26]
port 68 nsew signal input
rlabel metal2 s 22288 0 22344 400 6 mem_addr[27]
port 69 nsew signal input
rlabel metal2 s 22624 0 22680 400 6 mem_addr[28]
port 70 nsew signal input
rlabel metal2 s 22960 0 23016 400 6 mem_addr[29]
port 71 nsew signal input
rlabel metal2 s 13888 0 13944 400 6 mem_addr[2]
port 72 nsew signal input
rlabel metal2 s 23296 0 23352 400 6 mem_addr[30]
port 73 nsew signal input
rlabel metal2 s 23632 0 23688 400 6 mem_addr[31]
port 74 nsew signal input
rlabel metal2 s 14224 0 14280 400 6 mem_addr[3]
port 75 nsew signal input
rlabel metal2 s 14560 0 14616 400 6 mem_addr[4]
port 76 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 mem_addr[5]
port 77 nsew signal input
rlabel metal2 s 15232 0 15288 400 6 mem_addr[6]
port 78 nsew signal input
rlabel metal2 s 15568 0 15624 400 6 mem_addr[7]
port 79 nsew signal input
rlabel metal2 s 15904 0 15960 400 6 mem_addr[8]
port 80 nsew signal input
rlabel metal2 s 16240 0 16296 400 6 mem_addr[9]
port 81 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 mem_instr
port 82 nsew signal input
rlabel metal2 s 26320 0 26376 400 6 mem_rdata[0]
port 83 nsew signal output
rlabel metal2 s 29680 0 29736 400 6 mem_rdata[10]
port 84 nsew signal output
rlabel metal2 s 30016 0 30072 400 6 mem_rdata[11]
port 85 nsew signal output
rlabel metal2 s 30352 0 30408 400 6 mem_rdata[12]
port 86 nsew signal output
rlabel metal2 s 30688 0 30744 400 6 mem_rdata[13]
port 87 nsew signal output
rlabel metal2 s 31024 0 31080 400 6 mem_rdata[14]
port 88 nsew signal output
rlabel metal2 s 31360 0 31416 400 6 mem_rdata[15]
port 89 nsew signal output
rlabel metal2 s 31696 0 31752 400 6 mem_rdata[16]
port 90 nsew signal output
rlabel metal2 s 32032 0 32088 400 6 mem_rdata[17]
port 91 nsew signal output
rlabel metal2 s 32368 0 32424 400 6 mem_rdata[18]
port 92 nsew signal output
rlabel metal2 s 32704 0 32760 400 6 mem_rdata[19]
port 93 nsew signal output
rlabel metal2 s 26656 0 26712 400 6 mem_rdata[1]
port 94 nsew signal output
rlabel metal2 s 33040 0 33096 400 6 mem_rdata[20]
port 95 nsew signal output
rlabel metal2 s 33376 0 33432 400 6 mem_rdata[21]
port 96 nsew signal output
rlabel metal2 s 33712 0 33768 400 6 mem_rdata[22]
port 97 nsew signal output
rlabel metal2 s 34048 0 34104 400 6 mem_rdata[23]
port 98 nsew signal output
rlabel metal2 s 34384 0 34440 400 6 mem_rdata[24]
port 99 nsew signal output
rlabel metal2 s 34720 0 34776 400 6 mem_rdata[25]
port 100 nsew signal output
rlabel metal2 s 35056 0 35112 400 6 mem_rdata[26]
port 101 nsew signal output
rlabel metal2 s 35392 0 35448 400 6 mem_rdata[27]
port 102 nsew signal output
rlabel metal2 s 35728 0 35784 400 6 mem_rdata[28]
port 103 nsew signal output
rlabel metal2 s 36064 0 36120 400 6 mem_rdata[29]
port 104 nsew signal output
rlabel metal2 s 26992 0 27048 400 6 mem_rdata[2]
port 105 nsew signal output
rlabel metal2 s 36400 0 36456 400 6 mem_rdata[30]
port 106 nsew signal output
rlabel metal2 s 36736 0 36792 400 6 mem_rdata[31]
port 107 nsew signal output
rlabel metal2 s 27328 0 27384 400 6 mem_rdata[3]
port 108 nsew signal output
rlabel metal2 s 27664 0 27720 400 6 mem_rdata[4]
port 109 nsew signal output
rlabel metal2 s 28000 0 28056 400 6 mem_rdata[5]
port 110 nsew signal output
rlabel metal2 s 28336 0 28392 400 6 mem_rdata[6]
port 111 nsew signal output
rlabel metal2 s 28672 0 28728 400 6 mem_rdata[7]
port 112 nsew signal output
rlabel metal2 s 29008 0 29064 400 6 mem_rdata[8]
port 113 nsew signal output
rlabel metal2 s 29344 0 29400 400 6 mem_rdata[9]
port 114 nsew signal output
rlabel metal2 s 24640 0 24696 400 6 mem_ready
port 115 nsew signal output
rlabel metal2 s 23968 0 24024 400 6 mem_valid
port 116 nsew signal input
rlabel metal2 s 2464 0 2520 400 6 mem_wdata[0]
port 117 nsew signal input
rlabel metal2 s 5824 0 5880 400 6 mem_wdata[10]
port 118 nsew signal input
rlabel metal2 s 6160 0 6216 400 6 mem_wdata[11]
port 119 nsew signal input
rlabel metal2 s 6496 0 6552 400 6 mem_wdata[12]
port 120 nsew signal input
rlabel metal2 s 6832 0 6888 400 6 mem_wdata[13]
port 121 nsew signal input
rlabel metal2 s 7168 0 7224 400 6 mem_wdata[14]
port 122 nsew signal input
rlabel metal2 s 7504 0 7560 400 6 mem_wdata[15]
port 123 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 mem_wdata[16]
port 124 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 mem_wdata[17]
port 125 nsew signal input
rlabel metal2 s 8512 0 8568 400 6 mem_wdata[18]
port 126 nsew signal input
rlabel metal2 s 8848 0 8904 400 6 mem_wdata[19]
port 127 nsew signal input
rlabel metal2 s 2800 0 2856 400 6 mem_wdata[1]
port 128 nsew signal input
rlabel metal2 s 9184 0 9240 400 6 mem_wdata[20]
port 129 nsew signal input
rlabel metal2 s 9520 0 9576 400 6 mem_wdata[21]
port 130 nsew signal input
rlabel metal2 s 9856 0 9912 400 6 mem_wdata[22]
port 131 nsew signal input
rlabel metal2 s 10192 0 10248 400 6 mem_wdata[23]
port 132 nsew signal input
rlabel metal2 s 10528 0 10584 400 6 mem_wdata[24]
port 133 nsew signal input
rlabel metal2 s 10864 0 10920 400 6 mem_wdata[25]
port 134 nsew signal input
rlabel metal2 s 11200 0 11256 400 6 mem_wdata[26]
port 135 nsew signal input
rlabel metal2 s 11536 0 11592 400 6 mem_wdata[27]
port 136 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 mem_wdata[28]
port 137 nsew signal input
rlabel metal2 s 12208 0 12264 400 6 mem_wdata[29]
port 138 nsew signal input
rlabel metal2 s 3136 0 3192 400 6 mem_wdata[2]
port 139 nsew signal input
rlabel metal2 s 12544 0 12600 400 6 mem_wdata[30]
port 140 nsew signal input
rlabel metal2 s 12880 0 12936 400 6 mem_wdata[31]
port 141 nsew signal input
rlabel metal2 s 3472 0 3528 400 6 mem_wdata[3]
port 142 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 mem_wdata[4]
port 143 nsew signal input
rlabel metal2 s 4144 0 4200 400 6 mem_wdata[5]
port 144 nsew signal input
rlabel metal2 s 4480 0 4536 400 6 mem_wdata[6]
port 145 nsew signal input
rlabel metal2 s 4816 0 4872 400 6 mem_wdata[7]
port 146 nsew signal input
rlabel metal2 s 5152 0 5208 400 6 mem_wdata[8]
port 147 nsew signal input
rlabel metal2 s 5488 0 5544 400 6 mem_wdata[9]
port 148 nsew signal input
rlabel metal2 s 24976 0 25032 400 6 mem_wstrb[0]
port 149 nsew signal input
rlabel metal2 s 25312 0 25368 400 6 mem_wstrb[1]
port 150 nsew signal input
rlabel metal2 s 25648 0 25704 400 6 mem_wstrb[2]
port 151 nsew signal input
rlabel metal2 s 25984 0 26040 400 6 mem_wstrb[3]
port 152 nsew signal input
rlabel metal3 s 0 19040 400 19096 6 ram_gwenb[0]
port 153 nsew signal output
rlabel metal3 s 0 19600 400 19656 6 ram_gwenb[1]
port 154 nsew signal output
rlabel metal3 s 0 20160 400 20216 6 ram_gwenb[2]
port 155 nsew signal output
rlabel metal3 s 0 20720 400 20776 6 ram_gwenb[3]
port 156 nsew signal output
rlabel metal3 s 0 1120 400 1176 6 ram_rdata[0]
port 157 nsew signal input
rlabel metal3 s 0 6720 400 6776 6 ram_rdata[10]
port 158 nsew signal input
rlabel metal3 s 0 7280 400 7336 6 ram_rdata[11]
port 159 nsew signal input
rlabel metal3 s 0 7840 400 7896 6 ram_rdata[12]
port 160 nsew signal input
rlabel metal3 s 0 8400 400 8456 6 ram_rdata[13]
port 161 nsew signal input
rlabel metal3 s 0 8960 400 9016 6 ram_rdata[14]
port 162 nsew signal input
rlabel metal3 s 0 9520 400 9576 6 ram_rdata[15]
port 163 nsew signal input
rlabel metal3 s 0 10080 400 10136 6 ram_rdata[16]
port 164 nsew signal input
rlabel metal3 s 0 10640 400 10696 6 ram_rdata[17]
port 165 nsew signal input
rlabel metal3 s 0 11200 400 11256 6 ram_rdata[18]
port 166 nsew signal input
rlabel metal3 s 0 11760 400 11816 6 ram_rdata[19]
port 167 nsew signal input
rlabel metal3 s 0 1680 400 1736 6 ram_rdata[1]
port 168 nsew signal input
rlabel metal3 s 0 12320 400 12376 6 ram_rdata[20]
port 169 nsew signal input
rlabel metal3 s 0 12880 400 12936 6 ram_rdata[21]
port 170 nsew signal input
rlabel metal3 s 0 13440 400 13496 6 ram_rdata[22]
port 171 nsew signal input
rlabel metal3 s 0 14000 400 14056 6 ram_rdata[23]
port 172 nsew signal input
rlabel metal3 s 0 14560 400 14616 6 ram_rdata[24]
port 173 nsew signal input
rlabel metal3 s 0 15120 400 15176 6 ram_rdata[25]
port 174 nsew signal input
rlabel metal3 s 0 15680 400 15736 6 ram_rdata[26]
port 175 nsew signal input
rlabel metal3 s 0 16240 400 16296 6 ram_rdata[27]
port 176 nsew signal input
rlabel metal3 s 0 16800 400 16856 6 ram_rdata[28]
port 177 nsew signal input
rlabel metal3 s 0 17360 400 17416 6 ram_rdata[29]
port 178 nsew signal input
rlabel metal3 s 0 2240 400 2296 6 ram_rdata[2]
port 179 nsew signal input
rlabel metal3 s 0 17920 400 17976 6 ram_rdata[30]
port 180 nsew signal input
rlabel metal3 s 0 18480 400 18536 6 ram_rdata[31]
port 181 nsew signal input
rlabel metal3 s 0 2800 400 2856 6 ram_rdata[3]
port 182 nsew signal input
rlabel metal3 s 0 3360 400 3416 6 ram_rdata[4]
port 183 nsew signal input
rlabel metal3 s 0 3920 400 3976 6 ram_rdata[5]
port 184 nsew signal input
rlabel metal3 s 0 4480 400 4536 6 ram_rdata[6]
port 185 nsew signal input
rlabel metal3 s 0 5040 400 5096 6 ram_rdata[7]
port 186 nsew signal input
rlabel metal3 s 0 5600 400 5656 6 ram_rdata[8]
port 187 nsew signal input
rlabel metal3 s 0 6160 400 6216 6 ram_rdata[9]
port 188 nsew signal input
rlabel metal3 s 0 21280 400 21336 6 ram_wenb[0]
port 189 nsew signal output
rlabel metal3 s 0 26880 400 26936 6 ram_wenb[10]
port 190 nsew signal output
rlabel metal3 s 0 27440 400 27496 6 ram_wenb[11]
port 191 nsew signal output
rlabel metal3 s 0 28000 400 28056 6 ram_wenb[12]
port 192 nsew signal output
rlabel metal3 s 0 28560 400 28616 6 ram_wenb[13]
port 193 nsew signal output
rlabel metal3 s 0 29120 400 29176 6 ram_wenb[14]
port 194 nsew signal output
rlabel metal3 s 0 29680 400 29736 6 ram_wenb[15]
port 195 nsew signal output
rlabel metal3 s 0 30240 400 30296 6 ram_wenb[16]
port 196 nsew signal output
rlabel metal3 s 0 30800 400 30856 6 ram_wenb[17]
port 197 nsew signal output
rlabel metal3 s 0 31360 400 31416 6 ram_wenb[18]
port 198 nsew signal output
rlabel metal3 s 0 31920 400 31976 6 ram_wenb[19]
port 199 nsew signal output
rlabel metal3 s 0 21840 400 21896 6 ram_wenb[1]
port 200 nsew signal output
rlabel metal3 s 0 32480 400 32536 6 ram_wenb[20]
port 201 nsew signal output
rlabel metal3 s 0 33040 400 33096 6 ram_wenb[21]
port 202 nsew signal output
rlabel metal3 s 0 33600 400 33656 6 ram_wenb[22]
port 203 nsew signal output
rlabel metal3 s 0 34160 400 34216 6 ram_wenb[23]
port 204 nsew signal output
rlabel metal3 s 0 34720 400 34776 6 ram_wenb[24]
port 205 nsew signal output
rlabel metal3 s 0 35280 400 35336 6 ram_wenb[25]
port 206 nsew signal output
rlabel metal3 s 0 35840 400 35896 6 ram_wenb[26]
port 207 nsew signal output
rlabel metal3 s 0 36400 400 36456 6 ram_wenb[27]
port 208 nsew signal output
rlabel metal3 s 0 36960 400 37016 6 ram_wenb[28]
port 209 nsew signal output
rlabel metal3 s 0 37520 400 37576 6 ram_wenb[29]
port 210 nsew signal output
rlabel metal3 s 0 22400 400 22456 6 ram_wenb[2]
port 211 nsew signal output
rlabel metal3 s 0 38080 400 38136 6 ram_wenb[30]
port 212 nsew signal output
rlabel metal3 s 0 38640 400 38696 6 ram_wenb[31]
port 213 nsew signal output
rlabel metal3 s 0 22960 400 23016 6 ram_wenb[3]
port 214 nsew signal output
rlabel metal3 s 0 23520 400 23576 6 ram_wenb[4]
port 215 nsew signal output
rlabel metal3 s 0 24080 400 24136 6 ram_wenb[5]
port 216 nsew signal output
rlabel metal3 s 0 24640 400 24696 6 ram_wenb[6]
port 217 nsew signal output
rlabel metal3 s 0 25200 400 25256 6 ram_wenb[7]
port 218 nsew signal output
rlabel metal3 s 0 25760 400 25816 6 ram_wenb[8]
port 219 nsew signal output
rlabel metal3 s 0 26320 400 26376 6 ram_wenb[9]
port 220 nsew signal output
rlabel metal2 s 37408 0 37464 400 6 resetn
port 221 nsew signal input
rlabel metal3 s 39600 21056 40000 21112 6 simpleuart_dat_re
port 222 nsew signal output
rlabel metal3 s 39600 20496 40000 20552 6 simpleuart_dat_we
port 223 nsew signal output
rlabel metal3 s 39600 336 40000 392 6 simpleuart_div_we[0]
port 224 nsew signal output
rlabel metal3 s 39600 896 40000 952 6 simpleuart_div_we[1]
port 225 nsew signal output
rlabel metal3 s 39600 1456 40000 1512 6 simpleuart_div_we[2]
port 226 nsew signal output
rlabel metal3 s 39600 2016 40000 2072 6 simpleuart_div_we[3]
port 227 nsew signal output
rlabel metal3 s 39600 21616 40000 21672 6 simpleuart_reg_dat_do[0]
port 228 nsew signal input
rlabel metal3 s 39600 27216 40000 27272 6 simpleuart_reg_dat_do[10]
port 229 nsew signal input
rlabel metal3 s 39600 27776 40000 27832 6 simpleuart_reg_dat_do[11]
port 230 nsew signal input
rlabel metal3 s 39600 28336 40000 28392 6 simpleuart_reg_dat_do[12]
port 231 nsew signal input
rlabel metal3 s 39600 28896 40000 28952 6 simpleuart_reg_dat_do[13]
port 232 nsew signal input
rlabel metal3 s 39600 29456 40000 29512 6 simpleuart_reg_dat_do[14]
port 233 nsew signal input
rlabel metal3 s 39600 30016 40000 30072 6 simpleuart_reg_dat_do[15]
port 234 nsew signal input
rlabel metal3 s 39600 30576 40000 30632 6 simpleuart_reg_dat_do[16]
port 235 nsew signal input
rlabel metal3 s 39600 31136 40000 31192 6 simpleuart_reg_dat_do[17]
port 236 nsew signal input
rlabel metal3 s 39600 31696 40000 31752 6 simpleuart_reg_dat_do[18]
port 237 nsew signal input
rlabel metal3 s 39600 32256 40000 32312 6 simpleuart_reg_dat_do[19]
port 238 nsew signal input
rlabel metal3 s 39600 22176 40000 22232 6 simpleuart_reg_dat_do[1]
port 239 nsew signal input
rlabel metal3 s 39600 32816 40000 32872 6 simpleuart_reg_dat_do[20]
port 240 nsew signal input
rlabel metal3 s 39600 33376 40000 33432 6 simpleuart_reg_dat_do[21]
port 241 nsew signal input
rlabel metal3 s 39600 33936 40000 33992 6 simpleuart_reg_dat_do[22]
port 242 nsew signal input
rlabel metal3 s 39600 34496 40000 34552 6 simpleuart_reg_dat_do[23]
port 243 nsew signal input
rlabel metal3 s 39600 35056 40000 35112 6 simpleuart_reg_dat_do[24]
port 244 nsew signal input
rlabel metal3 s 39600 35616 40000 35672 6 simpleuart_reg_dat_do[25]
port 245 nsew signal input
rlabel metal3 s 39600 36176 40000 36232 6 simpleuart_reg_dat_do[26]
port 246 nsew signal input
rlabel metal3 s 39600 36736 40000 36792 6 simpleuart_reg_dat_do[27]
port 247 nsew signal input
rlabel metal3 s 39600 37296 40000 37352 6 simpleuart_reg_dat_do[28]
port 248 nsew signal input
rlabel metal3 s 39600 37856 40000 37912 6 simpleuart_reg_dat_do[29]
port 249 nsew signal input
rlabel metal3 s 39600 22736 40000 22792 6 simpleuart_reg_dat_do[2]
port 250 nsew signal input
rlabel metal3 s 39600 38416 40000 38472 6 simpleuart_reg_dat_do[30]
port 251 nsew signal input
rlabel metal3 s 39600 38976 40000 39032 6 simpleuart_reg_dat_do[31]
port 252 nsew signal input
rlabel metal3 s 39600 23296 40000 23352 6 simpleuart_reg_dat_do[3]
port 253 nsew signal input
rlabel metal3 s 39600 23856 40000 23912 6 simpleuart_reg_dat_do[4]
port 254 nsew signal input
rlabel metal3 s 39600 24416 40000 24472 6 simpleuart_reg_dat_do[5]
port 255 nsew signal input
rlabel metal3 s 39600 24976 40000 25032 6 simpleuart_reg_dat_do[6]
port 256 nsew signal input
rlabel metal3 s 39600 25536 40000 25592 6 simpleuart_reg_dat_do[7]
port 257 nsew signal input
rlabel metal3 s 39600 26096 40000 26152 6 simpleuart_reg_dat_do[8]
port 258 nsew signal input
rlabel metal3 s 39600 26656 40000 26712 6 simpleuart_reg_dat_do[9]
port 259 nsew signal input
rlabel metal3 s 39600 39536 40000 39592 6 simpleuart_reg_dat_wait
port 260 nsew signal input
rlabel metal3 s 39600 2576 40000 2632 6 simpleuart_reg_div_do[0]
port 261 nsew signal input
rlabel metal3 s 39600 8176 40000 8232 6 simpleuart_reg_div_do[10]
port 262 nsew signal input
rlabel metal3 s 39600 8736 40000 8792 6 simpleuart_reg_div_do[11]
port 263 nsew signal input
rlabel metal3 s 39600 9296 40000 9352 6 simpleuart_reg_div_do[12]
port 264 nsew signal input
rlabel metal3 s 39600 9856 40000 9912 6 simpleuart_reg_div_do[13]
port 265 nsew signal input
rlabel metal3 s 39600 10416 40000 10472 6 simpleuart_reg_div_do[14]
port 266 nsew signal input
rlabel metal3 s 39600 10976 40000 11032 6 simpleuart_reg_div_do[15]
port 267 nsew signal input
rlabel metal3 s 39600 11536 40000 11592 6 simpleuart_reg_div_do[16]
port 268 nsew signal input
rlabel metal3 s 39600 12096 40000 12152 6 simpleuart_reg_div_do[17]
port 269 nsew signal input
rlabel metal3 s 39600 12656 40000 12712 6 simpleuart_reg_div_do[18]
port 270 nsew signal input
rlabel metal3 s 39600 13216 40000 13272 6 simpleuart_reg_div_do[19]
port 271 nsew signal input
rlabel metal3 s 39600 3136 40000 3192 6 simpleuart_reg_div_do[1]
port 272 nsew signal input
rlabel metal3 s 39600 13776 40000 13832 6 simpleuart_reg_div_do[20]
port 273 nsew signal input
rlabel metal3 s 39600 14336 40000 14392 6 simpleuart_reg_div_do[21]
port 274 nsew signal input
rlabel metal3 s 39600 14896 40000 14952 6 simpleuart_reg_div_do[22]
port 275 nsew signal input
rlabel metal3 s 39600 15456 40000 15512 6 simpleuart_reg_div_do[23]
port 276 nsew signal input
rlabel metal3 s 39600 16016 40000 16072 6 simpleuart_reg_div_do[24]
port 277 nsew signal input
rlabel metal3 s 39600 16576 40000 16632 6 simpleuart_reg_div_do[25]
port 278 nsew signal input
rlabel metal3 s 39600 17136 40000 17192 6 simpleuart_reg_div_do[26]
port 279 nsew signal input
rlabel metal3 s 39600 17696 40000 17752 6 simpleuart_reg_div_do[27]
port 280 nsew signal input
rlabel metal3 s 39600 18256 40000 18312 6 simpleuart_reg_div_do[28]
port 281 nsew signal input
rlabel metal3 s 39600 18816 40000 18872 6 simpleuart_reg_div_do[29]
port 282 nsew signal input
rlabel metal3 s 39600 3696 40000 3752 6 simpleuart_reg_div_do[2]
port 283 nsew signal input
rlabel metal3 s 39600 19376 40000 19432 6 simpleuart_reg_div_do[30]
port 284 nsew signal input
rlabel metal3 s 39600 19936 40000 19992 6 simpleuart_reg_div_do[31]
port 285 nsew signal input
rlabel metal3 s 39600 4256 40000 4312 6 simpleuart_reg_div_do[3]
port 286 nsew signal input
rlabel metal3 s 39600 4816 40000 4872 6 simpleuart_reg_div_do[4]
port 287 nsew signal input
rlabel metal3 s 39600 5376 40000 5432 6 simpleuart_reg_div_do[5]
port 288 nsew signal input
rlabel metal3 s 39600 5936 40000 5992 6 simpleuart_reg_div_do[6]
port 289 nsew signal input
rlabel metal3 s 39600 6496 40000 6552 6 simpleuart_reg_div_do[7]
port 290 nsew signal input
rlabel metal3 s 39600 7056 40000 7112 6 simpleuart_reg_div_do[8]
port 291 nsew signal input
rlabel metal3 s 39600 7616 40000 7672 6 simpleuart_reg_div_do[9]
port 292 nsew signal input
rlabel metal2 s 17024 39600 17080 40000 6 spimem_rdata[0]
port 293 nsew signal input
rlabel metal2 s 20384 39600 20440 40000 6 spimem_rdata[10]
port 294 nsew signal input
rlabel metal2 s 20720 39600 20776 40000 6 spimem_rdata[11]
port 295 nsew signal input
rlabel metal2 s 21056 39600 21112 40000 6 spimem_rdata[12]
port 296 nsew signal input
rlabel metal2 s 21392 39600 21448 40000 6 spimem_rdata[13]
port 297 nsew signal input
rlabel metal2 s 21728 39600 21784 40000 6 spimem_rdata[14]
port 298 nsew signal input
rlabel metal2 s 22064 39600 22120 40000 6 spimem_rdata[15]
port 299 nsew signal input
rlabel metal2 s 22400 39600 22456 40000 6 spimem_rdata[16]
port 300 nsew signal input
rlabel metal2 s 22736 39600 22792 40000 6 spimem_rdata[17]
port 301 nsew signal input
rlabel metal2 s 23072 39600 23128 40000 6 spimem_rdata[18]
port 302 nsew signal input
rlabel metal2 s 23408 39600 23464 40000 6 spimem_rdata[19]
port 303 nsew signal input
rlabel metal2 s 17360 39600 17416 40000 6 spimem_rdata[1]
port 304 nsew signal input
rlabel metal2 s 23744 39600 23800 40000 6 spimem_rdata[20]
port 305 nsew signal input
rlabel metal2 s 24080 39600 24136 40000 6 spimem_rdata[21]
port 306 nsew signal input
rlabel metal2 s 24416 39600 24472 40000 6 spimem_rdata[22]
port 307 nsew signal input
rlabel metal2 s 24752 39600 24808 40000 6 spimem_rdata[23]
port 308 nsew signal input
rlabel metal2 s 25088 39600 25144 40000 6 spimem_rdata[24]
port 309 nsew signal input
rlabel metal2 s 25424 39600 25480 40000 6 spimem_rdata[25]
port 310 nsew signal input
rlabel metal2 s 25760 39600 25816 40000 6 spimem_rdata[26]
port 311 nsew signal input
rlabel metal2 s 26096 39600 26152 40000 6 spimem_rdata[27]
port 312 nsew signal input
rlabel metal2 s 26432 39600 26488 40000 6 spimem_rdata[28]
port 313 nsew signal input
rlabel metal2 s 26768 39600 26824 40000 6 spimem_rdata[29]
port 314 nsew signal input
rlabel metal2 s 17696 39600 17752 40000 6 spimem_rdata[2]
port 315 nsew signal input
rlabel metal2 s 27104 39600 27160 40000 6 spimem_rdata[30]
port 316 nsew signal input
rlabel metal2 s 27440 39600 27496 40000 6 spimem_rdata[31]
port 317 nsew signal input
rlabel metal2 s 18032 39600 18088 40000 6 spimem_rdata[3]
port 318 nsew signal input
rlabel metal2 s 18368 39600 18424 40000 6 spimem_rdata[4]
port 319 nsew signal input
rlabel metal2 s 18704 39600 18760 40000 6 spimem_rdata[5]
port 320 nsew signal input
rlabel metal2 s 19040 39600 19096 40000 6 spimem_rdata[6]
port 321 nsew signal input
rlabel metal2 s 19376 39600 19432 40000 6 spimem_rdata[7]
port 322 nsew signal input
rlabel metal2 s 19712 39600 19768 40000 6 spimem_rdata[8]
port 323 nsew signal input
rlabel metal2 s 20048 39600 20104 40000 6 spimem_rdata[9]
port 324 nsew signal input
rlabel metal2 s 16352 39600 16408 40000 6 spimem_ready
port 325 nsew signal input
rlabel metal2 s 16688 39600 16744 40000 6 spimem_valid
port 326 nsew signal output
rlabel metal2 s 29120 39600 29176 40000 6 spimemio_cfgreg_do[0]
port 327 nsew signal input
rlabel metal2 s 32480 39600 32536 40000 6 spimemio_cfgreg_do[10]
port 328 nsew signal input
rlabel metal2 s 32816 39600 32872 40000 6 spimemio_cfgreg_do[11]
port 329 nsew signal input
rlabel metal2 s 33152 39600 33208 40000 6 spimemio_cfgreg_do[12]
port 330 nsew signal input
rlabel metal2 s 33488 39600 33544 40000 6 spimemio_cfgreg_do[13]
port 331 nsew signal input
rlabel metal2 s 33824 39600 33880 40000 6 spimemio_cfgreg_do[14]
port 332 nsew signal input
rlabel metal2 s 34160 39600 34216 40000 6 spimemio_cfgreg_do[15]
port 333 nsew signal input
rlabel metal2 s 34496 39600 34552 40000 6 spimemio_cfgreg_do[16]
port 334 nsew signal input
rlabel metal2 s 34832 39600 34888 40000 6 spimemio_cfgreg_do[17]
port 335 nsew signal input
rlabel metal2 s 35168 39600 35224 40000 6 spimemio_cfgreg_do[18]
port 336 nsew signal input
rlabel metal2 s 35504 39600 35560 40000 6 spimemio_cfgreg_do[19]
port 337 nsew signal input
rlabel metal2 s 29456 39600 29512 40000 6 spimemio_cfgreg_do[1]
port 338 nsew signal input
rlabel metal2 s 35840 39600 35896 40000 6 spimemio_cfgreg_do[20]
port 339 nsew signal input
rlabel metal2 s 36176 39600 36232 40000 6 spimemio_cfgreg_do[21]
port 340 nsew signal input
rlabel metal2 s 36512 39600 36568 40000 6 spimemio_cfgreg_do[22]
port 341 nsew signal input
rlabel metal2 s 36848 39600 36904 40000 6 spimemio_cfgreg_do[23]
port 342 nsew signal input
rlabel metal2 s 37184 39600 37240 40000 6 spimemio_cfgreg_do[24]
port 343 nsew signal input
rlabel metal2 s 37520 39600 37576 40000 6 spimemio_cfgreg_do[25]
port 344 nsew signal input
rlabel metal2 s 37856 39600 37912 40000 6 spimemio_cfgreg_do[26]
port 345 nsew signal input
rlabel metal2 s 38192 39600 38248 40000 6 spimemio_cfgreg_do[27]
port 346 nsew signal input
rlabel metal2 s 38528 39600 38584 40000 6 spimemio_cfgreg_do[28]
port 347 nsew signal input
rlabel metal2 s 38864 39600 38920 40000 6 spimemio_cfgreg_do[29]
port 348 nsew signal input
rlabel metal2 s 29792 39600 29848 40000 6 spimemio_cfgreg_do[2]
port 349 nsew signal input
rlabel metal2 s 39200 39600 39256 40000 6 spimemio_cfgreg_do[30]
port 350 nsew signal input
rlabel metal2 s 39536 39600 39592 40000 6 spimemio_cfgreg_do[31]
port 351 nsew signal input
rlabel metal2 s 30128 39600 30184 40000 6 spimemio_cfgreg_do[3]
port 352 nsew signal input
rlabel metal2 s 30464 39600 30520 40000 6 spimemio_cfgreg_do[4]
port 353 nsew signal input
rlabel metal2 s 30800 39600 30856 40000 6 spimemio_cfgreg_do[5]
port 354 nsew signal input
rlabel metal2 s 31136 39600 31192 40000 6 spimemio_cfgreg_do[6]
port 355 nsew signal input
rlabel metal2 s 31472 39600 31528 40000 6 spimemio_cfgreg_do[7]
port 356 nsew signal input
rlabel metal2 s 31808 39600 31864 40000 6 spimemio_cfgreg_do[8]
port 357 nsew signal input
rlabel metal2 s 32144 39600 32200 40000 6 spimemio_cfgreg_do[9]
port 358 nsew signal input
rlabel metal2 s 27776 39600 27832 40000 6 spimemio_cfgreg_we[0]
port 359 nsew signal output
rlabel metal2 s 28112 39600 28168 40000 6 spimemio_cfgreg_we[1]
port 360 nsew signal output
rlabel metal2 s 28448 39600 28504 40000 6 spimemio_cfgreg_we[2]
port 361 nsew signal output
rlabel metal2 s 28784 39600 28840 40000 6 spimemio_cfgreg_we[3]
port 362 nsew signal output
rlabel metal4 s 2224 1538 2384 38446 6 vdd
port 363 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 38446 6 vdd
port 363 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 38446 6 vdd
port 363 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 38446 6 vss
port 364 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 38446 6 vss
port 364 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2445470
string GDS_FILE /home/luke/picosoc-w-approximation/openlane/simple_interconnect/runs/23_12_10_20_43/results/signoff/simple_interconnect.magic.gds
string GDS_START 200898
<< end >>


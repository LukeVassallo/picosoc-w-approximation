magic
tech gf180mcuD
magscale 1 10
timestamp 1702237379
<< metal1 >>
rect 16034 46734 16046 46786
rect 16098 46783 16110 46786
rect 17490 46783 17502 46786
rect 16098 46737 17502 46783
rect 16098 46734 16110 46737
rect 17490 46734 17502 46737
rect 17554 46734 17566 46786
rect 27570 46734 27582 46786
rect 27634 46783 27646 46786
rect 28578 46783 28590 46786
rect 27634 46737 28590 46783
rect 27634 46734 27646 46737
rect 28578 46734 28590 46737
rect 28642 46734 28654 46786
rect 19058 46510 19070 46562
rect 19122 46559 19134 46562
rect 19506 46559 19518 46562
rect 19122 46513 19518 46559
rect 19122 46510 19134 46513
rect 19506 46510 19518 46513
rect 19570 46559 19582 46562
rect 20066 46559 20078 46562
rect 19570 46513 20078 46559
rect 19570 46510 19582 46513
rect 20066 46510 20078 46513
rect 20130 46510 20142 46562
rect 18162 46398 18174 46450
rect 18226 46447 18238 46450
rect 21634 46447 21646 46450
rect 18226 46401 21646 46447
rect 18226 46398 18238 46401
rect 21634 46398 21646 46401
rect 21698 46398 21710 46450
rect 23762 46398 23774 46450
rect 23826 46447 23838 46450
rect 24882 46447 24894 46450
rect 23826 46401 24894 46447
rect 23826 46398 23838 46401
rect 24882 46398 24894 46401
rect 24946 46398 24958 46450
rect 26898 46398 26910 46450
rect 26962 46447 26974 46450
rect 27458 46447 27470 46450
rect 26962 46401 27470 46447
rect 26962 46398 26974 46401
rect 27458 46398 27470 46401
rect 27522 46398 27534 46450
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 17950 46114 18002 46126
rect 17950 46050 18002 46062
rect 25566 46114 25618 46126
rect 25566 46050 25618 46062
rect 30046 46114 30098 46126
rect 30046 46050 30098 46062
rect 36990 46114 37042 46126
rect 36990 46050 37042 46062
rect 41470 46114 41522 46126
rect 41470 46050 41522 46062
rect 44606 46114 44658 46126
rect 44606 46050 44658 46062
rect 8878 46002 8930 46014
rect 8878 45938 8930 45950
rect 13470 46002 13522 46014
rect 13470 45938 13522 45950
rect 22318 46002 22370 46014
rect 22318 45938 22370 45950
rect 35198 46002 35250 46014
rect 35198 45938 35250 45950
rect 9662 45890 9714 45902
rect 13694 45890 13746 45902
rect 16046 45890 16098 45902
rect 22990 45890 23042 45902
rect 27470 45890 27522 45902
rect 47406 45890 47458 45902
rect 10546 45838 10558 45890
rect 10610 45838 10622 45890
rect 11666 45838 11678 45890
rect 11730 45838 11742 45890
rect 12338 45838 12350 45890
rect 12402 45838 12414 45890
rect 14802 45838 14814 45890
rect 14866 45838 14878 45890
rect 15586 45838 15598 45890
rect 15650 45838 15662 45890
rect 17378 45838 17390 45890
rect 17442 45838 17454 45890
rect 20066 45838 20078 45890
rect 20130 45838 20142 45890
rect 20962 45838 20974 45890
rect 21026 45838 21038 45890
rect 21634 45838 21646 45890
rect 21698 45838 21710 45890
rect 23762 45838 23774 45890
rect 23826 45838 23838 45890
rect 24994 45838 25006 45890
rect 25058 45838 25070 45890
rect 28578 45838 28590 45890
rect 28642 45838 28654 45890
rect 29250 45838 29262 45890
rect 29314 45838 29326 45890
rect 32274 45838 32286 45890
rect 32338 45838 32350 45890
rect 32834 45838 32846 45890
rect 32898 45838 32910 45890
rect 35970 45838 35982 45890
rect 36034 45838 36046 45890
rect 40450 45838 40462 45890
rect 40514 45838 40526 45890
rect 43698 45838 43710 45890
rect 43762 45838 43774 45890
rect 9662 45826 9714 45838
rect 13694 45826 13746 45838
rect 16046 45826 16098 45838
rect 22990 45826 23042 45838
rect 27470 45826 27522 45838
rect 47406 45826 47458 45838
rect 22766 45778 22818 45790
rect 22766 45714 22818 45726
rect 38894 45778 38946 45790
rect 38894 45714 38946 45726
rect 39230 45778 39282 45790
rect 39230 45714 39282 45726
rect 39790 45778 39842 45790
rect 39790 45714 39842 45726
rect 40126 45778 40178 45790
rect 40126 45714 40178 45726
rect 9998 45666 10050 45678
rect 9998 45602 10050 45614
rect 10334 45666 10386 45678
rect 10334 45602 10386 45614
rect 11902 45666 11954 45678
rect 11902 45602 11954 45614
rect 12574 45666 12626 45678
rect 12574 45602 12626 45614
rect 14030 45666 14082 45678
rect 14030 45602 14082 45614
rect 15038 45666 15090 45678
rect 15038 45602 15090 45614
rect 15374 45666 15426 45678
rect 15374 45602 15426 45614
rect 16382 45666 16434 45678
rect 16382 45602 16434 45614
rect 19854 45666 19906 45678
rect 19854 45602 19906 45614
rect 20750 45666 20802 45678
rect 20750 45602 20802 45614
rect 21422 45666 21474 45678
rect 21422 45602 21474 45614
rect 23326 45666 23378 45678
rect 23326 45602 23378 45614
rect 23998 45666 24050 45678
rect 23998 45602 24050 45614
rect 27806 45666 27858 45678
rect 27806 45602 27858 45614
rect 28366 45666 28418 45678
rect 28366 45602 28418 45614
rect 32510 45666 32562 45678
rect 46846 45666 46898 45678
rect 46498 45614 46510 45666
rect 46562 45614 46574 45666
rect 32510 45602 32562 45614
rect 46846 45602 46898 45614
rect 47518 45666 47570 45678
rect 47518 45602 47570 45614
rect 47630 45666 47682 45678
rect 47630 45602 47682 45614
rect 47854 45666 47906 45678
rect 47854 45602 47906 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 10110 45330 10162 45342
rect 10110 45266 10162 45278
rect 12126 45330 12178 45342
rect 12126 45266 12178 45278
rect 12798 45330 12850 45342
rect 12798 45266 12850 45278
rect 14814 45330 14866 45342
rect 14814 45266 14866 45278
rect 15374 45330 15426 45342
rect 15374 45266 15426 45278
rect 15822 45330 15874 45342
rect 15822 45266 15874 45278
rect 16270 45330 16322 45342
rect 16270 45266 16322 45278
rect 29710 45330 29762 45342
rect 29710 45266 29762 45278
rect 42254 45330 42306 45342
rect 42254 45266 42306 45278
rect 47182 45330 47234 45342
rect 47182 45266 47234 45278
rect 16494 45218 16546 45230
rect 16494 45154 16546 45166
rect 16830 45218 16882 45230
rect 16830 45154 16882 45166
rect 24334 45218 24386 45230
rect 24334 45154 24386 45166
rect 28478 45218 28530 45230
rect 28478 45154 28530 45166
rect 28814 45218 28866 45230
rect 30830 45218 30882 45230
rect 31838 45218 31890 45230
rect 30482 45166 30494 45218
rect 30546 45166 30558 45218
rect 31154 45166 31166 45218
rect 31218 45166 31230 45218
rect 28814 45154 28866 45166
rect 30830 45154 30882 45166
rect 31838 45154 31890 45166
rect 32174 45218 32226 45230
rect 32174 45154 32226 45166
rect 32510 45218 32562 45230
rect 32510 45154 32562 45166
rect 33182 45218 33234 45230
rect 33182 45154 33234 45166
rect 33518 45218 33570 45230
rect 33518 45154 33570 45166
rect 33854 45218 33906 45230
rect 33854 45154 33906 45166
rect 29374 45106 29426 45118
rect 48078 45106 48130 45118
rect 17378 45054 17390 45106
rect 17442 45054 17454 45106
rect 21074 45054 21086 45106
rect 21138 45054 21150 45106
rect 24546 45054 24558 45106
rect 24610 45054 24622 45106
rect 25330 45054 25342 45106
rect 25394 45054 25406 45106
rect 30258 45054 30270 45106
rect 30322 45054 30334 45106
rect 31602 45054 31614 45106
rect 31666 45054 31678 45106
rect 34066 45054 34078 45106
rect 34130 45054 34142 45106
rect 36978 45054 36990 45106
rect 37042 45054 37054 45106
rect 37762 45054 37774 45106
rect 37826 45054 37838 45106
rect 41234 45054 41246 45106
rect 41298 45054 41310 45106
rect 44146 45054 44158 45106
rect 44210 45054 44222 45106
rect 29374 45042 29426 45054
rect 48078 45042 48130 45054
rect 47518 44994 47570 45006
rect 18162 44942 18174 44994
rect 18226 44942 18238 44994
rect 20290 44942 20302 44994
rect 20354 44942 20366 44994
rect 20514 44942 20526 44994
rect 20578 44991 20590 44994
rect 20738 44991 20750 44994
rect 20578 44945 20750 44991
rect 20578 44942 20590 44945
rect 20738 44942 20750 44945
rect 20802 44942 20814 44994
rect 21746 44942 21758 44994
rect 21810 44942 21822 44994
rect 23874 44942 23886 44994
rect 23938 44942 23950 44994
rect 26002 44942 26014 44994
rect 26066 44942 26078 44994
rect 28130 44942 28142 44994
rect 28194 44942 28206 44994
rect 45378 44942 45390 44994
rect 45442 44942 45454 44994
rect 47518 44930 47570 44942
rect 36430 44882 36482 44894
rect 36430 44818 36482 44830
rect 40126 44882 40178 44894
rect 40126 44818 40178 44830
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 36206 44546 36258 44558
rect 36206 44482 36258 44494
rect 41134 44546 41186 44558
rect 41134 44482 41186 44494
rect 45838 44546 45890 44558
rect 45838 44482 45890 44494
rect 18398 44434 18450 44446
rect 17042 44382 17054 44434
rect 17106 44382 17118 44434
rect 18398 44370 18450 44382
rect 19070 44434 19122 44446
rect 19070 44370 19122 44382
rect 21422 44434 21474 44446
rect 21422 44370 21474 44382
rect 21870 44434 21922 44446
rect 21870 44370 21922 44382
rect 24894 44434 24946 44446
rect 24894 44370 24946 44382
rect 27246 44434 27298 44446
rect 27246 44370 27298 44382
rect 28254 44434 28306 44446
rect 28254 44370 28306 44382
rect 30942 44434 30994 44446
rect 43810 44382 43822 44434
rect 43874 44382 43886 44434
rect 30942 44370 30994 44382
rect 18510 44322 18562 44334
rect 19742 44322 19794 44334
rect 20526 44322 20578 44334
rect 21310 44322 21362 44334
rect 14242 44270 14254 44322
rect 14306 44270 14318 44322
rect 19506 44270 19518 44322
rect 19570 44270 19582 44322
rect 20066 44270 20078 44322
rect 20130 44270 20142 44322
rect 20738 44270 20750 44322
rect 20802 44270 20814 44322
rect 18510 44258 18562 44270
rect 19742 44258 19794 44270
rect 20526 44258 20578 44270
rect 21310 44258 21362 44270
rect 31838 44322 31890 44334
rect 32610 44270 32622 44322
rect 32674 44270 32686 44322
rect 33842 44270 33854 44322
rect 33906 44270 33918 44322
rect 37538 44270 37550 44322
rect 37602 44270 37614 44322
rect 38210 44270 38222 44322
rect 38274 44270 38286 44322
rect 38770 44270 38782 44322
rect 38834 44270 38846 44322
rect 41682 44270 41694 44322
rect 41746 44270 41758 44322
rect 44818 44270 44830 44322
rect 44882 44270 44894 44322
rect 31838 44258 31890 44270
rect 19294 44210 19346 44222
rect 14914 44158 14926 44210
rect 14978 44158 14990 44210
rect 19294 44146 19346 44158
rect 19406 44210 19458 44222
rect 19406 44146 19458 44158
rect 20414 44210 20466 44222
rect 20414 44146 20466 44158
rect 23438 44210 23490 44222
rect 23438 44146 23490 44158
rect 32174 44210 32226 44222
rect 32174 44146 32226 44158
rect 32846 44210 32898 44222
rect 32846 44146 32898 44158
rect 37774 44210 37826 44222
rect 47742 44210 47794 44222
rect 38434 44158 38446 44210
rect 38498 44158 38510 44210
rect 37774 44146 37826 44158
rect 47742 44146 47794 44158
rect 18062 44098 18114 44110
rect 18062 44034 18114 44046
rect 18286 44098 18338 44110
rect 18286 44034 18338 44046
rect 23326 44098 23378 44110
rect 23326 44034 23378 44046
rect 29598 44098 29650 44110
rect 29598 44034 29650 44046
rect 29934 44098 29986 44110
rect 29934 44034 29986 44046
rect 30382 44098 30434 44110
rect 31502 44098 31554 44110
rect 31154 44046 31166 44098
rect 31218 44046 31230 44098
rect 30382 44034 30434 44046
rect 31502 44034 31554 44046
rect 33182 44098 33234 44110
rect 37102 44098 37154 44110
rect 33506 44046 33518 44098
rect 33570 44046 33582 44098
rect 33182 44034 33234 44046
rect 37102 44034 37154 44046
rect 48078 44098 48130 44110
rect 48078 44034 48130 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 18398 43762 18450 43774
rect 18398 43698 18450 43710
rect 22430 43762 22482 43774
rect 22430 43698 22482 43710
rect 22766 43762 22818 43774
rect 22766 43698 22818 43710
rect 24670 43762 24722 43774
rect 24670 43698 24722 43710
rect 25342 43762 25394 43774
rect 25342 43698 25394 43710
rect 27358 43762 27410 43774
rect 27358 43698 27410 43710
rect 27806 43762 27858 43774
rect 27806 43698 27858 43710
rect 28926 43762 28978 43774
rect 28926 43698 28978 43710
rect 17502 43650 17554 43662
rect 17502 43586 17554 43598
rect 18510 43650 18562 43662
rect 18510 43586 18562 43598
rect 19742 43650 19794 43662
rect 19742 43586 19794 43598
rect 20526 43650 20578 43662
rect 25230 43650 25282 43662
rect 21858 43598 21870 43650
rect 21922 43598 21934 43650
rect 24098 43598 24110 43650
rect 24162 43598 24174 43650
rect 20526 43586 20578 43598
rect 25230 43586 25282 43598
rect 25678 43650 25730 43662
rect 25678 43586 25730 43598
rect 26238 43650 26290 43662
rect 30382 43650 30434 43662
rect 32510 43650 32562 43662
rect 34526 43650 34578 43662
rect 26786 43598 26798 43650
rect 26850 43598 26862 43650
rect 31490 43598 31502 43650
rect 31554 43598 31566 43650
rect 33842 43598 33854 43650
rect 33906 43598 33918 43650
rect 26238 43586 26290 43598
rect 30382 43586 30434 43598
rect 32510 43586 32562 43598
rect 34526 43586 34578 43598
rect 41470 43650 41522 43662
rect 41470 43586 41522 43598
rect 4846 43538 4898 43550
rect 4274 43486 4286 43538
rect 4338 43486 4350 43538
rect 4846 43474 4898 43486
rect 10110 43538 10162 43550
rect 10110 43474 10162 43486
rect 10558 43538 10610 43550
rect 10558 43474 10610 43486
rect 10782 43538 10834 43550
rect 16718 43538 16770 43550
rect 16482 43486 16494 43538
rect 16546 43486 16558 43538
rect 10782 43474 10834 43486
rect 16718 43474 16770 43486
rect 17390 43538 17442 43550
rect 17390 43474 17442 43486
rect 17614 43538 17666 43550
rect 17614 43474 17666 43486
rect 18062 43538 18114 43550
rect 18062 43474 18114 43486
rect 21646 43538 21698 43550
rect 22990 43538 23042 43550
rect 22418 43486 22430 43538
rect 22482 43486 22494 43538
rect 21646 43474 21698 43486
rect 22990 43474 23042 43486
rect 23438 43538 23490 43550
rect 23438 43474 23490 43486
rect 23886 43538 23938 43550
rect 25454 43538 25506 43550
rect 24658 43486 24670 43538
rect 24722 43486 24734 43538
rect 23886 43474 23938 43486
rect 25454 43474 25506 43486
rect 26574 43538 26626 43550
rect 28030 43538 28082 43550
rect 28814 43538 28866 43550
rect 27122 43486 27134 43538
rect 27186 43486 27198 43538
rect 28354 43486 28366 43538
rect 28418 43486 28430 43538
rect 26574 43474 26626 43486
rect 28030 43474 28082 43486
rect 28814 43474 28866 43486
rect 30830 43538 30882 43550
rect 31714 43486 31726 43538
rect 31778 43486 31790 43538
rect 32274 43486 32286 43538
rect 32338 43486 32350 43538
rect 33618 43486 33630 43538
rect 33682 43486 33694 43538
rect 34290 43486 34302 43538
rect 34354 43486 34366 43538
rect 35074 43486 35086 43538
rect 35138 43486 35150 43538
rect 37762 43486 37774 43538
rect 37826 43486 37838 43538
rect 41234 43486 41246 43538
rect 41298 43486 41310 43538
rect 42914 43486 42926 43538
rect 42978 43486 42990 43538
rect 45826 43486 45838 43538
rect 45890 43486 45902 43538
rect 30830 43474 30882 43486
rect 10334 43426 10386 43438
rect 10334 43362 10386 43374
rect 16830 43426 16882 43438
rect 16830 43362 16882 43374
rect 18286 43426 18338 43438
rect 18286 43362 18338 43374
rect 22094 43426 22146 43438
rect 22094 43362 22146 43374
rect 22878 43426 22930 43438
rect 22878 43362 22930 43374
rect 27918 43426 27970 43438
rect 27918 43362 27970 43374
rect 31278 43426 31330 43438
rect 31278 43362 31330 43374
rect 33182 43426 33234 43438
rect 33182 43362 33234 43374
rect 42366 43426 42418 43438
rect 44930 43374 44942 43426
rect 44994 43374 45006 43426
rect 47842 43374 47854 43426
rect 47906 43374 47918 43426
rect 42366 43362 42418 43374
rect 1934 43314 1986 43326
rect 1934 43250 1986 43262
rect 19854 43314 19906 43326
rect 19854 43250 19906 43262
rect 24334 43314 24386 43326
rect 24334 43250 24386 43262
rect 26126 43314 26178 43326
rect 26126 43250 26178 43262
rect 27022 43314 27074 43326
rect 27022 43250 27074 43262
rect 28702 43314 28754 43326
rect 28702 43250 28754 43262
rect 37214 43314 37266 43326
rect 37214 43250 37266 43262
rect 40126 43314 40178 43326
rect 40126 43250 40178 43262
rect 41806 43314 41858 43326
rect 41806 43250 41858 43262
rect 42142 43314 42194 43326
rect 42142 43250 42194 43262
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 19854 42978 19906 42990
rect 19854 42914 19906 42926
rect 27134 42978 27186 42990
rect 27134 42914 27186 42926
rect 36206 42978 36258 42990
rect 36206 42914 36258 42926
rect 42814 42978 42866 42990
rect 42814 42914 42866 42926
rect 14478 42866 14530 42878
rect 2034 42814 2046 42866
rect 2098 42814 2110 42866
rect 8866 42814 8878 42866
rect 8930 42814 8942 42866
rect 10994 42814 11006 42866
rect 11058 42814 11070 42866
rect 14478 42802 14530 42814
rect 19518 42866 19570 42878
rect 19518 42802 19570 42814
rect 22542 42866 22594 42878
rect 22542 42802 22594 42814
rect 25006 42866 25058 42878
rect 25006 42802 25058 42814
rect 25566 42866 25618 42878
rect 43710 42866 43762 42878
rect 29138 42814 29150 42866
rect 29202 42814 29214 42866
rect 31266 42814 31278 42866
rect 31330 42814 31342 42866
rect 41906 42814 41918 42866
rect 41970 42814 41982 42866
rect 25566 42802 25618 42814
rect 43710 42802 43762 42814
rect 47966 42866 48018 42878
rect 47966 42802 48018 42814
rect 13582 42754 13634 42766
rect 4050 42702 4062 42754
rect 4114 42702 4126 42754
rect 8194 42702 8206 42754
rect 8258 42702 8270 42754
rect 13582 42690 13634 42702
rect 13806 42754 13858 42766
rect 13806 42690 13858 42702
rect 14142 42754 14194 42766
rect 14142 42690 14194 42702
rect 14366 42754 14418 42766
rect 14366 42690 14418 42702
rect 19406 42754 19458 42766
rect 25118 42754 25170 42766
rect 27470 42754 27522 42766
rect 37662 42754 37714 42766
rect 20066 42702 20078 42754
rect 20130 42702 20142 42754
rect 23202 42702 23214 42754
rect 23266 42702 23278 42754
rect 24770 42702 24782 42754
rect 24834 42702 24846 42754
rect 25778 42702 25790 42754
rect 25842 42702 25854 42754
rect 27122 42702 27134 42754
rect 27186 42702 27198 42754
rect 31938 42702 31950 42754
rect 32002 42702 32014 42754
rect 33282 42702 33294 42754
rect 33346 42702 33358 42754
rect 33842 42702 33854 42754
rect 33906 42702 33918 42754
rect 19406 42690 19458 42702
rect 25118 42690 25170 42702
rect 27470 42690 27522 42702
rect 37662 42690 37714 42702
rect 38334 42754 38386 42766
rect 42478 42754 42530 42766
rect 38994 42702 39006 42754
rect 39058 42702 39070 42754
rect 38334 42690 38386 42702
rect 42478 42690 42530 42702
rect 43486 42754 43538 42766
rect 45602 42702 45614 42754
rect 45666 42702 45678 42754
rect 43486 42690 43538 42702
rect 22430 42642 22482 42654
rect 19618 42590 19630 42642
rect 19682 42590 19694 42642
rect 22430 42578 22482 42590
rect 22654 42642 22706 42654
rect 22654 42578 22706 42590
rect 23550 42642 23602 42654
rect 23550 42578 23602 42590
rect 25454 42642 25506 42654
rect 25454 42578 25506 42590
rect 26798 42642 26850 42654
rect 26798 42578 26850 42590
rect 27582 42642 27634 42654
rect 27582 42578 27634 42590
rect 32510 42642 32562 42654
rect 32510 42578 32562 42590
rect 32846 42642 32898 42654
rect 32846 42578 32898 42590
rect 33518 42642 33570 42654
rect 33518 42578 33570 42590
rect 37998 42642 38050 42654
rect 42254 42642 42306 42654
rect 38658 42590 38670 42642
rect 38722 42590 38734 42642
rect 39778 42590 39790 42642
rect 39842 42590 39854 42642
rect 37998 42578 38050 42590
rect 42254 42578 42306 42590
rect 44830 42642 44882 42654
rect 44830 42578 44882 42590
rect 45166 42642 45218 42654
rect 45166 42578 45218 42590
rect 11454 42530 11506 42542
rect 11454 42466 11506 42478
rect 13918 42530 13970 42542
rect 13918 42466 13970 42478
rect 23438 42530 23490 42542
rect 23438 42466 23490 42478
rect 36990 42530 37042 42542
rect 44158 42530 44210 42542
rect 37314 42478 37326 42530
rect 37378 42478 37390 42530
rect 43138 42478 43150 42530
rect 43202 42478 43214 42530
rect 36990 42466 37042 42478
rect 44158 42466 44210 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 10110 42194 10162 42206
rect 10110 42130 10162 42142
rect 11006 42194 11058 42206
rect 15262 42194 15314 42206
rect 11890 42142 11902 42194
rect 11954 42142 11966 42194
rect 11006 42130 11058 42142
rect 15262 42130 15314 42142
rect 20078 42194 20130 42206
rect 35086 42194 35138 42206
rect 23202 42142 23214 42194
rect 23266 42142 23278 42194
rect 34738 42142 34750 42194
rect 34802 42142 34814 42194
rect 20078 42130 20130 42142
rect 35086 42130 35138 42142
rect 39230 42194 39282 42206
rect 39230 42130 39282 42142
rect 42030 42194 42082 42206
rect 42030 42130 42082 42142
rect 11118 42082 11170 42094
rect 15486 42082 15538 42094
rect 14130 42030 14142 42082
rect 14194 42030 14206 42082
rect 11118 42018 11170 42030
rect 15486 42018 15538 42030
rect 17390 42082 17442 42094
rect 39006 42082 39058 42094
rect 34066 42030 34078 42082
rect 34130 42030 34142 42082
rect 17390 42018 17442 42030
rect 39006 42018 39058 42030
rect 40350 42082 40402 42094
rect 40350 42018 40402 42030
rect 41806 42082 41858 42094
rect 41806 42018 41858 42030
rect 9998 41970 10050 41982
rect 4274 41918 4286 41970
rect 4338 41918 4350 41970
rect 5282 41918 5294 41970
rect 5346 41918 5358 41970
rect 9998 41906 10050 41918
rect 10894 41970 10946 41982
rect 10894 41906 10946 41918
rect 11566 41970 11618 41982
rect 15374 41970 15426 41982
rect 14802 41918 14814 41970
rect 14866 41918 14878 41970
rect 11566 41906 11618 41918
rect 15374 41906 15426 41918
rect 15934 41970 15986 41982
rect 15934 41906 15986 41918
rect 17614 41970 17666 41982
rect 17614 41906 17666 41918
rect 18062 41970 18114 41982
rect 18062 41906 18114 41918
rect 20302 41970 20354 41982
rect 20302 41906 20354 41918
rect 20638 41970 20690 41982
rect 20638 41906 20690 41918
rect 20750 41970 20802 41982
rect 21422 41970 21474 41982
rect 33742 41970 33794 41982
rect 21074 41918 21086 41970
rect 21138 41918 21150 41970
rect 23426 41918 23438 41970
rect 23490 41918 23502 41970
rect 20750 41906 20802 41918
rect 21422 41906 21474 41918
rect 33742 41906 33794 41918
rect 34414 41970 34466 41982
rect 34414 41906 34466 41918
rect 35422 41970 35474 41982
rect 39678 41970 39730 41982
rect 40910 41970 40962 41982
rect 35858 41918 35870 41970
rect 35922 41918 35934 41970
rect 40114 41918 40126 41970
rect 40178 41918 40190 41970
rect 35422 41906 35474 41918
rect 39678 41906 39730 41918
rect 40910 41906 40962 41918
rect 41022 41970 41074 41982
rect 41022 41906 41074 41918
rect 41246 41970 41298 41982
rect 41246 41906 41298 41918
rect 41358 41970 41410 41982
rect 41358 41906 41410 41918
rect 41918 41970 41970 41982
rect 42354 41918 42366 41970
rect 42418 41918 42430 41970
rect 42802 41918 42814 41970
rect 42866 41918 42878 41970
rect 45714 41918 45726 41970
rect 45778 41918 45790 41970
rect 41918 41906 41970 41918
rect 5742 41858 5794 41870
rect 5742 41794 5794 41806
rect 16270 41858 16322 41870
rect 16270 41794 16322 41806
rect 17502 41858 17554 41870
rect 17502 41794 17554 41806
rect 20190 41858 20242 41870
rect 20190 41794 20242 41806
rect 21310 41858 21362 41870
rect 21310 41794 21362 41806
rect 32174 41858 32226 41870
rect 32174 41794 32226 41806
rect 33182 41858 33234 41870
rect 39118 41858 39170 41870
rect 36530 41806 36542 41858
rect 36594 41806 36606 41858
rect 38658 41806 38670 41858
rect 38722 41806 38734 41858
rect 47618 41806 47630 41858
rect 47682 41806 47694 41858
rect 33182 41794 33234 41806
rect 39118 41794 39170 41806
rect 1934 41746 1986 41758
rect 1934 41682 1986 41694
rect 4958 41746 5010 41758
rect 4958 41682 5010 41694
rect 5294 41746 5346 41758
rect 5294 41682 5346 41694
rect 45054 41746 45106 41758
rect 45054 41682 45106 41694
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 21870 41410 21922 41422
rect 21870 41346 21922 41358
rect 26798 41410 26850 41422
rect 26798 41346 26850 41358
rect 41134 41410 41186 41422
rect 41134 41346 41186 41358
rect 44046 41410 44098 41422
rect 44046 41346 44098 41358
rect 48190 41410 48242 41422
rect 48190 41346 48242 41358
rect 14926 41298 14978 41310
rect 22206 41298 22258 41310
rect 27134 41298 27186 41310
rect 37102 41298 37154 41310
rect 4610 41246 4622 41298
rect 4674 41246 4686 41298
rect 6402 41246 6414 41298
rect 6466 41246 6478 41298
rect 8530 41246 8542 41298
rect 8594 41246 8606 41298
rect 16818 41246 16830 41298
rect 16882 41246 16894 41298
rect 18946 41246 18958 41298
rect 19010 41246 19022 41298
rect 26114 41246 26126 41298
rect 26178 41246 26190 41298
rect 34626 41246 34638 41298
rect 34690 41246 34702 41298
rect 47730 41246 47742 41298
rect 47794 41246 47806 41298
rect 14926 41234 14978 41246
rect 22206 41234 22258 41246
rect 27134 41234 27186 41246
rect 37102 41234 37154 41246
rect 22318 41186 22370 41198
rect 1698 41134 1710 41186
rect 1762 41134 1774 41186
rect 5730 41134 5742 41186
rect 5794 41134 5806 41186
rect 16034 41134 16046 41186
rect 16098 41134 16110 41186
rect 21522 41134 21534 41186
rect 21586 41134 21598 41186
rect 22318 41122 22370 41134
rect 25790 41186 25842 41198
rect 27582 41186 27634 41198
rect 26450 41134 26462 41186
rect 26514 41134 26526 41186
rect 27010 41134 27022 41186
rect 27074 41134 27086 41186
rect 25790 41122 25842 41134
rect 27582 41122 27634 41134
rect 30830 41186 30882 41198
rect 35086 41186 35138 41198
rect 31826 41134 31838 41186
rect 31890 41134 31902 41186
rect 30830 41122 30882 41134
rect 35086 41122 35138 41134
rect 35534 41186 35586 41198
rect 36878 41186 36930 41198
rect 36194 41134 36206 41186
rect 36258 41134 36270 41186
rect 35534 41122 35586 41134
rect 36878 41122 36930 41134
rect 37550 41186 37602 41198
rect 37550 41122 37602 41134
rect 38110 41186 38162 41198
rect 38770 41134 38782 41186
rect 38834 41134 38846 41186
rect 41682 41134 41694 41186
rect 41746 41134 41758 41186
rect 44930 41134 44942 41186
rect 44994 41134 45006 41186
rect 38110 41122 38162 41134
rect 23214 41074 23266 41086
rect 2482 41022 2494 41074
rect 2546 41022 2558 41074
rect 22082 41022 22094 41074
rect 22146 41022 22158 41074
rect 23214 41010 23266 41022
rect 23550 41074 23602 41086
rect 23550 41010 23602 41022
rect 25006 41074 25058 41086
rect 25006 41010 25058 41022
rect 25342 41074 25394 41086
rect 25342 41010 25394 41022
rect 27246 41074 27298 41086
rect 27246 41010 27298 41022
rect 28030 41074 28082 41086
rect 36430 41074 36482 41086
rect 32498 41022 32510 41074
rect 32562 41022 32574 41074
rect 28030 41010 28082 41022
rect 36430 41010 36482 41022
rect 37326 41074 37378 41086
rect 37326 41010 37378 41022
rect 38446 41074 38498 41086
rect 45602 41022 45614 41074
rect 45666 41022 45678 41074
rect 38446 41010 38498 41022
rect 5070 40962 5122 40974
rect 5070 40898 5122 40910
rect 8990 40962 9042 40974
rect 8990 40898 9042 40910
rect 23886 40962 23938 40974
rect 26014 40962 26066 40974
rect 24210 40910 24222 40962
rect 24274 40910 24286 40962
rect 23886 40898 23938 40910
rect 26014 40898 26066 40910
rect 27694 40962 27746 40974
rect 27694 40898 27746 40910
rect 27806 40962 27858 40974
rect 27806 40898 27858 40910
rect 35646 40962 35698 40974
rect 35646 40898 35698 40910
rect 35758 40962 35810 40974
rect 35758 40898 35810 40910
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 5742 40626 5794 40638
rect 5742 40562 5794 40574
rect 10222 40626 10274 40638
rect 10222 40562 10274 40574
rect 18958 40626 19010 40638
rect 22990 40626 23042 40638
rect 22642 40574 22654 40626
rect 22706 40574 22718 40626
rect 18958 40562 19010 40574
rect 22990 40562 23042 40574
rect 25230 40626 25282 40638
rect 27246 40626 27298 40638
rect 25554 40574 25566 40626
rect 25618 40574 25630 40626
rect 25230 40562 25282 40574
rect 27246 40562 27298 40574
rect 33742 40626 33794 40638
rect 41134 40626 41186 40638
rect 34066 40574 34078 40626
rect 34130 40574 34142 40626
rect 37090 40574 37102 40626
rect 37154 40574 37166 40626
rect 33742 40562 33794 40574
rect 41134 40562 41186 40574
rect 9774 40514 9826 40526
rect 4610 40462 4622 40514
rect 4674 40462 4686 40514
rect 5394 40462 5406 40514
rect 5458 40462 5470 40514
rect 6850 40462 6862 40514
rect 6914 40462 6926 40514
rect 9774 40450 9826 40462
rect 11230 40514 11282 40526
rect 11230 40450 11282 40462
rect 11454 40514 11506 40526
rect 11454 40450 11506 40462
rect 12126 40514 12178 40526
rect 12126 40450 12178 40462
rect 15150 40514 15202 40526
rect 15150 40450 15202 40462
rect 26462 40514 26514 40526
rect 26462 40450 26514 40462
rect 26574 40514 26626 40526
rect 34638 40514 34690 40526
rect 41470 40514 41522 40526
rect 29810 40462 29822 40514
rect 29874 40462 29886 40514
rect 36530 40462 36542 40514
rect 36594 40462 36606 40514
rect 39442 40462 39454 40514
rect 39506 40462 39518 40514
rect 26574 40450 26626 40462
rect 34638 40450 34690 40462
rect 41470 40450 41522 40462
rect 4958 40402 5010 40414
rect 9886 40402 9938 40414
rect 4274 40350 4286 40402
rect 4338 40350 4350 40402
rect 6178 40350 6190 40402
rect 6242 40350 6254 40402
rect 4958 40338 5010 40350
rect 9886 40338 9938 40350
rect 11006 40402 11058 40414
rect 11006 40338 11058 40350
rect 11566 40402 11618 40414
rect 23662 40402 23714 40414
rect 30942 40402 30994 40414
rect 35086 40402 35138 40414
rect 17378 40350 17390 40402
rect 17442 40350 17454 40402
rect 19506 40350 19518 40402
rect 19570 40350 19582 40402
rect 20178 40350 20190 40402
rect 20242 40350 20254 40402
rect 24210 40350 24222 40402
rect 24274 40350 24286 40402
rect 30594 40350 30606 40402
rect 30658 40350 30670 40402
rect 31378 40350 31390 40402
rect 31442 40350 31454 40402
rect 11566 40338 11618 40350
rect 23662 40338 23714 40350
rect 30942 40338 30994 40350
rect 35086 40338 35138 40350
rect 35310 40402 35362 40414
rect 35310 40338 35362 40350
rect 35422 40402 35474 40414
rect 35422 40338 35474 40350
rect 35646 40402 35698 40414
rect 35646 40338 35698 40350
rect 36206 40402 36258 40414
rect 36206 40338 36258 40350
rect 37438 40402 37490 40414
rect 40910 40402 40962 40414
rect 37762 40350 37774 40402
rect 37826 40350 37838 40402
rect 37438 40338 37490 40350
rect 40910 40338 40962 40350
rect 41246 40402 41298 40414
rect 42690 40350 42702 40402
rect 42754 40350 42766 40402
rect 45938 40350 45950 40402
rect 46002 40350 46014 40402
rect 41246 40338 41298 40350
rect 17614 40290 17666 40302
rect 8978 40238 8990 40290
rect 9042 40238 9054 40290
rect 10658 40238 10670 40290
rect 10722 40238 10734 40290
rect 17614 40226 17666 40238
rect 17726 40290 17778 40302
rect 17726 40226 17778 40238
rect 18734 40290 18786 40302
rect 23774 40290 23826 40302
rect 22306 40238 22318 40290
rect 22370 40238 22382 40290
rect 18734 40226 18786 40238
rect 23774 40226 23826 40238
rect 27022 40290 27074 40302
rect 42142 40290 42194 40302
rect 27346 40238 27358 40290
rect 27410 40238 27422 40290
rect 27682 40238 27694 40290
rect 27746 40238 27758 40290
rect 27022 40226 27074 40238
rect 42142 40226 42194 40238
rect 42366 40290 42418 40302
rect 47730 40238 47742 40290
rect 47794 40238 47806 40290
rect 42366 40226 42418 40238
rect 1934 40178 1986 40190
rect 1934 40114 1986 40126
rect 12238 40178 12290 40190
rect 12238 40114 12290 40126
rect 15262 40178 15314 40190
rect 15262 40114 15314 40126
rect 19070 40178 19122 40190
rect 19070 40114 19122 40126
rect 23998 40178 24050 40190
rect 23998 40114 24050 40126
rect 26462 40178 26514 40190
rect 26462 40114 26514 40126
rect 34414 40178 34466 40190
rect 34414 40114 34466 40126
rect 41806 40178 41858 40190
rect 41806 40114 41858 40126
rect 45054 40178 45106 40190
rect 45054 40114 45106 40126
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 26798 39842 26850 39854
rect 4386 39790 4398 39842
rect 4450 39790 4462 39842
rect 35970 39790 35982 39842
rect 36034 39839 36046 39842
rect 36530 39839 36542 39842
rect 36034 39793 36542 39839
rect 36034 39790 36046 39793
rect 36530 39790 36542 39793
rect 36594 39790 36606 39842
rect 43586 39790 43598 39842
rect 43650 39790 43662 39842
rect 26798 39778 26850 39790
rect 2494 39730 2546 39742
rect 5070 39730 5122 39742
rect 4274 39678 4286 39730
rect 4338 39678 4350 39730
rect 2494 39666 2546 39678
rect 5070 39666 5122 39678
rect 11566 39730 11618 39742
rect 20078 39730 20130 39742
rect 17602 39678 17614 39730
rect 17666 39678 17678 39730
rect 19394 39678 19406 39730
rect 19458 39727 19470 39730
rect 19618 39727 19630 39730
rect 19458 39681 19630 39727
rect 19458 39678 19470 39681
rect 19618 39678 19630 39681
rect 19682 39678 19694 39730
rect 11566 39666 11618 39678
rect 20078 39666 20130 39678
rect 26910 39730 26962 39742
rect 26910 39666 26962 39678
rect 34862 39730 34914 39742
rect 34862 39666 34914 39678
rect 35982 39730 36034 39742
rect 35982 39666 36034 39678
rect 36430 39730 36482 39742
rect 36430 39666 36482 39678
rect 37774 39730 37826 39742
rect 41010 39678 41022 39730
rect 41074 39678 41086 39730
rect 37774 39666 37826 39678
rect 10558 39618 10610 39630
rect 3714 39566 3726 39618
rect 3778 39566 3790 39618
rect 10098 39566 10110 39618
rect 10162 39566 10174 39618
rect 10558 39554 10610 39566
rect 11678 39618 11730 39630
rect 11678 39554 11730 39566
rect 12238 39618 12290 39630
rect 19182 39618 19234 39630
rect 14802 39566 14814 39618
rect 14866 39566 14878 39618
rect 12238 39554 12290 39566
rect 19182 39554 19234 39566
rect 19966 39618 20018 39630
rect 19966 39554 20018 39566
rect 20190 39618 20242 39630
rect 20190 39554 20242 39566
rect 24222 39618 24274 39630
rect 24222 39554 24274 39566
rect 36990 39618 37042 39630
rect 45166 39618 45218 39630
rect 38098 39566 38110 39618
rect 38162 39566 38174 39618
rect 41682 39566 41694 39618
rect 41746 39566 41758 39618
rect 48066 39566 48078 39618
rect 48130 39566 48142 39618
rect 36990 39554 37042 39566
rect 45166 39554 45218 39566
rect 2158 39506 2210 39518
rect 2158 39442 2210 39454
rect 2382 39506 2434 39518
rect 2382 39442 2434 39454
rect 7534 39506 7586 39518
rect 7534 39442 7586 39454
rect 11230 39506 11282 39518
rect 11230 39442 11282 39454
rect 12686 39506 12738 39518
rect 12686 39442 12738 39454
rect 12910 39506 12962 39518
rect 12910 39442 12962 39454
rect 13582 39506 13634 39518
rect 13582 39442 13634 39454
rect 13918 39506 13970 39518
rect 18174 39506 18226 39518
rect 15474 39454 15486 39506
rect 15538 39454 15550 39506
rect 13918 39442 13970 39454
rect 18174 39442 18226 39454
rect 18398 39506 18450 39518
rect 18398 39442 18450 39454
rect 18846 39506 18898 39518
rect 18846 39442 18898 39454
rect 34302 39506 34354 39518
rect 38882 39454 38894 39506
rect 38946 39454 38958 39506
rect 46610 39454 46622 39506
rect 46674 39454 46686 39506
rect 34302 39442 34354 39454
rect 2606 39394 2658 39406
rect 2606 39330 2658 39342
rect 3278 39394 3330 39406
rect 3278 39330 3330 39342
rect 8094 39394 8146 39406
rect 8094 39330 8146 39342
rect 9214 39394 9266 39406
rect 9214 39330 9266 39342
rect 11454 39394 11506 39406
rect 11454 39330 11506 39342
rect 12462 39394 12514 39406
rect 12462 39330 12514 39342
rect 13806 39394 13858 39406
rect 13806 39330 13858 39342
rect 14030 39394 14082 39406
rect 14030 39330 14082 39342
rect 17950 39394 18002 39406
rect 17950 39330 18002 39342
rect 18062 39394 18114 39406
rect 18062 39330 18114 39342
rect 19742 39394 19794 39406
rect 30606 39394 30658 39406
rect 23874 39342 23886 39394
rect 23938 39342 23950 39394
rect 19742 39330 19794 39342
rect 30606 39330 30658 39342
rect 31278 39394 31330 39406
rect 31278 39330 31330 39342
rect 31614 39394 31666 39406
rect 35310 39394 35362 39406
rect 44830 39394 44882 39406
rect 31938 39342 31950 39394
rect 32002 39342 32014 39394
rect 37314 39342 37326 39394
rect 37378 39342 37390 39394
rect 31614 39330 31666 39342
rect 35310 39330 35362 39342
rect 44830 39330 44882 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 7310 39058 7362 39070
rect 7310 38994 7362 39006
rect 10670 39058 10722 39070
rect 10670 38994 10722 39006
rect 15486 39058 15538 39070
rect 32510 39058 32562 39070
rect 18274 39006 18286 39058
rect 18338 39006 18350 39058
rect 19954 39006 19966 39058
rect 20018 39006 20030 39058
rect 23650 39006 23662 39058
rect 23714 39006 23726 39058
rect 15486 38994 15538 39006
rect 32510 38994 32562 39006
rect 34526 39058 34578 39070
rect 34526 38994 34578 39006
rect 36654 39058 36706 39070
rect 39454 39058 39506 39070
rect 38658 39006 38670 39058
rect 38722 39006 38734 39058
rect 36654 38994 36706 39006
rect 39454 38994 39506 39006
rect 40910 39058 40962 39070
rect 40910 38994 40962 39006
rect 41918 39058 41970 39070
rect 41918 38994 41970 39006
rect 3614 38946 3666 38958
rect 3614 38882 3666 38894
rect 3726 38946 3778 38958
rect 3726 38882 3778 38894
rect 4286 38946 4338 38958
rect 4286 38882 4338 38894
rect 4622 38946 4674 38958
rect 9550 38946 9602 38958
rect 8306 38894 8318 38946
rect 8370 38894 8382 38946
rect 4622 38882 4674 38894
rect 9550 38882 9602 38894
rect 11006 38946 11058 38958
rect 15934 38946 15986 38958
rect 12338 38894 12350 38946
rect 12402 38894 12414 38946
rect 11006 38882 11058 38894
rect 15934 38882 15986 38894
rect 33182 38946 33234 38958
rect 33182 38882 33234 38894
rect 33406 38946 33458 38958
rect 33406 38882 33458 38894
rect 33742 38946 33794 38958
rect 33742 38882 33794 38894
rect 33854 38946 33906 38958
rect 33854 38882 33906 38894
rect 33966 38946 34018 38958
rect 33966 38882 34018 38894
rect 36990 38946 37042 38958
rect 39342 38946 39394 38958
rect 37986 38894 37998 38946
rect 38050 38894 38062 38946
rect 36990 38882 37042 38894
rect 39342 38882 39394 38894
rect 41134 38946 41186 38958
rect 41134 38882 41186 38894
rect 41358 38946 41410 38958
rect 41358 38882 41410 38894
rect 42814 38946 42866 38958
rect 42814 38882 42866 38894
rect 47518 38946 47570 38958
rect 47518 38882 47570 38894
rect 48190 38946 48242 38958
rect 48190 38882 48242 38894
rect 2718 38834 2770 38846
rect 4398 38834 4450 38846
rect 3938 38782 3950 38834
rect 4002 38782 4014 38834
rect 2718 38770 2770 38782
rect 4398 38770 4450 38782
rect 4846 38834 4898 38846
rect 4846 38770 4898 38782
rect 6414 38834 6466 38846
rect 8990 38834 9042 38846
rect 6738 38782 6750 38834
rect 6802 38782 6814 38834
rect 7522 38782 7534 38834
rect 7586 38782 7598 38834
rect 7970 38782 7982 38834
rect 8034 38782 8046 38834
rect 6414 38770 6466 38782
rect 8990 38770 9042 38782
rect 9662 38834 9714 38846
rect 9662 38770 9714 38782
rect 10110 38834 10162 38846
rect 10110 38770 10162 38782
rect 11118 38834 11170 38846
rect 15262 38834 15314 38846
rect 11666 38782 11678 38834
rect 11730 38782 11742 38834
rect 11118 38770 11170 38782
rect 15262 38770 15314 38782
rect 15710 38834 15762 38846
rect 17950 38834 18002 38846
rect 17490 38782 17502 38834
rect 17554 38782 17566 38834
rect 15710 38770 15762 38782
rect 17950 38770 18002 38782
rect 18622 38834 18674 38846
rect 18622 38770 18674 38782
rect 20302 38834 20354 38846
rect 20302 38770 20354 38782
rect 23998 38834 24050 38846
rect 23998 38770 24050 38782
rect 24446 38834 24498 38846
rect 32398 38834 32450 38846
rect 29138 38782 29150 38834
rect 29202 38782 29214 38834
rect 24446 38770 24498 38782
rect 32398 38770 32450 38782
rect 37326 38834 37378 38846
rect 37326 38770 37378 38782
rect 37662 38834 37714 38846
rect 37662 38770 37714 38782
rect 38334 38834 38386 38846
rect 38334 38770 38386 38782
rect 39678 38834 39730 38846
rect 39678 38770 39730 38782
rect 39902 38834 39954 38846
rect 39902 38770 39954 38782
rect 41022 38834 41074 38846
rect 41022 38770 41074 38782
rect 42142 38834 42194 38846
rect 43038 38834 43090 38846
rect 46846 38834 46898 38846
rect 42466 38782 42478 38834
rect 42530 38782 42542 38834
rect 45826 38782 45838 38834
rect 45890 38782 45902 38834
rect 46498 38782 46510 38834
rect 46562 38782 46574 38834
rect 42142 38770 42194 38782
rect 43038 38770 43090 38782
rect 46846 38770 46898 38782
rect 47070 38834 47122 38846
rect 47070 38770 47122 38782
rect 47182 38834 47234 38846
rect 47182 38770 47234 38782
rect 47854 38834 47906 38846
rect 47854 38770 47906 38782
rect 2382 38722 2434 38734
rect 2382 38658 2434 38670
rect 2606 38722 2658 38734
rect 19070 38722 19122 38734
rect 40350 38722 40402 38734
rect 3154 38670 3166 38722
rect 3218 38670 3230 38722
rect 6626 38670 6638 38722
rect 6690 38670 6702 38722
rect 7858 38670 7870 38722
rect 7922 38670 7934 38722
rect 14466 38670 14478 38722
rect 14530 38670 14542 38722
rect 29810 38670 29822 38722
rect 29874 38670 29886 38722
rect 31938 38670 31950 38722
rect 32002 38670 32014 38722
rect 33058 38670 33070 38722
rect 33122 38670 33134 38722
rect 2606 38658 2658 38670
rect 19070 38658 19122 38670
rect 40350 38658 40402 38670
rect 42030 38722 42082 38734
rect 43698 38670 43710 38722
rect 43762 38670 43774 38722
rect 42030 38658 42082 38670
rect 2270 38610 2322 38622
rect 2270 38546 2322 38558
rect 43374 38610 43426 38622
rect 43374 38546 43426 38558
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 29934 38274 29986 38286
rect 29934 38210 29986 38222
rect 30270 38274 30322 38286
rect 43586 38222 43598 38274
rect 43650 38222 43662 38274
rect 30270 38210 30322 38222
rect 12014 38162 12066 38174
rect 36990 38162 37042 38174
rect 2482 38110 2494 38162
rect 2546 38110 2558 38162
rect 4610 38110 4622 38162
rect 4674 38110 4686 38162
rect 28354 38110 28366 38162
rect 28418 38110 28430 38162
rect 36082 38110 36094 38162
rect 36146 38110 36158 38162
rect 12014 38098 12066 38110
rect 36990 38098 37042 38110
rect 38110 38162 38162 38174
rect 38110 38098 38162 38110
rect 38558 38162 38610 38174
rect 38558 38098 38610 38110
rect 5630 38050 5682 38062
rect 1810 37998 1822 38050
rect 1874 37998 1886 38050
rect 5630 37986 5682 37998
rect 5966 38050 6018 38062
rect 5966 37986 6018 37998
rect 6414 38050 6466 38062
rect 9662 38050 9714 38062
rect 11454 38050 11506 38062
rect 23998 38050 24050 38062
rect 29262 38050 29314 38062
rect 41022 38050 41074 38062
rect 44830 38050 44882 38062
rect 7298 37998 7310 38050
rect 7362 37998 7374 38050
rect 8642 37998 8654 38050
rect 8706 37998 8718 38050
rect 10434 37998 10446 38050
rect 10498 37998 10510 38050
rect 20178 37998 20190 38050
rect 20242 37998 20254 38050
rect 23202 37998 23214 38050
rect 23266 37998 23278 38050
rect 24770 37998 24782 38050
rect 24834 37998 24846 38050
rect 25554 37998 25566 38050
rect 25618 37998 25630 38050
rect 33170 37998 33182 38050
rect 33234 37998 33246 38050
rect 39778 37998 39790 38050
rect 39842 37998 39854 38050
rect 41682 37998 41694 38050
rect 41746 37998 41758 38050
rect 46050 37998 46062 38050
rect 46114 37998 46126 38050
rect 6414 37986 6466 37998
rect 9662 37986 9714 37998
rect 11454 37986 11506 37998
rect 23998 37986 24050 37998
rect 29262 37986 29314 37998
rect 41022 37986 41074 37998
rect 44830 37986 44882 37998
rect 23774 37938 23826 37950
rect 40350 37938 40402 37950
rect 5730 37886 5742 37938
rect 5794 37886 5806 37938
rect 7522 37886 7534 37938
rect 7586 37886 7598 37938
rect 24994 37886 25006 37938
rect 25058 37886 25070 37938
rect 26226 37886 26238 37938
rect 26290 37886 26302 37938
rect 33954 37886 33966 37938
rect 34018 37886 34030 37938
rect 40002 37886 40014 37938
rect 40066 37886 40078 37938
rect 23774 37874 23826 37886
rect 40350 37874 40402 37886
rect 40686 37938 40738 37950
rect 40686 37874 40738 37886
rect 41358 37938 41410 37950
rect 45154 37886 45166 37938
rect 45218 37886 45230 37938
rect 47394 37886 47406 37938
rect 47458 37886 47470 37938
rect 41358 37874 41410 37886
rect 5070 37826 5122 37838
rect 5070 37762 5122 37774
rect 6638 37826 6690 37838
rect 6638 37762 6690 37774
rect 9550 37826 9602 37838
rect 9550 37762 9602 37774
rect 12462 37826 12514 37838
rect 12462 37762 12514 37774
rect 14030 37826 14082 37838
rect 14030 37762 14082 37774
rect 20414 37826 20466 37838
rect 30046 37826 30098 37838
rect 23426 37774 23438 37826
rect 23490 37774 23502 37826
rect 24322 37774 24334 37826
rect 24386 37774 24398 37826
rect 20414 37762 20466 37774
rect 30046 37762 30098 37774
rect 32174 37826 32226 37838
rect 32174 37762 32226 37774
rect 32846 37826 32898 37838
rect 32846 37762 32898 37774
rect 37102 37826 37154 37838
rect 37102 37762 37154 37774
rect 38894 37826 38946 37838
rect 38894 37762 38946 37774
rect 39454 37826 39506 37838
rect 39454 37762 39506 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 13134 37490 13186 37502
rect 4946 37438 4958 37490
rect 5010 37438 5022 37490
rect 13134 37426 13186 37438
rect 15598 37490 15650 37502
rect 18846 37490 18898 37502
rect 18498 37438 18510 37490
rect 18562 37438 18574 37490
rect 15598 37426 15650 37438
rect 18846 37426 18898 37438
rect 25342 37490 25394 37502
rect 25342 37426 25394 37438
rect 34974 37490 35026 37502
rect 34974 37426 35026 37438
rect 36094 37490 36146 37502
rect 36094 37426 36146 37438
rect 36206 37490 36258 37502
rect 36206 37426 36258 37438
rect 6638 37378 6690 37390
rect 13022 37378 13074 37390
rect 14926 37378 14978 37390
rect 7522 37326 7534 37378
rect 7586 37326 7598 37378
rect 11778 37326 11790 37378
rect 11842 37326 11854 37378
rect 14242 37326 14254 37378
rect 14306 37326 14318 37378
rect 6638 37314 6690 37326
rect 13022 37314 13074 37326
rect 14926 37314 14978 37326
rect 15710 37378 15762 37390
rect 15710 37314 15762 37326
rect 17838 37378 17890 37390
rect 17838 37314 17890 37326
rect 18174 37378 18226 37390
rect 25902 37378 25954 37390
rect 20514 37326 20526 37378
rect 20578 37326 20590 37378
rect 18174 37314 18226 37326
rect 25902 37314 25954 37326
rect 26014 37378 26066 37390
rect 26014 37314 26066 37326
rect 27694 37378 27746 37390
rect 27694 37314 27746 37326
rect 27806 37378 27858 37390
rect 27806 37314 27858 37326
rect 35422 37378 35474 37390
rect 35422 37314 35474 37326
rect 45278 37378 45330 37390
rect 45278 37314 45330 37326
rect 12910 37266 12962 37278
rect 14590 37266 14642 37278
rect 4274 37214 4286 37266
rect 4338 37214 4350 37266
rect 5170 37214 5182 37266
rect 5234 37214 5246 37266
rect 7074 37214 7086 37266
rect 7138 37214 7150 37266
rect 8082 37214 8094 37266
rect 8146 37214 8158 37266
rect 12562 37214 12574 37266
rect 12626 37214 12638 37266
rect 13346 37214 13358 37266
rect 13410 37214 13422 37266
rect 13570 37214 13582 37266
rect 13634 37214 13646 37266
rect 12910 37202 12962 37214
rect 14590 37202 14642 37214
rect 15262 37266 15314 37278
rect 15262 37202 15314 37214
rect 15934 37266 15986 37278
rect 25678 37266 25730 37278
rect 34862 37266 34914 37278
rect 19730 37214 19742 37266
rect 19794 37214 19806 37266
rect 26450 37214 26462 37266
rect 26514 37214 26526 37266
rect 15934 37202 15986 37214
rect 25678 37202 25730 37214
rect 34862 37202 34914 37214
rect 35086 37266 35138 37278
rect 35086 37202 35138 37214
rect 35982 37266 36034 37278
rect 35982 37202 36034 37214
rect 36654 37266 36706 37278
rect 44718 37266 44770 37278
rect 37202 37214 37214 37266
rect 37266 37214 37278 37266
rect 41010 37214 41022 37266
rect 41074 37214 41086 37266
rect 36654 37202 36706 37214
rect 44718 37202 44770 37214
rect 44942 37266 44994 37278
rect 45826 37214 45838 37266
rect 45890 37214 45902 37266
rect 44942 37202 44994 37214
rect 15038 37154 15090 37166
rect 44270 37154 44322 37166
rect 7746 37102 7758 37154
rect 7810 37102 7822 37154
rect 9650 37102 9662 37154
rect 9714 37102 9726 37154
rect 22642 37102 22654 37154
rect 22706 37102 22718 37154
rect 26002 37102 26014 37154
rect 26066 37102 26078 37154
rect 37986 37102 37998 37154
rect 38050 37102 38062 37154
rect 40114 37102 40126 37154
rect 40178 37102 40190 37154
rect 41682 37102 41694 37154
rect 41746 37102 41758 37154
rect 43810 37102 43822 37154
rect 43874 37102 43886 37154
rect 15038 37090 15090 37102
rect 44270 37090 44322 37102
rect 45166 37154 45218 37166
rect 47730 37102 47742 37154
rect 47794 37102 47806 37154
rect 45166 37090 45218 37102
rect 1934 37042 1986 37054
rect 44258 36990 44270 37042
rect 44322 37039 44334 37042
rect 44482 37039 44494 37042
rect 44322 36993 44494 37039
rect 44322 36990 44334 36993
rect 44482 36990 44494 36993
rect 44546 36990 44558 37042
rect 1934 36978 1986 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 4622 36706 4674 36718
rect 4622 36642 4674 36654
rect 10894 36706 10946 36718
rect 10894 36642 10946 36654
rect 13582 36706 13634 36718
rect 13582 36642 13634 36654
rect 19966 36706 20018 36718
rect 43038 36706 43090 36718
rect 20290 36654 20302 36706
rect 20354 36654 20366 36706
rect 40562 36654 40574 36706
rect 40626 36703 40638 36706
rect 41010 36703 41022 36706
rect 40626 36657 41022 36703
rect 40626 36654 40638 36657
rect 41010 36654 41022 36657
rect 41074 36654 41086 36706
rect 19966 36642 20018 36654
rect 43038 36642 43090 36654
rect 1934 36594 1986 36606
rect 9102 36594 9154 36606
rect 4946 36542 4958 36594
rect 5010 36542 5022 36594
rect 1934 36530 1986 36542
rect 9102 36530 9154 36542
rect 12798 36594 12850 36606
rect 18174 36594 18226 36606
rect 15586 36542 15598 36594
rect 15650 36542 15662 36594
rect 17714 36542 17726 36594
rect 17778 36542 17790 36594
rect 12798 36530 12850 36542
rect 18174 36530 18226 36542
rect 19742 36594 19794 36606
rect 19742 36530 19794 36542
rect 20750 36594 20802 36606
rect 29262 36594 29314 36606
rect 35646 36594 35698 36606
rect 25666 36542 25678 36594
rect 25730 36542 25742 36594
rect 32722 36542 32734 36594
rect 32786 36542 32798 36594
rect 20750 36530 20802 36542
rect 29262 36530 29314 36542
rect 35646 36530 35698 36542
rect 40014 36594 40066 36606
rect 40014 36530 40066 36542
rect 40574 36594 40626 36606
rect 40574 36530 40626 36542
rect 41806 36594 41858 36606
rect 41806 36530 41858 36542
rect 44158 36594 44210 36606
rect 44158 36530 44210 36542
rect 47966 36594 48018 36606
rect 47966 36530 48018 36542
rect 5742 36482 5794 36494
rect 4274 36430 4286 36482
rect 4338 36430 4350 36482
rect 5742 36418 5794 36430
rect 5854 36482 5906 36494
rect 5854 36418 5906 36430
rect 7198 36482 7250 36494
rect 7198 36418 7250 36430
rect 7646 36482 7698 36494
rect 7646 36418 7698 36430
rect 7870 36482 7922 36494
rect 7870 36418 7922 36430
rect 10782 36482 10834 36494
rect 10782 36418 10834 36430
rect 13470 36482 13522 36494
rect 18286 36482 18338 36494
rect 14802 36430 14814 36482
rect 14866 36430 14878 36482
rect 13470 36418 13522 36430
rect 18286 36418 18338 36430
rect 23774 36482 23826 36494
rect 24334 36482 24386 36494
rect 38110 36482 38162 36494
rect 24098 36430 24110 36482
rect 24162 36430 24174 36482
rect 28578 36430 28590 36482
rect 28642 36430 28654 36482
rect 29810 36430 29822 36482
rect 29874 36430 29886 36482
rect 23774 36418 23826 36430
rect 24334 36418 24386 36430
rect 38110 36418 38162 36430
rect 39342 36482 39394 36494
rect 39342 36418 39394 36430
rect 41582 36482 41634 36494
rect 41582 36418 41634 36430
rect 42142 36482 42194 36494
rect 42142 36418 42194 36430
rect 43598 36482 43650 36494
rect 45602 36430 45614 36482
rect 45666 36430 45678 36482
rect 43598 36418 43650 36430
rect 4846 36370 4898 36382
rect 4846 36306 4898 36318
rect 8318 36370 8370 36382
rect 8318 36306 8370 36318
rect 8430 36370 8482 36382
rect 8430 36306 8482 36318
rect 13582 36370 13634 36382
rect 13582 36306 13634 36318
rect 19294 36370 19346 36382
rect 19294 36306 19346 36318
rect 23326 36370 23378 36382
rect 35758 36370 35810 36382
rect 27794 36318 27806 36370
rect 27858 36318 27870 36370
rect 30594 36318 30606 36370
rect 30658 36318 30670 36370
rect 23326 36306 23378 36318
rect 35758 36306 35810 36318
rect 37774 36370 37826 36382
rect 37774 36306 37826 36318
rect 38334 36370 38386 36382
rect 38334 36306 38386 36318
rect 39230 36370 39282 36382
rect 39230 36306 39282 36318
rect 42030 36370 42082 36382
rect 42030 36306 42082 36318
rect 42814 36370 42866 36382
rect 45266 36318 45278 36370
rect 45330 36318 45342 36370
rect 42814 36306 42866 36318
rect 6302 36258 6354 36270
rect 6302 36194 6354 36206
rect 7758 36258 7810 36270
rect 7758 36194 7810 36206
rect 8654 36258 8706 36270
rect 8654 36194 8706 36206
rect 9214 36258 9266 36270
rect 9214 36194 9266 36206
rect 18062 36258 18114 36270
rect 18062 36194 18114 36206
rect 18510 36258 18562 36270
rect 18510 36194 18562 36206
rect 19182 36258 19234 36270
rect 19182 36194 19234 36206
rect 22430 36258 22482 36270
rect 22430 36194 22482 36206
rect 22654 36258 22706 36270
rect 22654 36194 22706 36206
rect 22766 36258 22818 36270
rect 22766 36194 22818 36206
rect 22878 36258 22930 36270
rect 22878 36194 22930 36206
rect 23438 36258 23490 36270
rect 23438 36194 23490 36206
rect 24222 36258 24274 36270
rect 24222 36194 24274 36206
rect 24446 36258 24498 36270
rect 24446 36194 24498 36206
rect 33182 36258 33234 36270
rect 33182 36194 33234 36206
rect 37998 36258 38050 36270
rect 37998 36194 38050 36206
rect 39118 36258 39170 36270
rect 39118 36194 39170 36206
rect 39566 36258 39618 36270
rect 39566 36194 39618 36206
rect 40126 36258 40178 36270
rect 40126 36194 40178 36206
rect 41022 36258 41074 36270
rect 44046 36258 44098 36270
rect 43362 36206 43374 36258
rect 43426 36206 43438 36258
rect 41022 36194 41074 36206
rect 44046 36194 44098 36206
rect 44270 36258 44322 36270
rect 44270 36194 44322 36206
rect 44942 36258 44994 36270
rect 44942 36194 44994 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 11566 35922 11618 35934
rect 10658 35870 10670 35922
rect 10722 35870 10734 35922
rect 10882 35870 10894 35922
rect 10946 35870 10958 35922
rect 11566 35858 11618 35870
rect 11790 35922 11842 35934
rect 14814 35922 14866 35934
rect 13794 35870 13806 35922
rect 13858 35870 13870 35922
rect 14466 35870 14478 35922
rect 14530 35870 14542 35922
rect 11790 35858 11842 35870
rect 14814 35858 14866 35870
rect 24670 35922 24722 35934
rect 24670 35858 24722 35870
rect 27022 35922 27074 35934
rect 27022 35858 27074 35870
rect 30606 35922 30658 35934
rect 30606 35858 30658 35870
rect 36878 35922 36930 35934
rect 36878 35858 36930 35870
rect 37102 35922 37154 35934
rect 37102 35858 37154 35870
rect 41582 35922 41634 35934
rect 41582 35858 41634 35870
rect 42926 35922 42978 35934
rect 44718 35922 44770 35934
rect 43250 35870 43262 35922
rect 43314 35870 43326 35922
rect 43586 35870 43598 35922
rect 43650 35870 43662 35922
rect 42926 35858 42978 35870
rect 44718 35858 44770 35870
rect 44830 35922 44882 35934
rect 44830 35858 44882 35870
rect 23214 35810 23266 35822
rect 9538 35758 9550 35810
rect 9602 35758 9614 35810
rect 19058 35758 19070 35810
rect 19122 35758 19134 35810
rect 22306 35758 22318 35810
rect 22370 35758 22382 35810
rect 22530 35758 22542 35810
rect 22594 35758 22606 35810
rect 23214 35746 23266 35758
rect 23326 35810 23378 35822
rect 23326 35746 23378 35758
rect 23774 35810 23826 35822
rect 23774 35746 23826 35758
rect 23998 35810 24050 35822
rect 23998 35746 24050 35758
rect 36654 35810 36706 35822
rect 36654 35746 36706 35758
rect 44494 35810 44546 35822
rect 46050 35758 46062 35810
rect 46114 35758 46126 35810
rect 44494 35746 44546 35758
rect 5518 35698 5570 35710
rect 8990 35698 9042 35710
rect 11902 35698 11954 35710
rect 25566 35698 25618 35710
rect 31166 35698 31218 35710
rect 42142 35698 42194 35710
rect 1810 35646 1822 35698
rect 1874 35646 1886 35698
rect 2482 35646 2494 35698
rect 2546 35646 2558 35698
rect 4946 35646 4958 35698
rect 5010 35646 5022 35698
rect 7522 35646 7534 35698
rect 7586 35646 7598 35698
rect 8754 35646 8766 35698
rect 8818 35646 8830 35698
rect 9986 35646 9998 35698
rect 10050 35646 10062 35698
rect 10546 35646 10558 35698
rect 10610 35646 10622 35698
rect 11330 35646 11342 35698
rect 11394 35646 11406 35698
rect 14018 35646 14030 35698
rect 14082 35646 14094 35698
rect 15810 35646 15822 35698
rect 15874 35646 15886 35698
rect 18386 35646 18398 35698
rect 18450 35646 18462 35698
rect 25778 35646 25790 35698
rect 25842 35646 25854 35698
rect 30370 35646 30382 35698
rect 30434 35646 30446 35698
rect 31714 35646 31726 35698
rect 31778 35646 31790 35698
rect 33394 35646 33406 35698
rect 33458 35646 33470 35698
rect 5518 35634 5570 35646
rect 8990 35634 9042 35646
rect 11902 35634 11954 35646
rect 25566 35634 25618 35646
rect 31166 35634 31218 35646
rect 42142 35634 42194 35646
rect 42590 35698 42642 35710
rect 42590 35634 42642 35646
rect 43934 35698 43986 35710
rect 43934 35634 43986 35646
rect 44942 35698 44994 35710
rect 45378 35646 45390 35698
rect 45442 35646 45454 35698
rect 44942 35634 44994 35646
rect 5182 35586 5234 35598
rect 4610 35534 4622 35586
rect 4674 35534 4686 35586
rect 5182 35522 5234 35534
rect 5966 35586 6018 35598
rect 11678 35586 11730 35598
rect 7970 35534 7982 35586
rect 8034 35534 8046 35586
rect 5966 35522 6018 35534
rect 11678 35522 11730 35534
rect 13470 35586 13522 35598
rect 13470 35522 13522 35534
rect 15262 35586 15314 35598
rect 17502 35586 17554 35598
rect 16258 35534 16270 35586
rect 16322 35534 16334 35586
rect 15262 35522 15314 35534
rect 17502 35522 17554 35534
rect 17950 35586 18002 35598
rect 26462 35586 26514 35598
rect 21186 35534 21198 35586
rect 21250 35534 21262 35586
rect 17950 35522 18002 35534
rect 26462 35522 26514 35534
rect 26798 35586 26850 35598
rect 30718 35586 30770 35598
rect 27122 35534 27134 35586
rect 27186 35534 27198 35586
rect 26798 35522 26850 35534
rect 30718 35522 30770 35534
rect 31054 35586 31106 35598
rect 31054 35522 31106 35534
rect 32510 35586 32562 35598
rect 36766 35586 36818 35598
rect 34178 35534 34190 35586
rect 34242 35534 34254 35586
rect 36306 35534 36318 35586
rect 36370 35534 36382 35586
rect 32510 35522 32562 35534
rect 36766 35522 36818 35534
rect 41134 35586 41186 35598
rect 48178 35534 48190 35586
rect 48242 35534 48254 35586
rect 41134 35522 41186 35534
rect 5406 35474 5458 35486
rect 15150 35474 15202 35486
rect 8306 35422 8318 35474
rect 8370 35422 8382 35474
rect 5406 35410 5458 35422
rect 15150 35410 15202 35422
rect 21646 35474 21698 35486
rect 21646 35410 21698 35422
rect 21982 35474 22034 35486
rect 21982 35410 22034 35422
rect 23326 35474 23378 35486
rect 23326 35410 23378 35422
rect 24334 35474 24386 35486
rect 24334 35410 24386 35422
rect 24558 35474 24610 35486
rect 24558 35410 24610 35422
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 11566 35138 11618 35150
rect 10770 35086 10782 35138
rect 10834 35086 10846 35138
rect 11566 35074 11618 35086
rect 22654 35138 22706 35150
rect 22654 35074 22706 35086
rect 22878 35138 22930 35150
rect 22878 35074 22930 35086
rect 23326 35138 23378 35150
rect 23326 35074 23378 35086
rect 41022 35138 41074 35150
rect 41022 35074 41074 35086
rect 43598 35138 43650 35150
rect 43598 35074 43650 35086
rect 1934 35026 1986 35038
rect 1934 34962 1986 34974
rect 15486 35026 15538 35038
rect 19742 35026 19794 35038
rect 16818 34974 16830 35026
rect 16882 34974 16894 35026
rect 15486 34962 15538 34974
rect 19742 34962 19794 34974
rect 22430 35026 22482 35038
rect 22430 34962 22482 34974
rect 26686 35026 26738 35038
rect 33742 35026 33794 35038
rect 32050 34974 32062 35026
rect 32114 34974 32126 35026
rect 26686 34962 26738 34974
rect 33742 34962 33794 34974
rect 34526 35026 34578 35038
rect 41470 35026 41522 35038
rect 40562 34974 40574 35026
rect 40626 34974 40638 35026
rect 34526 34962 34578 34974
rect 41470 34962 41522 34974
rect 42366 35026 42418 35038
rect 42366 34962 42418 34974
rect 42702 35026 42754 35038
rect 46946 34974 46958 35026
rect 47010 34974 47022 35026
rect 42702 34962 42754 34974
rect 4734 34914 4786 34926
rect 11790 34914 11842 34926
rect 4274 34862 4286 34914
rect 4338 34862 4350 34914
rect 8642 34862 8654 34914
rect 8706 34862 8718 34914
rect 9762 34862 9774 34914
rect 9826 34862 9838 34914
rect 11106 34862 11118 34914
rect 11170 34862 11182 34914
rect 4734 34850 4786 34862
rect 11790 34850 11842 34862
rect 12014 34914 12066 34926
rect 12014 34850 12066 34862
rect 14478 34914 14530 34926
rect 14478 34850 14530 34862
rect 14814 34914 14866 34926
rect 14814 34850 14866 34862
rect 15038 34914 15090 34926
rect 15038 34850 15090 34862
rect 15374 34914 15426 34926
rect 15374 34850 15426 34862
rect 16046 34914 16098 34926
rect 19854 34914 19906 34926
rect 25902 34914 25954 34926
rect 34638 34914 34690 34926
rect 18834 34862 18846 34914
rect 18898 34862 18910 34914
rect 24882 34862 24894 34914
rect 24946 34862 24958 34914
rect 29250 34862 29262 34914
rect 29314 34862 29326 34914
rect 32834 34862 32846 34914
rect 32898 34862 32910 34914
rect 16046 34850 16098 34862
rect 19854 34850 19906 34862
rect 25902 34850 25954 34862
rect 34638 34850 34690 34862
rect 34974 34914 35026 34926
rect 43150 34914 43202 34926
rect 37202 34862 37214 34914
rect 37266 34862 37278 34914
rect 37762 34862 37774 34914
rect 37826 34862 37838 34914
rect 34974 34850 35026 34862
rect 43150 34850 43202 34862
rect 43934 34914 43986 34926
rect 45042 34862 45054 34914
rect 45106 34862 45118 34914
rect 48066 34862 48078 34914
rect 48130 34862 48142 34914
rect 43934 34850 43986 34862
rect 12798 34802 12850 34814
rect 8754 34750 8766 34802
rect 8818 34750 8830 34802
rect 12798 34738 12850 34750
rect 12910 34802 12962 34814
rect 12910 34738 12962 34750
rect 13806 34802 13858 34814
rect 13806 34738 13858 34750
rect 24670 34802 24722 34814
rect 34414 34802 34466 34814
rect 40910 34802 40962 34814
rect 26226 34750 26238 34802
rect 26290 34750 26302 34802
rect 29922 34750 29934 34802
rect 29986 34750 29998 34802
rect 32610 34750 32622 34802
rect 32674 34750 32686 34802
rect 38434 34750 38446 34802
rect 38498 34750 38510 34802
rect 24670 34738 24722 34750
rect 34414 34738 34466 34750
rect 40910 34738 40962 34750
rect 43486 34802 43538 34814
rect 43486 34738 43538 34750
rect 44270 34802 44322 34814
rect 44270 34738 44322 34750
rect 45278 34802 45330 34814
rect 45278 34738 45330 34750
rect 12126 34690 12178 34702
rect 12126 34626 12178 34638
rect 12238 34690 12290 34702
rect 12238 34626 12290 34638
rect 12574 34690 12626 34702
rect 12574 34626 12626 34638
rect 13694 34690 13746 34702
rect 13694 34626 13746 34638
rect 14702 34690 14754 34702
rect 14702 34626 14754 34638
rect 15598 34690 15650 34702
rect 15598 34626 15650 34638
rect 19406 34690 19458 34702
rect 19406 34626 19458 34638
rect 19630 34690 19682 34702
rect 19630 34626 19682 34638
rect 20414 34690 20466 34702
rect 20414 34626 20466 34638
rect 20750 34690 20802 34702
rect 20750 34626 20802 34638
rect 33854 34690 33906 34702
rect 36978 34638 36990 34690
rect 37042 34638 37054 34690
rect 33854 34626 33906 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 2046 34354 2098 34366
rect 2046 34290 2098 34302
rect 2494 34354 2546 34366
rect 7310 34354 7362 34366
rect 20750 34354 20802 34366
rect 44718 34354 44770 34366
rect 6850 34302 6862 34354
rect 6914 34302 6926 34354
rect 7634 34302 7646 34354
rect 7698 34302 7710 34354
rect 37426 34302 37438 34354
rect 37490 34302 37502 34354
rect 2494 34290 2546 34302
rect 7310 34290 7362 34302
rect 20750 34290 20802 34302
rect 44718 34290 44770 34302
rect 45838 34354 45890 34366
rect 47842 34302 47854 34354
rect 47906 34302 47918 34354
rect 45838 34290 45890 34302
rect 1710 34242 1762 34254
rect 1710 34178 1762 34190
rect 10558 34242 10610 34254
rect 10558 34178 10610 34190
rect 11006 34242 11058 34254
rect 31054 34242 31106 34254
rect 47294 34242 47346 34254
rect 15138 34190 15150 34242
rect 15202 34190 15214 34242
rect 31714 34190 31726 34242
rect 31778 34190 31790 34242
rect 11006 34178 11058 34190
rect 31054 34178 31106 34190
rect 47294 34178 47346 34190
rect 10110 34130 10162 34142
rect 31390 34130 31442 34142
rect 3938 34078 3950 34130
rect 4002 34078 4014 34130
rect 10770 34078 10782 34130
rect 10834 34078 10846 34130
rect 12002 34078 12014 34130
rect 12066 34078 12078 34130
rect 13010 34078 13022 34130
rect 13074 34078 13086 34130
rect 13458 34078 13470 34130
rect 13522 34078 13534 34130
rect 13682 34078 13694 34130
rect 13746 34078 13758 34130
rect 16258 34078 16270 34130
rect 16322 34078 16334 34130
rect 18274 34078 18286 34130
rect 18338 34078 18350 34130
rect 10110 34066 10162 34078
rect 31390 34066 31442 34078
rect 32062 34130 32114 34142
rect 32062 34066 32114 34078
rect 33406 34130 33458 34142
rect 33406 34066 33458 34078
rect 33630 34130 33682 34142
rect 45726 34130 45778 34142
rect 37202 34078 37214 34130
rect 37266 34078 37278 34130
rect 37762 34078 37774 34130
rect 37826 34078 37838 34130
rect 41458 34078 41470 34130
rect 41522 34078 41534 34130
rect 44930 34078 44942 34130
rect 44994 34078 45006 34130
rect 45378 34078 45390 34130
rect 45442 34078 45454 34130
rect 33630 34066 33682 34078
rect 45726 34066 45778 34078
rect 45950 34130 46002 34142
rect 45950 34066 46002 34078
rect 46286 34130 46338 34142
rect 46286 34066 46338 34078
rect 46622 34130 46674 34142
rect 46622 34066 46674 34078
rect 46734 34130 46786 34142
rect 46734 34066 46786 34078
rect 47518 34130 47570 34142
rect 47518 34066 47570 34078
rect 8094 34018 8146 34030
rect 14926 34018 14978 34030
rect 33182 34018 33234 34030
rect 4610 33966 4622 34018
rect 4674 33966 4686 34018
rect 11106 33966 11118 34018
rect 11170 33966 11182 34018
rect 18834 33966 18846 34018
rect 18898 33966 18910 34018
rect 8094 33954 8146 33966
rect 14926 33954 14978 33966
rect 33182 33954 33234 33966
rect 36766 34018 36818 34030
rect 46398 34018 46450 34030
rect 40114 33966 40126 34018
rect 40178 33966 40190 34018
rect 42130 33966 42142 34018
rect 42194 33966 42206 34018
rect 44258 33966 44270 34018
rect 44322 33966 44334 34018
rect 36766 33954 36818 33966
rect 46398 33954 46450 33966
rect 10222 33906 10274 33918
rect 10222 33842 10274 33854
rect 34078 33906 34130 33918
rect 34078 33842 34130 33854
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 9214 33570 9266 33582
rect 9214 33506 9266 33518
rect 9886 33570 9938 33582
rect 9886 33506 9938 33518
rect 11454 33570 11506 33582
rect 11454 33506 11506 33518
rect 24558 33570 24610 33582
rect 24558 33506 24610 33518
rect 34414 33570 34466 33582
rect 34414 33506 34466 33518
rect 44942 33570 44994 33582
rect 44942 33506 44994 33518
rect 7422 33458 7474 33470
rect 7422 33394 7474 33406
rect 11230 33458 11282 33470
rect 20414 33458 20466 33470
rect 12898 33406 12910 33458
rect 12962 33406 12974 33458
rect 17154 33406 17166 33458
rect 17218 33406 17230 33458
rect 11230 33394 11282 33406
rect 20414 33394 20466 33406
rect 23102 33458 23154 33470
rect 26462 33458 26514 33470
rect 25890 33406 25902 33458
rect 25954 33406 25966 33458
rect 23102 33394 23154 33406
rect 26462 33394 26514 33406
rect 29598 33458 29650 33470
rect 37998 33458 38050 33470
rect 30930 33406 30942 33458
rect 30994 33406 31006 33458
rect 32498 33406 32510 33458
rect 32562 33406 32574 33458
rect 29598 33394 29650 33406
rect 37998 33394 38050 33406
rect 38446 33458 38498 33470
rect 42254 33458 42306 33470
rect 41570 33406 41582 33458
rect 41634 33406 41646 33458
rect 46050 33406 46062 33458
rect 46114 33406 46126 33458
rect 48178 33406 48190 33458
rect 48242 33406 48254 33458
rect 38446 33394 38498 33406
rect 42254 33394 42306 33406
rect 5742 33346 5794 33358
rect 8430 33346 8482 33358
rect 1810 33294 1822 33346
rect 1874 33294 1886 33346
rect 6290 33294 6302 33346
rect 6354 33294 6366 33346
rect 5742 33282 5794 33294
rect 8430 33282 8482 33294
rect 8766 33346 8818 33358
rect 8766 33282 8818 33294
rect 9102 33346 9154 33358
rect 9102 33282 9154 33294
rect 9998 33346 10050 33358
rect 9998 33282 10050 33294
rect 10222 33346 10274 33358
rect 10222 33282 10274 33294
rect 12126 33346 12178 33358
rect 12126 33282 12178 33294
rect 13694 33346 13746 33358
rect 13694 33282 13746 33294
rect 14366 33346 14418 33358
rect 19518 33346 19570 33358
rect 17938 33294 17950 33346
rect 18002 33294 18014 33346
rect 14366 33282 14418 33294
rect 19518 33282 19570 33294
rect 20078 33346 20130 33358
rect 27806 33346 27858 33358
rect 24098 33294 24110 33346
rect 24162 33294 24174 33346
rect 26002 33294 26014 33346
rect 26066 33294 26078 33346
rect 20078 33282 20130 33294
rect 27806 33282 27858 33294
rect 29150 33346 29202 33358
rect 29150 33282 29202 33294
rect 29486 33346 29538 33358
rect 34750 33346 34802 33358
rect 33618 33294 33630 33346
rect 33682 33294 33694 33346
rect 29486 33282 29538 33294
rect 34750 33282 34802 33294
rect 34974 33346 35026 33358
rect 34974 33282 35026 33294
rect 36318 33346 36370 33358
rect 36318 33282 36370 33294
rect 38222 33346 38274 33358
rect 38222 33282 38274 33294
rect 38670 33346 38722 33358
rect 42366 33346 42418 33358
rect 39218 33294 39230 33346
rect 39282 33294 39294 33346
rect 38670 33282 38722 33294
rect 42366 33282 42418 33294
rect 42702 33346 42754 33358
rect 42702 33282 42754 33294
rect 43374 33346 43426 33358
rect 43374 33282 43426 33294
rect 43486 33346 43538 33358
rect 43486 33282 43538 33294
rect 43934 33346 43986 33358
rect 43934 33282 43986 33294
rect 44830 33346 44882 33358
rect 45378 33294 45390 33346
rect 45442 33294 45454 33346
rect 44830 33282 44882 33294
rect 5630 33234 5682 33246
rect 2482 33182 2494 33234
rect 2546 33182 2558 33234
rect 5630 33170 5682 33182
rect 8206 33234 8258 33246
rect 8206 33170 8258 33182
rect 12350 33234 12402 33246
rect 12350 33170 12402 33182
rect 12462 33234 12514 33246
rect 13918 33234 13970 33246
rect 12562 33182 12574 33234
rect 12626 33182 12638 33234
rect 12462 33170 12514 33182
rect 13918 33170 13970 33182
rect 19630 33234 19682 33246
rect 19630 33170 19682 33182
rect 23214 33234 23266 33246
rect 23214 33170 23266 33182
rect 24558 33234 24610 33246
rect 24558 33170 24610 33182
rect 24670 33234 24722 33246
rect 25342 33234 25394 33246
rect 24994 33182 25006 33234
rect 25058 33182 25070 33234
rect 24670 33170 24722 33182
rect 25342 33170 25394 33182
rect 25678 33234 25730 33246
rect 29710 33234 29762 33246
rect 27122 33182 27134 33234
rect 27186 33182 27198 33234
rect 27458 33182 27470 33234
rect 27522 33182 27534 33234
rect 25678 33170 25730 33182
rect 29710 33170 29762 33182
rect 30606 33234 30658 33246
rect 30606 33170 30658 33182
rect 30830 33234 30882 33246
rect 30830 33170 30882 33182
rect 34302 33234 34354 33246
rect 34302 33170 34354 33182
rect 35310 33234 35362 33246
rect 35310 33170 35362 33182
rect 35534 33234 35586 33246
rect 35534 33170 35586 33182
rect 35870 33234 35922 33246
rect 35870 33170 35922 33182
rect 36206 33234 36258 33246
rect 36206 33170 36258 33182
rect 38894 33234 38946 33246
rect 38894 33170 38946 33182
rect 42142 33234 42194 33246
rect 42142 33170 42194 33182
rect 7310 33122 7362 33134
rect 4722 33070 4734 33122
rect 4786 33070 4798 33122
rect 7310 33058 7362 33070
rect 8654 33122 8706 33134
rect 8654 33058 8706 33070
rect 9886 33122 9938 33134
rect 9886 33058 9938 33070
rect 10894 33122 10946 33134
rect 14030 33122 14082 33134
rect 18398 33122 18450 33134
rect 11778 33070 11790 33122
rect 11842 33070 11854 33122
rect 14914 33070 14926 33122
rect 14978 33070 14990 33122
rect 10894 33058 10946 33070
rect 14030 33058 14082 33070
rect 18398 33058 18450 33070
rect 19182 33122 19234 33134
rect 19182 33058 19234 33070
rect 19406 33122 19458 33134
rect 19406 33058 19458 33070
rect 22990 33122 23042 33134
rect 22990 33058 23042 33070
rect 23550 33122 23602 33134
rect 23550 33058 23602 33070
rect 23662 33122 23714 33134
rect 23662 33058 23714 33070
rect 23774 33122 23826 33134
rect 23774 33058 23826 33070
rect 26350 33122 26402 33134
rect 26350 33058 26402 33070
rect 26798 33122 26850 33134
rect 26798 33058 26850 33070
rect 30270 33122 30322 33134
rect 30270 33058 30322 33070
rect 31054 33122 31106 33134
rect 31054 33058 31106 33070
rect 34526 33122 34578 33134
rect 34526 33058 34578 33070
rect 35758 33122 35810 33134
rect 35758 33058 35810 33070
rect 43262 33122 43314 33134
rect 43262 33058 43314 33070
rect 44270 33122 44322 33134
rect 44270 33058 44322 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 2942 32786 2994 32798
rect 7758 32786 7810 32798
rect 4946 32734 4958 32786
rect 5010 32734 5022 32786
rect 2942 32722 2994 32734
rect 7758 32722 7810 32734
rect 9886 32786 9938 32798
rect 9886 32722 9938 32734
rect 11006 32786 11058 32798
rect 11006 32722 11058 32734
rect 22206 32786 22258 32798
rect 22206 32722 22258 32734
rect 22430 32786 22482 32798
rect 22430 32722 22482 32734
rect 23774 32786 23826 32798
rect 27134 32786 27186 32798
rect 25778 32734 25790 32786
rect 25842 32734 25854 32786
rect 23774 32722 23826 32734
rect 27134 32722 27186 32734
rect 29710 32786 29762 32798
rect 29710 32722 29762 32734
rect 38222 32786 38274 32798
rect 38222 32722 38274 32734
rect 38894 32786 38946 32798
rect 39790 32786 39842 32798
rect 39218 32734 39230 32786
rect 39282 32734 39294 32786
rect 38894 32722 38946 32734
rect 39790 32722 39842 32734
rect 39902 32786 39954 32798
rect 39902 32722 39954 32734
rect 40014 32786 40066 32798
rect 40014 32722 40066 32734
rect 41806 32786 41858 32798
rect 44046 32786 44098 32798
rect 43698 32734 43710 32786
rect 43762 32734 43774 32786
rect 41806 32722 41858 32734
rect 44046 32722 44098 32734
rect 45614 32786 45666 32798
rect 45614 32722 45666 32734
rect 45950 32786 46002 32798
rect 45950 32722 46002 32734
rect 46174 32786 46226 32798
rect 46174 32722 46226 32734
rect 46846 32786 46898 32798
rect 46846 32722 46898 32734
rect 5854 32674 5906 32686
rect 5854 32610 5906 32622
rect 5966 32674 6018 32686
rect 8430 32674 8482 32686
rect 8194 32622 8206 32674
rect 8258 32622 8270 32674
rect 5966 32610 6018 32622
rect 8430 32610 8482 32622
rect 10446 32674 10498 32686
rect 10446 32610 10498 32622
rect 10782 32674 10834 32686
rect 14814 32674 14866 32686
rect 11778 32622 11790 32674
rect 11842 32622 11854 32674
rect 10782 32610 10834 32622
rect 14814 32610 14866 32622
rect 15934 32674 15986 32686
rect 15934 32610 15986 32622
rect 16606 32674 16658 32686
rect 23102 32674 23154 32686
rect 17378 32622 17390 32674
rect 17442 32622 17454 32674
rect 19282 32622 19294 32674
rect 19346 32622 19358 32674
rect 16606 32610 16658 32622
rect 23102 32610 23154 32622
rect 23662 32674 23714 32686
rect 40910 32674 40962 32686
rect 26786 32622 26798 32674
rect 26850 32622 26862 32674
rect 36978 32622 36990 32674
rect 37042 32622 37054 32674
rect 38546 32622 38558 32674
rect 38610 32622 38622 32674
rect 23662 32610 23714 32622
rect 40910 32610 40962 32622
rect 45502 32674 45554 32686
rect 45502 32610 45554 32622
rect 47630 32674 47682 32686
rect 47630 32610 47682 32622
rect 47966 32674 48018 32686
rect 47966 32610 48018 32622
rect 5294 32562 5346 32574
rect 7198 32562 7250 32574
rect 16718 32562 16770 32574
rect 22878 32562 22930 32574
rect 5618 32510 5630 32562
rect 5682 32510 5694 32562
rect 8642 32510 8654 32562
rect 8706 32510 8718 32562
rect 13234 32510 13246 32562
rect 13298 32510 13310 32562
rect 13682 32510 13694 32562
rect 13746 32510 13758 32562
rect 17602 32510 17614 32562
rect 17666 32510 17678 32562
rect 18610 32510 18622 32562
rect 18674 32510 18686 32562
rect 5294 32498 5346 32510
rect 7198 32498 7250 32510
rect 16718 32498 16770 32510
rect 22878 32498 22930 32510
rect 24110 32562 24162 32574
rect 24110 32498 24162 32510
rect 25230 32562 25282 32574
rect 25230 32498 25282 32510
rect 28478 32562 28530 32574
rect 33294 32562 33346 32574
rect 40462 32562 40514 32574
rect 29922 32510 29934 32562
rect 29986 32510 29998 32562
rect 33506 32510 33518 32562
rect 33570 32510 33582 32562
rect 37650 32510 37662 32562
rect 37714 32510 37726 32562
rect 28478 32498 28530 32510
rect 33294 32498 33346 32510
rect 40462 32498 40514 32510
rect 41134 32562 41186 32574
rect 41134 32498 41186 32510
rect 41358 32562 41410 32574
rect 41358 32498 41410 32510
rect 41918 32562 41970 32574
rect 41918 32498 41970 32510
rect 42030 32562 42082 32574
rect 42354 32510 42366 32562
rect 42418 32510 42430 32562
rect 46498 32510 46510 32562
rect 46562 32510 46574 32562
rect 47058 32510 47070 32562
rect 47122 32510 47134 32562
rect 42030 32498 42082 32510
rect 3166 32450 3218 32462
rect 2818 32398 2830 32450
rect 2882 32398 2894 32450
rect 3166 32386 3218 32398
rect 3614 32450 3666 32462
rect 3614 32386 3666 32398
rect 4622 32450 4674 32462
rect 4622 32386 4674 32398
rect 6414 32450 6466 32462
rect 6414 32386 6466 32398
rect 8094 32450 8146 32462
rect 13470 32450 13522 32462
rect 10210 32398 10222 32450
rect 10274 32398 10286 32450
rect 11106 32398 11118 32450
rect 11170 32398 11182 32450
rect 8094 32386 8146 32398
rect 13470 32386 13522 32398
rect 18174 32450 18226 32462
rect 22318 32450 22370 32462
rect 21410 32398 21422 32450
rect 21474 32398 21486 32450
rect 18174 32386 18226 32398
rect 22318 32386 22370 32398
rect 25454 32450 25506 32462
rect 25454 32386 25506 32398
rect 28814 32450 28866 32462
rect 33070 32450 33122 32462
rect 41022 32450 41074 32462
rect 31042 32398 31054 32450
rect 31106 32398 31118 32450
rect 34850 32398 34862 32450
rect 34914 32398 34926 32450
rect 28814 32386 28866 32398
rect 33070 32386 33122 32398
rect 41022 32386 41074 32398
rect 42702 32450 42754 32462
rect 42702 32386 42754 32398
rect 42814 32450 42866 32462
rect 42814 32386 42866 32398
rect 45166 32450 45218 32462
rect 45166 32386 45218 32398
rect 46062 32450 46114 32462
rect 46062 32386 46114 32398
rect 9102 32338 9154 32350
rect 9102 32274 9154 32286
rect 15822 32338 15874 32350
rect 15822 32274 15874 32286
rect 16158 32338 16210 32350
rect 16158 32274 16210 32286
rect 16606 32338 16658 32350
rect 16606 32274 16658 32286
rect 23214 32338 23266 32350
rect 23214 32274 23266 32286
rect 24334 32338 24386 32350
rect 29038 32338 29090 32350
rect 24658 32286 24670 32338
rect 24722 32286 24734 32338
rect 24334 32274 24386 32286
rect 29038 32274 29090 32286
rect 29262 32338 29314 32350
rect 29262 32274 29314 32286
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 19406 32002 19458 32014
rect 19406 31938 19458 31950
rect 19742 32002 19794 32014
rect 19742 31938 19794 31950
rect 31502 32002 31554 32014
rect 31502 31938 31554 31950
rect 3614 31890 3666 31902
rect 9214 31890 9266 31902
rect 30158 31890 30210 31902
rect 3266 31838 3278 31890
rect 3330 31838 3342 31890
rect 8530 31838 8542 31890
rect 8594 31838 8606 31890
rect 11106 31838 11118 31890
rect 11170 31838 11182 31890
rect 3614 31826 3666 31838
rect 9214 31826 9266 31838
rect 30158 31826 30210 31838
rect 34974 31890 35026 31902
rect 34974 31826 35026 31838
rect 37102 31890 37154 31902
rect 37102 31826 37154 31838
rect 38110 31890 38162 31902
rect 39890 31838 39902 31890
rect 39954 31838 39966 31890
rect 42018 31838 42030 31890
rect 42082 31838 42094 31890
rect 44146 31838 44158 31890
rect 44210 31838 44222 31890
rect 48178 31838 48190 31890
rect 48242 31838 48254 31890
rect 38110 31826 38162 31838
rect 9438 31778 9490 31790
rect 18510 31778 18562 31790
rect 5730 31726 5742 31778
rect 5794 31726 5806 31778
rect 8978 31726 8990 31778
rect 9042 31726 9054 31778
rect 10546 31726 10558 31778
rect 10610 31726 10622 31778
rect 13682 31726 13694 31778
rect 13746 31726 13758 31778
rect 14354 31726 14366 31778
rect 14418 31726 14430 31778
rect 18162 31726 18174 31778
rect 18226 31726 18238 31778
rect 9438 31714 9490 31726
rect 18510 31714 18562 31726
rect 19518 31778 19570 31790
rect 19518 31714 19570 31726
rect 19854 31778 19906 31790
rect 19854 31714 19906 31726
rect 20302 31778 20354 31790
rect 29710 31778 29762 31790
rect 31166 31778 31218 31790
rect 23202 31726 23214 31778
rect 23266 31726 23278 31778
rect 30594 31726 30606 31778
rect 30658 31726 30670 31778
rect 20302 31714 20354 31726
rect 29710 31714 29762 31726
rect 31166 31714 31218 31726
rect 31390 31778 31442 31790
rect 31390 31714 31442 31726
rect 31614 31778 31666 31790
rect 31614 31714 31666 31726
rect 33070 31778 33122 31790
rect 34078 31778 34130 31790
rect 33730 31726 33742 31778
rect 33794 31726 33806 31778
rect 33070 31714 33122 31726
rect 34078 31714 34130 31726
rect 35534 31778 35586 31790
rect 39106 31726 39118 31778
rect 39170 31726 39182 31778
rect 43810 31726 43822 31778
rect 43874 31726 43886 31778
rect 45378 31726 45390 31778
rect 45442 31726 45454 31778
rect 35534 31714 35586 31726
rect 19070 31666 19122 31678
rect 30942 31666 30994 31678
rect 33966 31666 34018 31678
rect 6402 31614 6414 31666
rect 6466 31614 6478 31666
rect 14466 31614 14478 31666
rect 14530 31614 14542 31666
rect 18050 31614 18062 31666
rect 18114 31614 18126 31666
rect 21298 31614 21310 31666
rect 21362 31614 21374 31666
rect 23314 31614 23326 31666
rect 23378 31614 23390 31666
rect 29026 31614 29038 31666
rect 29090 31663 29102 31666
rect 29250 31663 29262 31666
rect 29090 31617 29262 31663
rect 29090 31614 29102 31617
rect 29250 31614 29262 31617
rect 29314 31614 29326 31666
rect 32050 31614 32062 31666
rect 32114 31614 32126 31666
rect 32834 31614 32846 31666
rect 32898 31614 32910 31666
rect 19070 31602 19122 31614
rect 30942 31602 30994 31614
rect 33966 31602 34018 31614
rect 42590 31666 42642 31678
rect 42590 31602 42642 31614
rect 42926 31666 42978 31678
rect 42926 31602 42978 31614
rect 43262 31666 43314 31678
rect 46050 31614 46062 31666
rect 46114 31614 46126 31666
rect 43262 31602 43314 31614
rect 3390 31554 3442 31566
rect 3390 31490 3442 31502
rect 9102 31554 9154 31566
rect 9102 31490 9154 31502
rect 13694 31554 13746 31566
rect 21646 31554 21698 31566
rect 15362 31502 15374 31554
rect 15426 31502 15438 31554
rect 20626 31502 20638 31554
rect 20690 31502 20702 31554
rect 13694 31490 13746 31502
rect 21646 31490 21698 31502
rect 22094 31554 22146 31566
rect 29486 31554 29538 31566
rect 23650 31502 23662 31554
rect 23714 31502 23726 31554
rect 22094 31490 22146 31502
rect 29486 31490 29538 31502
rect 29598 31554 29650 31566
rect 29598 31490 29650 31502
rect 30046 31554 30098 31566
rect 30046 31490 30098 31502
rect 30270 31554 30322 31566
rect 34862 31554 34914 31566
rect 32498 31502 32510 31554
rect 32562 31502 32574 31554
rect 34514 31502 34526 31554
rect 34578 31502 34590 31554
rect 30270 31490 30322 31502
rect 34862 31490 34914 31502
rect 35086 31554 35138 31566
rect 35086 31490 35138 31502
rect 36318 31554 36370 31566
rect 36318 31490 36370 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 7198 31218 7250 31230
rect 7198 31154 7250 31166
rect 8430 31218 8482 31230
rect 8430 31154 8482 31166
rect 12910 31218 12962 31230
rect 12910 31154 12962 31166
rect 15262 31218 15314 31230
rect 15262 31154 15314 31166
rect 15374 31218 15426 31230
rect 15374 31154 15426 31166
rect 15598 31218 15650 31230
rect 15598 31154 15650 31166
rect 22654 31218 22706 31230
rect 22654 31154 22706 31166
rect 24558 31218 24610 31230
rect 24558 31154 24610 31166
rect 26238 31218 26290 31230
rect 29262 31218 29314 31230
rect 27122 31166 27134 31218
rect 27186 31166 27198 31218
rect 26238 31154 26290 31166
rect 29262 31154 29314 31166
rect 30158 31218 30210 31230
rect 30158 31154 30210 31166
rect 30830 31218 30882 31230
rect 30830 31154 30882 31166
rect 37886 31218 37938 31230
rect 37886 31154 37938 31166
rect 44718 31218 44770 31230
rect 44718 31154 44770 31166
rect 45726 31218 45778 31230
rect 45726 31154 45778 31166
rect 46622 31218 46674 31230
rect 46622 31154 46674 31166
rect 47070 31218 47122 31230
rect 47070 31154 47122 31166
rect 47518 31218 47570 31230
rect 47518 31154 47570 31166
rect 48190 31218 48242 31230
rect 48190 31154 48242 31166
rect 7422 31106 7474 31118
rect 7422 31042 7474 31054
rect 8766 31106 8818 31118
rect 8766 31042 8818 31054
rect 8990 31106 9042 31118
rect 15038 31106 15090 31118
rect 13570 31054 13582 31106
rect 13634 31054 13646 31106
rect 13794 31054 13806 31106
rect 13858 31054 13870 31106
rect 8990 31042 9042 31054
rect 15038 31042 15090 31054
rect 15486 31106 15538 31118
rect 15486 31042 15538 31054
rect 21758 31106 21810 31118
rect 21758 31042 21810 31054
rect 21982 31106 22034 31118
rect 21982 31042 22034 31054
rect 23326 31106 23378 31118
rect 23326 31042 23378 31054
rect 23886 31106 23938 31118
rect 23886 31042 23938 31054
rect 27470 31106 27522 31118
rect 27470 31042 27522 31054
rect 35758 31106 35810 31118
rect 35758 31042 35810 31054
rect 35982 31106 36034 31118
rect 35982 31042 36034 31054
rect 36094 31106 36146 31118
rect 36878 31106 36930 31118
rect 36642 31054 36654 31106
rect 36706 31054 36718 31106
rect 36094 31042 36146 31054
rect 36878 31042 36930 31054
rect 37998 31106 38050 31118
rect 45502 31106 45554 31118
rect 45042 31054 45054 31106
rect 45106 31054 45118 31106
rect 37998 31042 38050 31054
rect 45502 31042 45554 31054
rect 46062 31106 46114 31118
rect 46062 31042 46114 31054
rect 7534 30994 7586 31006
rect 20974 30994 21026 31006
rect 1810 30942 1822 30994
rect 1874 30942 1886 30994
rect 11890 30942 11902 30994
rect 11954 30942 11966 30994
rect 13346 30942 13358 30994
rect 13410 30942 13422 30994
rect 16594 30942 16606 30994
rect 16658 30942 16670 30994
rect 17602 30942 17614 30994
rect 17666 30942 17678 30994
rect 18722 30942 18734 30994
rect 18786 30942 18798 30994
rect 20738 30942 20750 30994
rect 20802 30942 20814 30994
rect 7534 30930 7586 30942
rect 20974 30930 21026 30942
rect 21422 30994 21474 31006
rect 21422 30930 21474 30942
rect 22318 30994 22370 31006
rect 22318 30930 22370 30942
rect 22878 30994 22930 31006
rect 22878 30930 22930 30942
rect 23438 30994 23490 31006
rect 24670 30994 24722 31006
rect 24210 30942 24222 30994
rect 24274 30942 24286 30994
rect 23438 30930 23490 30942
rect 24670 30930 24722 30942
rect 26574 30994 26626 31006
rect 29374 30994 29426 31006
rect 27682 30942 27694 30994
rect 27746 30942 27758 30994
rect 26574 30930 26626 30942
rect 29374 30930 29426 30942
rect 29934 30994 29986 31006
rect 29934 30930 29986 30942
rect 30382 30994 30434 31006
rect 37550 30994 37602 31006
rect 31042 30942 31054 30994
rect 31106 30942 31118 30994
rect 37090 30942 37102 30994
rect 37154 30942 37166 30994
rect 30382 30930 30434 30942
rect 37550 30930 37602 30942
rect 45726 30994 45778 31006
rect 45726 30930 45778 30942
rect 8878 30882 8930 30894
rect 14478 30882 14530 30894
rect 2482 30830 2494 30882
rect 2546 30830 2558 30882
rect 4610 30830 4622 30882
rect 4674 30830 4686 30882
rect 10098 30830 10110 30882
rect 10162 30830 10174 30882
rect 8878 30818 8930 30830
rect 14478 30818 14530 30830
rect 16158 30882 16210 30894
rect 16158 30818 16210 30830
rect 23102 30882 23154 30894
rect 26798 30882 26850 30894
rect 24098 30830 24110 30882
rect 24162 30830 24174 30882
rect 23102 30818 23154 30830
rect 26798 30818 26850 30830
rect 30270 30882 30322 30894
rect 30270 30818 30322 30830
rect 36542 30882 36594 30894
rect 36542 30818 36594 30830
rect 16718 30770 16770 30782
rect 22542 30770 22594 30782
rect 18050 30718 18062 30770
rect 18114 30718 18126 30770
rect 16718 30706 16770 30718
rect 22542 30706 22594 30718
rect 29262 30770 29314 30782
rect 29262 30706 29314 30718
rect 29710 30770 29762 30782
rect 29710 30706 29762 30718
rect 36094 30770 36146 30782
rect 36094 30706 36146 30718
rect 37774 30770 37826 30782
rect 37774 30706 37826 30718
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 2718 30434 2770 30446
rect 2718 30370 2770 30382
rect 2830 30434 2882 30446
rect 2830 30370 2882 30382
rect 3054 30434 3106 30446
rect 3054 30370 3106 30382
rect 4622 30434 4674 30446
rect 30382 30434 30434 30446
rect 35646 30434 35698 30446
rect 15026 30382 15038 30434
rect 15090 30382 15102 30434
rect 34178 30382 34190 30434
rect 34242 30382 34254 30434
rect 4622 30370 4674 30382
rect 30382 30370 30434 30382
rect 35646 30370 35698 30382
rect 13918 30322 13970 30334
rect 25342 30322 25394 30334
rect 12674 30270 12686 30322
rect 12738 30270 12750 30322
rect 14914 30270 14926 30322
rect 14978 30270 14990 30322
rect 16034 30270 16046 30322
rect 16098 30270 16110 30322
rect 22306 30270 22318 30322
rect 22370 30270 22382 30322
rect 24434 30270 24446 30322
rect 24498 30270 24510 30322
rect 13918 30258 13970 30270
rect 25342 30258 25394 30270
rect 33294 30322 33346 30334
rect 42130 30270 42142 30322
rect 42194 30270 42206 30322
rect 33294 30258 33346 30270
rect 4846 30210 4898 30222
rect 16942 30210 16994 30222
rect 3266 30158 3278 30210
rect 3330 30158 3342 30210
rect 9874 30158 9886 30210
rect 9938 30158 9950 30210
rect 14690 30158 14702 30210
rect 14754 30158 14766 30210
rect 15922 30158 15934 30210
rect 15986 30158 15998 30210
rect 4846 30146 4898 30158
rect 16942 30146 16994 30158
rect 17614 30210 17666 30222
rect 17614 30146 17666 30158
rect 18062 30210 18114 30222
rect 25118 30210 25170 30222
rect 30494 30210 30546 30222
rect 21634 30158 21646 30210
rect 21698 30158 21710 30210
rect 25666 30158 25678 30210
rect 25730 30158 25742 30210
rect 18062 30146 18114 30158
rect 25118 30146 25170 30158
rect 30494 30146 30546 30158
rect 32510 30210 32562 30222
rect 32510 30146 32562 30158
rect 32846 30210 32898 30222
rect 37214 30210 37266 30222
rect 33730 30158 33742 30210
rect 33794 30158 33806 30210
rect 35298 30158 35310 30210
rect 35362 30158 35374 30210
rect 36978 30158 36990 30210
rect 37042 30158 37054 30210
rect 38770 30158 38782 30210
rect 38834 30158 38846 30210
rect 32846 30146 32898 30158
rect 37214 30146 37266 30158
rect 13806 30098 13858 30110
rect 5954 30046 5966 30098
rect 6018 30046 6030 30098
rect 10546 30046 10558 30098
rect 10610 30046 10622 30098
rect 13806 30034 13858 30046
rect 14030 30098 14082 30110
rect 14030 30034 14082 30046
rect 17950 30098 18002 30110
rect 17950 30034 18002 30046
rect 18398 30098 18450 30110
rect 18398 30034 18450 30046
rect 18734 30098 18786 30110
rect 18734 30034 18786 30046
rect 19070 30098 19122 30110
rect 36094 30098 36146 30110
rect 31490 30046 31502 30098
rect 31554 30046 31566 30098
rect 32162 30046 32174 30098
rect 32226 30046 32238 30098
rect 34626 30046 34638 30098
rect 34690 30046 34702 30098
rect 35858 30046 35870 30098
rect 35922 30046 35934 30098
rect 19070 30034 19122 30046
rect 36094 30034 36146 30046
rect 37662 30098 37714 30110
rect 42254 30098 42306 30110
rect 39442 30046 39454 30098
rect 39506 30046 39518 30098
rect 37662 30034 37714 30046
rect 42254 30034 42306 30046
rect 42478 30098 42530 30110
rect 42478 30034 42530 30046
rect 5630 29986 5682 29998
rect 4274 29934 4286 29986
rect 4338 29934 4350 29986
rect 5630 29922 5682 29934
rect 9438 29986 9490 29998
rect 18510 29986 18562 29998
rect 17266 29934 17278 29986
rect 17330 29934 17342 29986
rect 9438 29922 9490 29934
rect 18510 29922 18562 29934
rect 19182 29986 19234 29998
rect 19182 29922 19234 29934
rect 19406 29986 19458 29998
rect 19406 29922 19458 29934
rect 19742 29986 19794 29998
rect 26574 29986 26626 29998
rect 26226 29934 26238 29986
rect 26290 29934 26302 29986
rect 19742 29922 19794 29934
rect 26574 29922 26626 29934
rect 30382 29986 30434 29998
rect 30382 29922 30434 29934
rect 31838 29986 31890 29998
rect 31838 29922 31890 29934
rect 35982 29986 36034 29998
rect 35982 29922 36034 29934
rect 37326 29986 37378 29998
rect 37326 29922 37378 29934
rect 37438 29986 37490 29998
rect 44158 29986 44210 29998
rect 41682 29934 41694 29986
rect 41746 29934 41758 29986
rect 37438 29922 37490 29934
rect 44158 29922 44210 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 10334 29650 10386 29662
rect 10334 29586 10386 29598
rect 12686 29650 12738 29662
rect 12686 29586 12738 29598
rect 13582 29650 13634 29662
rect 13582 29586 13634 29598
rect 14814 29650 14866 29662
rect 14814 29586 14866 29598
rect 15598 29650 15650 29662
rect 15598 29586 15650 29598
rect 17950 29650 18002 29662
rect 17950 29586 18002 29598
rect 32174 29650 32226 29662
rect 32174 29586 32226 29598
rect 33070 29650 33122 29662
rect 34862 29650 34914 29662
rect 34514 29598 34526 29650
rect 34578 29598 34590 29650
rect 33070 29586 33122 29598
rect 34862 29586 34914 29598
rect 38558 29650 38610 29662
rect 44034 29598 44046 29650
rect 44098 29598 44110 29650
rect 38558 29586 38610 29598
rect 17502 29538 17554 29550
rect 11442 29486 11454 29538
rect 11506 29486 11518 29538
rect 16146 29486 16158 29538
rect 16210 29486 16222 29538
rect 17502 29474 17554 29486
rect 18846 29538 18898 29550
rect 18846 29474 18898 29486
rect 20862 29538 20914 29550
rect 35646 29538 35698 29550
rect 27458 29486 27470 29538
rect 27522 29486 27534 29538
rect 20862 29474 20914 29486
rect 35646 29474 35698 29486
rect 38334 29538 38386 29550
rect 38334 29474 38386 29486
rect 41134 29538 41186 29550
rect 41134 29474 41186 29486
rect 42478 29538 42530 29550
rect 42478 29474 42530 29486
rect 10446 29426 10498 29438
rect 15262 29426 15314 29438
rect 2818 29374 2830 29426
rect 2882 29374 2894 29426
rect 10210 29374 10222 29426
rect 10274 29374 10286 29426
rect 11218 29374 11230 29426
rect 11282 29374 11294 29426
rect 10446 29362 10498 29374
rect 15262 29362 15314 29374
rect 15374 29426 15426 29438
rect 16494 29426 16546 29438
rect 15810 29374 15822 29426
rect 15874 29374 15886 29426
rect 15374 29362 15426 29374
rect 16494 29362 16546 29374
rect 18062 29426 18114 29438
rect 18062 29362 18114 29374
rect 18286 29426 18338 29438
rect 19518 29426 19570 29438
rect 18610 29374 18622 29426
rect 18674 29374 18686 29426
rect 18286 29362 18338 29374
rect 19518 29362 19570 29374
rect 19630 29426 19682 29438
rect 20302 29426 20354 29438
rect 19842 29374 19854 29426
rect 19906 29374 19918 29426
rect 19630 29362 19682 29374
rect 20302 29362 20354 29374
rect 20526 29426 20578 29438
rect 32286 29426 32338 29438
rect 38222 29426 38274 29438
rect 26786 29374 26798 29426
rect 26850 29374 26862 29426
rect 36082 29374 36094 29426
rect 36146 29374 36158 29426
rect 36754 29374 36766 29426
rect 36818 29374 36830 29426
rect 20526 29362 20578 29374
rect 32286 29362 32338 29374
rect 38222 29362 38274 29374
rect 38894 29426 38946 29438
rect 38894 29362 38946 29374
rect 41470 29426 41522 29438
rect 41470 29362 41522 29374
rect 42590 29426 42642 29438
rect 42590 29362 42642 29374
rect 42702 29426 42754 29438
rect 42702 29362 42754 29374
rect 43710 29426 43762 29438
rect 44606 29426 44658 29438
rect 44370 29374 44382 29426
rect 44434 29374 44446 29426
rect 45378 29374 45390 29426
rect 45442 29374 45454 29426
rect 43710 29362 43762 29374
rect 44606 29362 44658 29374
rect 2606 29314 2658 29326
rect 2606 29250 2658 29262
rect 3278 29314 3330 29326
rect 3278 29250 3330 29262
rect 10670 29314 10722 29326
rect 10670 29250 10722 29262
rect 11902 29314 11954 29326
rect 11902 29250 11954 29262
rect 13918 29314 13970 29326
rect 15486 29314 15538 29326
rect 19294 29314 19346 29326
rect 14354 29262 14366 29314
rect 14418 29262 14430 29314
rect 18834 29262 18846 29314
rect 18898 29262 18910 29314
rect 13918 29250 13970 29262
rect 15486 29250 15538 29262
rect 19294 29250 19346 29262
rect 21310 29314 21362 29326
rect 33182 29314 33234 29326
rect 40350 29314 40402 29326
rect 29586 29262 29598 29314
rect 29650 29262 29662 29314
rect 37090 29262 37102 29314
rect 37154 29262 37166 29314
rect 21310 29250 21362 29262
rect 33182 29250 33234 29262
rect 40350 29250 40402 29262
rect 43486 29314 43538 29326
rect 43486 29250 43538 29262
rect 44942 29314 44994 29326
rect 46050 29262 46062 29314
rect 46114 29262 46126 29314
rect 48178 29262 48190 29314
rect 48242 29262 48254 29314
rect 44942 29250 44994 29262
rect 2494 29202 2546 29214
rect 2494 29138 2546 29150
rect 5854 29202 5906 29214
rect 5854 29138 5906 29150
rect 5966 29202 6018 29214
rect 5966 29138 6018 29150
rect 6190 29202 6242 29214
rect 6190 29138 6242 29150
rect 6302 29202 6354 29214
rect 6302 29138 6354 29150
rect 17390 29202 17442 29214
rect 17390 29138 17442 29150
rect 32174 29202 32226 29214
rect 41246 29202 41298 29214
rect 36866 29150 36878 29202
rect 36930 29150 36942 29202
rect 32174 29138 32226 29150
rect 41246 29138 41298 29150
rect 41582 29202 41634 29214
rect 44830 29202 44882 29214
rect 42018 29150 42030 29202
rect 42082 29150 42094 29202
rect 41582 29138 41634 29150
rect 44830 29138 44882 29150
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 6638 28866 6690 28878
rect 13582 28866 13634 28878
rect 2482 28814 2494 28866
rect 2546 28814 2558 28866
rect 9874 28814 9886 28866
rect 9938 28814 9950 28866
rect 6638 28802 6690 28814
rect 13582 28802 13634 28814
rect 14926 28866 14978 28878
rect 43822 28866 43874 28878
rect 17826 28814 17838 28866
rect 17890 28814 17902 28866
rect 14926 28802 14978 28814
rect 43822 28802 43874 28814
rect 44158 28866 44210 28878
rect 44158 28802 44210 28814
rect 22094 28754 22146 28766
rect 45726 28754 45778 28766
rect 2930 28702 2942 28754
rect 2994 28702 3006 28754
rect 3714 28702 3726 28754
rect 3778 28702 3790 28754
rect 9762 28702 9774 28754
rect 9826 28702 9838 28754
rect 12562 28702 12574 28754
rect 12626 28702 12638 28754
rect 16370 28702 16382 28754
rect 16434 28702 16446 28754
rect 32050 28702 32062 28754
rect 32114 28702 32126 28754
rect 22094 28690 22146 28702
rect 45726 28690 45778 28702
rect 4174 28642 4226 28654
rect 3042 28590 3054 28642
rect 3106 28590 3118 28642
rect 4174 28578 4226 28590
rect 4398 28642 4450 28654
rect 4398 28578 4450 28590
rect 4622 28642 4674 28654
rect 4622 28578 4674 28590
rect 4846 28642 4898 28654
rect 4846 28578 4898 28590
rect 5070 28642 5122 28654
rect 5070 28578 5122 28590
rect 5630 28642 5682 28654
rect 5630 28578 5682 28590
rect 5966 28642 6018 28654
rect 5966 28578 6018 28590
rect 6414 28642 6466 28654
rect 6414 28578 6466 28590
rect 7198 28642 7250 28654
rect 8878 28642 8930 28654
rect 15038 28642 15090 28654
rect 18734 28642 18786 28654
rect 7634 28590 7646 28642
rect 7698 28590 7710 28642
rect 8642 28590 8654 28642
rect 8706 28590 8718 28642
rect 9650 28590 9662 28642
rect 9714 28590 9726 28642
rect 12338 28590 12350 28642
rect 12402 28590 12414 28642
rect 16818 28590 16830 28642
rect 16882 28590 16894 28642
rect 17378 28590 17390 28642
rect 17442 28590 17454 28642
rect 7198 28578 7250 28590
rect 8878 28578 8930 28590
rect 15038 28578 15090 28590
rect 18734 28578 18786 28590
rect 19070 28642 19122 28654
rect 24334 28642 24386 28654
rect 37102 28642 37154 28654
rect 37998 28642 38050 28654
rect 19394 28590 19406 28642
rect 19458 28590 19470 28642
rect 29138 28590 29150 28642
rect 29202 28590 29214 28642
rect 37426 28590 37438 28642
rect 37490 28590 37502 28642
rect 19070 28578 19122 28590
rect 24334 28578 24386 28590
rect 37102 28578 37154 28590
rect 37998 28578 38050 28590
rect 39566 28642 39618 28654
rect 44830 28642 44882 28654
rect 41682 28590 41694 28642
rect 41746 28590 41758 28642
rect 45266 28590 45278 28642
rect 45330 28590 45342 28642
rect 46162 28590 46174 28642
rect 46226 28590 46238 28642
rect 39566 28578 39618 28590
rect 44830 28578 44882 28590
rect 11678 28530 11730 28542
rect 5730 28478 5742 28530
rect 5794 28478 5806 28530
rect 11678 28466 11730 28478
rect 13694 28530 13746 28542
rect 13694 28466 13746 28478
rect 21422 28530 21474 28542
rect 21422 28466 21474 28478
rect 21534 28530 21586 28542
rect 21534 28466 21586 28478
rect 24222 28530 24274 28542
rect 44046 28530 44098 28542
rect 29922 28478 29934 28530
rect 29986 28478 29998 28530
rect 38658 28478 38670 28530
rect 38722 28478 38734 28530
rect 38994 28478 39006 28530
rect 39058 28478 39070 28530
rect 41458 28478 41470 28530
rect 41522 28478 41534 28530
rect 24222 28466 24274 28478
rect 44046 28466 44098 28478
rect 21758 28418 21810 28430
rect 21758 28354 21810 28366
rect 23998 28418 24050 28430
rect 39442 28366 39454 28418
rect 39506 28366 39518 28418
rect 23998 28354 24050 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 9998 28082 10050 28094
rect 16046 28082 16098 28094
rect 14018 28030 14030 28082
rect 14082 28030 14094 28082
rect 9998 28018 10050 28030
rect 16046 28018 16098 28030
rect 23774 28082 23826 28094
rect 23774 28018 23826 28030
rect 24110 28082 24162 28094
rect 24110 28018 24162 28030
rect 32398 28082 32450 28094
rect 32398 28018 32450 28030
rect 37550 28082 37602 28094
rect 37550 28018 37602 28030
rect 37998 28082 38050 28094
rect 37998 28018 38050 28030
rect 38222 28082 38274 28094
rect 38222 28018 38274 28030
rect 43486 28082 43538 28094
rect 43486 28018 43538 28030
rect 9774 27970 9826 27982
rect 2482 27918 2494 27970
rect 2546 27918 2558 27970
rect 6626 27918 6638 27970
rect 6690 27918 6702 27970
rect 9774 27906 9826 27918
rect 10222 27970 10274 27982
rect 10222 27906 10274 27918
rect 11790 27970 11842 27982
rect 11790 27906 11842 27918
rect 12014 27970 12066 27982
rect 12014 27906 12066 27918
rect 15822 27970 15874 27982
rect 18510 27970 18562 27982
rect 29934 27970 29986 27982
rect 37438 27970 37490 27982
rect 18274 27918 18286 27970
rect 18338 27918 18350 27970
rect 22194 27918 22206 27970
rect 22258 27918 22270 27970
rect 23426 27918 23438 27970
rect 23490 27918 23502 27970
rect 33842 27918 33854 27970
rect 33906 27918 33918 27970
rect 15822 27906 15874 27918
rect 18510 27906 18562 27918
rect 29934 27906 29986 27918
rect 37438 27906 37490 27918
rect 37886 27970 37938 27982
rect 37886 27906 37938 27918
rect 40014 27970 40066 27982
rect 40014 27906 40066 27918
rect 40126 27970 40178 27982
rect 40126 27906 40178 27918
rect 41358 27970 41410 27982
rect 41358 27906 41410 27918
rect 44830 27970 44882 27982
rect 44830 27906 44882 27918
rect 9886 27858 9938 27870
rect 1810 27806 1822 27858
rect 1874 27806 1886 27858
rect 5842 27806 5854 27858
rect 5906 27806 5918 27858
rect 9538 27806 9550 27858
rect 9602 27806 9614 27858
rect 9886 27794 9938 27806
rect 10446 27858 10498 27870
rect 10446 27794 10498 27806
rect 10782 27858 10834 27870
rect 10782 27794 10834 27806
rect 11006 27858 11058 27870
rect 11006 27794 11058 27806
rect 13694 27858 13746 27870
rect 13694 27794 13746 27806
rect 15374 27858 15426 27870
rect 15374 27794 15426 27806
rect 15598 27858 15650 27870
rect 15598 27794 15650 27806
rect 17950 27858 18002 27870
rect 17950 27794 18002 27806
rect 18734 27858 18786 27870
rect 18734 27794 18786 27806
rect 19070 27858 19122 27870
rect 41470 27858 41522 27870
rect 44270 27858 44322 27870
rect 19506 27806 19518 27858
rect 19570 27806 19582 27858
rect 22866 27806 22878 27858
rect 22930 27806 22942 27858
rect 25330 27806 25342 27858
rect 25394 27806 25406 27858
rect 28914 27806 28926 27858
rect 28978 27806 28990 27858
rect 32498 27806 32510 27858
rect 32562 27806 32574 27858
rect 33058 27806 33070 27858
rect 33122 27806 33134 27858
rect 39106 27806 39118 27858
rect 39170 27806 39182 27858
rect 39330 27806 39342 27858
rect 39394 27806 39406 27858
rect 43810 27806 43822 27858
rect 43874 27806 43886 27858
rect 45378 27806 45390 27858
rect 45442 27806 45454 27858
rect 19070 27794 19122 27806
rect 41470 27794 41522 27806
rect 44270 27794 44322 27806
rect 10670 27746 10722 27758
rect 4610 27694 4622 27746
rect 4674 27694 4686 27746
rect 8754 27694 8766 27746
rect 8818 27694 8830 27746
rect 10670 27682 10722 27694
rect 12462 27746 12514 27758
rect 12462 27682 12514 27694
rect 15934 27746 15986 27758
rect 30382 27746 30434 27758
rect 31390 27746 31442 27758
rect 44382 27746 44434 27758
rect 20066 27694 20078 27746
rect 20130 27694 20142 27746
rect 24546 27694 24558 27746
rect 24610 27694 24622 27746
rect 26002 27694 26014 27746
rect 26066 27694 26078 27746
rect 28130 27694 28142 27746
rect 28194 27694 28206 27746
rect 29138 27694 29150 27746
rect 29202 27694 29214 27746
rect 30818 27694 30830 27746
rect 30882 27694 30894 27746
rect 35970 27694 35982 27746
rect 36034 27694 36046 27746
rect 39554 27694 39566 27746
rect 39618 27694 39630 27746
rect 46050 27694 46062 27746
rect 46114 27694 46126 27746
rect 48178 27694 48190 27746
rect 48242 27694 48254 27746
rect 15934 27682 15986 27694
rect 30382 27682 30434 27694
rect 31390 27682 31442 27694
rect 44382 27682 44434 27694
rect 11678 27634 11730 27646
rect 11678 27570 11730 27582
rect 17726 27634 17778 27646
rect 30046 27634 30098 27646
rect 28578 27582 28590 27634
rect 28642 27582 28654 27634
rect 17726 27570 17778 27582
rect 30046 27570 30098 27582
rect 30270 27634 30322 27646
rect 30270 27570 30322 27582
rect 31166 27634 31218 27646
rect 31166 27570 31218 27582
rect 32062 27634 32114 27646
rect 32062 27570 32114 27582
rect 32286 27634 32338 27646
rect 40126 27634 40178 27646
rect 38658 27582 38670 27634
rect 38722 27582 38734 27634
rect 32286 27570 32338 27582
rect 40126 27570 40178 27582
rect 41358 27634 41410 27646
rect 41358 27570 41410 27582
rect 44046 27634 44098 27646
rect 44046 27570 44098 27582
rect 44718 27634 44770 27646
rect 44718 27570 44770 27582
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 9662 27298 9714 27310
rect 9662 27234 9714 27246
rect 26014 27298 26066 27310
rect 26014 27234 26066 27246
rect 30494 27298 30546 27310
rect 30494 27234 30546 27246
rect 32734 27298 32786 27310
rect 45166 27298 45218 27310
rect 43026 27246 43038 27298
rect 43090 27246 43102 27298
rect 32734 27234 32786 27246
rect 45166 27234 45218 27246
rect 7646 27186 7698 27198
rect 7646 27122 7698 27134
rect 9102 27186 9154 27198
rect 9102 27122 9154 27134
rect 9438 27186 9490 27198
rect 24894 27186 24946 27198
rect 10770 27134 10782 27186
rect 10834 27134 10846 27186
rect 12898 27134 12910 27186
rect 12962 27134 12974 27186
rect 9438 27122 9490 27134
rect 24894 27122 24946 27134
rect 25342 27186 25394 27198
rect 25342 27122 25394 27134
rect 25902 27186 25954 27198
rect 42590 27186 42642 27198
rect 30258 27134 30270 27186
rect 30322 27134 30334 27186
rect 25902 27122 25954 27134
rect 42590 27122 42642 27134
rect 43598 27186 43650 27198
rect 43598 27122 43650 27134
rect 44046 27186 44098 27198
rect 44818 27134 44830 27186
rect 44882 27134 44894 27186
rect 47842 27134 47854 27186
rect 47906 27134 47918 27186
rect 44046 27122 44098 27134
rect 15822 27074 15874 27086
rect 22542 27074 22594 27086
rect 10098 27022 10110 27074
rect 10162 27022 10174 27074
rect 13794 27022 13806 27074
rect 13858 27022 13870 27074
rect 14242 27022 14254 27074
rect 14306 27022 14318 27074
rect 14802 27022 14814 27074
rect 14866 27022 14878 27074
rect 16258 27022 16270 27074
rect 16322 27022 16334 27074
rect 17602 27022 17614 27074
rect 17666 27022 17678 27074
rect 18386 27022 18398 27074
rect 18450 27022 18462 27074
rect 21858 27022 21870 27074
rect 21922 27022 21934 27074
rect 15822 27010 15874 27022
rect 22542 27010 22594 27022
rect 23214 27074 23266 27086
rect 24110 27074 24162 27086
rect 23650 27022 23662 27074
rect 23714 27022 23726 27074
rect 23214 27010 23266 27022
rect 24110 27010 24162 27022
rect 29598 27074 29650 27086
rect 31614 27074 31666 27086
rect 30146 27022 30158 27074
rect 30210 27022 30222 27074
rect 29598 27010 29650 27022
rect 31614 27010 31666 27022
rect 35870 27074 35922 27086
rect 35870 27010 35922 27022
rect 36430 27074 36482 27086
rect 42254 27074 42306 27086
rect 38546 27022 38558 27074
rect 38610 27022 38622 27074
rect 39890 27022 39902 27074
rect 39954 27022 39966 27074
rect 40898 27022 40910 27074
rect 40962 27022 40974 27074
rect 36430 27010 36482 27022
rect 42254 27010 42306 27022
rect 42814 27074 42866 27086
rect 42814 27010 42866 27022
rect 43374 27074 43426 27086
rect 43374 27010 43426 27022
rect 43934 27074 43986 27086
rect 46050 27022 46062 27074
rect 46114 27022 46126 27074
rect 43934 27010 43986 27022
rect 8990 26962 9042 26974
rect 8990 26898 9042 26910
rect 9214 26962 9266 26974
rect 16494 26962 16546 26974
rect 25790 26962 25842 26974
rect 13458 26910 13470 26962
rect 13522 26910 13534 26962
rect 15362 26910 15374 26962
rect 15426 26910 15438 26962
rect 17266 26910 17278 26962
rect 17330 26910 17342 26962
rect 24434 26910 24446 26962
rect 24498 26910 24510 26962
rect 9214 26898 9266 26910
rect 16494 26898 16546 26910
rect 25790 26898 25842 26910
rect 32846 26962 32898 26974
rect 32846 26898 32898 26910
rect 33070 26962 33122 26974
rect 42366 26962 42418 26974
rect 41458 26910 41470 26962
rect 41522 26910 41534 26962
rect 33070 26898 33122 26910
rect 42366 26898 42418 26910
rect 44158 26962 44210 26974
rect 44158 26898 44210 26910
rect 44942 26962 44994 26974
rect 44942 26898 44994 26910
rect 18398 26850 18450 26862
rect 15138 26798 15150 26850
rect 15202 26798 15214 26850
rect 16594 26798 16606 26850
rect 16658 26798 16670 26850
rect 22082 26798 22094 26850
rect 22146 26798 22158 26850
rect 40562 26798 40574 26850
rect 40626 26798 40638 26850
rect 18398 26786 18450 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 7422 26514 7474 26526
rect 7422 26450 7474 26462
rect 17838 26514 17890 26526
rect 17838 26450 17890 26462
rect 22430 26514 22482 26526
rect 22430 26450 22482 26462
rect 22990 26514 23042 26526
rect 35422 26514 35474 26526
rect 33058 26462 33070 26514
rect 33122 26462 33134 26514
rect 22990 26450 23042 26462
rect 35422 26450 35474 26462
rect 39230 26514 39282 26526
rect 48066 26462 48078 26514
rect 48130 26462 48142 26514
rect 39230 26450 39282 26462
rect 8094 26402 8146 26414
rect 26462 26402 26514 26414
rect 7074 26350 7086 26402
rect 7138 26350 7150 26402
rect 15474 26350 15486 26402
rect 15538 26350 15550 26402
rect 8094 26338 8146 26350
rect 26462 26338 26514 26350
rect 33630 26402 33682 26414
rect 44270 26402 44322 26414
rect 35858 26350 35870 26402
rect 35922 26350 35934 26402
rect 33630 26338 33682 26350
rect 44270 26338 44322 26350
rect 4846 26290 4898 26302
rect 4846 26226 4898 26238
rect 5070 26290 5122 26302
rect 5966 26290 6018 26302
rect 5282 26238 5294 26290
rect 5346 26238 5358 26290
rect 5070 26226 5122 26238
rect 5966 26226 6018 26238
rect 15262 26290 15314 26302
rect 17614 26290 17666 26302
rect 15922 26238 15934 26290
rect 15986 26238 15998 26290
rect 16706 26238 16718 26290
rect 16770 26238 16782 26290
rect 17378 26238 17390 26290
rect 17442 26238 17454 26290
rect 15262 26226 15314 26238
rect 17614 26226 17666 26238
rect 17726 26290 17778 26302
rect 17726 26226 17778 26238
rect 17950 26290 18002 26302
rect 17950 26226 18002 26238
rect 18622 26290 18674 26302
rect 18622 26226 18674 26238
rect 18846 26290 18898 26302
rect 32174 26290 32226 26302
rect 33518 26290 33570 26302
rect 39342 26290 39394 26302
rect 19170 26238 19182 26290
rect 19234 26238 19246 26290
rect 19506 26238 19518 26290
rect 19570 26238 19582 26290
rect 26226 26238 26238 26290
rect 26290 26238 26302 26290
rect 32498 26238 32510 26290
rect 32562 26238 32574 26290
rect 33842 26238 33854 26290
rect 33906 26238 33918 26290
rect 36866 26238 36878 26290
rect 36930 26238 36942 26290
rect 38434 26238 38446 26290
rect 38498 26238 38510 26290
rect 38994 26238 39006 26290
rect 39058 26238 39070 26290
rect 18846 26226 18898 26238
rect 32174 26226 32226 26238
rect 33518 26226 33570 26238
rect 39342 26226 39394 26238
rect 39566 26290 39618 26302
rect 39566 26226 39618 26238
rect 39790 26290 39842 26302
rect 39790 26226 39842 26238
rect 39902 26290 39954 26302
rect 42590 26290 42642 26302
rect 41234 26238 41246 26290
rect 41298 26238 41310 26290
rect 41570 26238 41582 26290
rect 41634 26238 41646 26290
rect 42242 26238 42254 26290
rect 42306 26238 42318 26290
rect 39902 26226 39954 26238
rect 42590 26226 42642 26238
rect 42926 26290 42978 26302
rect 43138 26238 43150 26290
rect 43202 26238 43214 26290
rect 45154 26238 45166 26290
rect 45218 26238 45230 26290
rect 42926 26226 42978 26238
rect 6190 26178 6242 26190
rect 6190 26114 6242 26126
rect 8654 26178 8706 26190
rect 8654 26114 8706 26126
rect 20526 26178 20578 26190
rect 20526 26114 20578 26126
rect 21870 26178 21922 26190
rect 43922 26126 43934 26178
rect 43986 26126 43998 26178
rect 45826 26126 45838 26178
rect 45890 26126 45902 26178
rect 21870 26114 21922 26126
rect 4734 26066 4786 26078
rect 7870 26066 7922 26078
rect 5618 26014 5630 26066
rect 5682 26014 5694 26066
rect 4734 26002 4786 26014
rect 7870 26002 7922 26014
rect 8206 26066 8258 26078
rect 8206 26002 8258 26014
rect 15486 26066 15538 26078
rect 15486 26002 15538 26014
rect 19742 26066 19794 26078
rect 19742 26002 19794 26014
rect 19966 26066 20018 26078
rect 19966 26002 20018 26014
rect 20078 26066 20130 26078
rect 20078 26002 20130 26014
rect 32510 26066 32562 26078
rect 42130 26014 42142 26066
rect 42194 26014 42206 26066
rect 32510 26002 32562 26014
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 5630 25730 5682 25742
rect 5630 25666 5682 25678
rect 5966 25730 6018 25742
rect 5966 25666 6018 25678
rect 15262 25730 15314 25742
rect 15262 25666 15314 25678
rect 32622 25730 32674 25742
rect 32946 25678 32958 25730
rect 33010 25678 33022 25730
rect 32622 25666 32674 25678
rect 10558 25618 10610 25630
rect 2482 25566 2494 25618
rect 2546 25566 2558 25618
rect 4610 25566 4622 25618
rect 4674 25566 4686 25618
rect 8418 25566 8430 25618
rect 8482 25566 8494 25618
rect 10558 25554 10610 25566
rect 19182 25618 19234 25630
rect 19182 25554 19234 25566
rect 24670 25618 24722 25630
rect 32398 25618 32450 25630
rect 26450 25566 26462 25618
rect 26514 25566 26526 25618
rect 28578 25566 28590 25618
rect 28642 25566 28654 25618
rect 32050 25566 32062 25618
rect 32114 25566 32126 25618
rect 36418 25566 36430 25618
rect 36482 25566 36494 25618
rect 39106 25566 39118 25618
rect 39170 25566 39182 25618
rect 45602 25566 45614 25618
rect 45666 25566 45678 25618
rect 24670 25554 24722 25566
rect 32398 25554 32450 25566
rect 11342 25506 11394 25518
rect 1810 25454 1822 25506
rect 1874 25454 1886 25506
rect 7746 25454 7758 25506
rect 7810 25454 7822 25506
rect 11342 25442 11394 25454
rect 11566 25506 11618 25518
rect 15710 25506 15762 25518
rect 11778 25454 11790 25506
rect 11842 25454 11854 25506
rect 14914 25454 14926 25506
rect 14978 25454 14990 25506
rect 11566 25442 11618 25454
rect 15710 25442 15762 25454
rect 16494 25506 16546 25518
rect 25006 25506 25058 25518
rect 37326 25506 37378 25518
rect 38446 25506 38498 25518
rect 43598 25506 43650 25518
rect 16930 25454 16942 25506
rect 16994 25454 17006 25506
rect 17714 25454 17726 25506
rect 17778 25454 17790 25506
rect 25666 25454 25678 25506
rect 25730 25454 25742 25506
rect 29250 25454 29262 25506
rect 29314 25454 29326 25506
rect 33618 25454 33630 25506
rect 33682 25454 33694 25506
rect 38098 25454 38110 25506
rect 38162 25454 38174 25506
rect 39218 25454 39230 25506
rect 39282 25454 39294 25506
rect 41570 25454 41582 25506
rect 41634 25454 41646 25506
rect 41794 25454 41806 25506
rect 41858 25454 41870 25506
rect 43250 25454 43262 25506
rect 43314 25454 43326 25506
rect 44146 25454 44158 25506
rect 44210 25454 44222 25506
rect 45266 25454 45278 25506
rect 45330 25454 45342 25506
rect 45714 25454 45726 25506
rect 45778 25454 45790 25506
rect 16494 25442 16546 25454
rect 25006 25442 25058 25454
rect 37326 25442 37378 25454
rect 38446 25442 38498 25454
rect 43598 25442 43650 25454
rect 5742 25394 5794 25406
rect 22766 25394 22818 25406
rect 41918 25394 41970 25406
rect 46958 25394 47010 25406
rect 6626 25342 6638 25394
rect 6690 25342 6702 25394
rect 16034 25342 16046 25394
rect 16098 25342 16110 25394
rect 17938 25342 17950 25394
rect 18002 25342 18014 25394
rect 29922 25342 29934 25394
rect 29986 25342 29998 25394
rect 34290 25342 34302 25394
rect 34354 25342 34366 25394
rect 38770 25342 38782 25394
rect 38834 25342 38846 25394
rect 45826 25342 45838 25394
rect 45890 25342 45902 25394
rect 5742 25330 5794 25342
rect 22766 25330 22818 25342
rect 41918 25330 41970 25342
rect 46958 25330 47010 25342
rect 47518 25394 47570 25406
rect 47518 25330 47570 25342
rect 48190 25394 48242 25406
rect 48190 25330 48242 25342
rect 6302 25282 6354 25294
rect 6302 25218 6354 25230
rect 11230 25282 11282 25294
rect 11230 25218 11282 25230
rect 11454 25282 11506 25294
rect 11454 25218 11506 25230
rect 15150 25282 15202 25294
rect 23102 25282 23154 25294
rect 36990 25282 37042 25294
rect 16370 25230 16382 25282
rect 16434 25230 16446 25282
rect 25330 25230 25342 25282
rect 25394 25230 25406 25282
rect 15150 25218 15202 25230
rect 23102 25218 23154 25230
rect 36990 25218 37042 25230
rect 44158 25282 44210 25294
rect 44158 25218 44210 25230
rect 45054 25282 45106 25294
rect 45054 25218 45106 25230
rect 47182 25282 47234 25294
rect 47182 25218 47234 25230
rect 47854 25282 47906 25294
rect 47854 25218 47906 25230
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 22094 24946 22146 24958
rect 9538 24894 9550 24946
rect 9602 24894 9614 24946
rect 14690 24894 14702 24946
rect 14754 24894 14766 24946
rect 18610 24894 18622 24946
rect 18674 24894 18686 24946
rect 22094 24882 22146 24894
rect 38110 24946 38162 24958
rect 38110 24882 38162 24894
rect 38222 24946 38274 24958
rect 41134 24946 41186 24958
rect 38882 24894 38894 24946
rect 38946 24894 38958 24946
rect 38222 24882 38274 24894
rect 41134 24882 41186 24894
rect 41358 24946 41410 24958
rect 43710 24946 43762 24958
rect 42018 24894 42030 24946
rect 42082 24894 42094 24946
rect 42242 24894 42254 24946
rect 42306 24894 42318 24946
rect 41358 24882 41410 24894
rect 43710 24882 43762 24894
rect 46398 24946 46450 24958
rect 46398 24882 46450 24894
rect 47182 24946 47234 24958
rect 47182 24882 47234 24894
rect 30942 24834 30994 24846
rect 5954 24782 5966 24834
rect 6018 24782 6030 24834
rect 6738 24782 6750 24834
rect 6802 24782 6814 24834
rect 20850 24782 20862 24834
rect 20914 24782 20926 24834
rect 22642 24782 22654 24834
rect 22706 24782 22718 24834
rect 29810 24782 29822 24834
rect 29874 24782 29886 24834
rect 30942 24770 30994 24782
rect 33854 24834 33906 24846
rect 33854 24770 33906 24782
rect 37438 24834 37490 24846
rect 37438 24770 37490 24782
rect 37550 24834 37602 24846
rect 37550 24770 37602 24782
rect 37774 24834 37826 24846
rect 45614 24834 45666 24846
rect 39330 24782 39342 24834
rect 39394 24782 39406 24834
rect 42914 24782 42926 24834
rect 42978 24782 42990 24834
rect 37774 24770 37826 24782
rect 45614 24770 45666 24782
rect 47630 24834 47682 24846
rect 47630 24770 47682 24782
rect 9886 24722 9938 24734
rect 14366 24722 14418 24734
rect 4162 24670 4174 24722
rect 4226 24670 4238 24722
rect 6290 24670 6302 24722
rect 6354 24670 6366 24722
rect 6850 24670 6862 24722
rect 6914 24670 6926 24722
rect 11106 24670 11118 24722
rect 11170 24670 11182 24722
rect 9886 24658 9938 24670
rect 14366 24658 14418 24670
rect 15038 24722 15090 24734
rect 22318 24722 22370 24734
rect 15474 24670 15486 24722
rect 15538 24670 15550 24722
rect 16146 24670 16158 24722
rect 16210 24670 16222 24722
rect 21634 24670 21646 24722
rect 21698 24670 21710 24722
rect 15038 24658 15090 24670
rect 22318 24658 22370 24670
rect 22878 24722 22930 24734
rect 22878 24658 22930 24670
rect 24670 24722 24722 24734
rect 31054 24722 31106 24734
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 24670 24658 24722 24670
rect 31054 24658 31106 24670
rect 31390 24722 31442 24734
rect 33742 24722 33794 24734
rect 43822 24722 43874 24734
rect 31826 24670 31838 24722
rect 31890 24670 31902 24722
rect 33282 24670 33294 24722
rect 33346 24670 33358 24722
rect 38770 24670 38782 24722
rect 38834 24670 38846 24722
rect 39218 24670 39230 24722
rect 39282 24670 39294 24722
rect 40898 24670 40910 24722
rect 40962 24670 40974 24722
rect 41570 24670 41582 24722
rect 41634 24670 41646 24722
rect 42466 24670 42478 24722
rect 42530 24670 42542 24722
rect 43362 24670 43374 24722
rect 43426 24670 43438 24722
rect 31390 24658 31442 24670
rect 33742 24658 33794 24670
rect 43822 24658 43874 24670
rect 45838 24722 45890 24734
rect 45838 24658 45890 24670
rect 45950 24722 46002 24734
rect 45950 24658 46002 24670
rect 46174 24722 46226 24734
rect 46174 24658 46226 24670
rect 46510 24722 46562 24734
rect 46510 24658 46562 24670
rect 46846 24722 46898 24734
rect 46846 24658 46898 24670
rect 47294 24722 47346 24734
rect 47294 24658 47346 24670
rect 47406 24722 47458 24734
rect 47406 24658 47458 24670
rect 10334 24610 10386 24622
rect 23102 24610 23154 24622
rect 5618 24558 5630 24610
rect 5682 24558 5694 24610
rect 11890 24558 11902 24610
rect 11954 24558 11966 24610
rect 14018 24558 14030 24610
rect 14082 24558 14094 24610
rect 16370 24558 16382 24610
rect 16434 24558 16446 24610
rect 10334 24546 10386 24558
rect 23102 24546 23154 24558
rect 23550 24610 23602 24622
rect 48190 24610 48242 24622
rect 41010 24558 41022 24610
rect 41074 24558 41086 24610
rect 23550 24546 23602 24558
rect 48190 24546 48242 24558
rect 1934 24498 1986 24510
rect 31278 24498 31330 24510
rect 15474 24446 15486 24498
rect 15538 24446 15550 24498
rect 1934 24434 1986 24446
rect 31278 24434 31330 24446
rect 31838 24498 31890 24510
rect 31838 24434 31890 24446
rect 32174 24498 32226 24510
rect 32174 24434 32226 24446
rect 33518 24498 33570 24510
rect 33518 24434 33570 24446
rect 38334 24498 38386 24510
rect 38334 24434 38386 24446
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 11902 24162 11954 24174
rect 42926 24162 42978 24174
rect 26226 24110 26238 24162
rect 26290 24110 26302 24162
rect 11902 24098 11954 24110
rect 42926 24098 42978 24110
rect 7870 24050 7922 24062
rect 4610 23998 4622 24050
rect 4674 23998 4686 24050
rect 22866 23998 22878 24050
rect 22930 23998 22942 24050
rect 24994 23998 25006 24050
rect 25058 23998 25070 24050
rect 29922 23998 29934 24050
rect 29986 23998 29998 24050
rect 41122 23998 41134 24050
rect 41186 23998 41198 24050
rect 42018 23998 42030 24050
rect 42082 23998 42094 24050
rect 7870 23986 7922 23998
rect 5070 23938 5122 23950
rect 1810 23886 1822 23938
rect 1874 23886 1886 23938
rect 5070 23874 5122 23886
rect 5854 23938 5906 23950
rect 5854 23874 5906 23886
rect 6974 23938 7026 23950
rect 15934 23938 15986 23950
rect 20414 23938 20466 23950
rect 25678 23938 25730 23950
rect 7186 23886 7198 23938
rect 7250 23886 7262 23938
rect 12562 23886 12574 23938
rect 12626 23886 12638 23938
rect 19842 23886 19854 23938
rect 19906 23886 19918 23938
rect 22082 23886 22094 23938
rect 22146 23886 22158 23938
rect 25442 23886 25454 23938
rect 25506 23886 25518 23938
rect 6974 23874 7026 23886
rect 15934 23874 15986 23886
rect 20414 23874 20466 23886
rect 25678 23874 25730 23886
rect 26686 23938 26738 23950
rect 33518 23938 33570 23950
rect 28354 23886 28366 23938
rect 28418 23886 28430 23938
rect 29698 23886 29710 23938
rect 29762 23886 29774 23938
rect 26686 23874 26738 23886
rect 33518 23874 33570 23886
rect 33742 23938 33794 23950
rect 33742 23874 33794 23886
rect 41582 23938 41634 23950
rect 41582 23874 41634 23886
rect 42478 23938 42530 23950
rect 42478 23874 42530 23886
rect 45278 23938 45330 23950
rect 45278 23874 45330 23886
rect 46510 23938 46562 23950
rect 46510 23874 46562 23886
rect 46734 23938 46786 23950
rect 46734 23874 46786 23886
rect 47182 23938 47234 23950
rect 47182 23874 47234 23886
rect 47742 23938 47794 23950
rect 47742 23874 47794 23886
rect 48078 23938 48130 23950
rect 48078 23874 48130 23886
rect 5742 23826 5794 23838
rect 2482 23774 2494 23826
rect 2546 23774 2558 23826
rect 5742 23762 5794 23774
rect 8318 23826 8370 23838
rect 8318 23762 8370 23774
rect 12014 23826 12066 23838
rect 12014 23762 12066 23774
rect 25790 23826 25842 23838
rect 29150 23826 29202 23838
rect 28578 23774 28590 23826
rect 28642 23774 28654 23826
rect 25790 23762 25842 23774
rect 29150 23762 29202 23774
rect 33294 23826 33346 23838
rect 33294 23762 33346 23774
rect 43038 23826 43090 23838
rect 43038 23762 43090 23774
rect 46174 23826 46226 23838
rect 46174 23762 46226 23774
rect 5518 23714 5570 23726
rect 5518 23650 5570 23662
rect 8206 23714 8258 23726
rect 18398 23714 18450 23726
rect 33518 23714 33570 23726
rect 12338 23662 12350 23714
rect 12402 23662 12414 23714
rect 15586 23662 15598 23714
rect 15650 23662 15662 23714
rect 19618 23662 19630 23714
rect 19682 23662 19694 23714
rect 8206 23650 8258 23662
rect 18398 23650 18450 23662
rect 33518 23650 33570 23662
rect 38110 23714 38162 23726
rect 38110 23650 38162 23662
rect 45838 23714 45890 23726
rect 45838 23650 45890 23662
rect 46286 23714 46338 23726
rect 46286 23650 46338 23662
rect 47070 23714 47122 23726
rect 47070 23650 47122 23662
rect 47294 23714 47346 23726
rect 47294 23650 47346 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 3614 23378 3666 23390
rect 3614 23314 3666 23326
rect 18062 23378 18114 23390
rect 18062 23314 18114 23326
rect 18846 23378 18898 23390
rect 18846 23314 18898 23326
rect 19294 23378 19346 23390
rect 30718 23378 30770 23390
rect 29922 23326 29934 23378
rect 29986 23326 29998 23378
rect 19294 23314 19346 23326
rect 30718 23314 30770 23326
rect 38334 23378 38386 23390
rect 38334 23314 38386 23326
rect 39342 23378 39394 23390
rect 39342 23314 39394 23326
rect 44942 23378 44994 23390
rect 44942 23314 44994 23326
rect 2046 23266 2098 23278
rect 2046 23202 2098 23214
rect 2942 23266 2994 23278
rect 2942 23202 2994 23214
rect 6414 23266 6466 23278
rect 6414 23202 6466 23214
rect 17838 23266 17890 23278
rect 33518 23266 33570 23278
rect 18498 23214 18510 23266
rect 18562 23214 18574 23266
rect 31602 23214 31614 23266
rect 31666 23214 31678 23266
rect 17838 23202 17890 23214
rect 33518 23202 33570 23214
rect 39230 23266 39282 23278
rect 39230 23202 39282 23214
rect 43710 23266 43762 23278
rect 43710 23202 43762 23214
rect 44830 23266 44882 23278
rect 46050 23214 46062 23266
rect 46114 23214 46126 23266
rect 44830 23202 44882 23214
rect 1710 23154 1762 23166
rect 5518 23154 5570 23166
rect 31390 23154 31442 23166
rect 5282 23102 5294 23154
rect 5346 23102 5358 23154
rect 8866 23102 8878 23154
rect 8930 23102 8942 23154
rect 11330 23102 11342 23154
rect 11394 23102 11406 23154
rect 13906 23102 13918 23154
rect 13970 23102 13982 23154
rect 20514 23102 20526 23154
rect 20578 23102 20590 23154
rect 25330 23102 25342 23154
rect 25394 23102 25406 23154
rect 31154 23102 31166 23154
rect 31218 23102 31230 23154
rect 1710 23090 1762 23102
rect 5518 23090 5570 23102
rect 31390 23090 31442 23102
rect 33630 23154 33682 23166
rect 38222 23154 38274 23166
rect 33842 23102 33854 23154
rect 33906 23102 33918 23154
rect 34962 23102 34974 23154
rect 35026 23102 35038 23154
rect 33630 23090 33682 23102
rect 38222 23090 38274 23102
rect 38446 23154 38498 23166
rect 38446 23090 38498 23102
rect 38670 23154 38722 23166
rect 43598 23154 43650 23166
rect 42466 23102 42478 23154
rect 42530 23102 42542 23154
rect 42914 23102 42926 23154
rect 42978 23102 42990 23154
rect 45266 23102 45278 23154
rect 45330 23102 45342 23154
rect 38670 23090 38722 23102
rect 43598 23090 43650 23102
rect 2494 23042 2546 23054
rect 3166 23042 3218 23054
rect 2818 22990 2830 23042
rect 2882 22990 2894 23042
rect 2494 22978 2546 22990
rect 3166 22978 3218 22990
rect 4622 23042 4674 23054
rect 10558 23042 10610 23054
rect 8754 22990 8766 23042
rect 8818 22990 8830 23042
rect 4622 22978 4674 22990
rect 10558 22978 10610 22990
rect 10894 23042 10946 23054
rect 10894 22978 10946 22990
rect 11902 23042 11954 23054
rect 11902 22978 11954 22990
rect 12350 23042 12402 23054
rect 12350 22978 12402 22990
rect 12798 23042 12850 23054
rect 12798 22978 12850 22990
rect 13582 23042 13634 23054
rect 30494 23042 30546 23054
rect 14690 22990 14702 23042
rect 14754 22990 14766 23042
rect 16818 22990 16830 23042
rect 16882 22990 16894 23042
rect 21186 22990 21198 23042
rect 21250 22990 21262 23042
rect 23314 22990 23326 23042
rect 23378 22990 23390 23042
rect 26002 22990 26014 23042
rect 26066 22990 26078 23042
rect 28130 22990 28142 23042
rect 28194 22990 28206 23042
rect 13582 22978 13634 22990
rect 30494 22978 30546 22990
rect 31726 23042 31778 23054
rect 42254 23042 42306 23054
rect 35634 22990 35646 23042
rect 35698 22990 35710 23042
rect 37762 22990 37774 23042
rect 37826 22990 37838 23042
rect 31726 22978 31778 22990
rect 42254 22978 42306 22990
rect 44494 23042 44546 23054
rect 48178 22990 48190 23042
rect 48242 22990 48254 23042
rect 44494 22978 44546 22990
rect 6526 22930 6578 22942
rect 6526 22866 6578 22878
rect 8542 22930 8594 22942
rect 8542 22866 8594 22878
rect 11790 22930 11842 22942
rect 11790 22866 11842 22878
rect 18174 22930 18226 22942
rect 18174 22866 18226 22878
rect 30270 22930 30322 22942
rect 38894 22930 38946 22942
rect 33058 22878 33070 22930
rect 33122 22878 33134 22930
rect 30270 22866 30322 22878
rect 38894 22866 38946 22878
rect 39342 22930 39394 22942
rect 39342 22866 39394 22878
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 31614 22594 31666 22606
rect 34302 22594 34354 22606
rect 31938 22542 31950 22594
rect 32002 22542 32014 22594
rect 31614 22530 31666 22542
rect 34302 22530 34354 22542
rect 34638 22594 34690 22606
rect 34638 22530 34690 22542
rect 47966 22594 48018 22606
rect 47966 22530 48018 22542
rect 12462 22482 12514 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 11106 22430 11118 22482
rect 11170 22430 11182 22482
rect 12462 22418 12514 22430
rect 14478 22482 14530 22494
rect 22654 22482 22706 22494
rect 18274 22430 18286 22482
rect 18338 22430 18350 22482
rect 14478 22418 14530 22430
rect 22654 22418 22706 22430
rect 24446 22482 24498 22494
rect 24446 22418 24498 22430
rect 25678 22482 25730 22494
rect 31390 22482 31442 22494
rect 26898 22430 26910 22482
rect 26962 22430 26974 22482
rect 25678 22418 25730 22430
rect 31390 22418 31442 22430
rect 34414 22482 34466 22494
rect 34414 22418 34466 22430
rect 35086 22482 35138 22494
rect 42578 22430 42590 22482
rect 42642 22430 42654 22482
rect 44818 22430 44830 22482
rect 44882 22430 44894 22482
rect 35086 22418 35138 22430
rect 12126 22370 12178 22382
rect 1810 22318 1822 22370
rect 1874 22318 1886 22370
rect 8194 22318 8206 22370
rect 8258 22318 8270 22370
rect 12126 22306 12178 22318
rect 14030 22370 14082 22382
rect 22318 22370 22370 22382
rect 17602 22318 17614 22370
rect 17666 22318 17678 22370
rect 14030 22306 14082 22318
rect 22318 22306 22370 22318
rect 22542 22370 22594 22382
rect 22542 22306 22594 22318
rect 22878 22370 22930 22382
rect 22878 22306 22930 22318
rect 22990 22370 23042 22382
rect 24782 22370 24834 22382
rect 30158 22370 30210 22382
rect 23090 22318 23102 22370
rect 23154 22318 23166 22370
rect 25442 22318 25454 22370
rect 25506 22318 25518 22370
rect 27234 22318 27246 22370
rect 27298 22318 27310 22370
rect 28018 22318 28030 22370
rect 28082 22318 28094 22370
rect 22990 22306 23042 22318
rect 24782 22306 24834 22318
rect 30158 22306 30210 22318
rect 33406 22370 33458 22382
rect 34750 22370 34802 22382
rect 38782 22370 38834 22382
rect 43150 22370 43202 22382
rect 33842 22318 33854 22370
rect 33906 22318 33918 22370
rect 37986 22318 37998 22370
rect 38050 22318 38062 22370
rect 39666 22318 39678 22370
rect 39730 22318 39742 22370
rect 45826 22318 45838 22370
rect 45890 22318 45902 22370
rect 33406 22306 33458 22318
rect 34750 22306 34802 22318
rect 38782 22306 38834 22318
rect 43150 22306 43202 22318
rect 6190 22258 6242 22270
rect 12350 22258 12402 22270
rect 2482 22206 2494 22258
rect 2546 22206 2558 22258
rect 8978 22206 8990 22258
rect 9042 22206 9054 22258
rect 6190 22194 6242 22206
rect 12350 22194 12402 22206
rect 12686 22258 12738 22270
rect 12686 22194 12738 22206
rect 12910 22258 12962 22270
rect 12910 22194 12962 22206
rect 13582 22258 13634 22270
rect 13582 22194 13634 22206
rect 13918 22258 13970 22270
rect 13918 22194 13970 22206
rect 21982 22258 22034 22270
rect 21982 22194 22034 22206
rect 23774 22258 23826 22270
rect 23774 22194 23826 22206
rect 25790 22258 25842 22270
rect 25790 22194 25842 22206
rect 26574 22258 26626 22270
rect 26574 22194 26626 22206
rect 30494 22258 30546 22270
rect 30494 22194 30546 22206
rect 33182 22258 33234 22270
rect 33182 22194 33234 22206
rect 33294 22258 33346 22270
rect 33294 22194 33346 22206
rect 35310 22258 35362 22270
rect 35310 22194 35362 22206
rect 37774 22258 37826 22270
rect 37774 22194 37826 22206
rect 38446 22258 38498 22270
rect 43038 22258 43090 22270
rect 40450 22206 40462 22258
rect 40514 22206 40526 22258
rect 38446 22194 38498 22206
rect 43038 22194 43090 22206
rect 45166 22258 45218 22270
rect 45166 22194 45218 22206
rect 5070 22146 5122 22158
rect 5070 22082 5122 22094
rect 6302 22146 6354 22158
rect 6302 22082 6354 22094
rect 11454 22146 11506 22158
rect 11454 22082 11506 22094
rect 11566 22146 11618 22158
rect 11566 22082 11618 22094
rect 11678 22146 11730 22158
rect 11678 22082 11730 22094
rect 13806 22146 13858 22158
rect 22094 22146 22146 22158
rect 20514 22094 20526 22146
rect 20578 22094 20590 22146
rect 13806 22082 13858 22094
rect 22094 22082 22146 22094
rect 23662 22146 23714 22158
rect 35198 22146 35250 22158
rect 25106 22094 25118 22146
rect 25170 22094 25182 22146
rect 28242 22094 28254 22146
rect 28306 22094 28318 22146
rect 23662 22082 23714 22094
rect 35198 22082 35250 22094
rect 38558 22146 38610 22158
rect 38558 22082 38610 22094
rect 42814 22146 42866 22158
rect 42814 22082 42866 22094
rect 43598 22146 43650 22158
rect 43598 22082 43650 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 8318 21810 8370 21822
rect 8318 21746 8370 21758
rect 8654 21810 8706 21822
rect 8654 21746 8706 21758
rect 10334 21810 10386 21822
rect 12462 21810 12514 21822
rect 10994 21758 11006 21810
rect 11058 21758 11070 21810
rect 10334 21746 10386 21758
rect 12462 21746 12514 21758
rect 24558 21810 24610 21822
rect 24558 21746 24610 21758
rect 27806 21810 27858 21822
rect 27806 21746 27858 21758
rect 38894 21810 38946 21822
rect 38894 21746 38946 21758
rect 41022 21810 41074 21822
rect 41022 21746 41074 21758
rect 42030 21810 42082 21822
rect 42030 21746 42082 21758
rect 6862 21698 6914 21710
rect 6862 21634 6914 21646
rect 7198 21698 7250 21710
rect 7198 21634 7250 21646
rect 7534 21698 7586 21710
rect 7534 21634 7586 21646
rect 12014 21698 12066 21710
rect 12014 21634 12066 21646
rect 12574 21698 12626 21710
rect 12574 21634 12626 21646
rect 17390 21698 17442 21710
rect 17390 21634 17442 21646
rect 27918 21698 27970 21710
rect 27918 21634 27970 21646
rect 41246 21698 41298 21710
rect 41246 21634 41298 21646
rect 5742 21586 5794 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 5742 21522 5794 21534
rect 8430 21586 8482 21598
rect 10670 21586 10722 21598
rect 8866 21534 8878 21586
rect 8930 21534 8942 21586
rect 8430 21522 8482 21534
rect 10670 21522 10722 21534
rect 11566 21586 11618 21598
rect 11566 21522 11618 21534
rect 11678 21586 11730 21598
rect 11678 21522 11730 21534
rect 11902 21586 11954 21598
rect 34190 21586 34242 21598
rect 15138 21534 15150 21586
rect 15202 21534 15214 21586
rect 17826 21534 17838 21586
rect 17890 21534 17902 21586
rect 19282 21534 19294 21586
rect 19346 21534 19358 21586
rect 31378 21534 31390 21586
rect 31442 21534 31454 21586
rect 32050 21534 32062 21586
rect 32114 21534 32126 21586
rect 33954 21534 33966 21586
rect 34018 21534 34030 21586
rect 11902 21522 11954 21534
rect 34190 21522 34242 21534
rect 34414 21586 34466 21598
rect 34414 21522 34466 21534
rect 38782 21586 38834 21598
rect 38782 21522 38834 21534
rect 39006 21586 39058 21598
rect 39006 21522 39058 21534
rect 39454 21586 39506 21598
rect 39454 21522 39506 21534
rect 41806 21586 41858 21598
rect 42354 21534 42366 21586
rect 42418 21534 42430 21586
rect 43810 21534 43822 21586
rect 43874 21534 43886 21586
rect 45042 21534 45054 21586
rect 45106 21534 45118 21586
rect 46050 21534 46062 21586
rect 46114 21534 46126 21586
rect 41806 21522 41858 21534
rect 1934 21474 1986 21486
rect 1934 21410 1986 21422
rect 5966 21474 6018 21486
rect 5966 21410 6018 21422
rect 8542 21474 8594 21486
rect 8542 21410 8594 21422
rect 13134 21474 13186 21486
rect 13134 21410 13186 21422
rect 14926 21474 14978 21486
rect 23662 21474 23714 21486
rect 18274 21422 18286 21474
rect 18338 21422 18350 21474
rect 14926 21410 14978 21422
rect 23662 21410 23714 21422
rect 31166 21474 31218 21486
rect 31166 21410 31218 21422
rect 31838 21474 31890 21486
rect 31838 21410 31890 21422
rect 39230 21474 39282 21486
rect 39230 21410 39282 21422
rect 40350 21474 40402 21486
rect 41918 21474 41970 21486
rect 40898 21422 40910 21474
rect 40962 21422 40974 21474
rect 44034 21422 44046 21474
rect 44098 21422 44110 21474
rect 45154 21422 45166 21474
rect 45218 21422 45230 21474
rect 40350 21410 40402 21422
rect 41918 21410 41970 21422
rect 6414 21362 6466 21374
rect 5394 21310 5406 21362
rect 5458 21310 5470 21362
rect 6414 21298 6466 21310
rect 6526 21362 6578 21374
rect 6526 21298 6578 21310
rect 6750 21362 6802 21374
rect 6750 21298 6802 21310
rect 14814 21362 14866 21374
rect 14814 21298 14866 21310
rect 18734 21362 18786 21374
rect 18734 21298 18786 21310
rect 18846 21362 18898 21374
rect 18846 21298 18898 21310
rect 19070 21362 19122 21374
rect 19070 21298 19122 21310
rect 30830 21362 30882 21374
rect 30830 21298 30882 21310
rect 30942 21362 30994 21374
rect 30942 21298 30994 21310
rect 31726 21362 31778 21374
rect 31726 21298 31778 21310
rect 34526 21362 34578 21374
rect 47966 21362 48018 21374
rect 43922 21310 43934 21362
rect 43986 21310 43998 21362
rect 34526 21298 34578 21310
rect 47966 21298 48018 21310
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 4622 21026 4674 21038
rect 4622 20962 4674 20974
rect 4958 21026 5010 21038
rect 4958 20962 5010 20974
rect 14366 21026 14418 21038
rect 14366 20962 14418 20974
rect 14590 21026 14642 21038
rect 14590 20962 14642 20974
rect 21310 21026 21362 21038
rect 21310 20962 21362 20974
rect 22206 21026 22258 21038
rect 22206 20962 22258 20974
rect 2494 20914 2546 20926
rect 2494 20850 2546 20862
rect 10222 20914 10274 20926
rect 10222 20850 10274 20862
rect 14702 20914 14754 20926
rect 37662 20914 37714 20926
rect 15698 20862 15710 20914
rect 15762 20862 15774 20914
rect 14702 20850 14754 20862
rect 37662 20850 37714 20862
rect 37774 20914 37826 20926
rect 43598 20914 43650 20926
rect 38770 20862 38782 20914
rect 38834 20862 38846 20914
rect 41794 20862 41806 20914
rect 41858 20862 41870 20914
rect 48178 20862 48190 20914
rect 48242 20862 48254 20914
rect 37774 20850 37826 20862
rect 43598 20850 43650 20862
rect 1710 20802 1762 20814
rect 3726 20802 3778 20814
rect 3266 20750 3278 20802
rect 3330 20750 3342 20802
rect 1710 20738 1762 20750
rect 3726 20738 3778 20750
rect 4846 20802 4898 20814
rect 15150 20802 15202 20814
rect 5954 20750 5966 20802
rect 6018 20750 6030 20802
rect 7970 20750 7982 20802
rect 8034 20750 8046 20802
rect 4846 20738 4898 20750
rect 15150 20738 15202 20750
rect 15374 20802 15426 20814
rect 19630 20802 19682 20814
rect 16146 20750 16158 20802
rect 16210 20750 16222 20802
rect 17826 20750 17838 20802
rect 17890 20750 17902 20802
rect 15374 20738 15426 20750
rect 19630 20738 19682 20750
rect 19854 20802 19906 20814
rect 19854 20738 19906 20750
rect 19966 20802 20018 20814
rect 19966 20738 20018 20750
rect 20190 20802 20242 20814
rect 20190 20738 20242 20750
rect 22990 20802 23042 20814
rect 22990 20738 23042 20750
rect 23438 20802 23490 20814
rect 23438 20738 23490 20750
rect 23662 20802 23714 20814
rect 23662 20738 23714 20750
rect 24558 20802 24610 20814
rect 24558 20738 24610 20750
rect 24894 20802 24946 20814
rect 30382 20802 30434 20814
rect 29922 20750 29934 20802
rect 29986 20750 29998 20802
rect 24894 20738 24946 20750
rect 30382 20738 30434 20750
rect 30494 20802 30546 20814
rect 30494 20738 30546 20750
rect 30718 20802 30770 20814
rect 30718 20738 30770 20750
rect 31166 20802 31218 20814
rect 31166 20738 31218 20750
rect 37102 20802 37154 20814
rect 37102 20738 37154 20750
rect 38446 20802 38498 20814
rect 39118 20802 39170 20814
rect 38658 20750 38670 20802
rect 38722 20750 38734 20802
rect 38446 20738 38498 20750
rect 39118 20738 39170 20750
rect 39566 20802 39618 20814
rect 39566 20738 39618 20750
rect 40014 20802 40066 20814
rect 40014 20738 40066 20750
rect 40126 20802 40178 20814
rect 40126 20738 40178 20750
rect 40798 20802 40850 20814
rect 42814 20802 42866 20814
rect 41682 20750 41694 20802
rect 41746 20750 41758 20802
rect 42354 20750 42366 20802
rect 42418 20750 42430 20802
rect 40798 20738 40850 20750
rect 42814 20738 42866 20750
rect 43710 20802 43762 20814
rect 43710 20738 43762 20750
rect 43934 20802 43986 20814
rect 45266 20750 45278 20802
rect 45330 20750 45342 20802
rect 43934 20738 43986 20750
rect 2046 20690 2098 20702
rect 2046 20626 2098 20638
rect 2830 20690 2882 20702
rect 2830 20626 2882 20638
rect 4510 20690 4562 20702
rect 8542 20690 8594 20702
rect 6066 20638 6078 20690
rect 6130 20638 6142 20690
rect 4510 20626 4562 20638
rect 8542 20626 8594 20638
rect 14254 20690 14306 20702
rect 19518 20690 19570 20702
rect 16706 20638 16718 20690
rect 16770 20638 16782 20690
rect 17714 20638 17726 20690
rect 17778 20638 17790 20690
rect 14254 20626 14306 20638
rect 19518 20626 19570 20638
rect 21422 20690 21474 20702
rect 21422 20626 21474 20638
rect 22094 20690 22146 20702
rect 22094 20626 22146 20638
rect 23998 20690 24050 20702
rect 23998 20626 24050 20638
rect 25230 20690 25282 20702
rect 25230 20626 25282 20638
rect 29262 20690 29314 20702
rect 29262 20626 29314 20638
rect 29374 20690 29426 20702
rect 29374 20626 29426 20638
rect 29486 20690 29538 20702
rect 29486 20626 29538 20638
rect 30830 20690 30882 20702
rect 30830 20626 30882 20638
rect 36990 20690 37042 20702
rect 36990 20626 37042 20638
rect 38110 20690 38162 20702
rect 38110 20626 38162 20638
rect 38222 20690 38274 20702
rect 38222 20626 38274 20638
rect 39342 20690 39394 20702
rect 39342 20626 39394 20638
rect 39790 20690 39842 20702
rect 39790 20626 39842 20638
rect 40686 20690 40738 20702
rect 43486 20690 43538 20702
rect 41794 20638 41806 20690
rect 41858 20638 41870 20690
rect 40686 20626 40738 20638
rect 43486 20626 43538 20638
rect 44830 20690 44882 20702
rect 46050 20638 46062 20690
rect 46114 20638 46126 20690
rect 44830 20626 44882 20638
rect 10110 20578 10162 20590
rect 6962 20526 6974 20578
rect 7026 20526 7038 20578
rect 10110 20514 10162 20526
rect 11118 20578 11170 20590
rect 11118 20514 11170 20526
rect 22206 20578 22258 20590
rect 22206 20514 22258 20526
rect 23326 20578 23378 20590
rect 23326 20514 23378 20526
rect 23886 20578 23938 20590
rect 23886 20514 23938 20526
rect 24894 20578 24946 20590
rect 24894 20514 24946 20526
rect 31278 20578 31330 20590
rect 31278 20514 31330 20526
rect 31390 20578 31442 20590
rect 31390 20514 31442 20526
rect 38894 20578 38946 20590
rect 38894 20514 38946 20526
rect 40462 20578 40514 20590
rect 40462 20514 40514 20526
rect 44942 20578 44994 20590
rect 44942 20514 44994 20526
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 6414 20242 6466 20254
rect 6414 20178 6466 20190
rect 16830 20242 16882 20254
rect 16830 20178 16882 20190
rect 30382 20242 30434 20254
rect 30382 20178 30434 20190
rect 39118 20242 39170 20254
rect 39118 20178 39170 20190
rect 39230 20242 39282 20254
rect 39230 20178 39282 20190
rect 46846 20242 46898 20254
rect 46846 20178 46898 20190
rect 5630 20130 5682 20142
rect 5630 20066 5682 20078
rect 5742 20130 5794 20142
rect 5742 20066 5794 20078
rect 5854 20130 5906 20142
rect 5854 20066 5906 20078
rect 6190 20130 6242 20142
rect 6190 20066 6242 20078
rect 6750 20130 6802 20142
rect 6750 20066 6802 20078
rect 8654 20130 8706 20142
rect 8654 20066 8706 20078
rect 9886 20130 9938 20142
rect 9886 20066 9938 20078
rect 10782 20130 10834 20142
rect 37662 20130 37714 20142
rect 44270 20130 44322 20142
rect 12898 20078 12910 20130
rect 12962 20078 12974 20130
rect 18834 20078 18846 20130
rect 18898 20078 18910 20130
rect 23090 20078 23102 20130
rect 23154 20078 23166 20130
rect 24658 20078 24670 20130
rect 24722 20078 24734 20130
rect 34738 20078 34750 20130
rect 34802 20078 34814 20130
rect 41794 20078 41806 20130
rect 41858 20078 41870 20130
rect 10782 20066 10834 20078
rect 37662 20066 37714 20078
rect 44270 20066 44322 20078
rect 47854 20130 47906 20142
rect 47854 20066 47906 20078
rect 6526 20018 6578 20030
rect 1810 19966 1822 20018
rect 1874 19966 1886 20018
rect 6526 19954 6578 19966
rect 8542 20018 8594 20030
rect 8542 19954 8594 19966
rect 8878 20018 8930 20030
rect 8878 19954 8930 19966
rect 9102 20018 9154 20030
rect 9102 19954 9154 19966
rect 10334 20018 10386 20030
rect 10334 19954 10386 19966
rect 10558 20018 10610 20030
rect 10558 19954 10610 19966
rect 11006 20018 11058 20030
rect 15486 20018 15538 20030
rect 22542 20018 22594 20030
rect 24110 20018 24162 20030
rect 29038 20018 29090 20030
rect 12114 19966 12126 20018
rect 12178 19966 12190 20018
rect 18050 19966 18062 20018
rect 18114 19966 18126 20018
rect 22306 19966 22318 20018
rect 22370 19966 22382 20018
rect 22978 19966 22990 20018
rect 23042 19966 23054 20018
rect 25218 19966 25230 20018
rect 25282 19966 25294 20018
rect 11006 19954 11058 19966
rect 15486 19954 15538 19966
rect 22542 19954 22594 19966
rect 24110 19954 24162 19966
rect 29038 19954 29090 19966
rect 29486 20018 29538 20030
rect 29486 19954 29538 19966
rect 29598 20018 29650 20030
rect 29598 19954 29650 19966
rect 29710 20018 29762 20030
rect 29710 19954 29762 19966
rect 30046 20018 30098 20030
rect 30046 19954 30098 19966
rect 30382 20018 30434 20030
rect 30382 19954 30434 19966
rect 30718 20018 30770 20030
rect 30718 19954 30770 19966
rect 31166 20018 31218 20030
rect 31166 19954 31218 19966
rect 31390 20018 31442 20030
rect 37102 20018 37154 20030
rect 39006 20018 39058 20030
rect 43822 20018 43874 20030
rect 46622 20018 46674 20030
rect 31602 19966 31614 20018
rect 31666 19966 31678 20018
rect 33954 19966 33966 20018
rect 34018 19966 34030 20018
rect 37426 19966 37438 20018
rect 37490 19966 37502 20018
rect 43250 19966 43262 20018
rect 43314 19966 43326 20018
rect 45938 19966 45950 20018
rect 46002 19966 46014 20018
rect 31390 19954 31442 19966
rect 37102 19954 37154 19966
rect 39006 19954 39058 19966
rect 43822 19954 43874 19966
rect 46622 19954 46674 19966
rect 46958 20018 47010 20030
rect 46958 19954 47010 19966
rect 47182 20018 47234 20030
rect 48066 19966 48078 20018
rect 48130 19966 48142 20018
rect 47182 19954 47234 19966
rect 5070 19906 5122 19918
rect 2482 19854 2494 19906
rect 2546 19854 2558 19906
rect 4610 19854 4622 19906
rect 4674 19854 4686 19906
rect 5070 19842 5122 19854
rect 11118 19906 11170 19918
rect 16718 19906 16770 19918
rect 21646 19906 21698 19918
rect 37326 19906 37378 19918
rect 46398 19906 46450 19918
rect 15026 19854 15038 19906
rect 15090 19854 15102 19906
rect 20962 19854 20974 19906
rect 21026 19854 21038 19906
rect 24322 19854 24334 19906
rect 24386 19854 24398 19906
rect 26002 19854 26014 19906
rect 26066 19854 26078 19906
rect 28130 19854 28142 19906
rect 28194 19854 28206 19906
rect 36866 19854 36878 19906
rect 36930 19854 36942 19906
rect 43586 19854 43598 19906
rect 43650 19854 43662 19906
rect 11118 19842 11170 19854
rect 16718 19842 16770 19854
rect 21646 19842 21698 19854
rect 37326 19842 37378 19854
rect 46398 19842 46450 19854
rect 9662 19794 9714 19806
rect 9662 19730 9714 19742
rect 9998 19794 10050 19806
rect 9998 19730 10050 19742
rect 28814 19794 28866 19806
rect 28814 19730 28866 19742
rect 31054 19794 31106 19806
rect 31054 19730 31106 19742
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 2718 19458 2770 19470
rect 2718 19394 2770 19406
rect 3054 19458 3106 19470
rect 3054 19394 3106 19406
rect 8990 19458 9042 19470
rect 8990 19394 9042 19406
rect 9214 19458 9266 19470
rect 9214 19394 9266 19406
rect 11006 19458 11058 19470
rect 11006 19394 11058 19406
rect 11230 19458 11282 19470
rect 11230 19394 11282 19406
rect 20302 19458 20354 19470
rect 20302 19394 20354 19406
rect 25454 19458 25506 19470
rect 25454 19394 25506 19406
rect 25678 19458 25730 19470
rect 25678 19394 25730 19406
rect 3502 19346 3554 19358
rect 3502 19282 3554 19294
rect 12126 19346 12178 19358
rect 12126 19282 12178 19294
rect 15150 19346 15202 19358
rect 15150 19282 15202 19294
rect 17166 19346 17218 19358
rect 17166 19282 17218 19294
rect 19630 19346 19682 19358
rect 43934 19346 43986 19358
rect 31938 19294 31950 19346
rect 32002 19294 32014 19346
rect 34066 19294 34078 19346
rect 34130 19294 34142 19346
rect 39890 19294 39902 19346
rect 39954 19294 39966 19346
rect 42914 19294 42926 19346
rect 42978 19294 42990 19346
rect 19630 19282 19682 19294
rect 43934 19282 43986 19294
rect 44270 19346 44322 19358
rect 46734 19346 46786 19358
rect 44930 19294 44942 19346
rect 44994 19294 45006 19346
rect 44270 19282 44322 19294
rect 46734 19282 46786 19294
rect 5630 19234 5682 19246
rect 9774 19234 9826 19246
rect 8642 19182 8654 19234
rect 8706 19182 8718 19234
rect 5630 19170 5682 19182
rect 9774 19170 9826 19182
rect 10558 19234 10610 19246
rect 10558 19170 10610 19182
rect 12238 19234 12290 19246
rect 12238 19170 12290 19182
rect 13806 19234 13858 19246
rect 13806 19170 13858 19182
rect 13918 19234 13970 19246
rect 30158 19234 30210 19246
rect 14690 19182 14702 19234
rect 14754 19182 14766 19234
rect 19954 19182 19966 19234
rect 20018 19182 20030 19234
rect 25890 19182 25902 19234
rect 25954 19182 25966 19234
rect 27122 19182 27134 19234
rect 27186 19182 27198 19234
rect 13918 19170 13970 19182
rect 30158 19170 30210 19182
rect 30382 19234 30434 19246
rect 47294 19234 47346 19246
rect 31154 19182 31166 19234
rect 31218 19182 31230 19234
rect 38770 19182 38782 19234
rect 38834 19182 38846 19234
rect 42018 19182 42030 19234
rect 42082 19182 42094 19234
rect 43026 19182 43038 19234
rect 43090 19182 43102 19234
rect 45042 19182 45054 19234
rect 45106 19182 45118 19234
rect 46162 19182 46174 19234
rect 46226 19182 46238 19234
rect 30382 19170 30434 19182
rect 47294 19170 47346 19182
rect 2830 19122 2882 19134
rect 2830 19058 2882 19070
rect 10446 19122 10498 19134
rect 10446 19058 10498 19070
rect 11678 19122 11730 19134
rect 11678 19058 11730 19070
rect 11902 19122 11954 19134
rect 29934 19122 29986 19134
rect 26898 19070 26910 19122
rect 26962 19070 26974 19122
rect 42690 19070 42702 19122
rect 42754 19070 42766 19122
rect 45154 19070 45166 19122
rect 45218 19070 45230 19122
rect 11902 19058 11954 19070
rect 29934 19058 29986 19070
rect 5742 19010 5794 19022
rect 5742 18946 5794 18958
rect 8318 19010 8370 19022
rect 8318 18946 8370 18958
rect 8430 19010 8482 19022
rect 8430 18946 8482 18958
rect 8542 19010 8594 19022
rect 8542 18946 8594 18958
rect 9886 19010 9938 19022
rect 9886 18946 9938 18958
rect 10110 19010 10162 19022
rect 10110 18946 10162 18958
rect 11342 19010 11394 19022
rect 11342 18946 11394 18958
rect 17054 19010 17106 19022
rect 17054 18946 17106 18958
rect 20190 19010 20242 19022
rect 20190 18946 20242 18958
rect 25790 19010 25842 19022
rect 25790 18946 25842 18958
rect 30158 19010 30210 19022
rect 30158 18946 30210 18958
rect 37102 19010 37154 19022
rect 37102 18946 37154 18958
rect 38446 19010 38498 19022
rect 38446 18946 38498 18958
rect 41918 19010 41970 19022
rect 41918 18946 41970 18958
rect 46062 19010 46114 19022
rect 46062 18946 46114 18958
rect 46622 19010 46674 19022
rect 46622 18946 46674 18958
rect 46846 19010 46898 19022
rect 46846 18946 46898 18958
rect 47518 19010 47570 19022
rect 47842 18958 47854 19010
rect 47906 18958 47918 19010
rect 47518 18946 47570 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 6974 18674 7026 18686
rect 6974 18610 7026 18622
rect 7086 18674 7138 18686
rect 7086 18610 7138 18622
rect 8654 18674 8706 18686
rect 8654 18610 8706 18622
rect 8878 18674 8930 18686
rect 11454 18674 11506 18686
rect 40126 18674 40178 18686
rect 10434 18622 10446 18674
rect 10498 18622 10510 18674
rect 27122 18622 27134 18674
rect 27186 18622 27198 18674
rect 27346 18622 27358 18674
rect 27410 18622 27422 18674
rect 8878 18610 8930 18622
rect 11454 18610 11506 18622
rect 40126 18610 40178 18622
rect 8094 18562 8146 18574
rect 5954 18510 5966 18562
rect 6018 18510 6030 18562
rect 8094 18498 8146 18510
rect 11342 18562 11394 18574
rect 11342 18498 11394 18510
rect 13582 18562 13634 18574
rect 13582 18498 13634 18510
rect 17614 18562 17666 18574
rect 24334 18562 24386 18574
rect 33518 18562 33570 18574
rect 44606 18562 44658 18574
rect 20066 18510 20078 18562
rect 20130 18510 20142 18562
rect 28354 18510 28366 18562
rect 28418 18510 28430 18562
rect 41122 18510 41134 18562
rect 41186 18510 41198 18562
rect 44258 18510 44270 18562
rect 44322 18510 44334 18562
rect 17614 18498 17666 18510
rect 24334 18498 24386 18510
rect 33518 18498 33570 18510
rect 44606 18498 44658 18510
rect 45838 18562 45890 18574
rect 45838 18498 45890 18510
rect 47070 18562 47122 18574
rect 47070 18498 47122 18510
rect 7198 18450 7250 18462
rect 2818 18398 2830 18450
rect 2882 18398 2894 18450
rect 3490 18398 3502 18450
rect 3554 18398 3566 18450
rect 6178 18398 6190 18450
rect 6242 18398 6254 18450
rect 6738 18398 6750 18450
rect 6802 18398 6814 18450
rect 7198 18386 7250 18398
rect 7310 18450 7362 18462
rect 7310 18386 7362 18398
rect 7870 18450 7922 18462
rect 7870 18386 7922 18398
rect 8542 18450 8594 18462
rect 8542 18386 8594 18398
rect 9998 18450 10050 18462
rect 10558 18450 10610 18462
rect 10322 18398 10334 18450
rect 10386 18398 10398 18450
rect 9998 18386 10050 18398
rect 10558 18386 10610 18398
rect 10782 18450 10834 18462
rect 10782 18386 10834 18398
rect 11006 18450 11058 18462
rect 11006 18386 11058 18398
rect 11678 18450 11730 18462
rect 11678 18386 11730 18398
rect 13358 18450 13410 18462
rect 13358 18386 13410 18398
rect 14702 18450 14754 18462
rect 14702 18386 14754 18398
rect 17390 18450 17442 18462
rect 17390 18386 17442 18398
rect 17950 18450 18002 18462
rect 24110 18450 24162 18462
rect 19282 18398 19294 18450
rect 19346 18398 19358 18450
rect 22866 18398 22878 18450
rect 22930 18398 22942 18450
rect 17950 18386 18002 18398
rect 24110 18386 24162 18398
rect 25342 18450 25394 18462
rect 33854 18450 33906 18462
rect 41470 18450 41522 18462
rect 27570 18398 27582 18450
rect 27634 18398 27646 18450
rect 28242 18398 28254 18450
rect 28306 18398 28318 18450
rect 29698 18398 29710 18450
rect 29762 18398 29774 18450
rect 30370 18398 30382 18450
rect 30434 18398 30446 18450
rect 36866 18398 36878 18450
rect 36930 18398 36942 18450
rect 25342 18386 25394 18398
rect 33854 18386 33906 18398
rect 41470 18386 41522 18398
rect 41806 18450 41858 18462
rect 44718 18450 44770 18462
rect 42914 18398 42926 18450
rect 42978 18398 42990 18450
rect 43474 18398 43486 18450
rect 43538 18398 43550 18450
rect 44034 18398 44046 18450
rect 44098 18398 44110 18450
rect 41806 18386 41858 18398
rect 44718 18386 44770 18398
rect 44830 18450 44882 18462
rect 47294 18450 47346 18462
rect 45154 18398 45166 18450
rect 45218 18398 45230 18450
rect 45602 18398 45614 18450
rect 45666 18398 45678 18450
rect 46722 18398 46734 18450
rect 46786 18398 46798 18450
rect 48066 18398 48078 18450
rect 48130 18398 48142 18450
rect 44830 18386 44882 18398
rect 47294 18386 47346 18398
rect 17838 18338 17890 18350
rect 23886 18338 23938 18350
rect 5618 18286 5630 18338
rect 5682 18286 5694 18338
rect 8194 18286 8206 18338
rect 8258 18286 8270 18338
rect 13682 18286 13694 18338
rect 13746 18286 13758 18338
rect 22194 18286 22206 18338
rect 22258 18286 22270 18338
rect 23090 18286 23102 18338
rect 23154 18286 23166 18338
rect 17838 18274 17890 18286
rect 23886 18274 23938 18286
rect 24222 18338 24274 18350
rect 41918 18338 41970 18350
rect 32498 18286 32510 18338
rect 32562 18286 32574 18338
rect 37538 18286 37550 18338
rect 37602 18286 37614 18338
rect 39666 18286 39678 18338
rect 39730 18286 39742 18338
rect 24222 18274 24274 18286
rect 41918 18274 41970 18286
rect 42590 18338 42642 18350
rect 42590 18274 42642 18286
rect 46286 18338 46338 18350
rect 46286 18274 46338 18286
rect 47182 18338 47234 18350
rect 47182 18274 47234 18286
rect 47630 18338 47682 18350
rect 47630 18274 47682 18286
rect 13918 18226 13970 18238
rect 13918 18162 13970 18174
rect 14142 18226 14194 18238
rect 14142 18162 14194 18174
rect 23662 18226 23714 18238
rect 23662 18162 23714 18174
rect 25230 18226 25282 18238
rect 43138 18174 43150 18226
rect 43202 18174 43214 18226
rect 46050 18174 46062 18226
rect 46114 18223 46126 18226
rect 46498 18223 46510 18226
rect 46114 18177 46510 18223
rect 46114 18174 46126 18177
rect 46498 18174 46510 18177
rect 46562 18174 46574 18226
rect 25230 18162 25282 18174
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 1934 17890 1986 17902
rect 1934 17826 1986 17838
rect 15262 17890 15314 17902
rect 15262 17826 15314 17838
rect 22654 17890 22706 17902
rect 22654 17826 22706 17838
rect 26574 17890 26626 17902
rect 42702 17890 42754 17902
rect 30930 17838 30942 17890
rect 30994 17838 31006 17890
rect 26574 17826 26626 17838
rect 42702 17826 42754 17838
rect 6862 17778 6914 17790
rect 16270 17778 16322 17790
rect 34190 17778 34242 17790
rect 42254 17778 42306 17790
rect 11778 17726 11790 17778
rect 11842 17726 11854 17778
rect 14914 17726 14926 17778
rect 14978 17726 14990 17778
rect 19282 17726 19294 17778
rect 19346 17726 19358 17778
rect 29922 17726 29934 17778
rect 29986 17726 29998 17778
rect 36082 17726 36094 17778
rect 36146 17726 36158 17778
rect 40226 17726 40238 17778
rect 40290 17726 40302 17778
rect 6862 17714 6914 17726
rect 16270 17714 16322 17726
rect 34190 17714 34242 17726
rect 42254 17714 42306 17726
rect 44158 17778 44210 17790
rect 45602 17726 45614 17778
rect 45666 17726 45678 17778
rect 44158 17714 44210 17726
rect 6974 17666 7026 17678
rect 13582 17666 13634 17678
rect 4162 17614 4174 17666
rect 4226 17614 4238 17666
rect 6514 17614 6526 17666
rect 6578 17614 6590 17666
rect 10882 17614 10894 17666
rect 10946 17614 10958 17666
rect 6974 17602 7026 17614
rect 13582 17602 13634 17614
rect 14030 17666 14082 17678
rect 16046 17666 16098 17678
rect 15810 17614 15822 17666
rect 15874 17614 15886 17666
rect 14030 17602 14082 17614
rect 16046 17602 16098 17614
rect 17054 17666 17106 17678
rect 17054 17602 17106 17614
rect 17390 17666 17442 17678
rect 23662 17666 23714 17678
rect 20738 17614 20750 17666
rect 20802 17614 20814 17666
rect 17390 17602 17442 17614
rect 23662 17602 23714 17614
rect 23886 17666 23938 17678
rect 23886 17602 23938 17614
rect 23998 17666 24050 17678
rect 23998 17602 24050 17614
rect 25342 17666 25394 17678
rect 30494 17666 30546 17678
rect 34078 17666 34130 17678
rect 34750 17666 34802 17678
rect 43150 17666 43202 17678
rect 25890 17614 25902 17666
rect 25954 17614 25966 17666
rect 26786 17614 26798 17666
rect 26850 17614 26862 17666
rect 29362 17614 29374 17666
rect 29426 17614 29438 17666
rect 29586 17614 29598 17666
rect 29650 17614 29662 17666
rect 30706 17614 30718 17666
rect 30770 17614 30782 17666
rect 34402 17614 34414 17666
rect 34466 17614 34478 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 38210 17614 38222 17666
rect 38274 17614 38286 17666
rect 43026 17614 43038 17666
rect 43090 17614 43102 17666
rect 25342 17602 25394 17614
rect 30494 17602 30546 17614
rect 34078 17602 34130 17614
rect 34750 17602 34802 17614
rect 43150 17602 43202 17614
rect 44270 17666 44322 17678
rect 46622 17666 46674 17678
rect 44818 17614 44830 17666
rect 44882 17614 44894 17666
rect 45714 17614 45726 17666
rect 45778 17614 45790 17666
rect 44270 17602 44322 17614
rect 46622 17602 46674 17614
rect 46958 17666 47010 17678
rect 46958 17602 47010 17614
rect 47182 17666 47234 17678
rect 47842 17614 47854 17666
rect 47906 17614 47918 17666
rect 47182 17602 47234 17614
rect 7198 17554 7250 17566
rect 7198 17490 7250 17502
rect 15038 17554 15090 17566
rect 15038 17490 15090 17502
rect 15598 17554 15650 17566
rect 15598 17490 15650 17502
rect 16494 17554 16546 17566
rect 16494 17490 16546 17502
rect 16830 17554 16882 17566
rect 16830 17490 16882 17502
rect 22542 17554 22594 17566
rect 22542 17490 22594 17502
rect 24222 17554 24274 17566
rect 35758 17554 35810 17566
rect 25554 17502 25566 17554
rect 25618 17502 25630 17554
rect 24222 17490 24274 17502
rect 35758 17490 35810 17502
rect 36206 17554 36258 17566
rect 36206 17490 36258 17502
rect 36430 17554 36482 17566
rect 46050 17502 46062 17554
rect 46114 17502 46126 17554
rect 47618 17502 47630 17554
rect 47682 17502 47694 17554
rect 36430 17490 36482 17502
rect 5854 17442 5906 17454
rect 5854 17378 5906 17390
rect 6750 17442 6802 17454
rect 6750 17378 6802 17390
rect 14702 17442 14754 17454
rect 17166 17442 17218 17454
rect 15922 17390 15934 17442
rect 15986 17390 15998 17442
rect 14702 17378 14754 17390
rect 17166 17378 17218 17390
rect 17278 17442 17330 17454
rect 17278 17378 17330 17390
rect 21422 17442 21474 17454
rect 21422 17378 21474 17390
rect 21870 17442 21922 17454
rect 21870 17378 21922 17390
rect 23774 17442 23826 17454
rect 23774 17378 23826 17390
rect 34302 17442 34354 17454
rect 34302 17378 34354 17390
rect 37214 17442 37266 17454
rect 42366 17442 42418 17454
rect 37874 17390 37886 17442
rect 37938 17390 37950 17442
rect 37214 17378 37266 17390
rect 42366 17378 42418 17390
rect 43262 17442 43314 17454
rect 43262 17378 43314 17390
rect 43374 17442 43426 17454
rect 46734 17442 46786 17454
rect 44930 17390 44942 17442
rect 44994 17390 45006 17442
rect 43374 17378 43426 17390
rect 46734 17378 46786 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 5742 17106 5794 17118
rect 5742 17042 5794 17054
rect 16046 17106 16098 17118
rect 27134 17106 27186 17118
rect 39230 17106 39282 17118
rect 18050 17054 18062 17106
rect 18114 17054 18126 17106
rect 22754 17054 22766 17106
rect 22818 17054 22830 17106
rect 25554 17054 25566 17106
rect 25618 17054 25630 17106
rect 33506 17054 33518 17106
rect 33570 17054 33582 17106
rect 16046 17042 16098 17054
rect 27134 17042 27186 17054
rect 39230 17042 39282 17054
rect 40126 17106 40178 17118
rect 40126 17042 40178 17054
rect 43038 17106 43090 17118
rect 43038 17042 43090 17054
rect 44046 17106 44098 17118
rect 44046 17042 44098 17054
rect 44270 17106 44322 17118
rect 44270 17042 44322 17054
rect 44942 17106 44994 17118
rect 44942 17042 44994 17054
rect 6414 16994 6466 17006
rect 14366 16994 14418 17006
rect 6738 16942 6750 16994
rect 6802 16942 6814 16994
rect 6414 16930 6466 16942
rect 14366 16930 14418 16942
rect 15934 16994 15986 17006
rect 15934 16930 15986 16942
rect 16494 16994 16546 17006
rect 25454 16994 25506 17006
rect 28030 16994 28082 17006
rect 23650 16942 23662 16994
rect 23714 16942 23726 16994
rect 26562 16942 26574 16994
rect 26626 16942 26638 16994
rect 16494 16930 16546 16942
rect 25454 16930 25506 16942
rect 28030 16930 28082 16942
rect 29598 16994 29650 17006
rect 38782 16994 38834 17006
rect 43822 16994 43874 17006
rect 35410 16942 35422 16994
rect 35474 16942 35486 16994
rect 39778 16942 39790 16994
rect 39842 16942 39854 16994
rect 41010 16942 41022 16994
rect 41074 16942 41086 16994
rect 29598 16930 29650 16942
rect 38782 16930 38834 16942
rect 43822 16930 43874 16942
rect 8878 16882 8930 16894
rect 1810 16830 1822 16882
rect 1874 16830 1886 16882
rect 5282 16830 5294 16882
rect 5346 16830 5358 16882
rect 7410 16830 7422 16882
rect 7474 16830 7486 16882
rect 8418 16830 8430 16882
rect 8482 16830 8494 16882
rect 8878 16818 8930 16830
rect 10446 16882 10498 16894
rect 10446 16818 10498 16830
rect 10558 16882 10610 16894
rect 10558 16818 10610 16830
rect 10894 16882 10946 16894
rect 16158 16882 16210 16894
rect 17502 16882 17554 16894
rect 22430 16882 22482 16894
rect 27022 16882 27074 16894
rect 13570 16830 13582 16882
rect 13634 16830 13646 16882
rect 14914 16830 14926 16882
rect 14978 16830 14990 16882
rect 16818 16830 16830 16882
rect 16882 16830 16894 16882
rect 20962 16830 20974 16882
rect 21026 16830 21038 16882
rect 21410 16830 21422 16882
rect 21474 16830 21486 16882
rect 23090 16830 23102 16882
rect 23154 16830 23166 16882
rect 23874 16830 23886 16882
rect 23938 16830 23950 16882
rect 25666 16830 25678 16882
rect 25730 16830 25742 16882
rect 26114 16830 26126 16882
rect 26178 16830 26190 16882
rect 10894 16818 10946 16830
rect 16158 16818 16210 16830
rect 17502 16818 17554 16830
rect 22430 16818 22482 16830
rect 27022 16818 27074 16830
rect 27358 16882 27410 16894
rect 33854 16882 33906 16894
rect 28242 16830 28254 16882
rect 28306 16830 28318 16882
rect 28802 16830 28814 16882
rect 28866 16830 28878 16882
rect 30482 16830 30494 16882
rect 30546 16830 30558 16882
rect 31714 16830 31726 16882
rect 31778 16830 31790 16882
rect 27358 16818 27410 16830
rect 33854 16818 33906 16830
rect 34078 16882 34130 16894
rect 39006 16882 39058 16894
rect 34626 16830 34638 16882
rect 34690 16830 34702 16882
rect 34078 16818 34130 16830
rect 39006 16818 39058 16830
rect 39342 16882 39394 16894
rect 43262 16882 43314 16894
rect 44830 16882 44882 16894
rect 40898 16830 40910 16882
rect 40962 16830 40974 16882
rect 42130 16830 42142 16882
rect 42194 16830 42206 16882
rect 42354 16830 42366 16882
rect 42418 16830 42430 16882
rect 42802 16830 42814 16882
rect 42866 16830 42878 16882
rect 43474 16830 43486 16882
rect 43538 16830 43550 16882
rect 44482 16830 44494 16882
rect 44546 16830 44558 16882
rect 45602 16830 45614 16882
rect 45666 16830 45678 16882
rect 39342 16818 39394 16830
rect 43262 16818 43314 16830
rect 44830 16818 44882 16830
rect 5070 16770 5122 16782
rect 10782 16770 10834 16782
rect 15486 16770 15538 16782
rect 17726 16770 17778 16782
rect 27694 16770 27746 16782
rect 2482 16718 2494 16770
rect 2546 16718 2558 16770
rect 4610 16718 4622 16770
rect 4674 16718 4686 16770
rect 7634 16718 7646 16770
rect 7698 16718 7710 16770
rect 12562 16718 12574 16770
rect 12626 16718 12638 16770
rect 16706 16718 16718 16770
rect 16770 16718 16782 16770
rect 19842 16718 19854 16770
rect 19906 16718 19918 16770
rect 21746 16718 21758 16770
rect 21810 16718 21822 16770
rect 23986 16718 23998 16770
rect 24050 16718 24062 16770
rect 5070 16706 5122 16718
rect 10782 16706 10834 16718
rect 15486 16706 15538 16718
rect 17726 16706 17778 16718
rect 27694 16706 27746 16718
rect 28142 16770 28194 16782
rect 39118 16770 39170 16782
rect 37538 16718 37550 16770
rect 37602 16718 37614 16770
rect 41458 16718 41470 16770
rect 41522 16718 41534 16770
rect 43026 16718 43038 16770
rect 43090 16718 43102 16770
rect 44370 16718 44382 16770
rect 44434 16718 44446 16770
rect 28142 16706 28194 16718
rect 39118 16706 39170 16718
rect 4958 16658 5010 16670
rect 14478 16658 14530 16670
rect 8194 16606 8206 16658
rect 8258 16606 8270 16658
rect 4958 16594 5010 16606
rect 14478 16594 14530 16606
rect 14702 16658 14754 16670
rect 47966 16658 48018 16670
rect 28578 16606 28590 16658
rect 28642 16606 28654 16658
rect 14702 16594 14754 16606
rect 47966 16594 48018 16606
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 1934 16322 1986 16334
rect 1934 16258 1986 16270
rect 7310 16322 7362 16334
rect 7310 16258 7362 16270
rect 13470 16322 13522 16334
rect 13470 16258 13522 16270
rect 29934 16322 29986 16334
rect 29934 16258 29986 16270
rect 38110 16322 38162 16334
rect 38110 16258 38162 16270
rect 4958 16210 5010 16222
rect 16158 16210 16210 16222
rect 8194 16158 8206 16210
rect 8258 16158 8270 16210
rect 9762 16158 9774 16210
rect 9826 16158 9838 16210
rect 13794 16158 13806 16210
rect 13858 16158 13870 16210
rect 4958 16146 5010 16158
rect 16158 16146 16210 16158
rect 19070 16210 19122 16222
rect 25230 16210 25282 16222
rect 21746 16158 21758 16210
rect 21810 16158 21822 16210
rect 19070 16146 19122 16158
rect 25230 16146 25282 16158
rect 29598 16210 29650 16222
rect 34302 16210 34354 16222
rect 31154 16158 31166 16210
rect 31218 16158 31230 16210
rect 29598 16146 29650 16158
rect 34302 16146 34354 16158
rect 36430 16210 36482 16222
rect 36430 16146 36482 16158
rect 37998 16210 38050 16222
rect 37998 16146 38050 16158
rect 38558 16210 38610 16222
rect 42366 16210 42418 16222
rect 40898 16158 40910 16210
rect 40962 16158 40974 16210
rect 38558 16146 38610 16158
rect 42366 16146 42418 16158
rect 43486 16210 43538 16222
rect 45826 16158 45838 16210
rect 45890 16158 45902 16210
rect 48066 16158 48078 16210
rect 48130 16158 48142 16210
rect 43486 16146 43538 16158
rect 7198 16098 7250 16110
rect 7870 16098 7922 16110
rect 4050 16046 4062 16098
rect 4114 16046 4126 16098
rect 6402 16046 6414 16098
rect 6466 16046 6478 16098
rect 7634 16046 7646 16098
rect 7698 16046 7710 16098
rect 7198 16034 7250 16046
rect 7870 16034 7922 16046
rect 8094 16098 8146 16110
rect 8094 16034 8146 16046
rect 8766 16098 8818 16110
rect 19630 16098 19682 16110
rect 20526 16098 20578 16110
rect 9090 16046 9102 16098
rect 9154 16046 9166 16098
rect 10098 16046 10110 16098
rect 10162 16046 10174 16098
rect 11778 16046 11790 16098
rect 11842 16046 11854 16098
rect 12226 16046 12238 16098
rect 12290 16046 12302 16098
rect 15362 16046 15374 16098
rect 15426 16046 15438 16098
rect 16370 16046 16382 16098
rect 16434 16046 16446 16098
rect 18498 16046 18510 16098
rect 18562 16046 18574 16098
rect 20066 16046 20078 16098
rect 20130 16046 20142 16098
rect 8766 16034 8818 16046
rect 19630 16034 19682 16046
rect 20526 16034 20578 16046
rect 22094 16098 22146 16110
rect 22094 16034 22146 16046
rect 22878 16098 22930 16110
rect 22878 16034 22930 16046
rect 25118 16098 25170 16110
rect 25118 16034 25170 16046
rect 25342 16098 25394 16110
rect 25342 16034 25394 16046
rect 27582 16098 27634 16110
rect 27582 16034 27634 16046
rect 27918 16098 27970 16110
rect 27918 16034 27970 16046
rect 29710 16098 29762 16110
rect 36318 16098 36370 16110
rect 42478 16098 42530 16110
rect 32946 16046 32958 16098
rect 33010 16046 33022 16098
rect 35970 16046 35982 16098
rect 36034 16046 36046 16098
rect 40786 16046 40798 16098
rect 40850 16046 40862 16098
rect 41458 16046 41470 16098
rect 41522 16046 41534 16098
rect 41906 16046 41918 16098
rect 41970 16046 41982 16098
rect 29710 16034 29762 16046
rect 36318 16034 36370 16046
rect 42478 16034 42530 16046
rect 42814 16098 42866 16110
rect 45042 16046 45054 16098
rect 45106 16046 45118 16098
rect 42814 16034 42866 16046
rect 14254 15986 14306 15998
rect 17390 15986 17442 15998
rect 18062 15986 18114 15998
rect 6178 15934 6190 15986
rect 6242 15934 6254 15986
rect 9986 15934 9998 15986
rect 10050 15934 10062 15986
rect 11330 15934 11342 15986
rect 11394 15934 11406 15986
rect 12898 15928 12910 15980
rect 12962 15928 12974 15980
rect 14578 15934 14590 15986
rect 14642 15934 14654 15986
rect 15474 15934 15486 15986
rect 15538 15934 15550 15986
rect 16146 15934 16158 15986
rect 16210 15934 16222 15986
rect 17714 15934 17726 15986
rect 17778 15934 17790 15986
rect 14254 15922 14306 15934
rect 17390 15922 17442 15934
rect 18062 15922 18114 15934
rect 18734 15986 18786 15998
rect 18734 15922 18786 15934
rect 21422 15986 21474 15998
rect 21422 15922 21474 15934
rect 21646 15986 21698 15998
rect 21646 15922 21698 15934
rect 25566 15986 25618 15998
rect 25566 15922 25618 15934
rect 28478 15986 28530 15998
rect 28478 15922 28530 15934
rect 28590 15986 28642 15998
rect 28590 15922 28642 15934
rect 30270 15986 30322 15998
rect 30270 15922 30322 15934
rect 38446 15986 38498 15998
rect 42254 15986 42306 15998
rect 40450 15934 40462 15986
rect 40514 15934 40526 15986
rect 43810 15934 43822 15986
rect 43874 15934 43886 15986
rect 38446 15922 38498 15934
rect 42254 15922 42306 15934
rect 8206 15874 8258 15886
rect 13694 15874 13746 15886
rect 12786 15822 12798 15874
rect 12850 15822 12862 15874
rect 8206 15810 8258 15822
rect 13694 15810 13746 15822
rect 14926 15874 14978 15886
rect 27694 15874 27746 15886
rect 22418 15822 22430 15874
rect 22482 15822 22494 15874
rect 14926 15810 14978 15822
rect 27694 15810 27746 15822
rect 30046 15874 30098 15886
rect 30046 15810 30098 15822
rect 43374 15874 43426 15886
rect 43374 15810 43426 15822
rect 44158 15874 44210 15886
rect 44158 15810 44210 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 6302 15538 6354 15550
rect 6302 15474 6354 15486
rect 11454 15538 11506 15550
rect 11454 15474 11506 15486
rect 11566 15538 11618 15550
rect 11566 15474 11618 15486
rect 12686 15538 12738 15550
rect 16942 15538 16994 15550
rect 15138 15486 15150 15538
rect 15202 15486 15214 15538
rect 12686 15474 12738 15486
rect 16942 15474 16994 15486
rect 25678 15538 25730 15550
rect 25678 15474 25730 15486
rect 33294 15538 33346 15550
rect 33294 15474 33346 15486
rect 33406 15538 33458 15550
rect 33406 15474 33458 15486
rect 34190 15538 34242 15550
rect 34190 15474 34242 15486
rect 37102 15538 37154 15550
rect 37102 15474 37154 15486
rect 37438 15538 37490 15550
rect 37438 15474 37490 15486
rect 40798 15538 40850 15550
rect 40798 15474 40850 15486
rect 42030 15538 42082 15550
rect 42030 15474 42082 15486
rect 42254 15538 42306 15550
rect 42254 15474 42306 15486
rect 43038 15538 43090 15550
rect 45726 15538 45778 15550
rect 44258 15486 44270 15538
rect 44322 15486 44334 15538
rect 45154 15486 45166 15538
rect 45218 15486 45230 15538
rect 43038 15474 43090 15486
rect 45726 15474 45778 15486
rect 46398 15538 46450 15550
rect 47854 15538 47906 15550
rect 47506 15486 47518 15538
rect 47570 15486 47582 15538
rect 46398 15474 46450 15486
rect 47854 15474 47906 15486
rect 3390 15426 3442 15438
rect 3390 15362 3442 15374
rect 3838 15426 3890 15438
rect 3838 15362 3890 15374
rect 4174 15426 4226 15438
rect 4174 15362 4226 15374
rect 5182 15426 5234 15438
rect 5182 15362 5234 15374
rect 5294 15426 5346 15438
rect 5294 15362 5346 15374
rect 6190 15426 6242 15438
rect 6190 15362 6242 15374
rect 7086 15426 7138 15438
rect 7086 15362 7138 15374
rect 7758 15426 7810 15438
rect 14142 15426 14194 15438
rect 25230 15426 25282 15438
rect 8754 15374 8766 15426
rect 8818 15374 8830 15426
rect 21746 15374 21758 15426
rect 21810 15374 21822 15426
rect 7758 15362 7810 15374
rect 14142 15362 14194 15374
rect 25230 15362 25282 15374
rect 27358 15426 27410 15438
rect 32174 15426 32226 15438
rect 31042 15374 31054 15426
rect 31106 15374 31118 15426
rect 27358 15362 27410 15374
rect 32174 15362 32226 15374
rect 38222 15426 38274 15438
rect 38222 15362 38274 15374
rect 38558 15426 38610 15438
rect 38558 15362 38610 15374
rect 38894 15426 38946 15438
rect 41346 15374 41358 15426
rect 41410 15374 41422 15426
rect 41682 15374 41694 15426
rect 41746 15374 41758 15426
rect 43922 15374 43934 15426
rect 43986 15374 43998 15426
rect 38894 15362 38946 15374
rect 3278 15314 3330 15326
rect 2930 15262 2942 15314
rect 2994 15262 3006 15314
rect 3278 15250 3330 15262
rect 4398 15314 4450 15326
rect 6974 15314 7026 15326
rect 9998 15314 10050 15326
rect 5506 15262 5518 15314
rect 5570 15262 5582 15314
rect 7634 15262 7646 15314
rect 7698 15262 7710 15314
rect 8978 15262 8990 15314
rect 9042 15262 9054 15314
rect 4398 15250 4450 15262
rect 6974 15250 7026 15262
rect 9998 15250 10050 15262
rect 10222 15314 10274 15326
rect 10222 15250 10274 15262
rect 10446 15314 10498 15326
rect 10446 15250 10498 15262
rect 10670 15314 10722 15326
rect 10670 15250 10722 15262
rect 11006 15314 11058 15326
rect 11006 15250 11058 15262
rect 11678 15314 11730 15326
rect 11678 15250 11730 15262
rect 12238 15314 12290 15326
rect 12238 15250 12290 15262
rect 12462 15314 12514 15326
rect 12462 15250 12514 15262
rect 12910 15314 12962 15326
rect 12910 15250 12962 15262
rect 13694 15314 13746 15326
rect 13694 15250 13746 15262
rect 13806 15314 13858 15326
rect 13806 15250 13858 15262
rect 14254 15314 14306 15326
rect 14254 15250 14306 15262
rect 15486 15314 15538 15326
rect 15486 15250 15538 15262
rect 16158 15314 16210 15326
rect 25454 15314 25506 15326
rect 20178 15262 20190 15314
rect 20242 15262 20254 15314
rect 20962 15262 20974 15314
rect 21026 15262 21038 15314
rect 16158 15250 16210 15262
rect 25454 15250 25506 15262
rect 25790 15314 25842 15326
rect 25790 15250 25842 15262
rect 26126 15314 26178 15326
rect 26126 15250 26178 15262
rect 26462 15314 26514 15326
rect 26462 15250 26514 15262
rect 26686 15314 26738 15326
rect 26686 15250 26738 15262
rect 27470 15314 27522 15326
rect 33182 15314 33234 15326
rect 31826 15262 31838 15314
rect 31890 15262 31902 15314
rect 32386 15262 32398 15314
rect 32450 15262 32462 15314
rect 27470 15250 27522 15262
rect 33182 15250 33234 15262
rect 33854 15314 33906 15326
rect 33854 15250 33906 15262
rect 34078 15314 34130 15326
rect 34078 15250 34130 15262
rect 34414 15314 34466 15326
rect 34414 15250 34466 15262
rect 34638 15314 34690 15326
rect 39118 15314 39170 15326
rect 37426 15262 37438 15314
rect 37490 15262 37502 15314
rect 37986 15262 37998 15314
rect 38050 15262 38062 15314
rect 34638 15250 34690 15262
rect 39118 15250 39170 15262
rect 41022 15314 41074 15326
rect 41022 15250 41074 15262
rect 41806 15314 41858 15326
rect 41806 15250 41858 15262
rect 42366 15314 42418 15326
rect 43150 15314 43202 15326
rect 42802 15262 42814 15314
rect 42866 15262 42878 15314
rect 42366 15250 42418 15262
rect 43150 15250 43202 15262
rect 43262 15314 43314 15326
rect 43262 15250 43314 15262
rect 43374 15314 43426 15326
rect 45614 15314 45666 15326
rect 44370 15262 44382 15314
rect 44434 15262 44446 15314
rect 45266 15262 45278 15314
rect 45330 15262 45342 15314
rect 43374 15250 43426 15262
rect 45614 15250 45666 15262
rect 46958 15314 47010 15326
rect 46958 15250 47010 15262
rect 3950 15202 4002 15214
rect 10558 15202 10610 15214
rect 15710 15202 15762 15214
rect 25566 15202 25618 15214
rect 8306 15150 8318 15202
rect 8370 15150 8382 15202
rect 14690 15150 14702 15202
rect 14754 15150 14766 15202
rect 17378 15150 17390 15202
rect 17442 15150 17454 15202
rect 19506 15150 19518 15202
rect 19570 15150 19582 15202
rect 23874 15150 23886 15202
rect 23938 15150 23950 15202
rect 3950 15138 4002 15150
rect 10558 15138 10610 15150
rect 15710 15138 15762 15150
rect 25566 15138 25618 15150
rect 26350 15202 26402 15214
rect 38670 15202 38722 15214
rect 28914 15150 28926 15202
rect 28978 15150 28990 15202
rect 26350 15138 26402 15150
rect 38670 15138 38722 15150
rect 47070 15202 47122 15214
rect 47070 15138 47122 15150
rect 7086 15090 7138 15102
rect 4722 15038 4734 15090
rect 4786 15038 4798 15090
rect 7086 15026 7138 15038
rect 12350 15090 12402 15102
rect 12350 15026 12402 15038
rect 27358 15090 27410 15102
rect 27358 15026 27410 15038
rect 37774 15090 37826 15102
rect 37774 15026 37826 15038
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 4062 14754 4114 14766
rect 4062 14690 4114 14702
rect 11118 14754 11170 14766
rect 11118 14690 11170 14702
rect 11566 14754 11618 14766
rect 11566 14690 11618 14702
rect 12014 14754 12066 14766
rect 12014 14690 12066 14702
rect 17614 14754 17666 14766
rect 17614 14690 17666 14702
rect 18174 14754 18226 14766
rect 18174 14690 18226 14702
rect 18510 14754 18562 14766
rect 18510 14690 18562 14702
rect 25902 14754 25954 14766
rect 25902 14690 25954 14702
rect 27022 14754 27074 14766
rect 27022 14690 27074 14702
rect 15262 14642 15314 14654
rect 15262 14578 15314 14590
rect 21310 14642 21362 14654
rect 21310 14578 21362 14590
rect 24782 14642 24834 14654
rect 24782 14578 24834 14590
rect 26798 14642 26850 14654
rect 26798 14578 26850 14590
rect 29486 14642 29538 14654
rect 29486 14578 29538 14590
rect 32174 14642 32226 14654
rect 32174 14578 32226 14590
rect 35646 14642 35698 14654
rect 35646 14578 35698 14590
rect 44270 14642 44322 14654
rect 44270 14578 44322 14590
rect 3726 14530 3778 14542
rect 3726 14466 3778 14478
rect 3950 14530 4002 14542
rect 3950 14466 4002 14478
rect 5070 14530 5122 14542
rect 5070 14466 5122 14478
rect 6750 14530 6802 14542
rect 6750 14466 6802 14478
rect 8766 14530 8818 14542
rect 8766 14466 8818 14478
rect 11342 14530 11394 14542
rect 15486 14530 15538 14542
rect 18062 14530 18114 14542
rect 13458 14478 13470 14530
rect 13522 14478 13534 14530
rect 14802 14478 14814 14530
rect 14866 14478 14878 14530
rect 17602 14478 17614 14530
rect 17666 14478 17678 14530
rect 11342 14466 11394 14478
rect 15486 14466 15538 14478
rect 18062 14466 18114 14478
rect 18398 14530 18450 14542
rect 18398 14466 18450 14478
rect 19182 14530 19234 14542
rect 19182 14466 19234 14478
rect 19630 14530 19682 14542
rect 22206 14530 22258 14542
rect 21746 14478 21758 14530
rect 21810 14478 21822 14530
rect 19630 14466 19682 14478
rect 22206 14466 22258 14478
rect 26238 14530 26290 14542
rect 27694 14530 27746 14542
rect 27346 14478 27358 14530
rect 27410 14478 27422 14530
rect 26238 14466 26290 14478
rect 27694 14466 27746 14478
rect 29374 14530 29426 14542
rect 29374 14466 29426 14478
rect 29710 14530 29762 14542
rect 31278 14530 31330 14542
rect 31042 14478 31054 14530
rect 31106 14478 31118 14530
rect 29710 14466 29762 14478
rect 31278 14466 31330 14478
rect 31502 14530 31554 14542
rect 31502 14466 31554 14478
rect 33182 14530 33234 14542
rect 35422 14530 35474 14542
rect 35186 14478 35198 14530
rect 35250 14478 35262 14530
rect 33182 14466 33234 14478
rect 35422 14466 35474 14478
rect 38110 14530 38162 14542
rect 38110 14466 38162 14478
rect 38446 14530 38498 14542
rect 41570 14478 41582 14530
rect 41634 14478 41646 14530
rect 45042 14478 45054 14530
rect 45106 14478 45118 14530
rect 46274 14478 46286 14530
rect 46338 14478 46350 14530
rect 48066 14478 48078 14530
rect 48130 14478 48142 14530
rect 38446 14466 38498 14478
rect 3614 14418 3666 14430
rect 3614 14354 3666 14366
rect 4958 14418 5010 14430
rect 4958 14354 5010 14366
rect 5630 14418 5682 14430
rect 7870 14418 7922 14430
rect 5954 14366 5966 14418
rect 6018 14366 6030 14418
rect 5630 14354 5682 14366
rect 7870 14354 7922 14366
rect 9326 14418 9378 14430
rect 9326 14354 9378 14366
rect 10894 14418 10946 14430
rect 10894 14354 10946 14366
rect 12574 14418 12626 14430
rect 12574 14354 12626 14366
rect 12686 14418 12738 14430
rect 12686 14354 12738 14366
rect 13694 14418 13746 14430
rect 17278 14418 17330 14430
rect 14466 14366 14478 14418
rect 14530 14366 14542 14418
rect 13694 14354 13746 14366
rect 17278 14354 17330 14366
rect 25118 14418 25170 14430
rect 25118 14354 25170 14366
rect 25566 14418 25618 14430
rect 25566 14354 25618 14366
rect 26350 14418 26402 14430
rect 26350 14354 26402 14366
rect 29150 14418 29202 14430
rect 29150 14354 29202 14366
rect 31726 14418 31778 14430
rect 31726 14354 31778 14366
rect 32846 14418 32898 14430
rect 32846 14354 32898 14366
rect 32958 14418 33010 14430
rect 34862 14418 34914 14430
rect 34402 14366 34414 14418
rect 34466 14366 34478 14418
rect 32958 14354 33010 14366
rect 34862 14354 34914 14366
rect 34974 14418 35026 14430
rect 34974 14354 35026 14366
rect 35870 14418 35922 14430
rect 35870 14354 35922 14366
rect 36094 14418 36146 14430
rect 36094 14354 36146 14366
rect 38222 14418 38274 14430
rect 38222 14354 38274 14366
rect 41246 14418 41298 14430
rect 41246 14354 41298 14366
rect 44830 14418 44882 14430
rect 44830 14354 44882 14366
rect 45726 14418 45778 14430
rect 47854 14418 47906 14430
rect 47058 14366 47070 14418
rect 47122 14366 47134 14418
rect 45726 14354 45778 14366
rect 47854 14354 47906 14366
rect 4622 14306 4674 14318
rect 12350 14306 12402 14318
rect 24222 14306 24274 14318
rect 10322 14254 10334 14306
rect 10386 14254 10398 14306
rect 13794 14254 13806 14306
rect 13858 14254 13870 14306
rect 15810 14254 15822 14306
rect 15874 14254 15886 14306
rect 18834 14254 18846 14306
rect 18898 14254 18910 14306
rect 4622 14242 4674 14254
rect 12350 14242 12402 14254
rect 24222 14242 24274 14254
rect 25230 14306 25282 14318
rect 25230 14242 25282 14254
rect 25790 14306 25842 14318
rect 25790 14242 25842 14254
rect 27470 14306 27522 14318
rect 27470 14242 27522 14254
rect 27582 14306 27634 14318
rect 27582 14242 27634 14254
rect 29598 14306 29650 14318
rect 29598 14242 29650 14254
rect 31390 14306 31442 14318
rect 31390 14242 31442 14254
rect 41358 14306 41410 14318
rect 41358 14242 41410 14254
rect 42030 14306 42082 14318
rect 42030 14242 42082 14254
rect 45838 14306 45890 14318
rect 45838 14242 45890 14254
rect 45950 14306 46002 14318
rect 45950 14242 46002 14254
rect 46846 14306 46898 14318
rect 46846 14242 46898 14254
rect 47406 14306 47458 14318
rect 47406 14242 47458 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 7422 13970 7474 13982
rect 7422 13906 7474 13918
rect 14142 13970 14194 13982
rect 14142 13906 14194 13918
rect 17726 13970 17778 13982
rect 17726 13906 17778 13918
rect 28142 13970 28194 13982
rect 28142 13906 28194 13918
rect 32398 13970 32450 13982
rect 32398 13906 32450 13918
rect 34638 13970 34690 13982
rect 34638 13906 34690 13918
rect 35310 13970 35362 13982
rect 35310 13906 35362 13918
rect 36094 13970 36146 13982
rect 36094 13906 36146 13918
rect 36430 13970 36482 13982
rect 36430 13906 36482 13918
rect 37102 13970 37154 13982
rect 37102 13906 37154 13918
rect 37550 13970 37602 13982
rect 44382 13970 44434 13982
rect 40338 13918 40350 13970
rect 40402 13918 40414 13970
rect 37550 13906 37602 13918
rect 44382 13906 44434 13918
rect 45502 13970 45554 13982
rect 45502 13906 45554 13918
rect 46398 13970 46450 13982
rect 46398 13906 46450 13918
rect 46622 13970 46674 13982
rect 46622 13906 46674 13918
rect 7086 13858 7138 13870
rect 2482 13806 2494 13858
rect 2546 13806 2558 13858
rect 7086 13794 7138 13806
rect 8654 13858 8706 13870
rect 9886 13858 9938 13870
rect 27470 13858 27522 13870
rect 9650 13806 9662 13858
rect 9714 13806 9726 13858
rect 12226 13806 12238 13858
rect 12290 13806 12302 13858
rect 12898 13806 12910 13858
rect 12962 13806 12974 13858
rect 8654 13794 8706 13806
rect 9886 13794 9938 13806
rect 27470 13794 27522 13806
rect 29486 13858 29538 13870
rect 35086 13858 35138 13870
rect 39790 13858 39842 13870
rect 31042 13806 31054 13858
rect 31106 13806 31118 13858
rect 37874 13806 37886 13858
rect 37938 13855 37950 13858
rect 37938 13809 38271 13855
rect 37938 13806 37950 13809
rect 29486 13794 29538 13806
rect 35086 13794 35138 13806
rect 7310 13746 7362 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 7310 13682 7362 13694
rect 7534 13746 7586 13758
rect 8206 13746 8258 13758
rect 7746 13694 7758 13746
rect 7810 13694 7822 13746
rect 7534 13682 7586 13694
rect 8206 13682 8258 13694
rect 8318 13746 8370 13758
rect 8318 13682 8370 13694
rect 10334 13746 10386 13758
rect 27358 13746 27410 13758
rect 12002 13694 12014 13746
rect 12066 13694 12078 13746
rect 13010 13694 13022 13746
rect 13074 13694 13086 13746
rect 13570 13694 13582 13746
rect 13634 13694 13646 13746
rect 20178 13694 20190 13746
rect 20242 13694 20254 13746
rect 10334 13682 10386 13694
rect 27358 13682 27410 13694
rect 27918 13746 27970 13758
rect 27918 13682 27970 13694
rect 28926 13746 28978 13758
rect 31502 13746 31554 13758
rect 29250 13694 29262 13746
rect 29314 13694 29326 13746
rect 28926 13682 28978 13694
rect 31502 13682 31554 13694
rect 31614 13746 31666 13758
rect 33854 13746 33906 13758
rect 34302 13746 34354 13758
rect 34974 13746 35026 13758
rect 31826 13694 31838 13746
rect 31890 13694 31902 13746
rect 34066 13694 34078 13746
rect 34130 13694 34142 13746
rect 34402 13694 34414 13746
rect 34466 13694 34478 13746
rect 31614 13682 31666 13694
rect 33854 13682 33906 13694
rect 34302 13682 34354 13694
rect 34974 13682 35026 13694
rect 35982 13746 36034 13758
rect 35982 13682 36034 13694
rect 36206 13746 36258 13758
rect 38225 13746 38271 13809
rect 38658 13806 38670 13858
rect 38722 13806 38734 13858
rect 39790 13794 39842 13806
rect 39902 13858 39954 13870
rect 39902 13794 39954 13806
rect 41134 13858 41186 13870
rect 41134 13794 41186 13806
rect 46174 13858 46226 13870
rect 46174 13794 46226 13806
rect 47854 13858 47906 13870
rect 47854 13794 47906 13806
rect 39678 13746 39730 13758
rect 37762 13694 37774 13746
rect 37826 13694 37838 13746
rect 38210 13694 38222 13746
rect 38274 13694 38286 13746
rect 36206 13682 36258 13694
rect 39678 13682 39730 13694
rect 40910 13746 40962 13758
rect 40910 13682 40962 13694
rect 41246 13746 41298 13758
rect 41918 13746 41970 13758
rect 41458 13694 41470 13746
rect 41522 13694 41534 13746
rect 41246 13682 41298 13694
rect 41918 13682 41970 13694
rect 42478 13746 42530 13758
rect 48190 13746 48242 13758
rect 42690 13694 42702 13746
rect 42754 13694 42766 13746
rect 46946 13694 46958 13746
rect 47010 13694 47022 13746
rect 42478 13682 42530 13694
rect 48190 13682 48242 13694
rect 5070 13634 5122 13646
rect 4610 13582 4622 13634
rect 4674 13582 4686 13634
rect 5070 13570 5122 13582
rect 8542 13634 8594 13646
rect 8542 13570 8594 13582
rect 9550 13634 9602 13646
rect 18734 13634 18786 13646
rect 24558 13634 24610 13646
rect 18162 13582 18174 13634
rect 18226 13582 18238 13634
rect 20850 13582 20862 13634
rect 20914 13582 20926 13634
rect 22978 13582 22990 13634
rect 23042 13582 23054 13634
rect 9550 13570 9602 13582
rect 18734 13570 18786 13582
rect 24558 13570 24610 13582
rect 27134 13634 27186 13646
rect 38334 13634 38386 13646
rect 29474 13582 29486 13634
rect 29538 13582 29550 13634
rect 27134 13570 27186 13582
rect 38334 13570 38386 13582
rect 44718 13634 44770 13646
rect 44718 13570 44770 13582
rect 46510 13634 46562 13646
rect 46510 13570 46562 13582
rect 47518 13634 47570 13646
rect 47518 13570 47570 13582
rect 10558 13522 10610 13534
rect 10558 13458 10610 13470
rect 37438 13522 37490 13534
rect 37438 13458 37490 13470
rect 42142 13522 42194 13534
rect 42142 13458 42194 13470
rect 42254 13522 42306 13534
rect 42254 13458 42306 13470
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 10446 13186 10498 13198
rect 10446 13122 10498 13134
rect 13470 13186 13522 13198
rect 13470 13122 13522 13134
rect 29486 13186 29538 13198
rect 29486 13122 29538 13134
rect 29934 13186 29986 13198
rect 29934 13122 29986 13134
rect 22094 13074 22146 13086
rect 28254 13074 28306 13086
rect 4386 13022 4398 13074
rect 4450 13022 4462 13074
rect 26562 13022 26574 13074
rect 26626 13022 26638 13074
rect 22094 13010 22146 13022
rect 28254 13010 28306 13022
rect 32062 13074 32114 13086
rect 32062 13010 32114 13022
rect 41134 13074 41186 13086
rect 47966 13074 48018 13086
rect 42130 13022 42142 13074
rect 42194 13022 42206 13074
rect 44258 13022 44270 13074
rect 44322 13022 44334 13074
rect 41134 13010 41186 13022
rect 47966 13010 48018 13022
rect 6302 12962 6354 12974
rect 6302 12898 6354 12910
rect 6526 12962 6578 12974
rect 6526 12898 6578 12910
rect 9998 12962 10050 12974
rect 13582 12962 13634 12974
rect 10098 12910 10110 12962
rect 10162 12910 10174 12962
rect 9998 12898 10050 12910
rect 13582 12898 13634 12910
rect 14478 12962 14530 12974
rect 14478 12898 14530 12910
rect 14702 12962 14754 12974
rect 14702 12898 14754 12910
rect 14926 12962 14978 12974
rect 14926 12898 14978 12910
rect 15710 12962 15762 12974
rect 15710 12898 15762 12910
rect 15934 12962 15986 12974
rect 28366 12962 28418 12974
rect 17826 12910 17838 12962
rect 17890 12910 17902 12962
rect 23426 12910 23438 12962
rect 23490 12910 23502 12962
rect 24098 12910 24110 12962
rect 24162 12910 24174 12962
rect 25218 12910 25230 12962
rect 25282 12910 25294 12962
rect 25666 12910 25678 12962
rect 25730 12910 25742 12962
rect 26226 12910 26238 12962
rect 26290 12910 26302 12962
rect 27906 12910 27918 12962
rect 27970 12910 27982 12962
rect 15934 12898 15986 12910
rect 28366 12898 28418 12910
rect 29598 12962 29650 12974
rect 29598 12898 29650 12910
rect 29822 12962 29874 12974
rect 29822 12898 29874 12910
rect 32286 12962 32338 12974
rect 32286 12898 32338 12910
rect 40126 12962 40178 12974
rect 40126 12898 40178 12910
rect 40238 12962 40290 12974
rect 40238 12898 40290 12910
rect 40574 12962 40626 12974
rect 41346 12910 41358 12962
rect 41410 12910 41422 12962
rect 45042 12910 45054 12962
rect 45106 12910 45118 12962
rect 40574 12898 40626 12910
rect 4734 12850 4786 12862
rect 4734 12786 4786 12798
rect 6078 12850 6130 12862
rect 15150 12850 15202 12862
rect 8978 12798 8990 12850
rect 9042 12798 9054 12850
rect 6078 12786 6130 12798
rect 15150 12786 15202 12798
rect 15822 12850 15874 12862
rect 15822 12786 15874 12798
rect 18734 12850 18786 12862
rect 18734 12786 18786 12798
rect 18846 12850 18898 12862
rect 18846 12786 18898 12798
rect 18958 12850 19010 12862
rect 23326 12850 23378 12862
rect 31950 12850 32002 12862
rect 22418 12798 22430 12850
rect 22482 12798 22494 12850
rect 24322 12798 24334 12850
rect 24386 12798 24398 12850
rect 24882 12798 24894 12850
rect 24946 12798 24958 12850
rect 27010 12798 27022 12850
rect 27074 12798 27086 12850
rect 18958 12786 19010 12798
rect 23326 12786 23378 12798
rect 31950 12786 32002 12798
rect 32510 12850 32562 12862
rect 45826 12798 45838 12850
rect 45890 12798 45902 12850
rect 32510 12786 32562 12798
rect 6190 12738 6242 12750
rect 6190 12674 6242 12686
rect 9326 12738 9378 12750
rect 9326 12674 9378 12686
rect 9774 12738 9826 12750
rect 9774 12674 9826 12686
rect 9886 12738 9938 12750
rect 9886 12674 9938 12686
rect 15038 12738 15090 12750
rect 22766 12738 22818 12750
rect 27246 12738 27298 12750
rect 16370 12686 16382 12738
rect 16434 12686 16446 12738
rect 18050 12686 18062 12738
rect 18114 12686 18126 12738
rect 19394 12686 19406 12738
rect 19458 12686 19470 12738
rect 24210 12686 24222 12738
rect 24274 12686 24286 12738
rect 15038 12674 15090 12686
rect 22766 12674 22818 12686
rect 27246 12674 27298 12686
rect 28142 12738 28194 12750
rect 28142 12674 28194 12686
rect 28478 12738 28530 12750
rect 28478 12674 28530 12686
rect 40462 12738 40514 12750
rect 40462 12674 40514 12686
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 5294 12402 5346 12414
rect 5294 12338 5346 12350
rect 7310 12402 7362 12414
rect 7310 12338 7362 12350
rect 7758 12402 7810 12414
rect 7758 12338 7810 12350
rect 8878 12402 8930 12414
rect 8878 12338 8930 12350
rect 10558 12402 10610 12414
rect 10558 12338 10610 12350
rect 16158 12402 16210 12414
rect 16158 12338 16210 12350
rect 16270 12402 16322 12414
rect 16270 12338 16322 12350
rect 17502 12402 17554 12414
rect 17502 12338 17554 12350
rect 23998 12402 24050 12414
rect 23998 12338 24050 12350
rect 24558 12402 24610 12414
rect 24558 12338 24610 12350
rect 25454 12402 25506 12414
rect 25454 12338 25506 12350
rect 26238 12402 26290 12414
rect 34302 12402 34354 12414
rect 31378 12350 31390 12402
rect 31442 12350 31454 12402
rect 26238 12338 26290 12350
rect 34302 12338 34354 12350
rect 36094 12402 36146 12414
rect 36094 12338 36146 12350
rect 37998 12402 38050 12414
rect 37998 12338 38050 12350
rect 38110 12402 38162 12414
rect 38110 12338 38162 12350
rect 43374 12402 43426 12414
rect 43374 12338 43426 12350
rect 44942 12402 44994 12414
rect 44942 12338 44994 12350
rect 4846 12290 4898 12302
rect 4846 12226 4898 12238
rect 8654 12290 8706 12302
rect 21982 12290 22034 12302
rect 12674 12238 12686 12290
rect 12738 12238 12750 12290
rect 14578 12238 14590 12290
rect 14642 12238 14654 12290
rect 18610 12238 18622 12290
rect 18674 12238 18686 12290
rect 19618 12238 19630 12290
rect 19682 12238 19694 12290
rect 8654 12226 8706 12238
rect 21982 12226 22034 12238
rect 22206 12290 22258 12302
rect 23886 12290 23938 12302
rect 23426 12238 23438 12290
rect 23490 12238 23502 12290
rect 22206 12226 22258 12238
rect 23886 12226 23938 12238
rect 24670 12290 24722 12302
rect 24670 12226 24722 12238
rect 25230 12290 25282 12302
rect 31278 12290 31330 12302
rect 34190 12290 34242 12302
rect 28242 12238 28254 12290
rect 28306 12238 28318 12290
rect 29026 12238 29038 12290
rect 29090 12238 29102 12290
rect 30482 12238 30494 12290
rect 30546 12238 30558 12290
rect 32274 12238 32286 12290
rect 32338 12238 32350 12290
rect 25230 12226 25282 12238
rect 31278 12226 31330 12238
rect 34190 12226 34242 12238
rect 34862 12290 34914 12302
rect 34862 12226 34914 12238
rect 35870 12290 35922 12302
rect 35870 12226 35922 12238
rect 36990 12290 37042 12302
rect 43710 12290 43762 12302
rect 39106 12238 39118 12290
rect 39170 12238 39182 12290
rect 36990 12226 37042 12238
rect 43710 12226 43762 12238
rect 44270 12290 44322 12302
rect 44270 12226 44322 12238
rect 44382 12290 44434 12302
rect 44382 12226 44434 12238
rect 45054 12290 45106 12302
rect 45054 12226 45106 12238
rect 45278 12290 45330 12302
rect 45278 12226 45330 12238
rect 5854 12178 5906 12190
rect 6414 12178 6466 12190
rect 3826 12126 3838 12178
rect 3890 12126 3902 12178
rect 6178 12126 6190 12178
rect 6242 12126 6254 12178
rect 5854 12114 5906 12126
rect 6414 12114 6466 12126
rect 6638 12178 6690 12190
rect 6638 12114 6690 12126
rect 7198 12178 7250 12190
rect 9774 12178 9826 12190
rect 9538 12126 9550 12178
rect 9602 12126 9614 12178
rect 7198 12114 7250 12126
rect 9774 12114 9826 12126
rect 9998 12178 10050 12190
rect 15038 12178 15090 12190
rect 16046 12178 16098 12190
rect 21534 12178 21586 12190
rect 28478 12178 28530 12190
rect 33966 12178 34018 12190
rect 13010 12126 13022 12178
rect 13074 12126 13086 12178
rect 13682 12126 13694 12178
rect 13746 12126 13758 12178
rect 14018 12126 14030 12178
rect 14082 12126 14094 12178
rect 15810 12126 15822 12178
rect 15874 12126 15886 12178
rect 16482 12126 16494 12178
rect 16546 12126 16558 12178
rect 18162 12126 18174 12178
rect 18226 12126 18238 12178
rect 19730 12126 19742 12178
rect 19794 12126 19806 12178
rect 22866 12126 22878 12178
rect 22930 12126 22942 12178
rect 26450 12126 26462 12178
rect 26514 12126 26526 12178
rect 27234 12126 27246 12178
rect 27298 12126 27310 12178
rect 27458 12126 27470 12178
rect 27522 12126 27534 12178
rect 27906 12126 27918 12178
rect 27970 12126 27982 12178
rect 29474 12126 29486 12178
rect 29538 12126 29550 12178
rect 29922 12126 29934 12178
rect 29986 12126 29998 12178
rect 31042 12126 31054 12178
rect 31106 12126 31118 12178
rect 32498 12126 32510 12178
rect 32562 12126 32574 12178
rect 9998 12114 10050 12126
rect 15038 12114 15090 12126
rect 16046 12114 16098 12126
rect 21534 12114 21586 12126
rect 28478 12114 28530 12126
rect 33966 12114 34018 12126
rect 34414 12178 34466 12190
rect 34414 12114 34466 12126
rect 35422 12178 35474 12190
rect 35422 12114 35474 12126
rect 36206 12178 36258 12190
rect 36206 12114 36258 12126
rect 36430 12178 36482 12190
rect 37214 12178 37266 12190
rect 38222 12178 38274 12190
rect 38782 12178 38834 12190
rect 41134 12178 41186 12190
rect 36754 12126 36766 12178
rect 36818 12126 36830 12178
rect 37426 12126 37438 12178
rect 37490 12126 37502 12178
rect 37762 12126 37774 12178
rect 37826 12126 37838 12178
rect 38434 12126 38446 12178
rect 38498 12126 38510 12178
rect 40898 12126 40910 12178
rect 40962 12126 40974 12178
rect 36430 12114 36482 12126
rect 37214 12114 37266 12126
rect 38222 12114 38274 12126
rect 38782 12114 38834 12126
rect 41134 12114 41186 12126
rect 41358 12178 41410 12190
rect 41358 12114 41410 12126
rect 44718 12178 44770 12190
rect 46050 12126 46062 12178
rect 46114 12126 46126 12178
rect 44718 12114 44770 12126
rect 4286 12066 4338 12078
rect 3938 12014 3950 12066
rect 4002 12014 4014 12066
rect 4286 12002 4338 12014
rect 4622 12066 4674 12078
rect 4622 12002 4674 12014
rect 4734 12066 4786 12078
rect 21758 12066 21810 12078
rect 37102 12066 37154 12078
rect 8978 12014 8990 12066
rect 9042 12014 9054 12066
rect 14354 12014 14366 12066
rect 14418 12014 14430 12066
rect 21186 12014 21198 12066
rect 21250 12014 21262 12066
rect 25554 12014 25566 12066
rect 25618 12014 25630 12066
rect 30146 12014 30158 12066
rect 30210 12014 30222 12066
rect 4734 12002 4786 12014
rect 21758 12002 21810 12014
rect 37102 12002 37154 12014
rect 40350 12066 40402 12078
rect 40350 12002 40402 12014
rect 47966 12066 48018 12078
rect 47966 12002 48018 12014
rect 6750 11954 6802 11966
rect 6750 11890 6802 11902
rect 10110 11954 10162 11966
rect 10110 11890 10162 11902
rect 23326 11954 23378 11966
rect 23326 11890 23378 11902
rect 26126 11954 26178 11966
rect 26126 11890 26178 11902
rect 33742 11954 33794 11966
rect 33742 11890 33794 11902
rect 41470 11954 41522 11966
rect 41470 11890 41522 11902
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 13470 11618 13522 11630
rect 13470 11554 13522 11566
rect 21310 11618 21362 11630
rect 21310 11554 21362 11566
rect 21422 11618 21474 11630
rect 21422 11554 21474 11566
rect 21646 11618 21698 11630
rect 21646 11554 21698 11566
rect 27806 11618 27858 11630
rect 27806 11554 27858 11566
rect 30494 11618 30546 11630
rect 30494 11554 30546 11566
rect 34302 11618 34354 11630
rect 34302 11554 34354 11566
rect 37998 11618 38050 11630
rect 37998 11554 38050 11566
rect 16158 11506 16210 11518
rect 34414 11506 34466 11518
rect 47966 11506 48018 11518
rect 2482 11454 2494 11506
rect 2546 11454 2558 11506
rect 4610 11454 4622 11506
rect 4674 11454 4686 11506
rect 7410 11454 7422 11506
rect 7474 11454 7486 11506
rect 8866 11454 8878 11506
rect 8930 11454 8942 11506
rect 11666 11454 11678 11506
rect 11730 11454 11742 11506
rect 17938 11454 17950 11506
rect 18002 11454 18014 11506
rect 22530 11454 22542 11506
rect 22594 11454 22606 11506
rect 33506 11454 33518 11506
rect 33570 11454 33582 11506
rect 42018 11454 42030 11506
rect 42082 11454 42094 11506
rect 44146 11454 44158 11506
rect 44210 11454 44222 11506
rect 16158 11442 16210 11454
rect 34414 11442 34466 11454
rect 47966 11442 48018 11454
rect 10782 11394 10834 11406
rect 12238 11394 12290 11406
rect 1810 11342 1822 11394
rect 1874 11342 1886 11394
rect 7074 11342 7086 11394
rect 7138 11342 7150 11394
rect 11778 11342 11790 11394
rect 11842 11342 11854 11394
rect 10782 11330 10834 11342
rect 12238 11330 12290 11342
rect 12686 11394 12738 11406
rect 15486 11394 15538 11406
rect 13682 11342 13694 11394
rect 13746 11342 13758 11394
rect 14242 11342 14254 11394
rect 14306 11342 14318 11394
rect 15026 11342 15038 11394
rect 15090 11342 15102 11394
rect 12686 11330 12738 11342
rect 15486 11330 15538 11342
rect 15822 11394 15874 11406
rect 20862 11394 20914 11406
rect 17602 11342 17614 11394
rect 17666 11342 17678 11394
rect 18498 11342 18510 11394
rect 18562 11342 18574 11394
rect 15822 11330 15874 11342
rect 20862 11330 20914 11342
rect 21758 11394 21810 11406
rect 29486 11394 29538 11406
rect 23202 11342 23214 11394
rect 23266 11342 23278 11394
rect 25218 11342 25230 11394
rect 25282 11342 25294 11394
rect 21758 11330 21810 11342
rect 29486 11330 29538 11342
rect 29710 11394 29762 11406
rect 30718 11394 30770 11406
rect 30034 11342 30046 11394
rect 30098 11342 30110 11394
rect 29710 11330 29762 11342
rect 30718 11330 30770 11342
rect 30942 11394 30994 11406
rect 30942 11330 30994 11342
rect 31054 11394 31106 11406
rect 35646 11394 35698 11406
rect 37214 11394 37266 11406
rect 31714 11342 31726 11394
rect 31778 11342 31790 11394
rect 32722 11342 32734 11394
rect 32786 11342 32798 11394
rect 33618 11342 33630 11394
rect 33682 11342 33694 11394
rect 35858 11342 35870 11394
rect 35922 11342 35934 11394
rect 31054 11330 31106 11342
rect 35646 11330 35698 11342
rect 37214 11330 37266 11342
rect 40910 11394 40962 11406
rect 41234 11342 41246 11394
rect 41298 11342 41310 11394
rect 46050 11342 46062 11394
rect 46114 11342 46126 11394
rect 40910 11330 40962 11342
rect 9214 11282 9266 11294
rect 11118 11282 11170 11294
rect 9538 11230 9550 11282
rect 9602 11230 9614 11282
rect 9214 11218 9266 11230
rect 11118 11218 11170 11230
rect 12462 11282 12514 11294
rect 19630 11282 19682 11294
rect 13794 11230 13806 11282
rect 13858 11230 13870 11282
rect 18722 11230 18734 11282
rect 18786 11230 18798 11282
rect 18946 11230 18958 11282
rect 19010 11230 19022 11282
rect 12462 11218 12514 11230
rect 19630 11218 19682 11230
rect 22878 11282 22930 11294
rect 22878 11218 22930 11230
rect 24334 11282 24386 11294
rect 24334 11218 24386 11230
rect 25790 11282 25842 11294
rect 25790 11218 25842 11230
rect 27918 11282 27970 11294
rect 36878 11282 36930 11294
rect 33170 11230 33182 11282
rect 33234 11230 33246 11282
rect 33506 11230 33518 11282
rect 33570 11230 33582 11282
rect 27918 11218 27970 11230
rect 36878 11218 36930 11230
rect 38110 11282 38162 11294
rect 38110 11218 38162 11230
rect 5070 11170 5122 11182
rect 5070 11106 5122 11118
rect 5742 11170 5794 11182
rect 5742 11106 5794 11118
rect 9886 11170 9938 11182
rect 9886 11106 9938 11118
rect 10222 11170 10274 11182
rect 10222 11106 10274 11118
rect 11342 11170 11394 11182
rect 11342 11106 11394 11118
rect 11566 11170 11618 11182
rect 11566 11106 11618 11118
rect 12350 11170 12402 11182
rect 12350 11106 12402 11118
rect 12574 11170 12626 11182
rect 12574 11106 12626 11118
rect 15598 11170 15650 11182
rect 15598 11106 15650 11118
rect 22654 11170 22706 11182
rect 31166 11170 31218 11182
rect 26786 11118 26798 11170
rect 26850 11118 26862 11170
rect 22654 11106 22706 11118
rect 31166 11106 31218 11118
rect 35758 11170 35810 11182
rect 35758 11106 35810 11118
rect 37102 11170 37154 11182
rect 37102 11106 37154 11118
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 11790 10834 11842 10846
rect 11790 10770 11842 10782
rect 14702 10834 14754 10846
rect 16382 10834 16434 10846
rect 15586 10782 15598 10834
rect 15650 10782 15662 10834
rect 14702 10770 14754 10782
rect 16382 10770 16434 10782
rect 17502 10834 17554 10846
rect 17502 10770 17554 10782
rect 19294 10834 19346 10846
rect 19294 10770 19346 10782
rect 29150 10834 29202 10846
rect 29150 10770 29202 10782
rect 30718 10834 30770 10846
rect 30718 10770 30770 10782
rect 32062 10834 32114 10846
rect 32062 10770 32114 10782
rect 36878 10834 36930 10846
rect 39566 10834 39618 10846
rect 38434 10782 38446 10834
rect 38498 10782 38510 10834
rect 36878 10770 36930 10782
rect 39566 10770 39618 10782
rect 11902 10722 11954 10734
rect 14478 10722 14530 10734
rect 18286 10722 18338 10734
rect 4946 10670 4958 10722
rect 5010 10670 5022 10722
rect 12898 10670 12910 10722
rect 12962 10670 12974 10722
rect 15138 10670 15150 10722
rect 15202 10670 15214 10722
rect 23438 10722 23490 10734
rect 11902 10658 11954 10670
rect 14478 10658 14530 10670
rect 18286 10658 18338 10670
rect 19182 10666 19234 10678
rect 14366 10610 14418 10622
rect 17838 10610 17890 10622
rect 4274 10558 4286 10610
rect 4338 10558 4350 10610
rect 15698 10558 15710 10610
rect 15762 10558 15774 10610
rect 16034 10558 16046 10610
rect 16098 10558 16110 10610
rect 23438 10658 23490 10670
rect 23550 10722 23602 10734
rect 28926 10722 28978 10734
rect 36542 10722 36594 10734
rect 27570 10670 27582 10722
rect 27634 10670 27646 10722
rect 32386 10670 32398 10722
rect 32450 10670 32462 10722
rect 34738 10670 34750 10722
rect 34802 10670 34814 10722
rect 23550 10658 23602 10670
rect 28926 10658 28978 10670
rect 36542 10658 36594 10670
rect 43598 10722 43650 10734
rect 43598 10658 43650 10670
rect 43822 10722 43874 10734
rect 43822 10658 43874 10670
rect 47854 10722 47906 10734
rect 47854 10658 47906 10670
rect 48190 10722 48242 10734
rect 48190 10658 48242 10670
rect 19182 10602 19234 10614
rect 23774 10610 23826 10622
rect 14366 10546 14418 10558
rect 17838 10546 17890 10558
rect 23774 10546 23826 10558
rect 26686 10610 26738 10622
rect 28366 10610 28418 10622
rect 26898 10558 26910 10610
rect 26962 10558 26974 10610
rect 27794 10558 27806 10610
rect 27858 10558 27870 10610
rect 26686 10546 26738 10558
rect 28366 10546 28418 10558
rect 28814 10610 28866 10622
rect 34526 10610 34578 10622
rect 36766 10610 36818 10622
rect 30706 10558 30718 10610
rect 30770 10558 30782 10610
rect 35074 10558 35086 10610
rect 35138 10558 35150 10610
rect 35746 10558 35758 10610
rect 35810 10558 35822 10610
rect 28814 10546 28866 10558
rect 34526 10546 34578 10558
rect 36766 10546 36818 10558
rect 36990 10610 37042 10622
rect 37774 10610 37826 10622
rect 37202 10558 37214 10610
rect 37266 10558 37278 10610
rect 36990 10546 37042 10558
rect 37774 10546 37826 10558
rect 37886 10610 37938 10622
rect 37886 10546 37938 10558
rect 37998 10610 38050 10622
rect 37998 10546 38050 10558
rect 38782 10610 38834 10622
rect 38782 10546 38834 10558
rect 39118 10610 39170 10622
rect 39118 10546 39170 10558
rect 39230 10610 39282 10622
rect 44270 10610 44322 10622
rect 39330 10558 39342 10610
rect 39394 10558 39406 10610
rect 44482 10558 44494 10610
rect 44546 10558 44558 10610
rect 45266 10558 45278 10610
rect 45330 10558 45342 10610
rect 39230 10546 39282 10558
rect 44270 10546 44322 10558
rect 7534 10498 7586 10510
rect 7074 10446 7086 10498
rect 7138 10446 7150 10498
rect 7534 10434 7586 10446
rect 12574 10498 12626 10510
rect 12574 10434 12626 10446
rect 18846 10498 18898 10510
rect 18846 10434 18898 10446
rect 44046 10498 44098 10510
rect 47394 10446 47406 10498
rect 47458 10446 47470 10498
rect 44046 10434 44098 10446
rect 17950 10386 18002 10398
rect 17950 10322 18002 10334
rect 19294 10386 19346 10398
rect 35634 10334 35646 10386
rect 35698 10334 35710 10386
rect 19294 10322 19346 10334
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 44830 10050 44882 10062
rect 44830 9986 44882 9998
rect 27358 9938 27410 9950
rect 7970 9886 7982 9938
rect 8034 9886 8046 9938
rect 10098 9886 10110 9938
rect 10162 9886 10174 9938
rect 11890 9886 11902 9938
rect 11954 9886 11966 9938
rect 14354 9886 14366 9938
rect 14418 9886 14430 9938
rect 14914 9886 14926 9938
rect 14978 9886 14990 9938
rect 17826 9886 17838 9938
rect 17890 9886 17902 9938
rect 21634 9886 21646 9938
rect 21698 9886 21710 9938
rect 27358 9874 27410 9886
rect 28254 9938 28306 9950
rect 34414 9938 34466 9950
rect 43598 9938 43650 9950
rect 29922 9886 29934 9938
rect 29986 9886 29998 9938
rect 33618 9886 33630 9938
rect 33682 9886 33694 9938
rect 35522 9886 35534 9938
rect 35586 9886 35598 9938
rect 39218 9886 39230 9938
rect 39282 9886 39294 9938
rect 41346 9886 41358 9938
rect 41410 9886 41422 9938
rect 28254 9874 28306 9886
rect 34414 9874 34466 9886
rect 43598 9874 43650 9886
rect 44942 9938 44994 9950
rect 44942 9874 44994 9886
rect 47966 9938 48018 9950
rect 47966 9874 48018 9886
rect 12350 9826 12402 9838
rect 7298 9774 7310 9826
rect 7362 9774 7374 9826
rect 11554 9774 11566 9826
rect 11618 9774 11630 9826
rect 12350 9762 12402 9774
rect 12910 9826 12962 9838
rect 12910 9762 12962 9774
rect 13918 9826 13970 9838
rect 15038 9826 15090 9838
rect 27918 9826 27970 9838
rect 30942 9826 30994 9838
rect 33070 9826 33122 9838
rect 35310 9826 35362 9838
rect 38222 9826 38274 9838
rect 14466 9774 14478 9826
rect 14530 9774 14542 9826
rect 16370 9774 16382 9826
rect 16434 9774 16446 9826
rect 17266 9774 17278 9826
rect 17330 9774 17342 9826
rect 20626 9774 20638 9826
rect 20690 9774 20702 9826
rect 21970 9774 21982 9826
rect 22034 9774 22046 9826
rect 23202 9774 23214 9826
rect 23266 9774 23278 9826
rect 25218 9774 25230 9826
rect 25282 9774 25294 9826
rect 29586 9774 29598 9826
rect 29650 9774 29662 9826
rect 31826 9774 31838 9826
rect 31890 9774 31902 9826
rect 34178 9774 34190 9826
rect 34242 9774 34254 9826
rect 34514 9774 34526 9826
rect 34578 9774 34590 9826
rect 35746 9774 35758 9826
rect 35810 9774 35822 9826
rect 42018 9774 42030 9826
rect 42082 9774 42094 9826
rect 43138 9774 43150 9826
rect 43202 9774 43214 9826
rect 45602 9774 45614 9826
rect 45666 9774 45678 9826
rect 13918 9762 13970 9774
rect 15038 9762 15090 9774
rect 27918 9762 27970 9774
rect 30942 9762 30994 9774
rect 33070 9762 33122 9774
rect 35310 9762 35362 9774
rect 38222 9762 38274 9774
rect 14926 9714 14978 9726
rect 14926 9650 14978 9662
rect 15486 9714 15538 9726
rect 22430 9714 22482 9726
rect 17154 9662 17166 9714
rect 17218 9662 17230 9714
rect 19954 9662 19966 9714
rect 20018 9662 20030 9714
rect 15486 9650 15538 9662
rect 22430 9650 22482 9662
rect 24334 9714 24386 9726
rect 24334 9650 24386 9662
rect 25790 9714 25842 9726
rect 25790 9650 25842 9662
rect 28366 9714 28418 9726
rect 28366 9650 28418 9662
rect 30270 9714 30322 9726
rect 30270 9650 30322 9662
rect 31054 9714 31106 9726
rect 31054 9650 31106 9662
rect 32286 9714 32338 9726
rect 32286 9650 32338 9662
rect 32398 9714 32450 9726
rect 32398 9650 32450 9662
rect 32622 9714 32674 9726
rect 32622 9650 32674 9662
rect 32958 9714 33010 9726
rect 32958 9650 33010 9662
rect 33182 9714 33234 9726
rect 33182 9650 33234 9662
rect 33966 9714 34018 9726
rect 33966 9650 34018 9662
rect 35086 9714 35138 9726
rect 35086 9650 35138 9662
rect 35534 9714 35586 9726
rect 37886 9714 37938 9726
rect 37314 9662 37326 9714
rect 37378 9662 37390 9714
rect 35534 9650 35586 9662
rect 37886 9650 37938 9662
rect 37998 9714 38050 9726
rect 37998 9650 38050 9662
rect 10558 9602 10610 9614
rect 10558 9538 10610 9550
rect 14030 9602 14082 9614
rect 14030 9538 14082 9550
rect 14254 9602 14306 9614
rect 14254 9538 14306 9550
rect 15262 9602 15314 9614
rect 34750 9602 34802 9614
rect 15922 9550 15934 9602
rect 15986 9550 15998 9602
rect 16146 9550 16158 9602
rect 16210 9550 16222 9602
rect 26786 9550 26798 9602
rect 26850 9550 26862 9602
rect 31602 9550 31614 9602
rect 31666 9550 31678 9602
rect 15262 9538 15314 9550
rect 34750 9538 34802 9550
rect 36990 9602 37042 9614
rect 36990 9538 37042 9550
rect 38558 9602 38610 9614
rect 38558 9538 38610 9550
rect 42590 9602 42642 9614
rect 42590 9538 42642 9550
rect 44158 9602 44210 9614
rect 44158 9538 44210 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 7198 9266 7250 9278
rect 7198 9202 7250 9214
rect 12910 9266 12962 9278
rect 12910 9202 12962 9214
rect 14366 9266 14418 9278
rect 14366 9202 14418 9214
rect 15374 9266 15426 9278
rect 15374 9202 15426 9214
rect 19742 9266 19794 9278
rect 19742 9202 19794 9214
rect 24670 9266 24722 9278
rect 24670 9202 24722 9214
rect 27022 9266 27074 9278
rect 27022 9202 27074 9214
rect 27582 9266 27634 9278
rect 29486 9266 29538 9278
rect 28242 9214 28254 9266
rect 28306 9214 28318 9266
rect 27582 9202 27634 9214
rect 29486 9202 29538 9214
rect 34862 9266 34914 9278
rect 36990 9266 37042 9278
rect 35186 9214 35198 9266
rect 35250 9214 35262 9266
rect 34862 9202 34914 9214
rect 36990 9202 37042 9214
rect 41358 9266 41410 9278
rect 41358 9202 41410 9214
rect 47630 9266 47682 9278
rect 47630 9202 47682 9214
rect 14814 9154 14866 9166
rect 7522 9102 7534 9154
rect 7586 9102 7598 9154
rect 14814 9090 14866 9102
rect 18958 9154 19010 9166
rect 23886 9154 23938 9166
rect 26462 9154 26514 9166
rect 30158 9154 30210 9166
rect 19170 9102 19182 9154
rect 19234 9102 19246 9154
rect 24098 9102 24110 9154
rect 24162 9102 24174 9154
rect 28690 9102 28702 9154
rect 28754 9102 28766 9154
rect 18958 9090 19010 9102
rect 23886 9090 23938 9102
rect 26462 9090 26514 9102
rect 30158 9090 30210 9102
rect 33182 9154 33234 9166
rect 33182 9090 33234 9102
rect 47854 9154 47906 9166
rect 47854 9090 47906 9102
rect 14254 9042 14306 9054
rect 9650 8990 9662 9042
rect 9714 8990 9726 9042
rect 14254 8978 14306 8990
rect 14590 9042 14642 9054
rect 14590 8978 14642 8990
rect 15822 9042 15874 9054
rect 15822 8978 15874 8990
rect 15934 9042 15986 9054
rect 18286 9042 18338 9054
rect 17826 8990 17838 9042
rect 17890 8990 17902 9042
rect 15934 8978 15986 8990
rect 18286 8978 18338 8990
rect 19406 9042 19458 9054
rect 24334 9042 24386 9054
rect 48190 9042 48242 9054
rect 19506 8990 19518 9042
rect 19570 8990 19582 9042
rect 24658 8990 24670 9042
rect 24722 8990 24734 9042
rect 27570 8990 27582 9042
rect 27634 8990 27646 9042
rect 28466 8990 28478 9042
rect 28530 8990 28542 9042
rect 29810 8990 29822 9042
rect 29874 8990 29886 9042
rect 37650 8990 37662 9042
rect 37714 8990 37726 9042
rect 41682 8990 41694 9042
rect 41746 8990 41758 9042
rect 19406 8978 19458 8990
rect 24334 8978 24386 8990
rect 48190 8978 48242 8990
rect 15486 8930 15538 8942
rect 10322 8878 10334 8930
rect 10386 8878 10398 8930
rect 12450 8878 12462 8930
rect 12514 8878 12526 8930
rect 15486 8866 15538 8878
rect 17390 8930 17442 8942
rect 17390 8866 17442 8878
rect 20190 8930 20242 8942
rect 20190 8866 20242 8878
rect 23550 8930 23602 8942
rect 33070 8930 33122 8942
rect 29922 8878 29934 8930
rect 29986 8878 29998 8930
rect 23550 8866 23602 8878
rect 33070 8866 33122 8878
rect 33630 8930 33682 8942
rect 33630 8866 33682 8878
rect 36878 8930 36930 8942
rect 38334 8930 38386 8942
rect 37874 8878 37886 8930
rect 37938 8878 37950 8930
rect 42466 8878 42478 8930
rect 42530 8878 42542 8930
rect 44594 8878 44606 8930
rect 44658 8878 44670 8930
rect 36878 8866 36930 8878
rect 38334 8866 38386 8878
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 17726 8482 17778 8494
rect 17726 8418 17778 8430
rect 21870 8482 21922 8494
rect 21870 8418 21922 8430
rect 9998 8370 10050 8382
rect 9998 8306 10050 8318
rect 13582 8370 13634 8382
rect 13582 8306 13634 8318
rect 18174 8370 18226 8382
rect 22318 8370 22370 8382
rect 32510 8370 32562 8382
rect 41582 8370 41634 8382
rect 21522 8318 21534 8370
rect 21586 8318 21598 8370
rect 24882 8318 24894 8370
rect 24946 8318 24958 8370
rect 27010 8318 27022 8370
rect 27074 8318 27086 8370
rect 27906 8318 27918 8370
rect 27970 8318 27982 8370
rect 29922 8318 29934 8370
rect 29986 8318 29998 8370
rect 32050 8318 32062 8370
rect 32114 8318 32126 8370
rect 32834 8318 32846 8370
rect 32898 8318 32910 8370
rect 34962 8318 34974 8370
rect 35026 8318 35038 8370
rect 38210 8318 38222 8370
rect 38274 8318 38286 8370
rect 18174 8306 18226 8318
rect 22318 8306 22370 8318
rect 32510 8306 32562 8318
rect 41582 8306 41634 8318
rect 42030 8370 42082 8382
rect 42030 8306 42082 8318
rect 42590 8370 42642 8382
rect 42590 8306 42642 8318
rect 48302 8370 48354 8382
rect 48302 8306 48354 8318
rect 6974 8258 7026 8270
rect 6974 8194 7026 8206
rect 7198 8258 7250 8270
rect 7198 8194 7250 8206
rect 7646 8258 7698 8270
rect 7646 8194 7698 8206
rect 7870 8258 7922 8270
rect 7870 8194 7922 8206
rect 8318 8258 8370 8270
rect 8318 8194 8370 8206
rect 9550 8258 9602 8270
rect 9550 8194 9602 8206
rect 9774 8258 9826 8270
rect 9774 8194 9826 8206
rect 10222 8258 10274 8270
rect 10222 8194 10274 8206
rect 11454 8258 11506 8270
rect 42142 8258 42194 8270
rect 24210 8206 24222 8258
rect 24274 8206 24286 8258
rect 27682 8206 27694 8258
rect 27746 8206 27758 8258
rect 29138 8206 29150 8258
rect 29202 8206 29214 8258
rect 35746 8206 35758 8258
rect 35810 8206 35822 8258
rect 41122 8206 41134 8258
rect 41186 8206 41198 8258
rect 11454 8194 11506 8206
rect 42142 8194 42194 8206
rect 42366 8258 42418 8270
rect 42366 8194 42418 8206
rect 42814 8258 42866 8270
rect 42814 8194 42866 8206
rect 43262 8258 43314 8270
rect 43262 8194 43314 8206
rect 43934 8258 43986 8270
rect 45838 8258 45890 8270
rect 45378 8206 45390 8258
rect 45442 8206 45454 8258
rect 43934 8194 43986 8206
rect 45838 8194 45890 8206
rect 46622 8258 46674 8270
rect 46622 8194 46674 8206
rect 47070 8258 47122 8270
rect 47070 8194 47122 8206
rect 1710 8146 1762 8158
rect 1710 8082 1762 8094
rect 2046 8146 2098 8158
rect 2046 8082 2098 8094
rect 6862 8146 6914 8158
rect 6862 8082 6914 8094
rect 9438 8146 9490 8158
rect 9438 8082 9490 8094
rect 10446 8146 10498 8158
rect 10446 8082 10498 8094
rect 17502 8146 17554 8158
rect 17502 8082 17554 8094
rect 21646 8146 21698 8158
rect 43038 8146 43090 8158
rect 40338 8094 40350 8146
rect 40402 8094 40414 8146
rect 21646 8082 21698 8094
rect 43038 8082 43090 8094
rect 43822 8146 43874 8158
rect 45154 8094 45166 8146
rect 45218 8094 45230 8146
rect 46162 8094 46174 8146
rect 46226 8094 46238 8146
rect 43822 8082 43874 8094
rect 2494 8034 2546 8046
rect 2494 7970 2546 7982
rect 7422 8034 7474 8046
rect 7422 7970 7474 7982
rect 8206 8034 8258 8046
rect 8206 7970 8258 7982
rect 8430 8034 8482 8046
rect 8430 7970 8482 7982
rect 8654 8034 8706 8046
rect 8654 7970 8706 7982
rect 10782 8034 10834 8046
rect 10782 7970 10834 7982
rect 10894 8034 10946 8046
rect 10894 7970 10946 7982
rect 11006 8034 11058 8046
rect 11006 7970 11058 7982
rect 17614 8034 17666 8046
rect 17614 7970 17666 7982
rect 36206 8034 36258 8046
rect 36206 7970 36258 7982
rect 43710 8034 43762 8046
rect 43710 7970 43762 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 7422 7698 7474 7710
rect 8654 7698 8706 7710
rect 3938 7646 3950 7698
rect 4002 7646 4014 7698
rect 8306 7646 8318 7698
rect 8370 7646 8382 7698
rect 7422 7634 7474 7646
rect 8654 7634 8706 7646
rect 11902 7698 11954 7710
rect 11902 7634 11954 7646
rect 12350 7698 12402 7710
rect 12350 7634 12402 7646
rect 13582 7698 13634 7710
rect 13582 7634 13634 7646
rect 13806 7698 13858 7710
rect 16382 7698 16434 7710
rect 15138 7646 15150 7698
rect 15202 7646 15214 7698
rect 13806 7634 13858 7646
rect 16382 7634 16434 7646
rect 33406 7698 33458 7710
rect 33406 7634 33458 7646
rect 37438 7698 37490 7710
rect 37438 7634 37490 7646
rect 38894 7698 38946 7710
rect 38894 7634 38946 7646
rect 42926 7698 42978 7710
rect 42926 7634 42978 7646
rect 10670 7586 10722 7598
rect 6178 7534 6190 7586
rect 6242 7534 6254 7586
rect 10670 7522 10722 7534
rect 13022 7586 13074 7598
rect 13022 7522 13074 7534
rect 14030 7586 14082 7598
rect 38670 7586 38722 7598
rect 19506 7534 19518 7586
rect 19570 7534 19582 7586
rect 21410 7534 21422 7586
rect 21474 7534 21486 7586
rect 28466 7534 28478 7586
rect 28530 7534 28542 7586
rect 34178 7534 34190 7586
rect 34242 7534 34254 7586
rect 14030 7522 14082 7534
rect 38670 7522 38722 7534
rect 43150 7586 43202 7598
rect 43586 7534 43598 7586
rect 43650 7534 43662 7586
rect 43150 7522 43202 7534
rect 10334 7474 10386 7486
rect 6962 7422 6974 7474
rect 7026 7422 7038 7474
rect 10334 7410 10386 7422
rect 12686 7474 12738 7486
rect 12686 7410 12738 7422
rect 13134 7474 13186 7486
rect 13134 7410 13186 7422
rect 13694 7474 13746 7486
rect 13694 7410 13746 7422
rect 15486 7474 15538 7486
rect 24670 7474 24722 7486
rect 26126 7474 26178 7486
rect 20290 7422 20302 7474
rect 20354 7422 20366 7474
rect 20626 7422 20638 7474
rect 20690 7422 20702 7474
rect 25666 7422 25678 7474
rect 25730 7422 25742 7474
rect 15486 7410 15538 7422
rect 24670 7410 24722 7422
rect 26126 7410 26178 7422
rect 28030 7474 28082 7486
rect 33854 7474 33906 7486
rect 28690 7422 28702 7474
rect 28754 7422 28766 7474
rect 28030 7410 28082 7422
rect 33854 7410 33906 7422
rect 37550 7474 37602 7486
rect 37550 7410 37602 7422
rect 42702 7474 42754 7486
rect 42702 7410 42754 7422
rect 43934 7474 43986 7486
rect 43934 7410 43986 7422
rect 12238 7362 12290 7374
rect 12238 7298 12290 7310
rect 12798 7362 12850 7374
rect 24110 7362 24162 7374
rect 32510 7362 32562 7374
rect 15922 7310 15934 7362
rect 15986 7310 15998 7362
rect 17378 7310 17390 7362
rect 17442 7310 17454 7362
rect 23538 7310 23550 7362
rect 23602 7310 23614 7362
rect 27570 7310 27582 7362
rect 27634 7310 27646 7362
rect 12798 7298 12850 7310
rect 24110 7298 24162 7310
rect 32510 7298 32562 7310
rect 33518 7362 33570 7374
rect 33518 7298 33570 7310
rect 38446 7362 38498 7374
rect 42814 7362 42866 7374
rect 38994 7310 39006 7362
rect 39058 7310 39070 7362
rect 38446 7298 38498 7310
rect 42814 7298 42866 7310
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 19406 6914 19458 6926
rect 19406 6850 19458 6862
rect 26238 6802 26290 6814
rect 16370 6750 16382 6802
rect 16434 6750 16446 6802
rect 25778 6750 25790 6802
rect 25842 6750 25854 6802
rect 26238 6738 26290 6750
rect 32062 6802 32114 6814
rect 32062 6738 32114 6750
rect 35982 6802 36034 6814
rect 35982 6738 36034 6750
rect 6862 6690 6914 6702
rect 6862 6626 6914 6638
rect 7086 6690 7138 6702
rect 7086 6626 7138 6638
rect 8318 6690 8370 6702
rect 9886 6690 9938 6702
rect 8642 6638 8654 6690
rect 8706 6638 8718 6690
rect 8318 6626 8370 6638
rect 9886 6626 9938 6638
rect 10446 6690 10498 6702
rect 12910 6690 12962 6702
rect 17502 6690 17554 6702
rect 10882 6638 10894 6690
rect 10946 6638 10958 6690
rect 13570 6638 13582 6690
rect 13634 6638 13646 6690
rect 16818 6638 16830 6690
rect 16882 6638 16894 6690
rect 10446 6626 10498 6638
rect 12910 6626 12962 6638
rect 17502 6626 17554 6638
rect 18958 6690 19010 6702
rect 18958 6626 19010 6638
rect 19630 6690 19682 6702
rect 19630 6626 19682 6638
rect 19854 6690 19906 6702
rect 26126 6690 26178 6702
rect 22866 6638 22878 6690
rect 22930 6638 22942 6690
rect 19854 6626 19906 6638
rect 26126 6626 26178 6638
rect 26798 6690 26850 6702
rect 26798 6626 26850 6638
rect 27358 6690 27410 6702
rect 27358 6626 27410 6638
rect 28030 6690 28082 6702
rect 28030 6626 28082 6638
rect 29150 6690 29202 6702
rect 29150 6626 29202 6638
rect 29262 6690 29314 6702
rect 29262 6626 29314 6638
rect 30718 6690 30770 6702
rect 30718 6626 30770 6638
rect 31390 6690 31442 6702
rect 31390 6626 31442 6638
rect 32734 6690 32786 6702
rect 32734 6626 32786 6638
rect 34302 6690 34354 6702
rect 34302 6626 34354 6638
rect 36094 6690 36146 6702
rect 36094 6626 36146 6638
rect 36542 6690 36594 6702
rect 36542 6626 36594 6638
rect 41582 6690 41634 6702
rect 41582 6626 41634 6638
rect 41806 6690 41858 6702
rect 41806 6626 41858 6638
rect 42142 6690 42194 6702
rect 42142 6626 42194 6638
rect 42478 6690 42530 6702
rect 45602 6638 45614 6690
rect 45666 6638 45678 6690
rect 42478 6626 42530 6638
rect 6750 6578 6802 6590
rect 6750 6514 6802 6526
rect 7534 6578 7586 6590
rect 7534 6514 7586 6526
rect 7758 6578 7810 6590
rect 7758 6514 7810 6526
rect 8206 6578 8258 6590
rect 29598 6578 29650 6590
rect 33854 6578 33906 6590
rect 11442 6526 11454 6578
rect 11506 6526 11518 6578
rect 14242 6526 14254 6578
rect 14306 6526 14318 6578
rect 17042 6526 17054 6578
rect 17106 6526 17118 6578
rect 23650 6526 23662 6578
rect 23714 6526 23726 6578
rect 30146 6526 30158 6578
rect 30210 6526 30222 6578
rect 8206 6514 8258 6526
rect 29598 6514 29650 6526
rect 33854 6514 33906 6526
rect 35534 6578 35586 6590
rect 41470 6578 41522 6590
rect 37538 6526 37550 6578
rect 37602 6526 37614 6578
rect 47282 6526 47294 6578
rect 47346 6526 47358 6578
rect 35534 6514 35586 6526
rect 41470 6514 41522 6526
rect 7310 6466 7362 6478
rect 7310 6402 7362 6414
rect 8094 6466 8146 6478
rect 8094 6402 8146 6414
rect 9102 6466 9154 6478
rect 11790 6466 11842 6478
rect 11106 6414 11118 6466
rect 11170 6414 11182 6466
rect 9102 6402 9154 6414
rect 11790 6402 11842 6414
rect 12238 6466 12290 6478
rect 12238 6402 12290 6414
rect 20414 6466 20466 6478
rect 21646 6466 21698 6478
rect 21298 6414 21310 6466
rect 21362 6414 21374 6466
rect 20414 6402 20466 6414
rect 21646 6402 21698 6414
rect 26350 6466 26402 6478
rect 26350 6402 26402 6414
rect 27806 6466 27858 6478
rect 27806 6402 27858 6414
rect 27918 6466 27970 6478
rect 27918 6402 27970 6414
rect 28478 6466 28530 6478
rect 28478 6402 28530 6414
rect 29374 6466 29426 6478
rect 29374 6402 29426 6414
rect 30494 6466 30546 6478
rect 30494 6402 30546 6414
rect 31166 6466 31218 6478
rect 31166 6402 31218 6414
rect 31278 6466 31330 6478
rect 31278 6402 31330 6414
rect 33294 6466 33346 6478
rect 33294 6402 33346 6414
rect 34078 6466 34130 6478
rect 34078 6402 34130 6414
rect 34190 6466 34242 6478
rect 34190 6402 34242 6414
rect 34750 6466 34802 6478
rect 34750 6402 34802 6414
rect 35422 6466 35474 6478
rect 35422 6402 35474 6414
rect 35870 6466 35922 6478
rect 35870 6402 35922 6414
rect 37886 6466 37938 6478
rect 37886 6402 37938 6414
rect 42030 6466 42082 6478
rect 42030 6402 42082 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 8094 6130 8146 6142
rect 8094 6066 8146 6078
rect 8430 6130 8482 6142
rect 8430 6066 8482 6078
rect 9774 6130 9826 6142
rect 9774 6066 9826 6078
rect 10670 6130 10722 6142
rect 10670 6066 10722 6078
rect 20750 6130 20802 6142
rect 20750 6066 20802 6078
rect 23886 6130 23938 6142
rect 29262 6130 29314 6142
rect 28130 6078 28142 6130
rect 28194 6078 28206 6130
rect 23886 6066 23938 6078
rect 29262 6066 29314 6078
rect 31166 6130 31218 6142
rect 31166 6066 31218 6078
rect 33294 6130 33346 6142
rect 33294 6066 33346 6078
rect 38894 6130 38946 6142
rect 38894 6066 38946 6078
rect 40350 6130 40402 6142
rect 40350 6066 40402 6078
rect 9550 6018 9602 6030
rect 24334 6018 24386 6030
rect 27134 6018 27186 6030
rect 6514 5966 6526 6018
rect 6578 5966 6590 6018
rect 18162 5966 18174 6018
rect 18226 5966 18238 6018
rect 20290 5966 20302 6018
rect 20354 5966 20366 6018
rect 26786 5966 26798 6018
rect 26850 5966 26862 6018
rect 9550 5954 9602 5966
rect 24334 5954 24386 5966
rect 27134 5954 27186 5966
rect 29934 6018 29986 6030
rect 29934 5954 29986 5966
rect 34190 6018 34242 6030
rect 34190 5954 34242 5966
rect 34974 6018 35026 6030
rect 34974 5954 35026 5966
rect 35198 6018 35250 6030
rect 41682 5966 41694 6018
rect 41746 5966 41758 6018
rect 35198 5954 35250 5966
rect 19406 5906 19458 5918
rect 23438 5906 23490 5918
rect 7186 5854 7198 5906
rect 7250 5854 7262 5906
rect 10098 5854 10110 5906
rect 10162 5854 10174 5906
rect 10994 5854 11006 5906
rect 11058 5854 11070 5906
rect 20066 5854 20078 5906
rect 20130 5854 20142 5906
rect 19406 5842 19458 5854
rect 23438 5842 23490 5854
rect 23662 5906 23714 5918
rect 23662 5842 23714 5854
rect 24110 5906 24162 5918
rect 27470 5906 27522 5918
rect 26562 5854 26574 5906
rect 26626 5854 26638 5906
rect 24110 5842 24162 5854
rect 27470 5842 27522 5854
rect 27806 5906 27858 5918
rect 27806 5842 27858 5854
rect 30830 5906 30882 5918
rect 30830 5842 30882 5854
rect 31278 5906 31330 5918
rect 31278 5842 31330 5854
rect 31390 5906 31442 5918
rect 31390 5842 31442 5854
rect 33518 5906 33570 5918
rect 33518 5842 33570 5854
rect 33966 5906 34018 5918
rect 33966 5842 34018 5854
rect 34638 5906 34690 5918
rect 35634 5854 35646 5906
rect 35698 5854 35710 5906
rect 41010 5854 41022 5906
rect 41074 5854 41086 5906
rect 34638 5842 34690 5854
rect 9662 5794 9714 5806
rect 4386 5742 4398 5794
rect 4450 5742 4462 5794
rect 9662 5730 9714 5742
rect 18510 5794 18562 5806
rect 23326 5794 23378 5806
rect 18946 5742 18958 5794
rect 19010 5742 19022 5794
rect 18510 5730 18562 5742
rect 23326 5730 23378 5742
rect 25230 5794 25282 5806
rect 25230 5730 25282 5742
rect 25902 5794 25954 5806
rect 25902 5730 25954 5742
rect 28702 5794 28754 5806
rect 28702 5730 28754 5742
rect 31950 5794 32002 5806
rect 31950 5730 32002 5742
rect 32398 5794 32450 5806
rect 32398 5730 32450 5742
rect 33742 5794 33794 5806
rect 33742 5730 33794 5742
rect 34750 5794 34802 5806
rect 36306 5742 36318 5794
rect 36370 5742 36382 5794
rect 38434 5742 38446 5794
rect 38498 5742 38510 5794
rect 43810 5742 43822 5794
rect 43874 5742 43886 5794
rect 34750 5730 34802 5742
rect 12014 5682 12066 5694
rect 12014 5618 12066 5630
rect 25342 5682 25394 5694
rect 25342 5618 25394 5630
rect 28814 5682 28866 5694
rect 28814 5618 28866 5630
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 30270 5346 30322 5358
rect 30270 5282 30322 5294
rect 22318 5234 22370 5246
rect 25454 5234 25506 5246
rect 34862 5234 34914 5246
rect 10322 5182 10334 5234
rect 10386 5182 10398 5234
rect 15810 5182 15822 5234
rect 15874 5182 15886 5234
rect 16258 5182 16270 5234
rect 16322 5182 16334 5234
rect 23650 5182 23662 5234
rect 23714 5182 23726 5234
rect 31378 5182 31390 5234
rect 31442 5182 31454 5234
rect 33506 5182 33518 5234
rect 33570 5182 33582 5234
rect 22318 5170 22370 5182
rect 25454 5170 25506 5182
rect 34862 5170 34914 5182
rect 11118 5122 11170 5134
rect 7298 5070 7310 5122
rect 7362 5070 7374 5122
rect 11118 5058 11170 5070
rect 11454 5122 11506 5134
rect 11454 5058 11506 5070
rect 12462 5122 12514 5134
rect 12462 5058 12514 5070
rect 13022 5122 13074 5134
rect 19630 5122 19682 5134
rect 15586 5070 15598 5122
rect 15650 5070 15662 5122
rect 19170 5070 19182 5122
rect 19234 5070 19246 5122
rect 13022 5058 13074 5070
rect 19630 5058 19682 5070
rect 20190 5122 20242 5134
rect 20190 5058 20242 5070
rect 20302 5122 20354 5134
rect 20302 5058 20354 5070
rect 21758 5122 21810 5134
rect 21758 5058 21810 5070
rect 24110 5122 24162 5134
rect 27246 5122 27298 5134
rect 24546 5070 24558 5122
rect 24610 5070 24622 5122
rect 24110 5058 24162 5070
rect 27246 5058 27298 5070
rect 27694 5122 27746 5134
rect 27694 5058 27746 5070
rect 27918 5122 27970 5134
rect 29038 5122 29090 5134
rect 28466 5070 28478 5122
rect 28530 5070 28542 5122
rect 27918 5058 27970 5070
rect 29038 5058 29090 5070
rect 29374 5122 29426 5134
rect 29374 5058 29426 5070
rect 29598 5122 29650 5134
rect 30706 5070 30718 5122
rect 30770 5070 30782 5122
rect 33842 5070 33854 5122
rect 33906 5070 33918 5122
rect 29598 5058 29650 5070
rect 6862 5010 6914 5022
rect 12574 5010 12626 5022
rect 20414 5010 20466 5022
rect 8082 4958 8094 5010
rect 8146 4958 8158 5010
rect 11778 4958 11790 5010
rect 11842 4958 11854 5010
rect 18386 4958 18398 5010
rect 18450 4958 18462 5010
rect 6862 4946 6914 4958
rect 12574 4946 12626 4958
rect 20414 4946 20466 4958
rect 20638 5010 20690 5022
rect 20638 4946 20690 4958
rect 21422 5010 21474 5022
rect 21422 4946 21474 4958
rect 30158 5010 30210 5022
rect 30158 4946 30210 4958
rect 6974 4898 7026 4910
rect 12350 4898 12402 4910
rect 10770 4846 10782 4898
rect 10834 4846 10846 4898
rect 6974 4834 7026 4846
rect 12350 4834 12402 4846
rect 13694 4898 13746 4910
rect 13694 4834 13746 4846
rect 14814 4898 14866 4910
rect 19518 4898 19570 4910
rect 15138 4846 15150 4898
rect 15202 4846 15214 4898
rect 14814 4834 14866 4846
rect 19518 4834 19570 4846
rect 21310 4898 21362 4910
rect 21310 4834 21362 4846
rect 22206 4898 22258 4910
rect 22206 4834 22258 4846
rect 22430 4898 22482 4910
rect 22430 4834 22482 4846
rect 23326 4898 23378 4910
rect 23326 4834 23378 4846
rect 27582 4898 27634 4910
rect 27582 4834 27634 4846
rect 28254 4898 28306 4910
rect 28254 4834 28306 4846
rect 29374 4898 29426 4910
rect 29374 4834 29426 4846
rect 37214 4898 37266 4910
rect 37214 4834 37266 4846
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 8094 4562 8146 4574
rect 8094 4498 8146 4510
rect 10334 4562 10386 4574
rect 10334 4498 10386 4510
rect 14926 4562 14978 4574
rect 14926 4498 14978 4510
rect 19182 4562 19234 4574
rect 19182 4498 19234 4510
rect 19630 4562 19682 4574
rect 19630 4498 19682 4510
rect 32174 4562 32226 4574
rect 32174 4498 32226 4510
rect 33406 4562 33458 4574
rect 33406 4498 33458 4510
rect 37214 4562 37266 4574
rect 37214 4498 37266 4510
rect 8542 4450 8594 4462
rect 8542 4386 8594 4398
rect 9102 4450 9154 4462
rect 9102 4386 9154 4398
rect 9998 4450 10050 4462
rect 9998 4386 10050 4398
rect 11006 4450 11058 4462
rect 11006 4386 11058 4398
rect 11230 4450 11282 4462
rect 11230 4386 11282 4398
rect 19518 4450 19570 4462
rect 19518 4386 19570 4398
rect 19854 4450 19906 4462
rect 19854 4386 19906 4398
rect 20078 4450 20130 4462
rect 20078 4386 20130 4398
rect 20638 4450 20690 4462
rect 41246 4450 41298 4462
rect 27570 4398 27582 4450
rect 27634 4398 27646 4450
rect 29474 4398 29486 4450
rect 29538 4398 29550 4450
rect 34514 4398 34526 4450
rect 34578 4398 34590 4450
rect 20638 4386 20690 4398
rect 41246 4386 41298 4398
rect 7870 4338 7922 4350
rect 7870 4274 7922 4286
rect 8206 4338 8258 4350
rect 8206 4274 8258 4286
rect 9662 4338 9714 4350
rect 9662 4274 9714 4286
rect 10558 4338 10610 4350
rect 18846 4338 18898 4350
rect 11554 4286 11566 4338
rect 11618 4286 11630 4338
rect 10558 4274 10610 4286
rect 18846 4274 18898 4286
rect 20526 4338 20578 4350
rect 20526 4274 20578 4286
rect 21086 4338 21138 4350
rect 21410 4286 21422 4338
rect 21474 4286 21486 4338
rect 28354 4286 28366 4338
rect 28418 4286 28430 4338
rect 28802 4286 28814 4338
rect 28866 4286 28878 4338
rect 32386 4286 32398 4338
rect 32450 4286 32462 4338
rect 33730 4286 33742 4338
rect 33794 4286 33806 4338
rect 37426 4286 37438 4338
rect 37490 4286 37502 4338
rect 21086 4274 21138 4286
rect 7310 4226 7362 4238
rect 7310 4162 7362 4174
rect 7758 4226 7810 4238
rect 7758 4162 7810 4174
rect 9550 4226 9602 4238
rect 9550 4162 9602 4174
rect 10782 4226 10834 4238
rect 18174 4226 18226 4238
rect 12338 4174 12350 4226
rect 12402 4174 12414 4226
rect 14466 4174 14478 4226
rect 14530 4174 14542 4226
rect 10782 4162 10834 4174
rect 18174 4162 18226 4174
rect 18622 4226 18674 4238
rect 18622 4162 18674 4174
rect 20862 4226 20914 4238
rect 24222 4226 24274 4238
rect 22082 4174 22094 4226
rect 22146 4174 22158 4226
rect 20862 4162 20914 4174
rect 24222 4162 24274 4174
rect 25454 4226 25506 4238
rect 25454 4162 25506 4174
rect 31614 4226 31666 4238
rect 31614 4162 31666 4174
rect 33294 4226 33346 4238
rect 33294 4162 33346 4174
rect 36654 4226 36706 4238
rect 36654 4162 36706 4174
rect 37998 4226 38050 4238
rect 37998 4162 38050 4174
rect 42478 4226 42530 4238
rect 42478 4162 42530 4174
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 11566 3666 11618 3678
rect 29374 3666 29426 3678
rect 21858 3614 21870 3666
rect 21922 3614 21934 3666
rect 25554 3614 25566 3666
rect 25618 3614 25630 3666
rect 11566 3602 11618 3614
rect 29374 3602 29426 3614
rect 36990 3666 37042 3678
rect 36990 3602 37042 3614
rect 40798 3666 40850 3678
rect 40798 3602 40850 3614
rect 6862 3554 6914 3566
rect 6862 3490 6914 3502
rect 8430 3554 8482 3566
rect 8430 3490 8482 3502
rect 9326 3554 9378 3566
rect 19854 3554 19906 3566
rect 31614 3554 31666 3566
rect 35422 3554 35474 3566
rect 12114 3502 12126 3554
rect 12178 3502 12190 3554
rect 13346 3502 13358 3554
rect 13410 3502 13422 3554
rect 15922 3502 15934 3554
rect 15986 3502 15998 3554
rect 16930 3502 16942 3554
rect 16994 3502 17006 3554
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 23874 3502 23886 3554
rect 23938 3502 23950 3554
rect 24658 3502 24670 3554
rect 24722 3502 24734 3554
rect 27346 3502 27358 3554
rect 27410 3502 27422 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 32162 3502 32174 3554
rect 32226 3502 32238 3554
rect 36418 3502 36430 3554
rect 36482 3502 36494 3554
rect 39778 3502 39790 3554
rect 39842 3502 39854 3554
rect 42914 3502 42926 3554
rect 42978 3502 42990 3554
rect 9326 3490 9378 3502
rect 19854 3490 19906 3502
rect 31614 3490 31666 3502
rect 35422 3490 35474 3502
rect 6414 3442 6466 3454
rect 6414 3378 6466 3390
rect 7086 3442 7138 3454
rect 7086 3378 7138 3390
rect 7422 3442 7474 3454
rect 7422 3378 7474 3390
rect 7758 3442 7810 3454
rect 7758 3378 7810 3390
rect 8094 3442 8146 3454
rect 8094 3378 8146 3390
rect 8766 3442 8818 3454
rect 8766 3378 8818 3390
rect 9662 3442 9714 3454
rect 9662 3378 9714 3390
rect 13134 3442 13186 3454
rect 20190 3442 20242 3454
rect 14802 3390 14814 3442
rect 14866 3390 14878 3442
rect 18498 3390 18510 3442
rect 18562 3390 18574 3442
rect 13134 3378 13186 3390
rect 20190 3378 20242 3390
rect 23662 3442 23714 3454
rect 23662 3378 23714 3390
rect 24894 3442 24946 3454
rect 24894 3378 24946 3390
rect 31278 3442 31330 3454
rect 35086 3442 35138 3454
rect 33730 3390 33742 3442
rect 33794 3390 33806 3442
rect 31278 3378 31330 3390
rect 35086 3378 35138 3390
rect 42702 3442 42754 3454
rect 42702 3378 42754 3390
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
<< via1 >>
rect 16046 46734 16098 46786
rect 17502 46734 17554 46786
rect 27582 46734 27634 46786
rect 28590 46734 28642 46786
rect 19070 46510 19122 46562
rect 19518 46510 19570 46562
rect 20078 46510 20130 46562
rect 18174 46398 18226 46450
rect 21646 46398 21698 46450
rect 23774 46398 23826 46450
rect 24894 46398 24946 46450
rect 26910 46398 26962 46450
rect 27470 46398 27522 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 17950 46062 18002 46114
rect 25566 46062 25618 46114
rect 30046 46062 30098 46114
rect 36990 46062 37042 46114
rect 41470 46062 41522 46114
rect 44606 46062 44658 46114
rect 8878 45950 8930 46002
rect 13470 45950 13522 46002
rect 22318 45950 22370 46002
rect 35198 45950 35250 46002
rect 9662 45838 9714 45890
rect 10558 45838 10610 45890
rect 11678 45838 11730 45890
rect 12350 45838 12402 45890
rect 13694 45838 13746 45890
rect 14814 45838 14866 45890
rect 15598 45838 15650 45890
rect 16046 45838 16098 45890
rect 17390 45838 17442 45890
rect 20078 45838 20130 45890
rect 20974 45838 21026 45890
rect 21646 45838 21698 45890
rect 22990 45838 23042 45890
rect 23774 45838 23826 45890
rect 25006 45838 25058 45890
rect 27470 45838 27522 45890
rect 28590 45838 28642 45890
rect 29262 45838 29314 45890
rect 32286 45838 32338 45890
rect 32846 45838 32898 45890
rect 35982 45838 36034 45890
rect 40462 45838 40514 45890
rect 43710 45838 43762 45890
rect 47406 45838 47458 45890
rect 22766 45726 22818 45778
rect 38894 45726 38946 45778
rect 39230 45726 39282 45778
rect 39790 45726 39842 45778
rect 40126 45726 40178 45778
rect 9998 45614 10050 45666
rect 10334 45614 10386 45666
rect 11902 45614 11954 45666
rect 12574 45614 12626 45666
rect 14030 45614 14082 45666
rect 15038 45614 15090 45666
rect 15374 45614 15426 45666
rect 16382 45614 16434 45666
rect 19854 45614 19906 45666
rect 20750 45614 20802 45666
rect 21422 45614 21474 45666
rect 23326 45614 23378 45666
rect 23998 45614 24050 45666
rect 27806 45614 27858 45666
rect 28366 45614 28418 45666
rect 32510 45614 32562 45666
rect 46510 45614 46562 45666
rect 46846 45614 46898 45666
rect 47518 45614 47570 45666
rect 47630 45614 47682 45666
rect 47854 45614 47906 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 10110 45278 10162 45330
rect 12126 45278 12178 45330
rect 12798 45278 12850 45330
rect 14814 45278 14866 45330
rect 15374 45278 15426 45330
rect 15822 45278 15874 45330
rect 16270 45278 16322 45330
rect 29710 45278 29762 45330
rect 42254 45278 42306 45330
rect 47182 45278 47234 45330
rect 16494 45166 16546 45218
rect 16830 45166 16882 45218
rect 24334 45166 24386 45218
rect 28478 45166 28530 45218
rect 28814 45166 28866 45218
rect 30494 45166 30546 45218
rect 30830 45166 30882 45218
rect 31166 45166 31218 45218
rect 31838 45166 31890 45218
rect 32174 45166 32226 45218
rect 32510 45166 32562 45218
rect 33182 45166 33234 45218
rect 33518 45166 33570 45218
rect 33854 45166 33906 45218
rect 17390 45054 17442 45106
rect 21086 45054 21138 45106
rect 24558 45054 24610 45106
rect 25342 45054 25394 45106
rect 29374 45054 29426 45106
rect 30270 45054 30322 45106
rect 31614 45054 31666 45106
rect 34078 45054 34130 45106
rect 36990 45054 37042 45106
rect 37774 45054 37826 45106
rect 41246 45054 41298 45106
rect 44158 45054 44210 45106
rect 48078 45054 48130 45106
rect 18174 44942 18226 44994
rect 20302 44942 20354 44994
rect 20526 44942 20578 44994
rect 20750 44942 20802 44994
rect 21758 44942 21810 44994
rect 23886 44942 23938 44994
rect 26014 44942 26066 44994
rect 28142 44942 28194 44994
rect 45390 44942 45442 44994
rect 47518 44942 47570 44994
rect 36430 44830 36482 44882
rect 40126 44830 40178 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 36206 44494 36258 44546
rect 41134 44494 41186 44546
rect 45838 44494 45890 44546
rect 17054 44382 17106 44434
rect 18398 44382 18450 44434
rect 19070 44382 19122 44434
rect 21422 44382 21474 44434
rect 21870 44382 21922 44434
rect 24894 44382 24946 44434
rect 27246 44382 27298 44434
rect 28254 44382 28306 44434
rect 30942 44382 30994 44434
rect 43822 44382 43874 44434
rect 14254 44270 14306 44322
rect 18510 44270 18562 44322
rect 19518 44270 19570 44322
rect 19742 44270 19794 44322
rect 20078 44270 20130 44322
rect 20526 44270 20578 44322
rect 20750 44270 20802 44322
rect 21310 44270 21362 44322
rect 31838 44270 31890 44322
rect 32622 44270 32674 44322
rect 33854 44270 33906 44322
rect 37550 44270 37602 44322
rect 38222 44270 38274 44322
rect 38782 44270 38834 44322
rect 41694 44270 41746 44322
rect 44830 44270 44882 44322
rect 14926 44158 14978 44210
rect 19294 44158 19346 44210
rect 19406 44158 19458 44210
rect 20414 44158 20466 44210
rect 23438 44158 23490 44210
rect 32174 44158 32226 44210
rect 32846 44158 32898 44210
rect 37774 44158 37826 44210
rect 38446 44158 38498 44210
rect 47742 44158 47794 44210
rect 18062 44046 18114 44098
rect 18286 44046 18338 44098
rect 23326 44046 23378 44098
rect 29598 44046 29650 44098
rect 29934 44046 29986 44098
rect 30382 44046 30434 44098
rect 31166 44046 31218 44098
rect 31502 44046 31554 44098
rect 33182 44046 33234 44098
rect 33518 44046 33570 44098
rect 37102 44046 37154 44098
rect 48078 44046 48130 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 18398 43710 18450 43762
rect 22430 43710 22482 43762
rect 22766 43710 22818 43762
rect 24670 43710 24722 43762
rect 25342 43710 25394 43762
rect 27358 43710 27410 43762
rect 27806 43710 27858 43762
rect 28926 43710 28978 43762
rect 17502 43598 17554 43650
rect 18510 43598 18562 43650
rect 19742 43598 19794 43650
rect 20526 43598 20578 43650
rect 21870 43598 21922 43650
rect 24110 43598 24162 43650
rect 25230 43598 25282 43650
rect 25678 43598 25730 43650
rect 26238 43598 26290 43650
rect 26798 43598 26850 43650
rect 30382 43598 30434 43650
rect 31502 43598 31554 43650
rect 32510 43598 32562 43650
rect 33854 43598 33906 43650
rect 34526 43598 34578 43650
rect 41470 43598 41522 43650
rect 4286 43486 4338 43538
rect 4846 43486 4898 43538
rect 10110 43486 10162 43538
rect 10558 43486 10610 43538
rect 10782 43486 10834 43538
rect 16494 43486 16546 43538
rect 16718 43486 16770 43538
rect 17390 43486 17442 43538
rect 17614 43486 17666 43538
rect 18062 43486 18114 43538
rect 21646 43486 21698 43538
rect 22430 43486 22482 43538
rect 22990 43486 23042 43538
rect 23438 43486 23490 43538
rect 23886 43486 23938 43538
rect 24670 43486 24722 43538
rect 25454 43486 25506 43538
rect 26574 43486 26626 43538
rect 27134 43486 27186 43538
rect 28030 43486 28082 43538
rect 28366 43486 28418 43538
rect 28814 43486 28866 43538
rect 30830 43486 30882 43538
rect 31726 43486 31778 43538
rect 32286 43486 32338 43538
rect 33630 43486 33682 43538
rect 34302 43486 34354 43538
rect 35086 43486 35138 43538
rect 37774 43486 37826 43538
rect 41246 43486 41298 43538
rect 42926 43486 42978 43538
rect 45838 43486 45890 43538
rect 10334 43374 10386 43426
rect 16830 43374 16882 43426
rect 18286 43374 18338 43426
rect 22094 43374 22146 43426
rect 22878 43374 22930 43426
rect 27918 43374 27970 43426
rect 31278 43374 31330 43426
rect 33182 43374 33234 43426
rect 42366 43374 42418 43426
rect 44942 43374 44994 43426
rect 47854 43374 47906 43426
rect 1934 43262 1986 43314
rect 19854 43262 19906 43314
rect 24334 43262 24386 43314
rect 26126 43262 26178 43314
rect 27022 43262 27074 43314
rect 28702 43262 28754 43314
rect 37214 43262 37266 43314
rect 40126 43262 40178 43314
rect 41806 43262 41858 43314
rect 42142 43262 42194 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 19854 42926 19906 42978
rect 27134 42926 27186 42978
rect 36206 42926 36258 42978
rect 42814 42926 42866 42978
rect 2046 42814 2098 42866
rect 8878 42814 8930 42866
rect 11006 42814 11058 42866
rect 14478 42814 14530 42866
rect 19518 42814 19570 42866
rect 22542 42814 22594 42866
rect 25006 42814 25058 42866
rect 25566 42814 25618 42866
rect 29150 42814 29202 42866
rect 31278 42814 31330 42866
rect 41918 42814 41970 42866
rect 43710 42814 43762 42866
rect 47966 42814 48018 42866
rect 4062 42702 4114 42754
rect 8206 42702 8258 42754
rect 13582 42702 13634 42754
rect 13806 42702 13858 42754
rect 14142 42702 14194 42754
rect 14366 42702 14418 42754
rect 19406 42702 19458 42754
rect 20078 42702 20130 42754
rect 23214 42702 23266 42754
rect 24782 42702 24834 42754
rect 25118 42702 25170 42754
rect 25790 42702 25842 42754
rect 27134 42702 27186 42754
rect 27470 42702 27522 42754
rect 31950 42702 32002 42754
rect 33294 42702 33346 42754
rect 33854 42702 33906 42754
rect 37662 42702 37714 42754
rect 38334 42702 38386 42754
rect 39006 42702 39058 42754
rect 42478 42702 42530 42754
rect 43486 42702 43538 42754
rect 45614 42702 45666 42754
rect 19630 42590 19682 42642
rect 22430 42590 22482 42642
rect 22654 42590 22706 42642
rect 23550 42590 23602 42642
rect 25454 42590 25506 42642
rect 26798 42590 26850 42642
rect 27582 42590 27634 42642
rect 32510 42590 32562 42642
rect 32846 42590 32898 42642
rect 33518 42590 33570 42642
rect 37998 42590 38050 42642
rect 38670 42590 38722 42642
rect 39790 42590 39842 42642
rect 42254 42590 42306 42642
rect 44830 42590 44882 42642
rect 45166 42590 45218 42642
rect 11454 42478 11506 42530
rect 13918 42478 13970 42530
rect 23438 42478 23490 42530
rect 36990 42478 37042 42530
rect 37326 42478 37378 42530
rect 43150 42478 43202 42530
rect 44158 42478 44210 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 10110 42142 10162 42194
rect 11006 42142 11058 42194
rect 11902 42142 11954 42194
rect 15262 42142 15314 42194
rect 20078 42142 20130 42194
rect 23214 42142 23266 42194
rect 34750 42142 34802 42194
rect 35086 42142 35138 42194
rect 39230 42142 39282 42194
rect 42030 42142 42082 42194
rect 11118 42030 11170 42082
rect 14142 42030 14194 42082
rect 15486 42030 15538 42082
rect 17390 42030 17442 42082
rect 34078 42030 34130 42082
rect 39006 42030 39058 42082
rect 40350 42030 40402 42082
rect 41806 42030 41858 42082
rect 4286 41918 4338 41970
rect 5294 41918 5346 41970
rect 9998 41918 10050 41970
rect 10894 41918 10946 41970
rect 11566 41918 11618 41970
rect 14814 41918 14866 41970
rect 15374 41918 15426 41970
rect 15934 41918 15986 41970
rect 17614 41918 17666 41970
rect 18062 41918 18114 41970
rect 20302 41918 20354 41970
rect 20638 41918 20690 41970
rect 20750 41918 20802 41970
rect 21086 41918 21138 41970
rect 21422 41918 21474 41970
rect 23438 41918 23490 41970
rect 33742 41918 33794 41970
rect 34414 41918 34466 41970
rect 35422 41918 35474 41970
rect 35870 41918 35922 41970
rect 39678 41918 39730 41970
rect 40126 41918 40178 41970
rect 40910 41918 40962 41970
rect 41022 41918 41074 41970
rect 41246 41918 41298 41970
rect 41358 41918 41410 41970
rect 41918 41918 41970 41970
rect 42366 41918 42418 41970
rect 42814 41918 42866 41970
rect 45726 41918 45778 41970
rect 5742 41806 5794 41858
rect 16270 41806 16322 41858
rect 17502 41806 17554 41858
rect 20190 41806 20242 41858
rect 21310 41806 21362 41858
rect 32174 41806 32226 41858
rect 33182 41806 33234 41858
rect 36542 41806 36594 41858
rect 38670 41806 38722 41858
rect 39118 41806 39170 41858
rect 47630 41806 47682 41858
rect 1934 41694 1986 41746
rect 4958 41694 5010 41746
rect 5294 41694 5346 41746
rect 45054 41694 45106 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 21870 41358 21922 41410
rect 26798 41358 26850 41410
rect 41134 41358 41186 41410
rect 44046 41358 44098 41410
rect 48190 41358 48242 41410
rect 4622 41246 4674 41298
rect 6414 41246 6466 41298
rect 8542 41246 8594 41298
rect 14926 41246 14978 41298
rect 16830 41246 16882 41298
rect 18958 41246 19010 41298
rect 22206 41246 22258 41298
rect 26126 41246 26178 41298
rect 27134 41246 27186 41298
rect 34638 41246 34690 41298
rect 37102 41246 37154 41298
rect 47742 41246 47794 41298
rect 1710 41134 1762 41186
rect 5742 41134 5794 41186
rect 16046 41134 16098 41186
rect 21534 41134 21586 41186
rect 22318 41134 22370 41186
rect 25790 41134 25842 41186
rect 26462 41134 26514 41186
rect 27022 41134 27074 41186
rect 27582 41134 27634 41186
rect 30830 41134 30882 41186
rect 31838 41134 31890 41186
rect 35086 41134 35138 41186
rect 35534 41134 35586 41186
rect 36206 41134 36258 41186
rect 36878 41134 36930 41186
rect 37550 41134 37602 41186
rect 38110 41134 38162 41186
rect 38782 41134 38834 41186
rect 41694 41134 41746 41186
rect 44942 41134 44994 41186
rect 2494 41022 2546 41074
rect 22094 41022 22146 41074
rect 23214 41022 23266 41074
rect 23550 41022 23602 41074
rect 25006 41022 25058 41074
rect 25342 41022 25394 41074
rect 27246 41022 27298 41074
rect 28030 41022 28082 41074
rect 32510 41022 32562 41074
rect 36430 41022 36482 41074
rect 37326 41022 37378 41074
rect 38446 41022 38498 41074
rect 45614 41022 45666 41074
rect 5070 40910 5122 40962
rect 8990 40910 9042 40962
rect 23886 40910 23938 40962
rect 24222 40910 24274 40962
rect 26014 40910 26066 40962
rect 27694 40910 27746 40962
rect 27806 40910 27858 40962
rect 35646 40910 35698 40962
rect 35758 40910 35810 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 5742 40574 5794 40626
rect 10222 40574 10274 40626
rect 18958 40574 19010 40626
rect 22654 40574 22706 40626
rect 22990 40574 23042 40626
rect 25230 40574 25282 40626
rect 25566 40574 25618 40626
rect 27246 40574 27298 40626
rect 33742 40574 33794 40626
rect 34078 40574 34130 40626
rect 37102 40574 37154 40626
rect 41134 40574 41186 40626
rect 4622 40462 4674 40514
rect 5406 40462 5458 40514
rect 6862 40462 6914 40514
rect 9774 40462 9826 40514
rect 11230 40462 11282 40514
rect 11454 40462 11506 40514
rect 12126 40462 12178 40514
rect 15150 40462 15202 40514
rect 26462 40462 26514 40514
rect 26574 40462 26626 40514
rect 29822 40462 29874 40514
rect 34638 40462 34690 40514
rect 36542 40462 36594 40514
rect 39454 40462 39506 40514
rect 41470 40462 41522 40514
rect 4286 40350 4338 40402
rect 4958 40350 5010 40402
rect 6190 40350 6242 40402
rect 9886 40350 9938 40402
rect 11006 40350 11058 40402
rect 11566 40350 11618 40402
rect 17390 40350 17442 40402
rect 19518 40350 19570 40402
rect 20190 40350 20242 40402
rect 23662 40350 23714 40402
rect 24222 40350 24274 40402
rect 30606 40350 30658 40402
rect 30942 40350 30994 40402
rect 31390 40350 31442 40402
rect 35086 40350 35138 40402
rect 35310 40350 35362 40402
rect 35422 40350 35474 40402
rect 35646 40350 35698 40402
rect 36206 40350 36258 40402
rect 37438 40350 37490 40402
rect 37774 40350 37826 40402
rect 40910 40350 40962 40402
rect 41246 40350 41298 40402
rect 42702 40350 42754 40402
rect 45950 40350 46002 40402
rect 8990 40238 9042 40290
rect 10670 40238 10722 40290
rect 17614 40238 17666 40290
rect 17726 40238 17778 40290
rect 18734 40238 18786 40290
rect 22318 40238 22370 40290
rect 23774 40238 23826 40290
rect 27022 40238 27074 40290
rect 27358 40238 27410 40290
rect 27694 40238 27746 40290
rect 42142 40238 42194 40290
rect 42366 40238 42418 40290
rect 47742 40238 47794 40290
rect 1934 40126 1986 40178
rect 12238 40126 12290 40178
rect 15262 40126 15314 40178
rect 19070 40126 19122 40178
rect 23998 40126 24050 40178
rect 26462 40126 26514 40178
rect 34414 40126 34466 40178
rect 41806 40126 41858 40178
rect 45054 40126 45106 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 4398 39790 4450 39842
rect 26798 39790 26850 39842
rect 35982 39790 36034 39842
rect 36542 39790 36594 39842
rect 43598 39790 43650 39842
rect 2494 39678 2546 39730
rect 4286 39678 4338 39730
rect 5070 39678 5122 39730
rect 11566 39678 11618 39730
rect 17614 39678 17666 39730
rect 19406 39678 19458 39730
rect 19630 39678 19682 39730
rect 20078 39678 20130 39730
rect 26910 39678 26962 39730
rect 34862 39678 34914 39730
rect 35982 39678 36034 39730
rect 36430 39678 36482 39730
rect 37774 39678 37826 39730
rect 41022 39678 41074 39730
rect 3726 39566 3778 39618
rect 10110 39566 10162 39618
rect 10558 39566 10610 39618
rect 11678 39566 11730 39618
rect 12238 39566 12290 39618
rect 14814 39566 14866 39618
rect 19182 39566 19234 39618
rect 19966 39566 20018 39618
rect 20190 39566 20242 39618
rect 24222 39566 24274 39618
rect 36990 39566 37042 39618
rect 38110 39566 38162 39618
rect 41694 39566 41746 39618
rect 45166 39566 45218 39618
rect 48078 39566 48130 39618
rect 2158 39454 2210 39506
rect 2382 39454 2434 39506
rect 7534 39454 7586 39506
rect 11230 39454 11282 39506
rect 12686 39454 12738 39506
rect 12910 39454 12962 39506
rect 13582 39454 13634 39506
rect 13918 39454 13970 39506
rect 15486 39454 15538 39506
rect 18174 39454 18226 39506
rect 18398 39454 18450 39506
rect 18846 39454 18898 39506
rect 34302 39454 34354 39506
rect 38894 39454 38946 39506
rect 46622 39454 46674 39506
rect 2606 39342 2658 39394
rect 3278 39342 3330 39394
rect 8094 39342 8146 39394
rect 9214 39342 9266 39394
rect 11454 39342 11506 39394
rect 12462 39342 12514 39394
rect 13806 39342 13858 39394
rect 14030 39342 14082 39394
rect 17950 39342 18002 39394
rect 18062 39342 18114 39394
rect 19742 39342 19794 39394
rect 23886 39342 23938 39394
rect 30606 39342 30658 39394
rect 31278 39342 31330 39394
rect 31614 39342 31666 39394
rect 31950 39342 32002 39394
rect 35310 39342 35362 39394
rect 37326 39342 37378 39394
rect 44830 39342 44882 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 7310 39006 7362 39058
rect 10670 39006 10722 39058
rect 15486 39006 15538 39058
rect 18286 39006 18338 39058
rect 19966 39006 20018 39058
rect 23662 39006 23714 39058
rect 32510 39006 32562 39058
rect 34526 39006 34578 39058
rect 36654 39006 36706 39058
rect 38670 39006 38722 39058
rect 39454 39006 39506 39058
rect 40910 39006 40962 39058
rect 41918 39006 41970 39058
rect 3614 38894 3666 38946
rect 3726 38894 3778 38946
rect 4286 38894 4338 38946
rect 4622 38894 4674 38946
rect 8318 38894 8370 38946
rect 9550 38894 9602 38946
rect 11006 38894 11058 38946
rect 12350 38894 12402 38946
rect 15934 38894 15986 38946
rect 33182 38894 33234 38946
rect 33406 38894 33458 38946
rect 33742 38894 33794 38946
rect 33854 38894 33906 38946
rect 33966 38894 34018 38946
rect 36990 38894 37042 38946
rect 37998 38894 38050 38946
rect 39342 38894 39394 38946
rect 41134 38894 41186 38946
rect 41358 38894 41410 38946
rect 42814 38894 42866 38946
rect 47518 38894 47570 38946
rect 48190 38894 48242 38946
rect 2718 38782 2770 38834
rect 3950 38782 4002 38834
rect 4398 38782 4450 38834
rect 4846 38782 4898 38834
rect 6414 38782 6466 38834
rect 6750 38782 6802 38834
rect 7534 38782 7586 38834
rect 7982 38782 8034 38834
rect 8990 38782 9042 38834
rect 9662 38782 9714 38834
rect 10110 38782 10162 38834
rect 11118 38782 11170 38834
rect 11678 38782 11730 38834
rect 15262 38782 15314 38834
rect 15710 38782 15762 38834
rect 17502 38782 17554 38834
rect 17950 38782 18002 38834
rect 18622 38782 18674 38834
rect 20302 38782 20354 38834
rect 23998 38782 24050 38834
rect 24446 38782 24498 38834
rect 29150 38782 29202 38834
rect 32398 38782 32450 38834
rect 37326 38782 37378 38834
rect 37662 38782 37714 38834
rect 38334 38782 38386 38834
rect 39678 38782 39730 38834
rect 39902 38782 39954 38834
rect 41022 38782 41074 38834
rect 42142 38782 42194 38834
rect 42478 38782 42530 38834
rect 43038 38782 43090 38834
rect 45838 38782 45890 38834
rect 46510 38782 46562 38834
rect 46846 38782 46898 38834
rect 47070 38782 47122 38834
rect 47182 38782 47234 38834
rect 47854 38782 47906 38834
rect 2382 38670 2434 38722
rect 2606 38670 2658 38722
rect 3166 38670 3218 38722
rect 6638 38670 6690 38722
rect 7870 38670 7922 38722
rect 14478 38670 14530 38722
rect 19070 38670 19122 38722
rect 29822 38670 29874 38722
rect 31950 38670 32002 38722
rect 33070 38670 33122 38722
rect 40350 38670 40402 38722
rect 42030 38670 42082 38722
rect 43710 38670 43762 38722
rect 2270 38558 2322 38610
rect 43374 38558 43426 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 29934 38222 29986 38274
rect 30270 38222 30322 38274
rect 43598 38222 43650 38274
rect 2494 38110 2546 38162
rect 4622 38110 4674 38162
rect 12014 38110 12066 38162
rect 28366 38110 28418 38162
rect 36094 38110 36146 38162
rect 36990 38110 37042 38162
rect 38110 38110 38162 38162
rect 38558 38110 38610 38162
rect 1822 37998 1874 38050
rect 5630 37998 5682 38050
rect 5966 37998 6018 38050
rect 6414 37998 6466 38050
rect 7310 37998 7362 38050
rect 8654 37998 8706 38050
rect 9662 37998 9714 38050
rect 10446 37998 10498 38050
rect 11454 37998 11506 38050
rect 20190 37998 20242 38050
rect 23214 37998 23266 38050
rect 23998 37998 24050 38050
rect 24782 37998 24834 38050
rect 25566 37998 25618 38050
rect 29262 37998 29314 38050
rect 33182 37998 33234 38050
rect 39790 37998 39842 38050
rect 41022 37998 41074 38050
rect 41694 37998 41746 38050
rect 44830 37998 44882 38050
rect 46062 37998 46114 38050
rect 5742 37886 5794 37938
rect 7534 37886 7586 37938
rect 23774 37886 23826 37938
rect 25006 37886 25058 37938
rect 26238 37886 26290 37938
rect 33966 37886 34018 37938
rect 40014 37886 40066 37938
rect 40350 37886 40402 37938
rect 40686 37886 40738 37938
rect 41358 37886 41410 37938
rect 45166 37886 45218 37938
rect 47406 37886 47458 37938
rect 5070 37774 5122 37826
rect 6638 37774 6690 37826
rect 9550 37774 9602 37826
rect 12462 37774 12514 37826
rect 14030 37774 14082 37826
rect 20414 37774 20466 37826
rect 23438 37774 23490 37826
rect 24334 37774 24386 37826
rect 30046 37774 30098 37826
rect 32174 37774 32226 37826
rect 32846 37774 32898 37826
rect 37102 37774 37154 37826
rect 38894 37774 38946 37826
rect 39454 37774 39506 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 4958 37438 5010 37490
rect 13134 37438 13186 37490
rect 15598 37438 15650 37490
rect 18510 37438 18562 37490
rect 18846 37438 18898 37490
rect 25342 37438 25394 37490
rect 34974 37438 35026 37490
rect 36094 37438 36146 37490
rect 36206 37438 36258 37490
rect 6638 37326 6690 37378
rect 7534 37326 7586 37378
rect 11790 37326 11842 37378
rect 13022 37326 13074 37378
rect 14254 37326 14306 37378
rect 14926 37326 14978 37378
rect 15710 37326 15762 37378
rect 17838 37326 17890 37378
rect 18174 37326 18226 37378
rect 20526 37326 20578 37378
rect 25902 37326 25954 37378
rect 26014 37326 26066 37378
rect 27694 37326 27746 37378
rect 27806 37326 27858 37378
rect 35422 37326 35474 37378
rect 45278 37326 45330 37378
rect 4286 37214 4338 37266
rect 5182 37214 5234 37266
rect 7086 37214 7138 37266
rect 8094 37214 8146 37266
rect 12574 37214 12626 37266
rect 12910 37214 12962 37266
rect 13358 37214 13410 37266
rect 13582 37214 13634 37266
rect 14590 37214 14642 37266
rect 15262 37214 15314 37266
rect 15934 37214 15986 37266
rect 19742 37214 19794 37266
rect 25678 37214 25730 37266
rect 26462 37214 26514 37266
rect 34862 37214 34914 37266
rect 35086 37214 35138 37266
rect 35982 37214 36034 37266
rect 36654 37214 36706 37266
rect 37214 37214 37266 37266
rect 41022 37214 41074 37266
rect 44718 37214 44770 37266
rect 44942 37214 44994 37266
rect 45838 37214 45890 37266
rect 7758 37102 7810 37154
rect 9662 37102 9714 37154
rect 15038 37102 15090 37154
rect 22654 37102 22706 37154
rect 26014 37102 26066 37154
rect 37998 37102 38050 37154
rect 40126 37102 40178 37154
rect 41694 37102 41746 37154
rect 43822 37102 43874 37154
rect 44270 37102 44322 37154
rect 45166 37102 45218 37154
rect 47742 37102 47794 37154
rect 1934 36990 1986 37042
rect 44270 36990 44322 37042
rect 44494 36990 44546 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 4622 36654 4674 36706
rect 10894 36654 10946 36706
rect 13582 36654 13634 36706
rect 19966 36654 20018 36706
rect 20302 36654 20354 36706
rect 40574 36654 40626 36706
rect 41022 36654 41074 36706
rect 43038 36654 43090 36706
rect 1934 36542 1986 36594
rect 4958 36542 5010 36594
rect 9102 36542 9154 36594
rect 12798 36542 12850 36594
rect 15598 36542 15650 36594
rect 17726 36542 17778 36594
rect 18174 36542 18226 36594
rect 19742 36542 19794 36594
rect 20750 36542 20802 36594
rect 25678 36542 25730 36594
rect 29262 36542 29314 36594
rect 32734 36542 32786 36594
rect 35646 36542 35698 36594
rect 40014 36542 40066 36594
rect 40574 36542 40626 36594
rect 41806 36542 41858 36594
rect 44158 36542 44210 36594
rect 47966 36542 48018 36594
rect 4286 36430 4338 36482
rect 5742 36430 5794 36482
rect 5854 36430 5906 36482
rect 7198 36430 7250 36482
rect 7646 36430 7698 36482
rect 7870 36430 7922 36482
rect 10782 36430 10834 36482
rect 13470 36430 13522 36482
rect 14814 36430 14866 36482
rect 18286 36430 18338 36482
rect 23774 36430 23826 36482
rect 24110 36430 24162 36482
rect 24334 36430 24386 36482
rect 28590 36430 28642 36482
rect 29822 36430 29874 36482
rect 38110 36430 38162 36482
rect 39342 36430 39394 36482
rect 41582 36430 41634 36482
rect 42142 36430 42194 36482
rect 43598 36430 43650 36482
rect 45614 36430 45666 36482
rect 4846 36318 4898 36370
rect 8318 36318 8370 36370
rect 8430 36318 8482 36370
rect 13582 36318 13634 36370
rect 19294 36318 19346 36370
rect 23326 36318 23378 36370
rect 27806 36318 27858 36370
rect 30606 36318 30658 36370
rect 35758 36318 35810 36370
rect 37774 36318 37826 36370
rect 38334 36318 38386 36370
rect 39230 36318 39282 36370
rect 42030 36318 42082 36370
rect 42814 36318 42866 36370
rect 45278 36318 45330 36370
rect 6302 36206 6354 36258
rect 7758 36206 7810 36258
rect 8654 36206 8706 36258
rect 9214 36206 9266 36258
rect 18062 36206 18114 36258
rect 18510 36206 18562 36258
rect 19182 36206 19234 36258
rect 22430 36206 22482 36258
rect 22654 36206 22706 36258
rect 22766 36206 22818 36258
rect 22878 36206 22930 36258
rect 23438 36206 23490 36258
rect 24222 36206 24274 36258
rect 24446 36206 24498 36258
rect 33182 36206 33234 36258
rect 37998 36206 38050 36258
rect 39118 36206 39170 36258
rect 39566 36206 39618 36258
rect 40126 36206 40178 36258
rect 41022 36206 41074 36258
rect 43374 36206 43426 36258
rect 44046 36206 44098 36258
rect 44270 36206 44322 36258
rect 44942 36206 44994 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 10670 35870 10722 35922
rect 10894 35870 10946 35922
rect 11566 35870 11618 35922
rect 11790 35870 11842 35922
rect 13806 35870 13858 35922
rect 14478 35870 14530 35922
rect 14814 35870 14866 35922
rect 24670 35870 24722 35922
rect 27022 35870 27074 35922
rect 30606 35870 30658 35922
rect 36878 35870 36930 35922
rect 37102 35870 37154 35922
rect 41582 35870 41634 35922
rect 42926 35870 42978 35922
rect 43262 35870 43314 35922
rect 43598 35870 43650 35922
rect 44718 35870 44770 35922
rect 44830 35870 44882 35922
rect 9550 35758 9602 35810
rect 19070 35758 19122 35810
rect 22318 35758 22370 35810
rect 22542 35758 22594 35810
rect 23214 35758 23266 35810
rect 23326 35758 23378 35810
rect 23774 35758 23826 35810
rect 23998 35758 24050 35810
rect 36654 35758 36706 35810
rect 44494 35758 44546 35810
rect 46062 35758 46114 35810
rect 1822 35646 1874 35698
rect 2494 35646 2546 35698
rect 4958 35646 5010 35698
rect 5518 35646 5570 35698
rect 7534 35646 7586 35698
rect 8766 35646 8818 35698
rect 8990 35646 9042 35698
rect 9998 35646 10050 35698
rect 10558 35646 10610 35698
rect 11342 35646 11394 35698
rect 11902 35646 11954 35698
rect 14030 35646 14082 35698
rect 15822 35646 15874 35698
rect 18398 35646 18450 35698
rect 25566 35646 25618 35698
rect 25790 35646 25842 35698
rect 30382 35646 30434 35698
rect 31166 35646 31218 35698
rect 31726 35646 31778 35698
rect 33406 35646 33458 35698
rect 42142 35646 42194 35698
rect 42590 35646 42642 35698
rect 43934 35646 43986 35698
rect 44942 35646 44994 35698
rect 45390 35646 45442 35698
rect 4622 35534 4674 35586
rect 5182 35534 5234 35586
rect 5966 35534 6018 35586
rect 7982 35534 8034 35586
rect 11678 35534 11730 35586
rect 13470 35534 13522 35586
rect 15262 35534 15314 35586
rect 16270 35534 16322 35586
rect 17502 35534 17554 35586
rect 17950 35534 18002 35586
rect 21198 35534 21250 35586
rect 26462 35534 26514 35586
rect 26798 35534 26850 35586
rect 27134 35534 27186 35586
rect 30718 35534 30770 35586
rect 31054 35534 31106 35586
rect 32510 35534 32562 35586
rect 34190 35534 34242 35586
rect 36318 35534 36370 35586
rect 36766 35534 36818 35586
rect 41134 35534 41186 35586
rect 48190 35534 48242 35586
rect 5406 35422 5458 35474
rect 8318 35422 8370 35474
rect 15150 35422 15202 35474
rect 21646 35422 21698 35474
rect 21982 35422 22034 35474
rect 23326 35422 23378 35474
rect 24334 35422 24386 35474
rect 24558 35422 24610 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 10782 35086 10834 35138
rect 11566 35086 11618 35138
rect 22654 35086 22706 35138
rect 22878 35086 22930 35138
rect 23326 35086 23378 35138
rect 41022 35086 41074 35138
rect 43598 35086 43650 35138
rect 1934 34974 1986 35026
rect 15486 34974 15538 35026
rect 16830 34974 16882 35026
rect 19742 34974 19794 35026
rect 22430 34974 22482 35026
rect 26686 34974 26738 35026
rect 32062 34974 32114 35026
rect 33742 34974 33794 35026
rect 34526 34974 34578 35026
rect 40574 34974 40626 35026
rect 41470 34974 41522 35026
rect 42366 34974 42418 35026
rect 42702 34974 42754 35026
rect 46958 34974 47010 35026
rect 4286 34862 4338 34914
rect 4734 34862 4786 34914
rect 8654 34862 8706 34914
rect 9774 34862 9826 34914
rect 11118 34862 11170 34914
rect 11790 34862 11842 34914
rect 12014 34862 12066 34914
rect 14478 34862 14530 34914
rect 14814 34862 14866 34914
rect 15038 34862 15090 34914
rect 15374 34862 15426 34914
rect 16046 34862 16098 34914
rect 18846 34862 18898 34914
rect 19854 34862 19906 34914
rect 24894 34862 24946 34914
rect 25902 34862 25954 34914
rect 29262 34862 29314 34914
rect 32846 34862 32898 34914
rect 34638 34862 34690 34914
rect 34974 34862 35026 34914
rect 37214 34862 37266 34914
rect 37774 34862 37826 34914
rect 43150 34862 43202 34914
rect 43934 34862 43986 34914
rect 45054 34862 45106 34914
rect 48078 34862 48130 34914
rect 8766 34750 8818 34802
rect 12798 34750 12850 34802
rect 12910 34750 12962 34802
rect 13806 34750 13858 34802
rect 24670 34750 24722 34802
rect 26238 34750 26290 34802
rect 29934 34750 29986 34802
rect 32622 34750 32674 34802
rect 34414 34750 34466 34802
rect 38446 34750 38498 34802
rect 40910 34750 40962 34802
rect 43486 34750 43538 34802
rect 44270 34750 44322 34802
rect 45278 34750 45330 34802
rect 12126 34638 12178 34690
rect 12238 34638 12290 34690
rect 12574 34638 12626 34690
rect 13694 34638 13746 34690
rect 14702 34638 14754 34690
rect 15598 34638 15650 34690
rect 19406 34638 19458 34690
rect 19630 34638 19682 34690
rect 20414 34638 20466 34690
rect 20750 34638 20802 34690
rect 33854 34638 33906 34690
rect 36990 34638 37042 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 2046 34302 2098 34354
rect 2494 34302 2546 34354
rect 6862 34302 6914 34354
rect 7310 34302 7362 34354
rect 7646 34302 7698 34354
rect 20750 34302 20802 34354
rect 37438 34302 37490 34354
rect 44718 34302 44770 34354
rect 45838 34302 45890 34354
rect 47854 34302 47906 34354
rect 1710 34190 1762 34242
rect 10558 34190 10610 34242
rect 11006 34190 11058 34242
rect 15150 34190 15202 34242
rect 31054 34190 31106 34242
rect 31726 34190 31778 34242
rect 47294 34190 47346 34242
rect 3950 34078 4002 34130
rect 10110 34078 10162 34130
rect 10782 34078 10834 34130
rect 12014 34078 12066 34130
rect 13022 34078 13074 34130
rect 13470 34078 13522 34130
rect 13694 34078 13746 34130
rect 16270 34078 16322 34130
rect 18286 34078 18338 34130
rect 31390 34078 31442 34130
rect 32062 34078 32114 34130
rect 33406 34078 33458 34130
rect 33630 34078 33682 34130
rect 37214 34078 37266 34130
rect 37774 34078 37826 34130
rect 41470 34078 41522 34130
rect 44942 34078 44994 34130
rect 45390 34078 45442 34130
rect 45726 34078 45778 34130
rect 45950 34078 46002 34130
rect 46286 34078 46338 34130
rect 46622 34078 46674 34130
rect 46734 34078 46786 34130
rect 47518 34078 47570 34130
rect 4622 33966 4674 34018
rect 8094 33966 8146 34018
rect 11118 33966 11170 34018
rect 14926 33966 14978 34018
rect 18846 33966 18898 34018
rect 33182 33966 33234 34018
rect 36766 33966 36818 34018
rect 40126 33966 40178 34018
rect 42142 33966 42194 34018
rect 44270 33966 44322 34018
rect 46398 33966 46450 34018
rect 10222 33854 10274 33906
rect 34078 33854 34130 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 9214 33518 9266 33570
rect 9886 33518 9938 33570
rect 11454 33518 11506 33570
rect 24558 33518 24610 33570
rect 34414 33518 34466 33570
rect 44942 33518 44994 33570
rect 7422 33406 7474 33458
rect 11230 33406 11282 33458
rect 12910 33406 12962 33458
rect 17166 33406 17218 33458
rect 20414 33406 20466 33458
rect 23102 33406 23154 33458
rect 25902 33406 25954 33458
rect 26462 33406 26514 33458
rect 29598 33406 29650 33458
rect 30942 33406 30994 33458
rect 32510 33406 32562 33458
rect 37998 33406 38050 33458
rect 38446 33406 38498 33458
rect 41582 33406 41634 33458
rect 42254 33406 42306 33458
rect 46062 33406 46114 33458
rect 48190 33406 48242 33458
rect 1822 33294 1874 33346
rect 5742 33294 5794 33346
rect 6302 33294 6354 33346
rect 8430 33294 8482 33346
rect 8766 33294 8818 33346
rect 9102 33294 9154 33346
rect 9998 33294 10050 33346
rect 10222 33294 10274 33346
rect 12126 33294 12178 33346
rect 13694 33294 13746 33346
rect 14366 33294 14418 33346
rect 17950 33294 18002 33346
rect 19518 33294 19570 33346
rect 20078 33294 20130 33346
rect 24110 33294 24162 33346
rect 26014 33294 26066 33346
rect 27806 33294 27858 33346
rect 29150 33294 29202 33346
rect 29486 33294 29538 33346
rect 33630 33294 33682 33346
rect 34750 33294 34802 33346
rect 34974 33294 35026 33346
rect 36318 33294 36370 33346
rect 38222 33294 38274 33346
rect 38670 33294 38722 33346
rect 39230 33294 39282 33346
rect 42366 33294 42418 33346
rect 42702 33294 42754 33346
rect 43374 33294 43426 33346
rect 43486 33294 43538 33346
rect 43934 33294 43986 33346
rect 44830 33294 44882 33346
rect 45390 33294 45442 33346
rect 2494 33182 2546 33234
rect 5630 33182 5682 33234
rect 8206 33182 8258 33234
rect 12350 33182 12402 33234
rect 12462 33182 12514 33234
rect 12574 33182 12626 33234
rect 13918 33182 13970 33234
rect 19630 33182 19682 33234
rect 23214 33182 23266 33234
rect 24558 33182 24610 33234
rect 24670 33182 24722 33234
rect 25006 33182 25058 33234
rect 25342 33182 25394 33234
rect 25678 33182 25730 33234
rect 27134 33182 27186 33234
rect 27470 33182 27522 33234
rect 29710 33182 29762 33234
rect 30606 33182 30658 33234
rect 30830 33182 30882 33234
rect 34302 33182 34354 33234
rect 35310 33182 35362 33234
rect 35534 33182 35586 33234
rect 35870 33182 35922 33234
rect 36206 33182 36258 33234
rect 38894 33182 38946 33234
rect 42142 33182 42194 33234
rect 4734 33070 4786 33122
rect 7310 33070 7362 33122
rect 8654 33070 8706 33122
rect 9886 33070 9938 33122
rect 10894 33070 10946 33122
rect 11790 33070 11842 33122
rect 14030 33070 14082 33122
rect 14926 33070 14978 33122
rect 18398 33070 18450 33122
rect 19182 33070 19234 33122
rect 19406 33070 19458 33122
rect 22990 33070 23042 33122
rect 23550 33070 23602 33122
rect 23662 33070 23714 33122
rect 23774 33070 23826 33122
rect 26350 33070 26402 33122
rect 26798 33070 26850 33122
rect 30270 33070 30322 33122
rect 31054 33070 31106 33122
rect 34526 33070 34578 33122
rect 35758 33070 35810 33122
rect 43262 33070 43314 33122
rect 44270 33070 44322 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 2942 32734 2994 32786
rect 4958 32734 5010 32786
rect 7758 32734 7810 32786
rect 9886 32734 9938 32786
rect 11006 32734 11058 32786
rect 22206 32734 22258 32786
rect 22430 32734 22482 32786
rect 23774 32734 23826 32786
rect 25790 32734 25842 32786
rect 27134 32734 27186 32786
rect 29710 32734 29762 32786
rect 38222 32734 38274 32786
rect 38894 32734 38946 32786
rect 39230 32734 39282 32786
rect 39790 32734 39842 32786
rect 39902 32734 39954 32786
rect 40014 32734 40066 32786
rect 41806 32734 41858 32786
rect 43710 32734 43762 32786
rect 44046 32734 44098 32786
rect 45614 32734 45666 32786
rect 45950 32734 46002 32786
rect 46174 32734 46226 32786
rect 46846 32734 46898 32786
rect 5854 32622 5906 32674
rect 5966 32622 6018 32674
rect 8206 32622 8258 32674
rect 8430 32622 8482 32674
rect 10446 32622 10498 32674
rect 10782 32622 10834 32674
rect 11790 32622 11842 32674
rect 14814 32622 14866 32674
rect 15934 32622 15986 32674
rect 16606 32622 16658 32674
rect 17390 32622 17442 32674
rect 19294 32622 19346 32674
rect 23102 32622 23154 32674
rect 23662 32622 23714 32674
rect 26798 32622 26850 32674
rect 36990 32622 37042 32674
rect 38558 32622 38610 32674
rect 40910 32622 40962 32674
rect 45502 32622 45554 32674
rect 47630 32622 47682 32674
rect 47966 32622 48018 32674
rect 5294 32510 5346 32562
rect 5630 32510 5682 32562
rect 7198 32510 7250 32562
rect 8654 32510 8706 32562
rect 13246 32510 13298 32562
rect 13694 32510 13746 32562
rect 16718 32510 16770 32562
rect 17614 32510 17666 32562
rect 18622 32510 18674 32562
rect 22878 32510 22930 32562
rect 24110 32510 24162 32562
rect 25230 32510 25282 32562
rect 28478 32510 28530 32562
rect 29934 32510 29986 32562
rect 33294 32510 33346 32562
rect 33518 32510 33570 32562
rect 37662 32510 37714 32562
rect 40462 32510 40514 32562
rect 41134 32510 41186 32562
rect 41358 32510 41410 32562
rect 41918 32510 41970 32562
rect 42030 32510 42082 32562
rect 42366 32510 42418 32562
rect 46510 32510 46562 32562
rect 47070 32510 47122 32562
rect 2830 32398 2882 32450
rect 3166 32398 3218 32450
rect 3614 32398 3666 32450
rect 4622 32398 4674 32450
rect 6414 32398 6466 32450
rect 8094 32398 8146 32450
rect 10222 32398 10274 32450
rect 11118 32398 11170 32450
rect 13470 32398 13522 32450
rect 18174 32398 18226 32450
rect 21422 32398 21474 32450
rect 22318 32398 22370 32450
rect 25454 32398 25506 32450
rect 28814 32398 28866 32450
rect 31054 32398 31106 32450
rect 33070 32398 33122 32450
rect 34862 32398 34914 32450
rect 41022 32398 41074 32450
rect 42702 32398 42754 32450
rect 42814 32398 42866 32450
rect 45166 32398 45218 32450
rect 46062 32398 46114 32450
rect 9102 32286 9154 32338
rect 15822 32286 15874 32338
rect 16158 32286 16210 32338
rect 16606 32286 16658 32338
rect 23214 32286 23266 32338
rect 24334 32286 24386 32338
rect 24670 32286 24722 32338
rect 29038 32286 29090 32338
rect 29262 32286 29314 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19406 31950 19458 32002
rect 19742 31950 19794 32002
rect 31502 31950 31554 32002
rect 3278 31838 3330 31890
rect 3614 31838 3666 31890
rect 8542 31838 8594 31890
rect 9214 31838 9266 31890
rect 11118 31838 11170 31890
rect 30158 31838 30210 31890
rect 34974 31838 35026 31890
rect 37102 31838 37154 31890
rect 38110 31838 38162 31890
rect 39902 31838 39954 31890
rect 42030 31838 42082 31890
rect 44158 31838 44210 31890
rect 48190 31838 48242 31890
rect 5742 31726 5794 31778
rect 8990 31726 9042 31778
rect 9438 31726 9490 31778
rect 10558 31726 10610 31778
rect 13694 31726 13746 31778
rect 14366 31726 14418 31778
rect 18174 31726 18226 31778
rect 18510 31726 18562 31778
rect 19518 31726 19570 31778
rect 19854 31726 19906 31778
rect 20302 31726 20354 31778
rect 23214 31726 23266 31778
rect 29710 31726 29762 31778
rect 30606 31726 30658 31778
rect 31166 31726 31218 31778
rect 31390 31726 31442 31778
rect 31614 31726 31666 31778
rect 33070 31726 33122 31778
rect 33742 31726 33794 31778
rect 34078 31726 34130 31778
rect 35534 31726 35586 31778
rect 39118 31726 39170 31778
rect 43822 31726 43874 31778
rect 45390 31726 45442 31778
rect 6414 31614 6466 31666
rect 14478 31614 14530 31666
rect 18062 31614 18114 31666
rect 19070 31614 19122 31666
rect 21310 31614 21362 31666
rect 23326 31614 23378 31666
rect 29038 31614 29090 31666
rect 29262 31614 29314 31666
rect 30942 31614 30994 31666
rect 32062 31614 32114 31666
rect 32846 31614 32898 31666
rect 33966 31614 34018 31666
rect 42590 31614 42642 31666
rect 42926 31614 42978 31666
rect 43262 31614 43314 31666
rect 46062 31614 46114 31666
rect 3390 31502 3442 31554
rect 9102 31502 9154 31554
rect 13694 31502 13746 31554
rect 15374 31502 15426 31554
rect 20638 31502 20690 31554
rect 21646 31502 21698 31554
rect 22094 31502 22146 31554
rect 23662 31502 23714 31554
rect 29486 31502 29538 31554
rect 29598 31502 29650 31554
rect 30046 31502 30098 31554
rect 30270 31502 30322 31554
rect 32510 31502 32562 31554
rect 34526 31502 34578 31554
rect 34862 31502 34914 31554
rect 35086 31502 35138 31554
rect 36318 31502 36370 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 7198 31166 7250 31218
rect 8430 31166 8482 31218
rect 12910 31166 12962 31218
rect 15262 31166 15314 31218
rect 15374 31166 15426 31218
rect 15598 31166 15650 31218
rect 22654 31166 22706 31218
rect 24558 31166 24610 31218
rect 26238 31166 26290 31218
rect 27134 31166 27186 31218
rect 29262 31166 29314 31218
rect 30158 31166 30210 31218
rect 30830 31166 30882 31218
rect 37886 31166 37938 31218
rect 44718 31166 44770 31218
rect 45726 31166 45778 31218
rect 46622 31166 46674 31218
rect 47070 31166 47122 31218
rect 47518 31166 47570 31218
rect 48190 31166 48242 31218
rect 7422 31054 7474 31106
rect 8766 31054 8818 31106
rect 8990 31054 9042 31106
rect 13582 31054 13634 31106
rect 13806 31054 13858 31106
rect 15038 31054 15090 31106
rect 15486 31054 15538 31106
rect 21758 31054 21810 31106
rect 21982 31054 22034 31106
rect 23326 31054 23378 31106
rect 23886 31054 23938 31106
rect 27470 31054 27522 31106
rect 35758 31054 35810 31106
rect 35982 31054 36034 31106
rect 36094 31054 36146 31106
rect 36654 31054 36706 31106
rect 36878 31054 36930 31106
rect 37998 31054 38050 31106
rect 45054 31054 45106 31106
rect 45502 31054 45554 31106
rect 46062 31054 46114 31106
rect 1822 30942 1874 30994
rect 7534 30942 7586 30994
rect 11902 30942 11954 30994
rect 13358 30942 13410 30994
rect 16606 30942 16658 30994
rect 17614 30942 17666 30994
rect 18734 30942 18786 30994
rect 20750 30942 20802 30994
rect 20974 30942 21026 30994
rect 21422 30942 21474 30994
rect 22318 30942 22370 30994
rect 22878 30942 22930 30994
rect 23438 30942 23490 30994
rect 24222 30942 24274 30994
rect 24670 30942 24722 30994
rect 26574 30942 26626 30994
rect 27694 30942 27746 30994
rect 29374 30942 29426 30994
rect 29934 30942 29986 30994
rect 30382 30942 30434 30994
rect 31054 30942 31106 30994
rect 37102 30942 37154 30994
rect 37550 30942 37602 30994
rect 45726 30942 45778 30994
rect 2494 30830 2546 30882
rect 4622 30830 4674 30882
rect 8878 30830 8930 30882
rect 10110 30830 10162 30882
rect 14478 30830 14530 30882
rect 16158 30830 16210 30882
rect 23102 30830 23154 30882
rect 24110 30830 24162 30882
rect 26798 30830 26850 30882
rect 30270 30830 30322 30882
rect 36542 30830 36594 30882
rect 16718 30718 16770 30770
rect 18062 30718 18114 30770
rect 22542 30718 22594 30770
rect 29262 30718 29314 30770
rect 29710 30718 29762 30770
rect 36094 30718 36146 30770
rect 37774 30718 37826 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 2718 30382 2770 30434
rect 2830 30382 2882 30434
rect 3054 30382 3106 30434
rect 4622 30382 4674 30434
rect 15038 30382 15090 30434
rect 30382 30382 30434 30434
rect 34190 30382 34242 30434
rect 35646 30382 35698 30434
rect 12686 30270 12738 30322
rect 13918 30270 13970 30322
rect 14926 30270 14978 30322
rect 16046 30270 16098 30322
rect 22318 30270 22370 30322
rect 24446 30270 24498 30322
rect 25342 30270 25394 30322
rect 33294 30270 33346 30322
rect 42142 30270 42194 30322
rect 3278 30158 3330 30210
rect 4846 30158 4898 30210
rect 9886 30158 9938 30210
rect 14702 30158 14754 30210
rect 15934 30158 15986 30210
rect 16942 30158 16994 30210
rect 17614 30158 17666 30210
rect 18062 30158 18114 30210
rect 21646 30158 21698 30210
rect 25118 30158 25170 30210
rect 25678 30158 25730 30210
rect 30494 30158 30546 30210
rect 32510 30158 32562 30210
rect 32846 30158 32898 30210
rect 33742 30158 33794 30210
rect 35310 30158 35362 30210
rect 36990 30158 37042 30210
rect 37214 30158 37266 30210
rect 38782 30158 38834 30210
rect 5966 30046 6018 30098
rect 10558 30046 10610 30098
rect 13806 30046 13858 30098
rect 14030 30046 14082 30098
rect 17950 30046 18002 30098
rect 18398 30046 18450 30098
rect 18734 30046 18786 30098
rect 19070 30046 19122 30098
rect 31502 30046 31554 30098
rect 32174 30046 32226 30098
rect 34638 30046 34690 30098
rect 35870 30046 35922 30098
rect 36094 30046 36146 30098
rect 37662 30046 37714 30098
rect 39454 30046 39506 30098
rect 42254 30046 42306 30098
rect 42478 30046 42530 30098
rect 4286 29934 4338 29986
rect 5630 29934 5682 29986
rect 9438 29934 9490 29986
rect 17278 29934 17330 29986
rect 18510 29934 18562 29986
rect 19182 29934 19234 29986
rect 19406 29934 19458 29986
rect 19742 29934 19794 29986
rect 26238 29934 26290 29986
rect 26574 29934 26626 29986
rect 30382 29934 30434 29986
rect 31838 29934 31890 29986
rect 35982 29934 36034 29986
rect 37326 29934 37378 29986
rect 37438 29934 37490 29986
rect 41694 29934 41746 29986
rect 44158 29934 44210 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 10334 29598 10386 29650
rect 12686 29598 12738 29650
rect 13582 29598 13634 29650
rect 14814 29598 14866 29650
rect 15598 29598 15650 29650
rect 17950 29598 18002 29650
rect 32174 29598 32226 29650
rect 33070 29598 33122 29650
rect 34526 29598 34578 29650
rect 34862 29598 34914 29650
rect 38558 29598 38610 29650
rect 44046 29598 44098 29650
rect 11454 29486 11506 29538
rect 16158 29486 16210 29538
rect 17502 29486 17554 29538
rect 18846 29486 18898 29538
rect 20862 29486 20914 29538
rect 27470 29486 27522 29538
rect 35646 29486 35698 29538
rect 38334 29486 38386 29538
rect 41134 29486 41186 29538
rect 42478 29486 42530 29538
rect 2830 29374 2882 29426
rect 10222 29374 10274 29426
rect 10446 29374 10498 29426
rect 11230 29374 11282 29426
rect 15262 29374 15314 29426
rect 15374 29374 15426 29426
rect 15822 29374 15874 29426
rect 16494 29374 16546 29426
rect 18062 29374 18114 29426
rect 18286 29374 18338 29426
rect 18622 29374 18674 29426
rect 19518 29374 19570 29426
rect 19630 29374 19682 29426
rect 19854 29374 19906 29426
rect 20302 29374 20354 29426
rect 20526 29374 20578 29426
rect 26798 29374 26850 29426
rect 32286 29374 32338 29426
rect 36094 29374 36146 29426
rect 36766 29374 36818 29426
rect 38222 29374 38274 29426
rect 38894 29374 38946 29426
rect 41470 29374 41522 29426
rect 42590 29374 42642 29426
rect 42702 29374 42754 29426
rect 43710 29374 43762 29426
rect 44382 29374 44434 29426
rect 44606 29374 44658 29426
rect 45390 29374 45442 29426
rect 2606 29262 2658 29314
rect 3278 29262 3330 29314
rect 10670 29262 10722 29314
rect 11902 29262 11954 29314
rect 13918 29262 13970 29314
rect 14366 29262 14418 29314
rect 15486 29262 15538 29314
rect 18846 29262 18898 29314
rect 19294 29262 19346 29314
rect 21310 29262 21362 29314
rect 29598 29262 29650 29314
rect 33182 29262 33234 29314
rect 37102 29262 37154 29314
rect 40350 29262 40402 29314
rect 43486 29262 43538 29314
rect 44942 29262 44994 29314
rect 46062 29262 46114 29314
rect 48190 29262 48242 29314
rect 2494 29150 2546 29202
rect 5854 29150 5906 29202
rect 5966 29150 6018 29202
rect 6190 29150 6242 29202
rect 6302 29150 6354 29202
rect 17390 29150 17442 29202
rect 32174 29150 32226 29202
rect 36878 29150 36930 29202
rect 41246 29150 41298 29202
rect 41582 29150 41634 29202
rect 42030 29150 42082 29202
rect 44830 29150 44882 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 2494 28814 2546 28866
rect 6638 28814 6690 28866
rect 9886 28814 9938 28866
rect 13582 28814 13634 28866
rect 14926 28814 14978 28866
rect 17838 28814 17890 28866
rect 43822 28814 43874 28866
rect 44158 28814 44210 28866
rect 2942 28702 2994 28754
rect 3726 28702 3778 28754
rect 9774 28702 9826 28754
rect 12574 28702 12626 28754
rect 16382 28702 16434 28754
rect 22094 28702 22146 28754
rect 32062 28702 32114 28754
rect 45726 28702 45778 28754
rect 3054 28590 3106 28642
rect 4174 28590 4226 28642
rect 4398 28590 4450 28642
rect 4622 28590 4674 28642
rect 4846 28590 4898 28642
rect 5070 28590 5122 28642
rect 5630 28590 5682 28642
rect 5966 28590 6018 28642
rect 6414 28590 6466 28642
rect 7198 28590 7250 28642
rect 7646 28590 7698 28642
rect 8654 28590 8706 28642
rect 8878 28590 8930 28642
rect 9662 28590 9714 28642
rect 12350 28590 12402 28642
rect 15038 28590 15090 28642
rect 16830 28590 16882 28642
rect 17390 28590 17442 28642
rect 18734 28590 18786 28642
rect 19070 28590 19122 28642
rect 19406 28590 19458 28642
rect 24334 28590 24386 28642
rect 29150 28590 29202 28642
rect 37102 28590 37154 28642
rect 37438 28590 37490 28642
rect 37998 28590 38050 28642
rect 39566 28590 39618 28642
rect 41694 28590 41746 28642
rect 44830 28590 44882 28642
rect 45278 28590 45330 28642
rect 46174 28590 46226 28642
rect 5742 28478 5794 28530
rect 11678 28478 11730 28530
rect 13694 28478 13746 28530
rect 21422 28478 21474 28530
rect 21534 28478 21586 28530
rect 24222 28478 24274 28530
rect 29934 28478 29986 28530
rect 38670 28478 38722 28530
rect 39006 28478 39058 28530
rect 41470 28478 41522 28530
rect 44046 28478 44098 28530
rect 21758 28366 21810 28418
rect 23998 28366 24050 28418
rect 39454 28366 39506 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 9998 28030 10050 28082
rect 14030 28030 14082 28082
rect 16046 28030 16098 28082
rect 23774 28030 23826 28082
rect 24110 28030 24162 28082
rect 32398 28030 32450 28082
rect 37550 28030 37602 28082
rect 37998 28030 38050 28082
rect 38222 28030 38274 28082
rect 43486 28030 43538 28082
rect 2494 27918 2546 27970
rect 6638 27918 6690 27970
rect 9774 27918 9826 27970
rect 10222 27918 10274 27970
rect 11790 27918 11842 27970
rect 12014 27918 12066 27970
rect 15822 27918 15874 27970
rect 18286 27918 18338 27970
rect 18510 27918 18562 27970
rect 22206 27918 22258 27970
rect 23438 27918 23490 27970
rect 29934 27918 29986 27970
rect 33854 27918 33906 27970
rect 37438 27918 37490 27970
rect 37886 27918 37938 27970
rect 40014 27918 40066 27970
rect 40126 27918 40178 27970
rect 41358 27918 41410 27970
rect 44830 27918 44882 27970
rect 1822 27806 1874 27858
rect 5854 27806 5906 27858
rect 9550 27806 9602 27858
rect 9886 27806 9938 27858
rect 10446 27806 10498 27858
rect 10782 27806 10834 27858
rect 11006 27806 11058 27858
rect 13694 27806 13746 27858
rect 15374 27806 15426 27858
rect 15598 27806 15650 27858
rect 17950 27806 18002 27858
rect 18734 27806 18786 27858
rect 19070 27806 19122 27858
rect 19518 27806 19570 27858
rect 22878 27806 22930 27858
rect 25342 27806 25394 27858
rect 28926 27806 28978 27858
rect 32510 27806 32562 27858
rect 33070 27806 33122 27858
rect 39118 27806 39170 27858
rect 39342 27806 39394 27858
rect 41470 27806 41522 27858
rect 43822 27806 43874 27858
rect 44270 27806 44322 27858
rect 45390 27806 45442 27858
rect 4622 27694 4674 27746
rect 8766 27694 8818 27746
rect 10670 27694 10722 27746
rect 12462 27694 12514 27746
rect 15934 27694 15986 27746
rect 20078 27694 20130 27746
rect 24558 27694 24610 27746
rect 26014 27694 26066 27746
rect 28142 27694 28194 27746
rect 29150 27694 29202 27746
rect 30382 27694 30434 27746
rect 30830 27694 30882 27746
rect 31390 27694 31442 27746
rect 35982 27694 36034 27746
rect 39566 27694 39618 27746
rect 44382 27694 44434 27746
rect 46062 27694 46114 27746
rect 48190 27694 48242 27746
rect 11678 27582 11730 27634
rect 17726 27582 17778 27634
rect 28590 27582 28642 27634
rect 30046 27582 30098 27634
rect 30270 27582 30322 27634
rect 31166 27582 31218 27634
rect 32062 27582 32114 27634
rect 32286 27582 32338 27634
rect 38670 27582 38722 27634
rect 40126 27582 40178 27634
rect 41358 27582 41410 27634
rect 44046 27582 44098 27634
rect 44718 27582 44770 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 9662 27246 9714 27298
rect 26014 27246 26066 27298
rect 30494 27246 30546 27298
rect 32734 27246 32786 27298
rect 43038 27246 43090 27298
rect 45166 27246 45218 27298
rect 7646 27134 7698 27186
rect 9102 27134 9154 27186
rect 9438 27134 9490 27186
rect 10782 27134 10834 27186
rect 12910 27134 12962 27186
rect 24894 27134 24946 27186
rect 25342 27134 25394 27186
rect 25902 27134 25954 27186
rect 30270 27134 30322 27186
rect 42590 27134 42642 27186
rect 43598 27134 43650 27186
rect 44046 27134 44098 27186
rect 44830 27134 44882 27186
rect 47854 27134 47906 27186
rect 10110 27022 10162 27074
rect 13806 27022 13858 27074
rect 14254 27022 14306 27074
rect 14814 27022 14866 27074
rect 15822 27022 15874 27074
rect 16270 27022 16322 27074
rect 17614 27022 17666 27074
rect 18398 27022 18450 27074
rect 21870 27022 21922 27074
rect 22542 27022 22594 27074
rect 23214 27022 23266 27074
rect 23662 27022 23714 27074
rect 24110 27022 24162 27074
rect 29598 27022 29650 27074
rect 30158 27022 30210 27074
rect 31614 27022 31666 27074
rect 35870 27022 35922 27074
rect 36430 27022 36482 27074
rect 38558 27022 38610 27074
rect 39902 27022 39954 27074
rect 40910 27022 40962 27074
rect 42254 27022 42306 27074
rect 42814 27022 42866 27074
rect 43374 27022 43426 27074
rect 43934 27022 43986 27074
rect 46062 27022 46114 27074
rect 8990 26910 9042 26962
rect 9214 26910 9266 26962
rect 13470 26910 13522 26962
rect 15374 26910 15426 26962
rect 16494 26910 16546 26962
rect 17278 26910 17330 26962
rect 24446 26910 24498 26962
rect 25790 26910 25842 26962
rect 32846 26910 32898 26962
rect 33070 26910 33122 26962
rect 41470 26910 41522 26962
rect 42366 26910 42418 26962
rect 44158 26910 44210 26962
rect 44942 26910 44994 26962
rect 15150 26798 15202 26850
rect 16606 26798 16658 26850
rect 18398 26798 18450 26850
rect 22094 26798 22146 26850
rect 40574 26798 40626 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 7422 26462 7474 26514
rect 17838 26462 17890 26514
rect 22430 26462 22482 26514
rect 22990 26462 23042 26514
rect 33070 26462 33122 26514
rect 35422 26462 35474 26514
rect 39230 26462 39282 26514
rect 48078 26462 48130 26514
rect 7086 26350 7138 26402
rect 8094 26350 8146 26402
rect 15486 26350 15538 26402
rect 26462 26350 26514 26402
rect 33630 26350 33682 26402
rect 35870 26350 35922 26402
rect 44270 26350 44322 26402
rect 4846 26238 4898 26290
rect 5070 26238 5122 26290
rect 5294 26238 5346 26290
rect 5966 26238 6018 26290
rect 15262 26238 15314 26290
rect 15934 26238 15986 26290
rect 16718 26238 16770 26290
rect 17390 26238 17442 26290
rect 17614 26238 17666 26290
rect 17726 26238 17778 26290
rect 17950 26238 18002 26290
rect 18622 26238 18674 26290
rect 18846 26238 18898 26290
rect 19182 26238 19234 26290
rect 19518 26238 19570 26290
rect 26238 26238 26290 26290
rect 32174 26238 32226 26290
rect 32510 26238 32562 26290
rect 33518 26238 33570 26290
rect 33854 26238 33906 26290
rect 36878 26238 36930 26290
rect 38446 26238 38498 26290
rect 39006 26238 39058 26290
rect 39342 26238 39394 26290
rect 39566 26238 39618 26290
rect 39790 26238 39842 26290
rect 39902 26238 39954 26290
rect 41246 26238 41298 26290
rect 41582 26238 41634 26290
rect 42254 26238 42306 26290
rect 42590 26238 42642 26290
rect 42926 26238 42978 26290
rect 43150 26238 43202 26290
rect 45166 26238 45218 26290
rect 6190 26126 6242 26178
rect 8654 26126 8706 26178
rect 20526 26126 20578 26178
rect 21870 26126 21922 26178
rect 43934 26126 43986 26178
rect 45838 26126 45890 26178
rect 4734 26014 4786 26066
rect 5630 26014 5682 26066
rect 7870 26014 7922 26066
rect 8206 26014 8258 26066
rect 15486 26014 15538 26066
rect 19742 26014 19794 26066
rect 19966 26014 20018 26066
rect 20078 26014 20130 26066
rect 32510 26014 32562 26066
rect 42142 26014 42194 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 5630 25678 5682 25730
rect 5966 25678 6018 25730
rect 15262 25678 15314 25730
rect 32622 25678 32674 25730
rect 32958 25678 33010 25730
rect 2494 25566 2546 25618
rect 4622 25566 4674 25618
rect 8430 25566 8482 25618
rect 10558 25566 10610 25618
rect 19182 25566 19234 25618
rect 24670 25566 24722 25618
rect 26462 25566 26514 25618
rect 28590 25566 28642 25618
rect 32062 25566 32114 25618
rect 32398 25566 32450 25618
rect 36430 25566 36482 25618
rect 39118 25566 39170 25618
rect 45614 25566 45666 25618
rect 1822 25454 1874 25506
rect 7758 25454 7810 25506
rect 11342 25454 11394 25506
rect 11566 25454 11618 25506
rect 11790 25454 11842 25506
rect 14926 25454 14978 25506
rect 15710 25454 15762 25506
rect 16494 25454 16546 25506
rect 16942 25454 16994 25506
rect 17726 25454 17778 25506
rect 25006 25454 25058 25506
rect 25678 25454 25730 25506
rect 29262 25454 29314 25506
rect 33630 25454 33682 25506
rect 37326 25454 37378 25506
rect 38110 25454 38162 25506
rect 38446 25454 38498 25506
rect 39230 25454 39282 25506
rect 41582 25454 41634 25506
rect 41806 25454 41858 25506
rect 43262 25454 43314 25506
rect 43598 25454 43650 25506
rect 44158 25454 44210 25506
rect 45278 25454 45330 25506
rect 45726 25454 45778 25506
rect 5742 25342 5794 25394
rect 6638 25342 6690 25394
rect 16046 25342 16098 25394
rect 17950 25342 18002 25394
rect 22766 25342 22818 25394
rect 29934 25342 29986 25394
rect 34302 25342 34354 25394
rect 38782 25342 38834 25394
rect 41918 25342 41970 25394
rect 45838 25342 45890 25394
rect 46958 25342 47010 25394
rect 47518 25342 47570 25394
rect 48190 25342 48242 25394
rect 6302 25230 6354 25282
rect 11230 25230 11282 25282
rect 11454 25230 11506 25282
rect 15150 25230 15202 25282
rect 16382 25230 16434 25282
rect 23102 25230 23154 25282
rect 25342 25230 25394 25282
rect 36990 25230 37042 25282
rect 44158 25230 44210 25282
rect 45054 25230 45106 25282
rect 47182 25230 47234 25282
rect 47854 25230 47906 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 9550 24894 9602 24946
rect 14702 24894 14754 24946
rect 18622 24894 18674 24946
rect 22094 24894 22146 24946
rect 38110 24894 38162 24946
rect 38222 24894 38274 24946
rect 38894 24894 38946 24946
rect 41134 24894 41186 24946
rect 41358 24894 41410 24946
rect 42030 24894 42082 24946
rect 42254 24894 42306 24946
rect 43710 24894 43762 24946
rect 46398 24894 46450 24946
rect 47182 24894 47234 24946
rect 5966 24782 6018 24834
rect 6750 24782 6802 24834
rect 20862 24782 20914 24834
rect 22654 24782 22706 24834
rect 29822 24782 29874 24834
rect 30942 24782 30994 24834
rect 33854 24782 33906 24834
rect 37438 24782 37490 24834
rect 37550 24782 37602 24834
rect 37774 24782 37826 24834
rect 39342 24782 39394 24834
rect 42926 24782 42978 24834
rect 45614 24782 45666 24834
rect 47630 24782 47682 24834
rect 4174 24670 4226 24722
rect 6302 24670 6354 24722
rect 6862 24670 6914 24722
rect 9886 24670 9938 24722
rect 11118 24670 11170 24722
rect 14366 24670 14418 24722
rect 15038 24670 15090 24722
rect 15486 24670 15538 24722
rect 16158 24670 16210 24722
rect 21646 24670 21698 24722
rect 22318 24670 22370 24722
rect 22878 24670 22930 24722
rect 24670 24670 24722 24722
rect 25230 24670 25282 24722
rect 31054 24670 31106 24722
rect 31390 24670 31442 24722
rect 31838 24670 31890 24722
rect 33294 24670 33346 24722
rect 33742 24670 33794 24722
rect 38782 24670 38834 24722
rect 39230 24670 39282 24722
rect 40910 24670 40962 24722
rect 41582 24670 41634 24722
rect 42478 24670 42530 24722
rect 43374 24670 43426 24722
rect 43822 24670 43874 24722
rect 45838 24670 45890 24722
rect 45950 24670 46002 24722
rect 46174 24670 46226 24722
rect 46510 24670 46562 24722
rect 46846 24670 46898 24722
rect 47294 24670 47346 24722
rect 47406 24670 47458 24722
rect 5630 24558 5682 24610
rect 10334 24558 10386 24610
rect 11902 24558 11954 24610
rect 14030 24558 14082 24610
rect 16382 24558 16434 24610
rect 23102 24558 23154 24610
rect 23550 24558 23602 24610
rect 41022 24558 41074 24610
rect 48190 24558 48242 24610
rect 1934 24446 1986 24498
rect 15486 24446 15538 24498
rect 31278 24446 31330 24498
rect 31838 24446 31890 24498
rect 32174 24446 32226 24498
rect 33518 24446 33570 24498
rect 38334 24446 38386 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 11902 24110 11954 24162
rect 26238 24110 26290 24162
rect 42926 24110 42978 24162
rect 4622 23998 4674 24050
rect 7870 23998 7922 24050
rect 22878 23998 22930 24050
rect 25006 23998 25058 24050
rect 29934 23998 29986 24050
rect 41134 23998 41186 24050
rect 42030 23998 42082 24050
rect 1822 23886 1874 23938
rect 5070 23886 5122 23938
rect 5854 23886 5906 23938
rect 6974 23886 7026 23938
rect 7198 23886 7250 23938
rect 12574 23886 12626 23938
rect 15934 23886 15986 23938
rect 19854 23886 19906 23938
rect 20414 23886 20466 23938
rect 22094 23886 22146 23938
rect 25454 23886 25506 23938
rect 25678 23886 25730 23938
rect 26686 23886 26738 23938
rect 28366 23886 28418 23938
rect 29710 23886 29762 23938
rect 33518 23886 33570 23938
rect 33742 23886 33794 23938
rect 41582 23886 41634 23938
rect 42478 23886 42530 23938
rect 45278 23886 45330 23938
rect 46510 23886 46562 23938
rect 46734 23886 46786 23938
rect 47182 23886 47234 23938
rect 47742 23886 47794 23938
rect 48078 23886 48130 23938
rect 2494 23774 2546 23826
rect 5742 23774 5794 23826
rect 8318 23774 8370 23826
rect 12014 23774 12066 23826
rect 25790 23774 25842 23826
rect 28590 23774 28642 23826
rect 29150 23774 29202 23826
rect 33294 23774 33346 23826
rect 43038 23774 43090 23826
rect 46174 23774 46226 23826
rect 5518 23662 5570 23714
rect 8206 23662 8258 23714
rect 12350 23662 12402 23714
rect 15598 23662 15650 23714
rect 18398 23662 18450 23714
rect 19630 23662 19682 23714
rect 33518 23662 33570 23714
rect 38110 23662 38162 23714
rect 45838 23662 45890 23714
rect 46286 23662 46338 23714
rect 47070 23662 47122 23714
rect 47294 23662 47346 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 3614 23326 3666 23378
rect 18062 23326 18114 23378
rect 18846 23326 18898 23378
rect 19294 23326 19346 23378
rect 29934 23326 29986 23378
rect 30718 23326 30770 23378
rect 38334 23326 38386 23378
rect 39342 23326 39394 23378
rect 44942 23326 44994 23378
rect 2046 23214 2098 23266
rect 2942 23214 2994 23266
rect 6414 23214 6466 23266
rect 17838 23214 17890 23266
rect 18510 23214 18562 23266
rect 31614 23214 31666 23266
rect 33518 23214 33570 23266
rect 39230 23214 39282 23266
rect 43710 23214 43762 23266
rect 44830 23214 44882 23266
rect 46062 23214 46114 23266
rect 1710 23102 1762 23154
rect 5294 23102 5346 23154
rect 5518 23102 5570 23154
rect 8878 23102 8930 23154
rect 11342 23102 11394 23154
rect 13918 23102 13970 23154
rect 20526 23102 20578 23154
rect 25342 23102 25394 23154
rect 31166 23102 31218 23154
rect 31390 23102 31442 23154
rect 33630 23102 33682 23154
rect 33854 23102 33906 23154
rect 34974 23102 35026 23154
rect 38222 23102 38274 23154
rect 38446 23102 38498 23154
rect 38670 23102 38722 23154
rect 42478 23102 42530 23154
rect 42926 23102 42978 23154
rect 43598 23102 43650 23154
rect 45278 23102 45330 23154
rect 2494 22990 2546 23042
rect 2830 22990 2882 23042
rect 3166 22990 3218 23042
rect 4622 22990 4674 23042
rect 8766 22990 8818 23042
rect 10558 22990 10610 23042
rect 10894 22990 10946 23042
rect 11902 22990 11954 23042
rect 12350 22990 12402 23042
rect 12798 22990 12850 23042
rect 13582 22990 13634 23042
rect 14702 22990 14754 23042
rect 16830 22990 16882 23042
rect 21198 22990 21250 23042
rect 23326 22990 23378 23042
rect 26014 22990 26066 23042
rect 28142 22990 28194 23042
rect 30494 22990 30546 23042
rect 31726 22990 31778 23042
rect 35646 22990 35698 23042
rect 37774 22990 37826 23042
rect 42254 22990 42306 23042
rect 44494 22990 44546 23042
rect 48190 22990 48242 23042
rect 6526 22878 6578 22930
rect 8542 22878 8594 22930
rect 11790 22878 11842 22930
rect 18174 22878 18226 22930
rect 30270 22878 30322 22930
rect 33070 22878 33122 22930
rect 38894 22878 38946 22930
rect 39342 22878 39394 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 31614 22542 31666 22594
rect 31950 22542 32002 22594
rect 34302 22542 34354 22594
rect 34638 22542 34690 22594
rect 47966 22542 48018 22594
rect 4622 22430 4674 22482
rect 11118 22430 11170 22482
rect 12462 22430 12514 22482
rect 14478 22430 14530 22482
rect 18286 22430 18338 22482
rect 22654 22430 22706 22482
rect 24446 22430 24498 22482
rect 25678 22430 25730 22482
rect 26910 22430 26962 22482
rect 31390 22430 31442 22482
rect 34414 22430 34466 22482
rect 35086 22430 35138 22482
rect 42590 22430 42642 22482
rect 44830 22430 44882 22482
rect 1822 22318 1874 22370
rect 8206 22318 8258 22370
rect 12126 22318 12178 22370
rect 14030 22318 14082 22370
rect 17614 22318 17666 22370
rect 22318 22318 22370 22370
rect 22542 22318 22594 22370
rect 22878 22318 22930 22370
rect 22990 22318 23042 22370
rect 23102 22318 23154 22370
rect 24782 22318 24834 22370
rect 25454 22318 25506 22370
rect 27246 22318 27298 22370
rect 28030 22318 28082 22370
rect 30158 22318 30210 22370
rect 33406 22318 33458 22370
rect 33854 22318 33906 22370
rect 34750 22318 34802 22370
rect 37998 22318 38050 22370
rect 38782 22318 38834 22370
rect 39678 22318 39730 22370
rect 43150 22318 43202 22370
rect 45838 22318 45890 22370
rect 2494 22206 2546 22258
rect 6190 22206 6242 22258
rect 8990 22206 9042 22258
rect 12350 22206 12402 22258
rect 12686 22206 12738 22258
rect 12910 22206 12962 22258
rect 13582 22206 13634 22258
rect 13918 22206 13970 22258
rect 21982 22206 22034 22258
rect 23774 22206 23826 22258
rect 25790 22206 25842 22258
rect 26574 22206 26626 22258
rect 30494 22206 30546 22258
rect 33182 22206 33234 22258
rect 33294 22206 33346 22258
rect 35310 22206 35362 22258
rect 37774 22206 37826 22258
rect 38446 22206 38498 22258
rect 40462 22206 40514 22258
rect 43038 22206 43090 22258
rect 45166 22206 45218 22258
rect 5070 22094 5122 22146
rect 6302 22094 6354 22146
rect 11454 22094 11506 22146
rect 11566 22094 11618 22146
rect 11678 22094 11730 22146
rect 13806 22094 13858 22146
rect 20526 22094 20578 22146
rect 22094 22094 22146 22146
rect 23662 22094 23714 22146
rect 25118 22094 25170 22146
rect 28254 22094 28306 22146
rect 35198 22094 35250 22146
rect 38558 22094 38610 22146
rect 42814 22094 42866 22146
rect 43598 22094 43650 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 8318 21758 8370 21810
rect 8654 21758 8706 21810
rect 10334 21758 10386 21810
rect 11006 21758 11058 21810
rect 12462 21758 12514 21810
rect 24558 21758 24610 21810
rect 27806 21758 27858 21810
rect 38894 21758 38946 21810
rect 41022 21758 41074 21810
rect 42030 21758 42082 21810
rect 6862 21646 6914 21698
rect 7198 21646 7250 21698
rect 7534 21646 7586 21698
rect 12014 21646 12066 21698
rect 12574 21646 12626 21698
rect 17390 21646 17442 21698
rect 27918 21646 27970 21698
rect 41246 21646 41298 21698
rect 4286 21534 4338 21586
rect 5742 21534 5794 21586
rect 8430 21534 8482 21586
rect 8878 21534 8930 21586
rect 10670 21534 10722 21586
rect 11566 21534 11618 21586
rect 11678 21534 11730 21586
rect 11902 21534 11954 21586
rect 15150 21534 15202 21586
rect 17838 21534 17890 21586
rect 19294 21534 19346 21586
rect 31390 21534 31442 21586
rect 32062 21534 32114 21586
rect 33966 21534 34018 21586
rect 34190 21534 34242 21586
rect 34414 21534 34466 21586
rect 38782 21534 38834 21586
rect 39006 21534 39058 21586
rect 39454 21534 39506 21586
rect 41806 21534 41858 21586
rect 42366 21534 42418 21586
rect 43822 21534 43874 21586
rect 45054 21534 45106 21586
rect 46062 21534 46114 21586
rect 1934 21422 1986 21474
rect 5966 21422 6018 21474
rect 8542 21422 8594 21474
rect 13134 21422 13186 21474
rect 14926 21422 14978 21474
rect 18286 21422 18338 21474
rect 23662 21422 23714 21474
rect 31166 21422 31218 21474
rect 31838 21422 31890 21474
rect 39230 21422 39282 21474
rect 40350 21422 40402 21474
rect 40910 21422 40962 21474
rect 41918 21422 41970 21474
rect 44046 21422 44098 21474
rect 45166 21422 45218 21474
rect 5406 21310 5458 21362
rect 6414 21310 6466 21362
rect 6526 21310 6578 21362
rect 6750 21310 6802 21362
rect 14814 21310 14866 21362
rect 18734 21310 18786 21362
rect 18846 21310 18898 21362
rect 19070 21310 19122 21362
rect 30830 21310 30882 21362
rect 30942 21310 30994 21362
rect 31726 21310 31778 21362
rect 34526 21310 34578 21362
rect 43934 21310 43986 21362
rect 47966 21310 48018 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 4622 20974 4674 21026
rect 4958 20974 5010 21026
rect 14366 20974 14418 21026
rect 14590 20974 14642 21026
rect 21310 20974 21362 21026
rect 22206 20974 22258 21026
rect 2494 20862 2546 20914
rect 10222 20862 10274 20914
rect 14702 20862 14754 20914
rect 15710 20862 15762 20914
rect 37662 20862 37714 20914
rect 37774 20862 37826 20914
rect 38782 20862 38834 20914
rect 41806 20862 41858 20914
rect 43598 20862 43650 20914
rect 48190 20862 48242 20914
rect 1710 20750 1762 20802
rect 3278 20750 3330 20802
rect 3726 20750 3778 20802
rect 4846 20750 4898 20802
rect 5966 20750 6018 20802
rect 7982 20750 8034 20802
rect 15150 20750 15202 20802
rect 15374 20750 15426 20802
rect 16158 20750 16210 20802
rect 17838 20750 17890 20802
rect 19630 20750 19682 20802
rect 19854 20750 19906 20802
rect 19966 20750 20018 20802
rect 20190 20750 20242 20802
rect 22990 20750 23042 20802
rect 23438 20750 23490 20802
rect 23662 20750 23714 20802
rect 24558 20750 24610 20802
rect 24894 20750 24946 20802
rect 29934 20750 29986 20802
rect 30382 20750 30434 20802
rect 30494 20750 30546 20802
rect 30718 20750 30770 20802
rect 31166 20750 31218 20802
rect 37102 20750 37154 20802
rect 38446 20750 38498 20802
rect 38670 20750 38722 20802
rect 39118 20750 39170 20802
rect 39566 20750 39618 20802
rect 40014 20750 40066 20802
rect 40126 20750 40178 20802
rect 40798 20750 40850 20802
rect 41694 20750 41746 20802
rect 42366 20750 42418 20802
rect 42814 20750 42866 20802
rect 43710 20750 43762 20802
rect 43934 20750 43986 20802
rect 45278 20750 45330 20802
rect 2046 20638 2098 20690
rect 2830 20638 2882 20690
rect 4510 20638 4562 20690
rect 6078 20638 6130 20690
rect 8542 20638 8594 20690
rect 14254 20638 14306 20690
rect 16718 20638 16770 20690
rect 17726 20638 17778 20690
rect 19518 20638 19570 20690
rect 21422 20638 21474 20690
rect 22094 20638 22146 20690
rect 23998 20638 24050 20690
rect 25230 20638 25282 20690
rect 29262 20638 29314 20690
rect 29374 20638 29426 20690
rect 29486 20638 29538 20690
rect 30830 20638 30882 20690
rect 36990 20638 37042 20690
rect 38110 20638 38162 20690
rect 38222 20638 38274 20690
rect 39342 20638 39394 20690
rect 39790 20638 39842 20690
rect 40686 20638 40738 20690
rect 41806 20638 41858 20690
rect 43486 20638 43538 20690
rect 44830 20638 44882 20690
rect 46062 20638 46114 20690
rect 6974 20526 7026 20578
rect 10110 20526 10162 20578
rect 11118 20526 11170 20578
rect 22206 20526 22258 20578
rect 23326 20526 23378 20578
rect 23886 20526 23938 20578
rect 24894 20526 24946 20578
rect 31278 20526 31330 20578
rect 31390 20526 31442 20578
rect 38894 20526 38946 20578
rect 40462 20526 40514 20578
rect 44942 20526 44994 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 6414 20190 6466 20242
rect 16830 20190 16882 20242
rect 30382 20190 30434 20242
rect 39118 20190 39170 20242
rect 39230 20190 39282 20242
rect 46846 20190 46898 20242
rect 5630 20078 5682 20130
rect 5742 20078 5794 20130
rect 5854 20078 5906 20130
rect 6190 20078 6242 20130
rect 6750 20078 6802 20130
rect 8654 20078 8706 20130
rect 9886 20078 9938 20130
rect 10782 20078 10834 20130
rect 12910 20078 12962 20130
rect 18846 20078 18898 20130
rect 23102 20078 23154 20130
rect 24670 20078 24722 20130
rect 34750 20078 34802 20130
rect 37662 20078 37714 20130
rect 41806 20078 41858 20130
rect 44270 20078 44322 20130
rect 47854 20078 47906 20130
rect 1822 19966 1874 20018
rect 6526 19966 6578 20018
rect 8542 19966 8594 20018
rect 8878 19966 8930 20018
rect 9102 19966 9154 20018
rect 10334 19966 10386 20018
rect 10558 19966 10610 20018
rect 11006 19966 11058 20018
rect 12126 19966 12178 20018
rect 15486 19966 15538 20018
rect 18062 19966 18114 20018
rect 22318 19966 22370 20018
rect 22542 19966 22594 20018
rect 22990 19966 23042 20018
rect 24110 19966 24162 20018
rect 25230 19966 25282 20018
rect 29038 19966 29090 20018
rect 29486 19966 29538 20018
rect 29598 19966 29650 20018
rect 29710 19966 29762 20018
rect 30046 19966 30098 20018
rect 30382 19966 30434 20018
rect 30718 19966 30770 20018
rect 31166 19966 31218 20018
rect 31390 19966 31442 20018
rect 31614 19966 31666 20018
rect 33966 19966 34018 20018
rect 37102 19966 37154 20018
rect 37438 19966 37490 20018
rect 39006 19966 39058 20018
rect 43262 19966 43314 20018
rect 43822 19966 43874 20018
rect 45950 19966 46002 20018
rect 46622 19966 46674 20018
rect 46958 19966 47010 20018
rect 47182 19966 47234 20018
rect 48078 19966 48130 20018
rect 2494 19854 2546 19906
rect 4622 19854 4674 19906
rect 5070 19854 5122 19906
rect 11118 19854 11170 19906
rect 15038 19854 15090 19906
rect 16718 19854 16770 19906
rect 20974 19854 21026 19906
rect 21646 19854 21698 19906
rect 24334 19854 24386 19906
rect 26014 19854 26066 19906
rect 28142 19854 28194 19906
rect 36878 19854 36930 19906
rect 37326 19854 37378 19906
rect 43598 19854 43650 19906
rect 46398 19854 46450 19906
rect 9662 19742 9714 19794
rect 9998 19742 10050 19794
rect 28814 19742 28866 19794
rect 31054 19742 31106 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 2718 19406 2770 19458
rect 3054 19406 3106 19458
rect 8990 19406 9042 19458
rect 9214 19406 9266 19458
rect 11006 19406 11058 19458
rect 11230 19406 11282 19458
rect 20302 19406 20354 19458
rect 25454 19406 25506 19458
rect 25678 19406 25730 19458
rect 3502 19294 3554 19346
rect 12126 19294 12178 19346
rect 15150 19294 15202 19346
rect 17166 19294 17218 19346
rect 19630 19294 19682 19346
rect 31950 19294 32002 19346
rect 34078 19294 34130 19346
rect 39902 19294 39954 19346
rect 42926 19294 42978 19346
rect 43934 19294 43986 19346
rect 44270 19294 44322 19346
rect 44942 19294 44994 19346
rect 46734 19294 46786 19346
rect 5630 19182 5682 19234
rect 8654 19182 8706 19234
rect 9774 19182 9826 19234
rect 10558 19182 10610 19234
rect 12238 19182 12290 19234
rect 13806 19182 13858 19234
rect 13918 19182 13970 19234
rect 14702 19182 14754 19234
rect 19966 19182 20018 19234
rect 25902 19182 25954 19234
rect 27134 19182 27186 19234
rect 30158 19182 30210 19234
rect 30382 19182 30434 19234
rect 31166 19182 31218 19234
rect 38782 19182 38834 19234
rect 42030 19182 42082 19234
rect 43038 19182 43090 19234
rect 45054 19182 45106 19234
rect 46174 19182 46226 19234
rect 47294 19182 47346 19234
rect 2830 19070 2882 19122
rect 10446 19070 10498 19122
rect 11678 19070 11730 19122
rect 11902 19070 11954 19122
rect 26910 19070 26962 19122
rect 29934 19070 29986 19122
rect 42702 19070 42754 19122
rect 45166 19070 45218 19122
rect 5742 18958 5794 19010
rect 8318 18958 8370 19010
rect 8430 18958 8482 19010
rect 8542 18958 8594 19010
rect 9886 18958 9938 19010
rect 10110 18958 10162 19010
rect 11342 18958 11394 19010
rect 17054 18958 17106 19010
rect 20190 18958 20242 19010
rect 25790 18958 25842 19010
rect 30158 18958 30210 19010
rect 37102 18958 37154 19010
rect 38446 18958 38498 19010
rect 41918 18958 41970 19010
rect 46062 18958 46114 19010
rect 46622 18958 46674 19010
rect 46846 18958 46898 19010
rect 47518 18958 47570 19010
rect 47854 18958 47906 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 6974 18622 7026 18674
rect 7086 18622 7138 18674
rect 8654 18622 8706 18674
rect 8878 18622 8930 18674
rect 10446 18622 10498 18674
rect 11454 18622 11506 18674
rect 27134 18622 27186 18674
rect 27358 18622 27410 18674
rect 40126 18622 40178 18674
rect 5966 18510 6018 18562
rect 8094 18510 8146 18562
rect 11342 18510 11394 18562
rect 13582 18510 13634 18562
rect 17614 18510 17666 18562
rect 20078 18510 20130 18562
rect 24334 18510 24386 18562
rect 28366 18510 28418 18562
rect 33518 18510 33570 18562
rect 41134 18510 41186 18562
rect 44270 18510 44322 18562
rect 44606 18510 44658 18562
rect 45838 18510 45890 18562
rect 47070 18510 47122 18562
rect 2830 18398 2882 18450
rect 3502 18398 3554 18450
rect 6190 18398 6242 18450
rect 6750 18398 6802 18450
rect 7198 18398 7250 18450
rect 7310 18398 7362 18450
rect 7870 18398 7922 18450
rect 8542 18398 8594 18450
rect 9998 18398 10050 18450
rect 10334 18398 10386 18450
rect 10558 18398 10610 18450
rect 10782 18398 10834 18450
rect 11006 18398 11058 18450
rect 11678 18398 11730 18450
rect 13358 18398 13410 18450
rect 14702 18398 14754 18450
rect 17390 18398 17442 18450
rect 17950 18398 18002 18450
rect 19294 18398 19346 18450
rect 22878 18398 22930 18450
rect 24110 18398 24162 18450
rect 25342 18398 25394 18450
rect 27582 18398 27634 18450
rect 28254 18398 28306 18450
rect 29710 18398 29762 18450
rect 30382 18398 30434 18450
rect 33854 18398 33906 18450
rect 36878 18398 36930 18450
rect 41470 18398 41522 18450
rect 41806 18398 41858 18450
rect 42926 18398 42978 18450
rect 43486 18398 43538 18450
rect 44046 18398 44098 18450
rect 44718 18398 44770 18450
rect 44830 18398 44882 18450
rect 45166 18398 45218 18450
rect 45614 18398 45666 18450
rect 46734 18398 46786 18450
rect 47294 18398 47346 18450
rect 48078 18398 48130 18450
rect 5630 18286 5682 18338
rect 8206 18286 8258 18338
rect 13694 18286 13746 18338
rect 17838 18286 17890 18338
rect 22206 18286 22258 18338
rect 23102 18286 23154 18338
rect 23886 18286 23938 18338
rect 24222 18286 24274 18338
rect 32510 18286 32562 18338
rect 37550 18286 37602 18338
rect 39678 18286 39730 18338
rect 41918 18286 41970 18338
rect 42590 18286 42642 18338
rect 46286 18286 46338 18338
rect 47182 18286 47234 18338
rect 47630 18286 47682 18338
rect 13918 18174 13970 18226
rect 14142 18174 14194 18226
rect 23662 18174 23714 18226
rect 25230 18174 25282 18226
rect 43150 18174 43202 18226
rect 46062 18174 46114 18226
rect 46510 18174 46562 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 1934 17838 1986 17890
rect 15262 17838 15314 17890
rect 22654 17838 22706 17890
rect 26574 17838 26626 17890
rect 30942 17838 30994 17890
rect 42702 17838 42754 17890
rect 6862 17726 6914 17778
rect 11790 17726 11842 17778
rect 14926 17726 14978 17778
rect 16270 17726 16322 17778
rect 19294 17726 19346 17778
rect 29934 17726 29986 17778
rect 34190 17726 34242 17778
rect 36094 17726 36146 17778
rect 40238 17726 40290 17778
rect 42254 17726 42306 17778
rect 44158 17726 44210 17778
rect 45614 17726 45666 17778
rect 4174 17614 4226 17666
rect 6526 17614 6578 17666
rect 6974 17614 7026 17666
rect 10894 17614 10946 17666
rect 13582 17614 13634 17666
rect 14030 17614 14082 17666
rect 15822 17614 15874 17666
rect 16046 17614 16098 17666
rect 17054 17614 17106 17666
rect 17390 17614 17442 17666
rect 20750 17614 20802 17666
rect 23662 17614 23714 17666
rect 23886 17614 23938 17666
rect 23998 17614 24050 17666
rect 25342 17614 25394 17666
rect 25902 17614 25954 17666
rect 26798 17614 26850 17666
rect 29374 17614 29426 17666
rect 29598 17614 29650 17666
rect 30494 17614 30546 17666
rect 30718 17614 30770 17666
rect 34078 17614 34130 17666
rect 34414 17614 34466 17666
rect 34750 17614 34802 17666
rect 37662 17614 37714 17666
rect 38222 17614 38274 17666
rect 43038 17614 43090 17666
rect 43150 17614 43202 17666
rect 44270 17614 44322 17666
rect 44830 17614 44882 17666
rect 45726 17614 45778 17666
rect 46622 17614 46674 17666
rect 46958 17614 47010 17666
rect 47182 17614 47234 17666
rect 47854 17614 47906 17666
rect 7198 17502 7250 17554
rect 15038 17502 15090 17554
rect 15598 17502 15650 17554
rect 16494 17502 16546 17554
rect 16830 17502 16882 17554
rect 22542 17502 22594 17554
rect 24222 17502 24274 17554
rect 25566 17502 25618 17554
rect 35758 17502 35810 17554
rect 36206 17502 36258 17554
rect 36430 17502 36482 17554
rect 46062 17502 46114 17554
rect 47630 17502 47682 17554
rect 5854 17390 5906 17442
rect 6750 17390 6802 17442
rect 14702 17390 14754 17442
rect 15934 17390 15986 17442
rect 17166 17390 17218 17442
rect 17278 17390 17330 17442
rect 21422 17390 21474 17442
rect 21870 17390 21922 17442
rect 23774 17390 23826 17442
rect 34302 17390 34354 17442
rect 37214 17390 37266 17442
rect 37886 17390 37938 17442
rect 42366 17390 42418 17442
rect 43262 17390 43314 17442
rect 43374 17390 43426 17442
rect 44942 17390 44994 17442
rect 46734 17390 46786 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 5742 17054 5794 17106
rect 16046 17054 16098 17106
rect 18062 17054 18114 17106
rect 22766 17054 22818 17106
rect 25566 17054 25618 17106
rect 27134 17054 27186 17106
rect 33518 17054 33570 17106
rect 39230 17054 39282 17106
rect 40126 17054 40178 17106
rect 43038 17054 43090 17106
rect 44046 17054 44098 17106
rect 44270 17054 44322 17106
rect 44942 17054 44994 17106
rect 6414 16942 6466 16994
rect 6750 16942 6802 16994
rect 14366 16942 14418 16994
rect 15934 16942 15986 16994
rect 16494 16942 16546 16994
rect 23662 16942 23714 16994
rect 25454 16942 25506 16994
rect 26574 16942 26626 16994
rect 28030 16942 28082 16994
rect 29598 16942 29650 16994
rect 35422 16942 35474 16994
rect 38782 16942 38834 16994
rect 39790 16942 39842 16994
rect 41022 16942 41074 16994
rect 43822 16942 43874 16994
rect 1822 16830 1874 16882
rect 5294 16830 5346 16882
rect 7422 16830 7474 16882
rect 8430 16830 8482 16882
rect 8878 16830 8930 16882
rect 10446 16830 10498 16882
rect 10558 16830 10610 16882
rect 10894 16830 10946 16882
rect 13582 16830 13634 16882
rect 14926 16830 14978 16882
rect 16158 16830 16210 16882
rect 16830 16830 16882 16882
rect 17502 16830 17554 16882
rect 20974 16830 21026 16882
rect 21422 16830 21474 16882
rect 22430 16830 22482 16882
rect 23102 16830 23154 16882
rect 23886 16830 23938 16882
rect 25678 16830 25730 16882
rect 26126 16830 26178 16882
rect 27022 16830 27074 16882
rect 27358 16830 27410 16882
rect 28254 16830 28306 16882
rect 28814 16830 28866 16882
rect 30494 16830 30546 16882
rect 31726 16830 31778 16882
rect 33854 16830 33906 16882
rect 34078 16830 34130 16882
rect 34638 16830 34690 16882
rect 39006 16830 39058 16882
rect 39342 16830 39394 16882
rect 40910 16830 40962 16882
rect 42142 16830 42194 16882
rect 42366 16830 42418 16882
rect 42814 16830 42866 16882
rect 43262 16830 43314 16882
rect 43486 16830 43538 16882
rect 44494 16830 44546 16882
rect 44830 16830 44882 16882
rect 45614 16830 45666 16882
rect 2494 16718 2546 16770
rect 4622 16718 4674 16770
rect 5070 16718 5122 16770
rect 7646 16718 7698 16770
rect 10782 16718 10834 16770
rect 12574 16718 12626 16770
rect 15486 16718 15538 16770
rect 16718 16718 16770 16770
rect 17726 16718 17778 16770
rect 19854 16718 19906 16770
rect 21758 16718 21810 16770
rect 23998 16718 24050 16770
rect 27694 16718 27746 16770
rect 28142 16718 28194 16770
rect 37550 16718 37602 16770
rect 39118 16718 39170 16770
rect 41470 16718 41522 16770
rect 43038 16718 43090 16770
rect 44382 16718 44434 16770
rect 4958 16606 5010 16658
rect 8206 16606 8258 16658
rect 14478 16606 14530 16658
rect 14702 16606 14754 16658
rect 28590 16606 28642 16658
rect 47966 16606 48018 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 1934 16270 1986 16322
rect 7310 16270 7362 16322
rect 13470 16270 13522 16322
rect 29934 16270 29986 16322
rect 38110 16270 38162 16322
rect 4958 16158 5010 16210
rect 8206 16158 8258 16210
rect 9774 16158 9826 16210
rect 13806 16158 13858 16210
rect 16158 16158 16210 16210
rect 19070 16158 19122 16210
rect 21758 16158 21810 16210
rect 25230 16158 25282 16210
rect 29598 16158 29650 16210
rect 31166 16158 31218 16210
rect 34302 16158 34354 16210
rect 36430 16158 36482 16210
rect 37998 16158 38050 16210
rect 38558 16158 38610 16210
rect 40910 16158 40962 16210
rect 42366 16158 42418 16210
rect 43486 16158 43538 16210
rect 45838 16158 45890 16210
rect 48078 16158 48130 16210
rect 4062 16046 4114 16098
rect 6414 16046 6466 16098
rect 7198 16046 7250 16098
rect 7646 16046 7698 16098
rect 7870 16046 7922 16098
rect 8094 16046 8146 16098
rect 8766 16046 8818 16098
rect 9102 16046 9154 16098
rect 10110 16046 10162 16098
rect 11790 16046 11842 16098
rect 12238 16046 12290 16098
rect 15374 16046 15426 16098
rect 16382 16046 16434 16098
rect 18510 16046 18562 16098
rect 19630 16046 19682 16098
rect 20078 16046 20130 16098
rect 20526 16046 20578 16098
rect 22094 16046 22146 16098
rect 22878 16046 22930 16098
rect 25118 16046 25170 16098
rect 25342 16046 25394 16098
rect 27582 16046 27634 16098
rect 27918 16046 27970 16098
rect 29710 16046 29762 16098
rect 32958 16046 33010 16098
rect 35982 16046 36034 16098
rect 36318 16046 36370 16098
rect 40798 16046 40850 16098
rect 41470 16046 41522 16098
rect 41918 16046 41970 16098
rect 42478 16046 42530 16098
rect 42814 16046 42866 16098
rect 45054 16046 45106 16098
rect 6190 15934 6242 15986
rect 9998 15934 10050 15986
rect 11342 15934 11394 15986
rect 12910 15928 12962 15980
rect 14254 15934 14306 15986
rect 14590 15934 14642 15986
rect 15486 15934 15538 15986
rect 16158 15934 16210 15986
rect 17390 15934 17442 15986
rect 17726 15934 17778 15986
rect 18062 15934 18114 15986
rect 18734 15934 18786 15986
rect 21422 15934 21474 15986
rect 21646 15934 21698 15986
rect 25566 15934 25618 15986
rect 28478 15934 28530 15986
rect 28590 15934 28642 15986
rect 30270 15934 30322 15986
rect 38446 15934 38498 15986
rect 40462 15934 40514 15986
rect 42254 15934 42306 15986
rect 43822 15934 43874 15986
rect 8206 15822 8258 15874
rect 12798 15822 12850 15874
rect 13694 15822 13746 15874
rect 14926 15822 14978 15874
rect 22430 15822 22482 15874
rect 27694 15822 27746 15874
rect 30046 15822 30098 15874
rect 43374 15822 43426 15874
rect 44158 15822 44210 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 6302 15486 6354 15538
rect 11454 15486 11506 15538
rect 11566 15486 11618 15538
rect 12686 15486 12738 15538
rect 15150 15486 15202 15538
rect 16942 15486 16994 15538
rect 25678 15486 25730 15538
rect 33294 15486 33346 15538
rect 33406 15486 33458 15538
rect 34190 15486 34242 15538
rect 37102 15486 37154 15538
rect 37438 15486 37490 15538
rect 40798 15486 40850 15538
rect 42030 15486 42082 15538
rect 42254 15486 42306 15538
rect 43038 15486 43090 15538
rect 44270 15486 44322 15538
rect 45166 15486 45218 15538
rect 45726 15486 45778 15538
rect 46398 15486 46450 15538
rect 47518 15486 47570 15538
rect 47854 15486 47906 15538
rect 3390 15374 3442 15426
rect 3838 15374 3890 15426
rect 4174 15374 4226 15426
rect 5182 15374 5234 15426
rect 5294 15374 5346 15426
rect 6190 15374 6242 15426
rect 7086 15374 7138 15426
rect 7758 15374 7810 15426
rect 8766 15374 8818 15426
rect 14142 15374 14194 15426
rect 21758 15374 21810 15426
rect 25230 15374 25282 15426
rect 27358 15374 27410 15426
rect 31054 15374 31106 15426
rect 32174 15374 32226 15426
rect 38222 15374 38274 15426
rect 38558 15374 38610 15426
rect 38894 15374 38946 15426
rect 41358 15374 41410 15426
rect 41694 15374 41746 15426
rect 43934 15374 43986 15426
rect 2942 15262 2994 15314
rect 3278 15262 3330 15314
rect 4398 15262 4450 15314
rect 5518 15262 5570 15314
rect 6974 15262 7026 15314
rect 7646 15262 7698 15314
rect 8990 15262 9042 15314
rect 9998 15262 10050 15314
rect 10222 15262 10274 15314
rect 10446 15262 10498 15314
rect 10670 15262 10722 15314
rect 11006 15262 11058 15314
rect 11678 15262 11730 15314
rect 12238 15262 12290 15314
rect 12462 15262 12514 15314
rect 12910 15262 12962 15314
rect 13694 15262 13746 15314
rect 13806 15262 13858 15314
rect 14254 15262 14306 15314
rect 15486 15262 15538 15314
rect 16158 15262 16210 15314
rect 20190 15262 20242 15314
rect 20974 15262 21026 15314
rect 25454 15262 25506 15314
rect 25790 15262 25842 15314
rect 26126 15262 26178 15314
rect 26462 15262 26514 15314
rect 26686 15262 26738 15314
rect 27470 15262 27522 15314
rect 31838 15262 31890 15314
rect 32398 15262 32450 15314
rect 33182 15262 33234 15314
rect 33854 15262 33906 15314
rect 34078 15262 34130 15314
rect 34414 15262 34466 15314
rect 34638 15262 34690 15314
rect 37438 15262 37490 15314
rect 37998 15262 38050 15314
rect 39118 15262 39170 15314
rect 41022 15262 41074 15314
rect 41806 15262 41858 15314
rect 42366 15262 42418 15314
rect 42814 15262 42866 15314
rect 43150 15262 43202 15314
rect 43262 15262 43314 15314
rect 43374 15262 43426 15314
rect 44382 15262 44434 15314
rect 45278 15262 45330 15314
rect 45614 15262 45666 15314
rect 46958 15262 47010 15314
rect 3950 15150 4002 15202
rect 8318 15150 8370 15202
rect 10558 15150 10610 15202
rect 14702 15150 14754 15202
rect 15710 15150 15762 15202
rect 17390 15150 17442 15202
rect 19518 15150 19570 15202
rect 23886 15150 23938 15202
rect 25566 15150 25618 15202
rect 26350 15150 26402 15202
rect 28926 15150 28978 15202
rect 38670 15150 38722 15202
rect 47070 15150 47122 15202
rect 4734 15038 4786 15090
rect 7086 15038 7138 15090
rect 12350 15038 12402 15090
rect 27358 15038 27410 15090
rect 37774 15038 37826 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 4062 14702 4114 14754
rect 11118 14702 11170 14754
rect 11566 14702 11618 14754
rect 12014 14702 12066 14754
rect 17614 14702 17666 14754
rect 18174 14702 18226 14754
rect 18510 14702 18562 14754
rect 25902 14702 25954 14754
rect 27022 14702 27074 14754
rect 15262 14590 15314 14642
rect 21310 14590 21362 14642
rect 24782 14590 24834 14642
rect 26798 14590 26850 14642
rect 29486 14590 29538 14642
rect 32174 14590 32226 14642
rect 35646 14590 35698 14642
rect 44270 14590 44322 14642
rect 3726 14478 3778 14530
rect 3950 14478 4002 14530
rect 5070 14478 5122 14530
rect 6750 14478 6802 14530
rect 8766 14478 8818 14530
rect 11342 14478 11394 14530
rect 13470 14478 13522 14530
rect 14814 14478 14866 14530
rect 15486 14478 15538 14530
rect 17614 14478 17666 14530
rect 18062 14478 18114 14530
rect 18398 14478 18450 14530
rect 19182 14478 19234 14530
rect 19630 14478 19682 14530
rect 21758 14478 21810 14530
rect 22206 14478 22258 14530
rect 26238 14478 26290 14530
rect 27358 14478 27410 14530
rect 27694 14478 27746 14530
rect 29374 14478 29426 14530
rect 29710 14478 29762 14530
rect 31054 14478 31106 14530
rect 31278 14478 31330 14530
rect 31502 14478 31554 14530
rect 33182 14478 33234 14530
rect 35198 14478 35250 14530
rect 35422 14478 35474 14530
rect 38110 14478 38162 14530
rect 38446 14478 38498 14530
rect 41582 14478 41634 14530
rect 45054 14478 45106 14530
rect 46286 14478 46338 14530
rect 48078 14478 48130 14530
rect 3614 14366 3666 14418
rect 4958 14366 5010 14418
rect 5630 14366 5682 14418
rect 5966 14366 6018 14418
rect 7870 14366 7922 14418
rect 9326 14366 9378 14418
rect 10894 14366 10946 14418
rect 12574 14366 12626 14418
rect 12686 14366 12738 14418
rect 13694 14366 13746 14418
rect 14478 14366 14530 14418
rect 17278 14366 17330 14418
rect 25118 14366 25170 14418
rect 25566 14366 25618 14418
rect 26350 14366 26402 14418
rect 29150 14366 29202 14418
rect 31726 14366 31778 14418
rect 32846 14366 32898 14418
rect 32958 14366 33010 14418
rect 34414 14366 34466 14418
rect 34862 14366 34914 14418
rect 34974 14366 35026 14418
rect 35870 14366 35922 14418
rect 36094 14366 36146 14418
rect 38222 14366 38274 14418
rect 41246 14366 41298 14418
rect 44830 14366 44882 14418
rect 45726 14366 45778 14418
rect 47070 14366 47122 14418
rect 47854 14366 47906 14418
rect 4622 14254 4674 14306
rect 10334 14254 10386 14306
rect 12350 14254 12402 14306
rect 13806 14254 13858 14306
rect 15822 14254 15874 14306
rect 18846 14254 18898 14306
rect 24222 14254 24274 14306
rect 25230 14254 25282 14306
rect 25790 14254 25842 14306
rect 27470 14254 27522 14306
rect 27582 14254 27634 14306
rect 29598 14254 29650 14306
rect 31390 14254 31442 14306
rect 41358 14254 41410 14306
rect 42030 14254 42082 14306
rect 45838 14254 45890 14306
rect 45950 14254 46002 14306
rect 46846 14254 46898 14306
rect 47406 14254 47458 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 7422 13918 7474 13970
rect 14142 13918 14194 13970
rect 17726 13918 17778 13970
rect 28142 13918 28194 13970
rect 32398 13918 32450 13970
rect 34638 13918 34690 13970
rect 35310 13918 35362 13970
rect 36094 13918 36146 13970
rect 36430 13918 36482 13970
rect 37102 13918 37154 13970
rect 37550 13918 37602 13970
rect 40350 13918 40402 13970
rect 44382 13918 44434 13970
rect 45502 13918 45554 13970
rect 46398 13918 46450 13970
rect 46622 13918 46674 13970
rect 2494 13806 2546 13858
rect 7086 13806 7138 13858
rect 8654 13806 8706 13858
rect 9662 13806 9714 13858
rect 9886 13806 9938 13858
rect 12238 13806 12290 13858
rect 12910 13806 12962 13858
rect 27470 13806 27522 13858
rect 29486 13806 29538 13858
rect 31054 13806 31106 13858
rect 35086 13806 35138 13858
rect 37886 13806 37938 13858
rect 1822 13694 1874 13746
rect 7310 13694 7362 13746
rect 7534 13694 7586 13746
rect 7758 13694 7810 13746
rect 8206 13694 8258 13746
rect 8318 13694 8370 13746
rect 10334 13694 10386 13746
rect 12014 13694 12066 13746
rect 13022 13694 13074 13746
rect 13582 13694 13634 13746
rect 20190 13694 20242 13746
rect 27358 13694 27410 13746
rect 27918 13694 27970 13746
rect 28926 13694 28978 13746
rect 29262 13694 29314 13746
rect 31502 13694 31554 13746
rect 31614 13694 31666 13746
rect 31838 13694 31890 13746
rect 33854 13694 33906 13746
rect 34078 13694 34130 13746
rect 34302 13694 34354 13746
rect 34414 13694 34466 13746
rect 34974 13694 35026 13746
rect 35982 13694 36034 13746
rect 38670 13806 38722 13858
rect 39790 13806 39842 13858
rect 39902 13806 39954 13858
rect 41134 13806 41186 13858
rect 46174 13806 46226 13858
rect 47854 13806 47906 13858
rect 36206 13694 36258 13746
rect 37774 13694 37826 13746
rect 38222 13694 38274 13746
rect 39678 13694 39730 13746
rect 40910 13694 40962 13746
rect 41246 13694 41298 13746
rect 41470 13694 41522 13746
rect 41918 13694 41970 13746
rect 42478 13694 42530 13746
rect 42702 13694 42754 13746
rect 46958 13694 47010 13746
rect 48190 13694 48242 13746
rect 4622 13582 4674 13634
rect 5070 13582 5122 13634
rect 8542 13582 8594 13634
rect 9550 13582 9602 13634
rect 18174 13582 18226 13634
rect 18734 13582 18786 13634
rect 20862 13582 20914 13634
rect 22990 13582 23042 13634
rect 24558 13582 24610 13634
rect 27134 13582 27186 13634
rect 29486 13582 29538 13634
rect 38334 13582 38386 13634
rect 44718 13582 44770 13634
rect 46510 13582 46562 13634
rect 47518 13582 47570 13634
rect 10558 13470 10610 13522
rect 37438 13470 37490 13522
rect 42142 13470 42194 13522
rect 42254 13470 42306 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 10446 13134 10498 13186
rect 13470 13134 13522 13186
rect 29486 13134 29538 13186
rect 29934 13134 29986 13186
rect 4398 13022 4450 13074
rect 22094 13022 22146 13074
rect 26574 13022 26626 13074
rect 28254 13022 28306 13074
rect 32062 13022 32114 13074
rect 41134 13022 41186 13074
rect 42142 13022 42194 13074
rect 44270 13022 44322 13074
rect 47966 13022 48018 13074
rect 6302 12910 6354 12962
rect 6526 12910 6578 12962
rect 9998 12910 10050 12962
rect 10110 12910 10162 12962
rect 13582 12910 13634 12962
rect 14478 12910 14530 12962
rect 14702 12910 14754 12962
rect 14926 12910 14978 12962
rect 15710 12910 15762 12962
rect 15934 12910 15986 12962
rect 17838 12910 17890 12962
rect 23438 12910 23490 12962
rect 24110 12910 24162 12962
rect 25230 12910 25282 12962
rect 25678 12910 25730 12962
rect 26238 12910 26290 12962
rect 27918 12910 27970 12962
rect 28366 12910 28418 12962
rect 29598 12910 29650 12962
rect 29822 12910 29874 12962
rect 32286 12910 32338 12962
rect 40126 12910 40178 12962
rect 40238 12910 40290 12962
rect 40574 12910 40626 12962
rect 41358 12910 41410 12962
rect 45054 12910 45106 12962
rect 4734 12798 4786 12850
rect 6078 12798 6130 12850
rect 8990 12798 9042 12850
rect 15150 12798 15202 12850
rect 15822 12798 15874 12850
rect 18734 12798 18786 12850
rect 18846 12798 18898 12850
rect 18958 12798 19010 12850
rect 22430 12798 22482 12850
rect 23326 12798 23378 12850
rect 24334 12798 24386 12850
rect 24894 12798 24946 12850
rect 27022 12798 27074 12850
rect 31950 12798 32002 12850
rect 32510 12798 32562 12850
rect 45838 12798 45890 12850
rect 6190 12686 6242 12738
rect 9326 12686 9378 12738
rect 9774 12686 9826 12738
rect 9886 12686 9938 12738
rect 15038 12686 15090 12738
rect 16382 12686 16434 12738
rect 18062 12686 18114 12738
rect 19406 12686 19458 12738
rect 22766 12686 22818 12738
rect 24222 12686 24274 12738
rect 27246 12686 27298 12738
rect 28142 12686 28194 12738
rect 28478 12686 28530 12738
rect 40462 12686 40514 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 5294 12350 5346 12402
rect 7310 12350 7362 12402
rect 7758 12350 7810 12402
rect 8878 12350 8930 12402
rect 10558 12350 10610 12402
rect 16158 12350 16210 12402
rect 16270 12350 16322 12402
rect 17502 12350 17554 12402
rect 23998 12350 24050 12402
rect 24558 12350 24610 12402
rect 25454 12350 25506 12402
rect 26238 12350 26290 12402
rect 31390 12350 31442 12402
rect 34302 12350 34354 12402
rect 36094 12350 36146 12402
rect 37998 12350 38050 12402
rect 38110 12350 38162 12402
rect 43374 12350 43426 12402
rect 44942 12350 44994 12402
rect 4846 12238 4898 12290
rect 8654 12238 8706 12290
rect 12686 12238 12738 12290
rect 14590 12238 14642 12290
rect 18622 12238 18674 12290
rect 19630 12238 19682 12290
rect 21982 12238 22034 12290
rect 22206 12238 22258 12290
rect 23438 12238 23490 12290
rect 23886 12238 23938 12290
rect 24670 12238 24722 12290
rect 25230 12238 25282 12290
rect 28254 12238 28306 12290
rect 29038 12238 29090 12290
rect 30494 12238 30546 12290
rect 31278 12238 31330 12290
rect 32286 12238 32338 12290
rect 34190 12238 34242 12290
rect 34862 12238 34914 12290
rect 35870 12238 35922 12290
rect 36990 12238 37042 12290
rect 39118 12238 39170 12290
rect 43710 12238 43762 12290
rect 44270 12238 44322 12290
rect 44382 12238 44434 12290
rect 45054 12238 45106 12290
rect 45278 12238 45330 12290
rect 3838 12126 3890 12178
rect 5854 12126 5906 12178
rect 6190 12126 6242 12178
rect 6414 12126 6466 12178
rect 6638 12126 6690 12178
rect 7198 12126 7250 12178
rect 9550 12126 9602 12178
rect 9774 12126 9826 12178
rect 9998 12126 10050 12178
rect 13022 12126 13074 12178
rect 13694 12126 13746 12178
rect 14030 12126 14082 12178
rect 15038 12126 15090 12178
rect 15822 12126 15874 12178
rect 16046 12126 16098 12178
rect 16494 12126 16546 12178
rect 18174 12126 18226 12178
rect 19742 12126 19794 12178
rect 21534 12126 21586 12178
rect 22878 12126 22930 12178
rect 26462 12126 26514 12178
rect 27246 12126 27298 12178
rect 27470 12126 27522 12178
rect 27918 12126 27970 12178
rect 28478 12126 28530 12178
rect 29486 12126 29538 12178
rect 29934 12126 29986 12178
rect 31054 12126 31106 12178
rect 32510 12126 32562 12178
rect 33966 12126 34018 12178
rect 34414 12126 34466 12178
rect 35422 12126 35474 12178
rect 36206 12126 36258 12178
rect 36430 12126 36482 12178
rect 36766 12126 36818 12178
rect 37214 12126 37266 12178
rect 37438 12126 37490 12178
rect 37774 12126 37826 12178
rect 38222 12126 38274 12178
rect 38446 12126 38498 12178
rect 38782 12126 38834 12178
rect 40910 12126 40962 12178
rect 41134 12126 41186 12178
rect 41358 12126 41410 12178
rect 44718 12126 44770 12178
rect 46062 12126 46114 12178
rect 3950 12014 4002 12066
rect 4286 12014 4338 12066
rect 4622 12014 4674 12066
rect 4734 12014 4786 12066
rect 8990 12014 9042 12066
rect 14366 12014 14418 12066
rect 21198 12014 21250 12066
rect 21758 12014 21810 12066
rect 25566 12014 25618 12066
rect 30158 12014 30210 12066
rect 37102 12014 37154 12066
rect 40350 12014 40402 12066
rect 47966 12014 48018 12066
rect 6750 11902 6802 11954
rect 10110 11902 10162 11954
rect 23326 11902 23378 11954
rect 26126 11902 26178 11954
rect 33742 11902 33794 11954
rect 41470 11902 41522 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 13470 11566 13522 11618
rect 21310 11566 21362 11618
rect 21422 11566 21474 11618
rect 21646 11566 21698 11618
rect 27806 11566 27858 11618
rect 30494 11566 30546 11618
rect 34302 11566 34354 11618
rect 37998 11566 38050 11618
rect 2494 11454 2546 11506
rect 4622 11454 4674 11506
rect 7422 11454 7474 11506
rect 8878 11454 8930 11506
rect 11678 11454 11730 11506
rect 16158 11454 16210 11506
rect 17950 11454 18002 11506
rect 22542 11454 22594 11506
rect 33518 11454 33570 11506
rect 34414 11454 34466 11506
rect 42030 11454 42082 11506
rect 44158 11454 44210 11506
rect 47966 11454 48018 11506
rect 1822 11342 1874 11394
rect 7086 11342 7138 11394
rect 10782 11342 10834 11394
rect 11790 11342 11842 11394
rect 12238 11342 12290 11394
rect 12686 11342 12738 11394
rect 13694 11342 13746 11394
rect 14254 11342 14306 11394
rect 15038 11342 15090 11394
rect 15486 11342 15538 11394
rect 15822 11342 15874 11394
rect 17614 11342 17666 11394
rect 18510 11342 18562 11394
rect 20862 11342 20914 11394
rect 21758 11342 21810 11394
rect 23214 11342 23266 11394
rect 25230 11342 25282 11394
rect 29486 11342 29538 11394
rect 29710 11342 29762 11394
rect 30046 11342 30098 11394
rect 30718 11342 30770 11394
rect 30942 11342 30994 11394
rect 31054 11342 31106 11394
rect 31726 11342 31778 11394
rect 32734 11342 32786 11394
rect 33630 11342 33682 11394
rect 35646 11342 35698 11394
rect 35870 11342 35922 11394
rect 37214 11342 37266 11394
rect 40910 11342 40962 11394
rect 41246 11342 41298 11394
rect 46062 11342 46114 11394
rect 9214 11230 9266 11282
rect 9550 11230 9602 11282
rect 11118 11230 11170 11282
rect 12462 11230 12514 11282
rect 13806 11230 13858 11282
rect 18734 11230 18786 11282
rect 18958 11230 19010 11282
rect 19630 11230 19682 11282
rect 22878 11230 22930 11282
rect 24334 11230 24386 11282
rect 25790 11230 25842 11282
rect 27918 11230 27970 11282
rect 33182 11230 33234 11282
rect 33518 11230 33570 11282
rect 36878 11230 36930 11282
rect 38110 11230 38162 11282
rect 5070 11118 5122 11170
rect 5742 11118 5794 11170
rect 9886 11118 9938 11170
rect 10222 11118 10274 11170
rect 11342 11118 11394 11170
rect 11566 11118 11618 11170
rect 12350 11118 12402 11170
rect 12574 11118 12626 11170
rect 15598 11118 15650 11170
rect 22654 11118 22706 11170
rect 26798 11118 26850 11170
rect 31166 11118 31218 11170
rect 35758 11118 35810 11170
rect 37102 11118 37154 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 11790 10782 11842 10834
rect 14702 10782 14754 10834
rect 15598 10782 15650 10834
rect 16382 10782 16434 10834
rect 17502 10782 17554 10834
rect 19294 10782 19346 10834
rect 29150 10782 29202 10834
rect 30718 10782 30770 10834
rect 32062 10782 32114 10834
rect 36878 10782 36930 10834
rect 38446 10782 38498 10834
rect 39566 10782 39618 10834
rect 4958 10670 5010 10722
rect 11902 10670 11954 10722
rect 12910 10670 12962 10722
rect 14478 10670 14530 10722
rect 15150 10670 15202 10722
rect 18286 10670 18338 10722
rect 4286 10558 4338 10610
rect 14366 10558 14418 10610
rect 15710 10558 15762 10610
rect 16046 10558 16098 10610
rect 17838 10558 17890 10610
rect 19182 10614 19234 10666
rect 23438 10670 23490 10722
rect 23550 10670 23602 10722
rect 27582 10670 27634 10722
rect 28926 10670 28978 10722
rect 32398 10670 32450 10722
rect 34750 10670 34802 10722
rect 36542 10670 36594 10722
rect 43598 10670 43650 10722
rect 43822 10670 43874 10722
rect 47854 10670 47906 10722
rect 48190 10670 48242 10722
rect 23774 10558 23826 10610
rect 26686 10558 26738 10610
rect 26910 10558 26962 10610
rect 27806 10558 27858 10610
rect 28366 10558 28418 10610
rect 28814 10558 28866 10610
rect 30718 10558 30770 10610
rect 34526 10558 34578 10610
rect 35086 10558 35138 10610
rect 35758 10558 35810 10610
rect 36766 10558 36818 10610
rect 36990 10558 37042 10610
rect 37214 10558 37266 10610
rect 37774 10558 37826 10610
rect 37886 10558 37938 10610
rect 37998 10558 38050 10610
rect 38782 10558 38834 10610
rect 39118 10558 39170 10610
rect 39230 10558 39282 10610
rect 39342 10558 39394 10610
rect 44270 10558 44322 10610
rect 44494 10558 44546 10610
rect 45278 10558 45330 10610
rect 7086 10446 7138 10498
rect 7534 10446 7586 10498
rect 12574 10446 12626 10498
rect 18846 10446 18898 10498
rect 44046 10446 44098 10498
rect 47406 10446 47458 10498
rect 17950 10334 18002 10386
rect 19294 10334 19346 10386
rect 35646 10334 35698 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 44830 9998 44882 10050
rect 7982 9886 8034 9938
rect 10110 9886 10162 9938
rect 11902 9886 11954 9938
rect 14366 9886 14418 9938
rect 14926 9886 14978 9938
rect 17838 9886 17890 9938
rect 21646 9886 21698 9938
rect 27358 9886 27410 9938
rect 28254 9886 28306 9938
rect 29934 9886 29986 9938
rect 33630 9886 33682 9938
rect 34414 9886 34466 9938
rect 35534 9886 35586 9938
rect 39230 9886 39282 9938
rect 41358 9886 41410 9938
rect 43598 9886 43650 9938
rect 44942 9886 44994 9938
rect 47966 9886 48018 9938
rect 7310 9774 7362 9826
rect 11566 9774 11618 9826
rect 12350 9774 12402 9826
rect 12910 9774 12962 9826
rect 13918 9774 13970 9826
rect 14478 9774 14530 9826
rect 15038 9774 15090 9826
rect 16382 9774 16434 9826
rect 17278 9774 17330 9826
rect 20638 9774 20690 9826
rect 21982 9774 22034 9826
rect 23214 9774 23266 9826
rect 25230 9774 25282 9826
rect 27918 9774 27970 9826
rect 29598 9774 29650 9826
rect 30942 9774 30994 9826
rect 31838 9774 31890 9826
rect 33070 9774 33122 9826
rect 34190 9774 34242 9826
rect 34526 9774 34578 9826
rect 35310 9774 35362 9826
rect 35758 9774 35810 9826
rect 38222 9774 38274 9826
rect 42030 9774 42082 9826
rect 43150 9774 43202 9826
rect 45614 9774 45666 9826
rect 14926 9662 14978 9714
rect 15486 9662 15538 9714
rect 17166 9662 17218 9714
rect 19966 9662 20018 9714
rect 22430 9662 22482 9714
rect 24334 9662 24386 9714
rect 25790 9662 25842 9714
rect 28366 9662 28418 9714
rect 30270 9662 30322 9714
rect 31054 9662 31106 9714
rect 32286 9662 32338 9714
rect 32398 9662 32450 9714
rect 32622 9662 32674 9714
rect 32958 9662 33010 9714
rect 33182 9662 33234 9714
rect 33966 9662 34018 9714
rect 35086 9662 35138 9714
rect 35534 9662 35586 9714
rect 37326 9662 37378 9714
rect 37886 9662 37938 9714
rect 37998 9662 38050 9714
rect 10558 9550 10610 9602
rect 14030 9550 14082 9602
rect 14254 9550 14306 9602
rect 15262 9550 15314 9602
rect 15934 9550 15986 9602
rect 16158 9550 16210 9602
rect 26798 9550 26850 9602
rect 31614 9550 31666 9602
rect 34750 9550 34802 9602
rect 36990 9550 37042 9602
rect 38558 9550 38610 9602
rect 42590 9550 42642 9602
rect 44158 9550 44210 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 7198 9214 7250 9266
rect 12910 9214 12962 9266
rect 14366 9214 14418 9266
rect 15374 9214 15426 9266
rect 19742 9214 19794 9266
rect 24670 9214 24722 9266
rect 27022 9214 27074 9266
rect 27582 9214 27634 9266
rect 28254 9214 28306 9266
rect 29486 9214 29538 9266
rect 34862 9214 34914 9266
rect 35198 9214 35250 9266
rect 36990 9214 37042 9266
rect 41358 9214 41410 9266
rect 47630 9214 47682 9266
rect 7534 9102 7586 9154
rect 14814 9102 14866 9154
rect 18958 9102 19010 9154
rect 19182 9102 19234 9154
rect 23886 9102 23938 9154
rect 24110 9102 24162 9154
rect 26462 9102 26514 9154
rect 28702 9102 28754 9154
rect 30158 9102 30210 9154
rect 33182 9102 33234 9154
rect 47854 9102 47906 9154
rect 9662 8990 9714 9042
rect 14254 8990 14306 9042
rect 14590 8990 14642 9042
rect 15822 8990 15874 9042
rect 15934 8990 15986 9042
rect 17838 8990 17890 9042
rect 18286 8990 18338 9042
rect 19406 8990 19458 9042
rect 19518 8990 19570 9042
rect 24334 8990 24386 9042
rect 24670 8990 24722 9042
rect 27582 8990 27634 9042
rect 28478 8990 28530 9042
rect 29822 8990 29874 9042
rect 37662 8990 37714 9042
rect 41694 8990 41746 9042
rect 48190 8990 48242 9042
rect 10334 8878 10386 8930
rect 12462 8878 12514 8930
rect 15486 8878 15538 8930
rect 17390 8878 17442 8930
rect 20190 8878 20242 8930
rect 23550 8878 23602 8930
rect 29934 8878 29986 8930
rect 33070 8878 33122 8930
rect 33630 8878 33682 8930
rect 36878 8878 36930 8930
rect 37886 8878 37938 8930
rect 38334 8878 38386 8930
rect 42478 8878 42530 8930
rect 44606 8878 44658 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 17726 8430 17778 8482
rect 21870 8430 21922 8482
rect 9998 8318 10050 8370
rect 13582 8318 13634 8370
rect 18174 8318 18226 8370
rect 21534 8318 21586 8370
rect 22318 8318 22370 8370
rect 24894 8318 24946 8370
rect 27022 8318 27074 8370
rect 27918 8318 27970 8370
rect 29934 8318 29986 8370
rect 32062 8318 32114 8370
rect 32510 8318 32562 8370
rect 32846 8318 32898 8370
rect 34974 8318 35026 8370
rect 38222 8318 38274 8370
rect 41582 8318 41634 8370
rect 42030 8318 42082 8370
rect 42590 8318 42642 8370
rect 48302 8318 48354 8370
rect 6974 8206 7026 8258
rect 7198 8206 7250 8258
rect 7646 8206 7698 8258
rect 7870 8206 7922 8258
rect 8318 8206 8370 8258
rect 9550 8206 9602 8258
rect 9774 8206 9826 8258
rect 10222 8206 10274 8258
rect 11454 8206 11506 8258
rect 24222 8206 24274 8258
rect 27694 8206 27746 8258
rect 29150 8206 29202 8258
rect 35758 8206 35810 8258
rect 41134 8206 41186 8258
rect 42142 8206 42194 8258
rect 42366 8206 42418 8258
rect 42814 8206 42866 8258
rect 43262 8206 43314 8258
rect 43934 8206 43986 8258
rect 45390 8206 45442 8258
rect 45838 8206 45890 8258
rect 46622 8206 46674 8258
rect 47070 8206 47122 8258
rect 1710 8094 1762 8146
rect 2046 8094 2098 8146
rect 6862 8094 6914 8146
rect 9438 8094 9490 8146
rect 10446 8094 10498 8146
rect 17502 8094 17554 8146
rect 21646 8094 21698 8146
rect 40350 8094 40402 8146
rect 43038 8094 43090 8146
rect 43822 8094 43874 8146
rect 45166 8094 45218 8146
rect 46174 8094 46226 8146
rect 2494 7982 2546 8034
rect 7422 7982 7474 8034
rect 8206 7982 8258 8034
rect 8430 7982 8482 8034
rect 8654 7982 8706 8034
rect 10782 7982 10834 8034
rect 10894 7982 10946 8034
rect 11006 7982 11058 8034
rect 17614 7982 17666 8034
rect 36206 7982 36258 8034
rect 43710 7982 43762 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 3950 7646 4002 7698
rect 7422 7646 7474 7698
rect 8318 7646 8370 7698
rect 8654 7646 8706 7698
rect 11902 7646 11954 7698
rect 12350 7646 12402 7698
rect 13582 7646 13634 7698
rect 13806 7646 13858 7698
rect 15150 7646 15202 7698
rect 16382 7646 16434 7698
rect 33406 7646 33458 7698
rect 37438 7646 37490 7698
rect 38894 7646 38946 7698
rect 42926 7646 42978 7698
rect 6190 7534 6242 7586
rect 10670 7534 10722 7586
rect 13022 7534 13074 7586
rect 14030 7534 14082 7586
rect 19518 7534 19570 7586
rect 21422 7534 21474 7586
rect 28478 7534 28530 7586
rect 34190 7534 34242 7586
rect 38670 7534 38722 7586
rect 43150 7534 43202 7586
rect 43598 7534 43650 7586
rect 6974 7422 7026 7474
rect 10334 7422 10386 7474
rect 12686 7422 12738 7474
rect 13134 7422 13186 7474
rect 13694 7422 13746 7474
rect 15486 7422 15538 7474
rect 20302 7422 20354 7474
rect 20638 7422 20690 7474
rect 24670 7422 24722 7474
rect 25678 7422 25730 7474
rect 26126 7422 26178 7474
rect 28030 7422 28082 7474
rect 28702 7422 28754 7474
rect 33854 7422 33906 7474
rect 37550 7422 37602 7474
rect 42702 7422 42754 7474
rect 43934 7422 43986 7474
rect 12238 7310 12290 7362
rect 12798 7310 12850 7362
rect 15934 7310 15986 7362
rect 17390 7310 17442 7362
rect 23550 7310 23602 7362
rect 24110 7310 24162 7362
rect 27582 7310 27634 7362
rect 32510 7310 32562 7362
rect 33518 7310 33570 7362
rect 38446 7310 38498 7362
rect 39006 7310 39058 7362
rect 42814 7310 42866 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19406 6862 19458 6914
rect 16382 6750 16434 6802
rect 25790 6750 25842 6802
rect 26238 6750 26290 6802
rect 32062 6750 32114 6802
rect 35982 6750 36034 6802
rect 6862 6638 6914 6690
rect 7086 6638 7138 6690
rect 8318 6638 8370 6690
rect 8654 6638 8706 6690
rect 9886 6638 9938 6690
rect 10446 6638 10498 6690
rect 10894 6638 10946 6690
rect 12910 6638 12962 6690
rect 13582 6638 13634 6690
rect 16830 6638 16882 6690
rect 17502 6638 17554 6690
rect 18958 6638 19010 6690
rect 19630 6638 19682 6690
rect 19854 6638 19906 6690
rect 22878 6638 22930 6690
rect 26126 6638 26178 6690
rect 26798 6638 26850 6690
rect 27358 6638 27410 6690
rect 28030 6638 28082 6690
rect 29150 6638 29202 6690
rect 29262 6638 29314 6690
rect 30718 6638 30770 6690
rect 31390 6638 31442 6690
rect 32734 6638 32786 6690
rect 34302 6638 34354 6690
rect 36094 6638 36146 6690
rect 36542 6638 36594 6690
rect 41582 6638 41634 6690
rect 41806 6638 41858 6690
rect 42142 6638 42194 6690
rect 42478 6638 42530 6690
rect 45614 6638 45666 6690
rect 6750 6526 6802 6578
rect 7534 6526 7586 6578
rect 7758 6526 7810 6578
rect 8206 6526 8258 6578
rect 11454 6526 11506 6578
rect 14254 6526 14306 6578
rect 17054 6526 17106 6578
rect 23662 6526 23714 6578
rect 29598 6526 29650 6578
rect 30158 6526 30210 6578
rect 33854 6526 33906 6578
rect 35534 6526 35586 6578
rect 37550 6526 37602 6578
rect 41470 6526 41522 6578
rect 47294 6526 47346 6578
rect 7310 6414 7362 6466
rect 8094 6414 8146 6466
rect 9102 6414 9154 6466
rect 11118 6414 11170 6466
rect 11790 6414 11842 6466
rect 12238 6414 12290 6466
rect 20414 6414 20466 6466
rect 21310 6414 21362 6466
rect 21646 6414 21698 6466
rect 26350 6414 26402 6466
rect 27806 6414 27858 6466
rect 27918 6414 27970 6466
rect 28478 6414 28530 6466
rect 29374 6414 29426 6466
rect 30494 6414 30546 6466
rect 31166 6414 31218 6466
rect 31278 6414 31330 6466
rect 33294 6414 33346 6466
rect 34078 6414 34130 6466
rect 34190 6414 34242 6466
rect 34750 6414 34802 6466
rect 35422 6414 35474 6466
rect 35870 6414 35922 6466
rect 37886 6414 37938 6466
rect 42030 6414 42082 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 8094 6078 8146 6130
rect 8430 6078 8482 6130
rect 9774 6078 9826 6130
rect 10670 6078 10722 6130
rect 20750 6078 20802 6130
rect 23886 6078 23938 6130
rect 28142 6078 28194 6130
rect 29262 6078 29314 6130
rect 31166 6078 31218 6130
rect 33294 6078 33346 6130
rect 38894 6078 38946 6130
rect 40350 6078 40402 6130
rect 6526 5966 6578 6018
rect 9550 5966 9602 6018
rect 18174 5966 18226 6018
rect 20302 5966 20354 6018
rect 24334 5966 24386 6018
rect 26798 5966 26850 6018
rect 27134 5966 27186 6018
rect 29934 5966 29986 6018
rect 34190 5966 34242 6018
rect 34974 5966 35026 6018
rect 35198 5966 35250 6018
rect 41694 5966 41746 6018
rect 7198 5854 7250 5906
rect 10110 5854 10162 5906
rect 11006 5854 11058 5906
rect 19406 5854 19458 5906
rect 20078 5854 20130 5906
rect 23438 5854 23490 5906
rect 23662 5854 23714 5906
rect 24110 5854 24162 5906
rect 26574 5854 26626 5906
rect 27470 5854 27522 5906
rect 27806 5854 27858 5906
rect 30830 5854 30882 5906
rect 31278 5854 31330 5906
rect 31390 5854 31442 5906
rect 33518 5854 33570 5906
rect 33966 5854 34018 5906
rect 34638 5854 34690 5906
rect 35646 5854 35698 5906
rect 41022 5854 41074 5906
rect 4398 5742 4450 5794
rect 9662 5742 9714 5794
rect 18510 5742 18562 5794
rect 18958 5742 19010 5794
rect 23326 5742 23378 5794
rect 25230 5742 25282 5794
rect 25902 5742 25954 5794
rect 28702 5742 28754 5794
rect 31950 5742 32002 5794
rect 32398 5742 32450 5794
rect 33742 5742 33794 5794
rect 34750 5742 34802 5794
rect 36318 5742 36370 5794
rect 38446 5742 38498 5794
rect 43822 5742 43874 5794
rect 12014 5630 12066 5682
rect 25342 5630 25394 5682
rect 28814 5630 28866 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 30270 5294 30322 5346
rect 10334 5182 10386 5234
rect 15822 5182 15874 5234
rect 16270 5182 16322 5234
rect 22318 5182 22370 5234
rect 23662 5182 23714 5234
rect 25454 5182 25506 5234
rect 31390 5182 31442 5234
rect 33518 5182 33570 5234
rect 34862 5182 34914 5234
rect 7310 5070 7362 5122
rect 11118 5070 11170 5122
rect 11454 5070 11506 5122
rect 12462 5070 12514 5122
rect 13022 5070 13074 5122
rect 15598 5070 15650 5122
rect 19182 5070 19234 5122
rect 19630 5070 19682 5122
rect 20190 5070 20242 5122
rect 20302 5070 20354 5122
rect 21758 5070 21810 5122
rect 24110 5070 24162 5122
rect 24558 5070 24610 5122
rect 27246 5070 27298 5122
rect 27694 5070 27746 5122
rect 27918 5070 27970 5122
rect 28478 5070 28530 5122
rect 29038 5070 29090 5122
rect 29374 5070 29426 5122
rect 29598 5070 29650 5122
rect 30718 5070 30770 5122
rect 33854 5070 33906 5122
rect 6862 4958 6914 5010
rect 8094 4958 8146 5010
rect 11790 4958 11842 5010
rect 12574 4958 12626 5010
rect 18398 4958 18450 5010
rect 20414 4958 20466 5010
rect 20638 4958 20690 5010
rect 21422 4958 21474 5010
rect 30158 4958 30210 5010
rect 6974 4846 7026 4898
rect 10782 4846 10834 4898
rect 12350 4846 12402 4898
rect 13694 4846 13746 4898
rect 14814 4846 14866 4898
rect 15150 4846 15202 4898
rect 19518 4846 19570 4898
rect 21310 4846 21362 4898
rect 22206 4846 22258 4898
rect 22430 4846 22482 4898
rect 23326 4846 23378 4898
rect 27582 4846 27634 4898
rect 28254 4846 28306 4898
rect 29374 4846 29426 4898
rect 37214 4846 37266 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 8094 4510 8146 4562
rect 10334 4510 10386 4562
rect 14926 4510 14978 4562
rect 19182 4510 19234 4562
rect 19630 4510 19682 4562
rect 32174 4510 32226 4562
rect 33406 4510 33458 4562
rect 37214 4510 37266 4562
rect 8542 4398 8594 4450
rect 9102 4398 9154 4450
rect 9998 4398 10050 4450
rect 11006 4398 11058 4450
rect 11230 4398 11282 4450
rect 19518 4398 19570 4450
rect 19854 4398 19906 4450
rect 20078 4398 20130 4450
rect 20638 4398 20690 4450
rect 27582 4398 27634 4450
rect 29486 4398 29538 4450
rect 34526 4398 34578 4450
rect 41246 4398 41298 4450
rect 7870 4286 7922 4338
rect 8206 4286 8258 4338
rect 9662 4286 9714 4338
rect 10558 4286 10610 4338
rect 11566 4286 11618 4338
rect 18846 4286 18898 4338
rect 20526 4286 20578 4338
rect 21086 4286 21138 4338
rect 21422 4286 21474 4338
rect 28366 4286 28418 4338
rect 28814 4286 28866 4338
rect 32398 4286 32450 4338
rect 33742 4286 33794 4338
rect 37438 4286 37490 4338
rect 7310 4174 7362 4226
rect 7758 4174 7810 4226
rect 9550 4174 9602 4226
rect 10782 4174 10834 4226
rect 12350 4174 12402 4226
rect 14478 4174 14530 4226
rect 18174 4174 18226 4226
rect 18622 4174 18674 4226
rect 20862 4174 20914 4226
rect 22094 4174 22146 4226
rect 24222 4174 24274 4226
rect 25454 4174 25506 4226
rect 31614 4174 31666 4226
rect 33294 4174 33346 4226
rect 36654 4174 36706 4226
rect 37998 4174 38050 4226
rect 42478 4174 42530 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 11566 3614 11618 3666
rect 21870 3614 21922 3666
rect 25566 3614 25618 3666
rect 29374 3614 29426 3666
rect 36990 3614 37042 3666
rect 40798 3614 40850 3666
rect 6862 3502 6914 3554
rect 8430 3502 8482 3554
rect 9326 3502 9378 3554
rect 12126 3502 12178 3554
rect 13358 3502 13410 3554
rect 15934 3502 15986 3554
rect 16942 3502 16994 3554
rect 19854 3502 19906 3554
rect 20750 3502 20802 3554
rect 23886 3502 23938 3554
rect 24670 3502 24722 3554
rect 27358 3502 27410 3554
rect 28590 3502 28642 3554
rect 31614 3502 31666 3554
rect 32174 3502 32226 3554
rect 35422 3502 35474 3554
rect 36430 3502 36482 3554
rect 39790 3502 39842 3554
rect 42926 3502 42978 3554
rect 6414 3390 6466 3442
rect 7086 3390 7138 3442
rect 7422 3390 7474 3442
rect 7758 3390 7810 3442
rect 8094 3390 8146 3442
rect 8766 3390 8818 3442
rect 9662 3390 9714 3442
rect 13134 3390 13186 3442
rect 14814 3390 14866 3442
rect 18510 3390 18562 3442
rect 20190 3390 20242 3442
rect 23662 3390 23714 3442
rect 24894 3390 24946 3442
rect 31278 3390 31330 3442
rect 33742 3390 33794 3442
rect 35086 3390 35138 3442
rect 42702 3390 42754 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 9408 49200 9520 50000
rect 10080 49200 10192 50000
rect 12096 49200 12208 50000
rect 12768 49200 12880 50000
rect 13440 49200 13552 50000
rect 14784 49200 14896 50000
rect 15456 49200 15568 50000
rect 16128 49200 16240 50000
rect 16800 49200 16912 50000
rect 17472 49200 17584 50000
rect 18144 49200 18256 50000
rect 18816 49200 18928 50000
rect 19488 49200 19600 50000
rect 22848 49200 22960 50000
rect 23520 49200 23632 50000
rect 24192 49200 24304 50000
rect 24864 49200 24976 50000
rect 26880 49200 26992 50000
rect 27552 49200 27664 50000
rect 28224 49200 28336 50000
rect 28896 49200 29008 50000
rect 32928 49200 33040 50000
rect 33600 49200 33712 50000
rect 34944 49200 35056 50000
rect 40320 49200 40432 50000
rect 40992 49200 41104 50000
rect 41664 49200 41776 50000
rect 42336 49200 42448 50000
rect 43008 49200 43120 50000
rect 43680 49200 43792 50000
rect 44352 49200 44464 50000
rect 44716 49812 44772 49822
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 8876 46004 8932 46014
rect 9436 46004 9492 49200
rect 8876 46002 9492 46004
rect 8876 45950 8878 46002
rect 8930 45950 9492 46002
rect 8876 45948 9492 45950
rect 8876 45938 8932 45948
rect 9436 45892 9492 45948
rect 10108 46788 10164 49200
rect 12124 46788 12180 49200
rect 10108 46732 10612 46788
rect 9660 45892 9716 45902
rect 9436 45890 9716 45892
rect 9436 45838 9662 45890
rect 9714 45838 9716 45890
rect 9436 45836 9716 45838
rect 9660 45826 9716 45836
rect 9996 45668 10052 45678
rect 9772 45666 10052 45668
rect 9772 45614 9998 45666
rect 10050 45614 10052 45666
rect 9772 45612 10052 45614
rect 4172 45108 4228 45118
rect 1932 43314 1988 43326
rect 1932 43262 1934 43314
rect 1986 43262 1988 43314
rect 1932 42420 1988 43262
rect 1932 42354 1988 42364
rect 2044 42866 2100 42878
rect 2044 42814 2046 42866
rect 2098 42814 2100 42866
rect 1932 41746 1988 41758
rect 1932 41694 1934 41746
rect 1986 41694 1988 41746
rect 1708 41186 1764 41198
rect 1708 41134 1710 41186
rect 1762 41134 1764 41186
rect 1708 40964 1764 41134
rect 1708 40898 1764 40908
rect 1932 40404 1988 41694
rect 2044 41748 2100 42814
rect 2044 41682 2100 41692
rect 4060 42754 4116 42766
rect 4060 42702 4062 42754
rect 4114 42702 4116 42754
rect 1932 40338 1988 40348
rect 2492 41074 2548 41086
rect 2492 41022 2494 41074
rect 2546 41022 2548 41074
rect 1932 40178 1988 40190
rect 1932 40126 1934 40178
rect 1986 40126 1988 40178
rect 1932 39732 1988 40126
rect 1932 39666 1988 39676
rect 2492 39730 2548 41022
rect 2492 39678 2494 39730
rect 2546 39678 2548 39730
rect 2492 39666 2548 39678
rect 3724 39618 3780 39630
rect 3724 39566 3726 39618
rect 3778 39566 3780 39618
rect 2156 39508 2212 39518
rect 2380 39508 2436 39518
rect 2492 39508 2548 39518
rect 2156 39506 2492 39508
rect 2156 39454 2158 39506
rect 2210 39454 2382 39506
rect 2434 39454 2492 39506
rect 2156 39452 2492 39454
rect 2156 39442 2212 39452
rect 2380 39442 2436 39452
rect 2380 39060 2436 39070
rect 2380 38722 2436 39004
rect 2380 38670 2382 38722
rect 2434 38670 2436 38722
rect 2268 38610 2324 38622
rect 2268 38558 2270 38610
rect 2322 38558 2324 38610
rect 2268 38276 2324 38558
rect 2380 38388 2436 38670
rect 2492 38500 2548 39452
rect 2604 39394 2660 39406
rect 2604 39342 2606 39394
rect 2658 39342 2660 39394
rect 2604 38948 2660 39342
rect 3276 39394 3332 39406
rect 3276 39342 3278 39394
rect 3330 39342 3332 39394
rect 3164 39060 3220 39070
rect 3276 39060 3332 39342
rect 3220 39004 3332 39060
rect 3724 39060 3780 39566
rect 4060 39396 4116 42702
rect 4060 39330 4116 39340
rect 3164 38994 3220 39004
rect 2604 38882 2660 38892
rect 3612 38948 3668 38958
rect 3612 38854 3668 38892
rect 3724 38946 3780 39004
rect 3724 38894 3726 38946
rect 3778 38894 3780 38946
rect 3724 38882 3780 38894
rect 2716 38836 2772 38846
rect 2716 38742 2772 38780
rect 3948 38834 4004 38846
rect 3948 38782 3950 38834
rect 4002 38782 4004 38834
rect 2604 38722 2660 38734
rect 2604 38670 2606 38722
rect 2658 38670 2660 38722
rect 2604 38612 2660 38670
rect 3164 38722 3220 38734
rect 3164 38670 3166 38722
rect 3218 38670 3220 38722
rect 3164 38612 3220 38670
rect 3948 38724 4004 38782
rect 3948 38658 4004 38668
rect 2604 38556 3220 38612
rect 2492 38444 3108 38500
rect 2380 38332 2660 38388
rect 2268 38220 2548 38276
rect 2492 38162 2548 38220
rect 2492 38110 2494 38162
rect 2546 38110 2548 38162
rect 2492 38098 2548 38110
rect 1820 38050 1876 38062
rect 1820 37998 1822 38050
rect 1874 37998 1876 38050
rect 1820 35698 1876 37998
rect 2604 37492 2660 38332
rect 2380 37436 2660 37492
rect 1932 37044 1988 37054
rect 1932 36950 1988 36988
rect 1932 36596 1988 36606
rect 1932 36502 1988 36540
rect 1820 35646 1822 35698
rect 1874 35646 1876 35698
rect 1820 35588 1876 35646
rect 1820 35522 1876 35532
rect 1932 35026 1988 35038
rect 1932 34974 1934 35026
rect 1986 34974 1988 35026
rect 1708 34356 1764 34366
rect 1708 34242 1764 34300
rect 1708 34190 1710 34242
rect 1762 34190 1764 34242
rect 1708 34178 1764 34190
rect 1932 33684 1988 34974
rect 2044 34468 2100 34478
rect 2044 34354 2100 34412
rect 2044 34302 2046 34354
rect 2098 34302 2100 34354
rect 2044 34290 2100 34302
rect 1932 33618 1988 33628
rect 1820 33348 1876 33358
rect 1820 33254 1876 33292
rect 1820 30994 1876 31006
rect 1820 30942 1822 30994
rect 1874 30942 1876 30994
rect 1820 27860 1876 30942
rect 1820 25506 1876 27804
rect 2380 27636 2436 37436
rect 2492 35700 2548 35710
rect 2492 35606 2548 35644
rect 2492 34356 2548 34366
rect 2492 34262 2548 34300
rect 2492 33236 2548 33246
rect 2492 33234 2884 33236
rect 2492 33182 2494 33234
rect 2546 33182 2884 33234
rect 2492 33180 2884 33182
rect 2492 33170 2548 33180
rect 2828 32450 2884 33180
rect 2940 32788 2996 32798
rect 2940 32694 2996 32732
rect 2828 32398 2830 32450
rect 2882 32398 2884 32450
rect 2828 32386 2884 32398
rect 3052 31948 3108 38444
rect 3164 37044 3220 38556
rect 3164 36978 3220 36988
rect 3948 35364 4004 35374
rect 3948 34130 4004 35308
rect 3948 34078 3950 34130
rect 4002 34078 4004 34130
rect 3948 33348 4004 34078
rect 3164 32452 3220 32462
rect 3612 32452 3668 32462
rect 3164 32450 3668 32452
rect 3164 32398 3166 32450
rect 3218 32398 3614 32450
rect 3666 32398 3668 32450
rect 3164 32396 3668 32398
rect 3164 32386 3220 32396
rect 3612 32340 3668 32396
rect 3948 32452 4004 33292
rect 3948 32386 4004 32396
rect 3612 32274 3668 32284
rect 3052 31892 3220 31948
rect 2492 30882 2548 30894
rect 2492 30830 2494 30882
rect 2546 30830 2548 30882
rect 2492 30436 2548 30830
rect 2828 30772 2884 30782
rect 2716 30436 2772 30446
rect 2492 30434 2772 30436
rect 2492 30382 2718 30434
rect 2770 30382 2772 30434
rect 2492 30380 2772 30382
rect 2716 30370 2772 30380
rect 2828 30434 2884 30716
rect 3052 30436 3108 30446
rect 2828 30382 2830 30434
rect 2882 30382 2884 30434
rect 2828 30370 2884 30382
rect 2940 30434 3108 30436
rect 2940 30382 3054 30434
rect 3106 30382 3108 30434
rect 2940 30380 3108 30382
rect 2828 29426 2884 29438
rect 2828 29374 2830 29426
rect 2882 29374 2884 29426
rect 2604 29314 2660 29326
rect 2604 29262 2606 29314
rect 2658 29262 2660 29314
rect 2492 29202 2548 29214
rect 2492 29150 2494 29202
rect 2546 29150 2548 29202
rect 2492 28866 2548 29150
rect 2492 28814 2494 28866
rect 2546 28814 2548 28866
rect 2492 28802 2548 28814
rect 2492 27972 2548 27982
rect 2604 27972 2660 29262
rect 2828 29316 2884 29374
rect 2828 29250 2884 29260
rect 2940 28756 2996 30380
rect 3052 30370 3108 30380
rect 3164 29316 3220 31892
rect 3276 31890 3332 31902
rect 3276 31838 3278 31890
rect 3330 31838 3332 31890
rect 3276 30210 3332 31838
rect 3612 31892 3668 31902
rect 3612 31798 3668 31836
rect 3388 31554 3444 31566
rect 3388 31502 3390 31554
rect 3442 31502 3444 31554
rect 3388 30436 3444 31502
rect 3388 30370 3444 30380
rect 3276 30158 3278 30210
rect 3330 30158 3332 30210
rect 3276 30146 3332 30158
rect 3948 29988 4004 29998
rect 3276 29316 3332 29326
rect 3164 29260 3276 29316
rect 3276 29222 3332 29260
rect 2940 28662 2996 28700
rect 3052 28868 3108 28878
rect 3052 28642 3108 28812
rect 3724 28868 3780 28878
rect 3724 28754 3780 28812
rect 3724 28702 3726 28754
rect 3778 28702 3780 28754
rect 3724 28690 3780 28702
rect 3948 28756 4004 29932
rect 4172 29764 4228 45052
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4284 43540 4340 43550
rect 4844 43540 4900 43550
rect 4284 43538 4844 43540
rect 4284 43486 4286 43538
rect 4338 43486 4844 43538
rect 4284 43484 4844 43486
rect 4284 43474 4340 43484
rect 4844 43446 4900 43484
rect 8764 43540 8820 43550
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 8204 42754 8260 42766
rect 8204 42702 8206 42754
rect 8258 42702 8260 42754
rect 8204 42084 8260 42702
rect 8204 42018 8260 42028
rect 4284 41970 4340 41982
rect 4284 41918 4286 41970
rect 4338 41918 4340 41970
rect 4284 40740 4340 41918
rect 5292 41972 5348 41982
rect 6188 41972 6244 41982
rect 5292 41970 5460 41972
rect 5292 41918 5294 41970
rect 5346 41918 5460 41970
rect 5292 41916 5460 41918
rect 5292 41906 5348 41916
rect 5404 41860 5460 41916
rect 5740 41860 5796 41870
rect 5404 41858 5796 41860
rect 5404 41806 5742 41858
rect 5794 41806 5796 41858
rect 5404 41804 5796 41806
rect 4956 41748 5012 41758
rect 4956 41654 5012 41692
rect 5292 41748 5348 41758
rect 5292 41654 5348 41692
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 5404 41524 5460 41804
rect 5740 41794 5796 41804
rect 4476 41514 4740 41524
rect 5292 41468 5460 41524
rect 4620 41300 4676 41310
rect 4620 41298 5012 41300
rect 4620 41246 4622 41298
rect 4674 41246 5012 41298
rect 4620 41244 5012 41246
rect 4620 41234 4676 41244
rect 4284 40674 4340 40684
rect 4284 40516 4340 40526
rect 4284 40402 4340 40460
rect 4284 40350 4286 40402
rect 4338 40350 4340 40402
rect 4284 40338 4340 40350
rect 4620 40514 4676 40526
rect 4620 40462 4622 40514
rect 4674 40462 4676 40514
rect 4620 40180 4676 40462
rect 4284 40124 4676 40180
rect 4956 40402 5012 41244
rect 5068 40964 5124 40974
rect 5124 40908 5236 40964
rect 5068 40870 5124 40908
rect 4956 40350 4958 40402
rect 5010 40350 5012 40402
rect 4284 39730 4340 40124
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4396 39844 4452 39854
rect 4396 39750 4452 39788
rect 4284 39678 4286 39730
rect 4338 39678 4340 39730
rect 4284 38948 4340 39678
rect 4284 38854 4340 38892
rect 4620 38948 4676 38958
rect 4620 38854 4676 38892
rect 4396 38836 4452 38846
rect 4396 38742 4452 38780
rect 4844 38836 4900 38846
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4620 38164 4676 38174
rect 4620 38070 4676 38108
rect 4844 37492 4900 38780
rect 4956 38052 5012 40350
rect 5068 40516 5124 40526
rect 5068 39730 5124 40460
rect 5068 39678 5070 39730
rect 5122 39678 5124 39730
rect 5068 39666 5124 39678
rect 5180 40404 5236 40908
rect 5180 38668 5236 40348
rect 5292 39508 5348 41468
rect 5740 41188 5796 41198
rect 6188 41188 6244 41916
rect 6300 41748 6356 41758
rect 6356 41692 6468 41748
rect 6300 41682 6356 41692
rect 6412 41298 6468 41692
rect 6412 41246 6414 41298
rect 6466 41246 6468 41298
rect 6412 41234 6468 41246
rect 8540 41298 8596 41310
rect 8540 41246 8542 41298
rect 8594 41246 8596 41298
rect 5740 41186 6244 41188
rect 5740 41134 5742 41186
rect 5794 41134 6244 41186
rect 5740 41132 6244 41134
rect 5740 41122 5796 41132
rect 5740 40628 5796 40638
rect 5796 40572 6020 40628
rect 5740 40534 5796 40572
rect 5292 39442 5348 39452
rect 5404 40514 5460 40526
rect 5404 40462 5406 40514
rect 5458 40462 5460 40514
rect 5404 38948 5460 40462
rect 5404 38882 5460 38892
rect 4956 37986 5012 37996
rect 5068 38612 5236 38668
rect 5068 37826 5124 38612
rect 5068 37774 5070 37826
rect 5122 37774 5124 37826
rect 4956 37492 5012 37502
rect 4844 37490 5012 37492
rect 4844 37438 4958 37490
rect 5010 37438 5012 37490
rect 4844 37436 5012 37438
rect 4956 37426 5012 37436
rect 4284 37268 4340 37278
rect 4284 37174 4340 37212
rect 4284 37044 4340 37054
rect 4284 36708 4340 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4620 36708 4676 36718
rect 4284 36706 4676 36708
rect 4284 36654 4622 36706
rect 4674 36654 4676 36706
rect 4284 36652 4676 36654
rect 4620 36642 4676 36652
rect 4956 36594 5012 36606
rect 4956 36542 4958 36594
rect 5010 36542 5012 36594
rect 4284 36482 4340 36494
rect 4284 36430 4286 36482
rect 4338 36430 4340 36482
rect 4284 36260 4340 36430
rect 4844 36484 4900 36494
rect 4844 36372 4900 36428
rect 4284 36194 4340 36204
rect 4620 36370 4900 36372
rect 4620 36318 4846 36370
rect 4898 36318 4900 36370
rect 4620 36316 4900 36318
rect 4620 35586 4676 36316
rect 4844 36306 4900 36316
rect 4956 35698 5012 36542
rect 4956 35646 4958 35698
rect 5010 35646 5012 35698
rect 4956 35634 5012 35646
rect 4620 35534 4622 35586
rect 4674 35534 4676 35586
rect 4620 35522 4676 35534
rect 5068 35476 5124 37774
rect 5180 38164 5236 38174
rect 5180 37266 5236 38108
rect 5740 38164 5796 38174
rect 5628 38050 5684 38062
rect 5628 37998 5630 38050
rect 5682 37998 5684 38050
rect 5516 37828 5572 37838
rect 5180 37214 5182 37266
rect 5234 37214 5236 37266
rect 5180 37202 5236 37214
rect 5292 37772 5516 37828
rect 5068 35410 5124 35420
rect 5180 35588 5236 35598
rect 5292 35588 5348 37772
rect 5516 37762 5572 37772
rect 5628 36484 5684 37998
rect 5740 37938 5796 38108
rect 5964 38050 6020 40572
rect 6076 40516 6132 40526
rect 6076 38668 6132 40460
rect 6188 40404 6244 41132
rect 7196 40628 7252 40638
rect 7084 40572 7196 40628
rect 6860 40516 6916 40526
rect 6860 40422 6916 40460
rect 6188 40310 6244 40348
rect 7084 39060 7140 40572
rect 7196 40562 7252 40572
rect 8540 40628 8596 41246
rect 8540 40562 8596 40572
rect 7532 39506 7588 39518
rect 7532 39454 7534 39506
rect 7586 39454 7588 39506
rect 7308 39060 7364 39070
rect 7084 39058 7364 39060
rect 7084 39006 7310 39058
rect 7362 39006 7364 39058
rect 7084 39004 7364 39006
rect 7308 38994 7364 39004
rect 6412 38836 6468 38846
rect 6412 38742 6468 38780
rect 6748 38834 6804 38846
rect 7532 38836 7588 39454
rect 8092 39396 8148 39406
rect 8092 39394 8260 39396
rect 8092 39342 8094 39394
rect 8146 39342 8260 39394
rect 8092 39340 8260 39342
rect 8092 39330 8148 39340
rect 6748 38782 6750 38834
rect 6802 38782 6804 38834
rect 6636 38722 6692 38734
rect 6636 38670 6638 38722
rect 6690 38670 6692 38722
rect 6076 38612 6244 38668
rect 5964 37998 5966 38050
rect 6018 37998 6020 38050
rect 5964 37986 6020 37998
rect 5740 37886 5742 37938
rect 5794 37886 5796 37938
rect 5740 37874 5796 37886
rect 5740 36484 5796 36494
rect 5684 36482 5796 36484
rect 5684 36430 5742 36482
rect 5794 36430 5796 36482
rect 5684 36428 5796 36430
rect 5628 36390 5684 36428
rect 5740 36418 5796 36428
rect 5852 36484 5908 36494
rect 5852 36390 5908 36428
rect 5516 35700 5572 35710
rect 5516 35606 5572 35644
rect 5180 35586 5348 35588
rect 5180 35534 5182 35586
rect 5234 35534 5348 35586
rect 5180 35532 5348 35534
rect 5964 35586 6020 35598
rect 5964 35534 5966 35586
rect 6018 35534 6020 35586
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4284 34916 4340 34926
rect 4732 34916 4788 34926
rect 4284 34914 4788 34916
rect 4284 34862 4286 34914
rect 4338 34862 4734 34914
rect 4786 34862 4788 34914
rect 4284 34860 4788 34862
rect 4284 33012 4340 34860
rect 4732 34850 4788 34860
rect 4620 34020 4676 34030
rect 4620 34018 4900 34020
rect 4620 33966 4622 34018
rect 4674 33966 4900 34018
rect 4620 33964 4900 33966
rect 4620 33954 4676 33964
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4284 32946 4340 32956
rect 4732 33122 4788 33134
rect 4732 33070 4734 33122
rect 4786 33070 4788 33122
rect 4732 32564 4788 33070
rect 4844 32676 4900 33964
rect 4956 32788 5012 32798
rect 4956 32694 5012 32732
rect 4844 32610 4900 32620
rect 4732 32498 4788 32508
rect 4620 32452 4676 32462
rect 4620 32340 4676 32396
rect 4620 32284 4900 32340
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4844 32004 4900 32284
rect 4844 31938 4900 31948
rect 4396 31892 4452 31902
rect 4284 31836 4396 31892
rect 4284 30436 4340 31836
rect 4396 31826 4452 31836
rect 5180 31892 5236 35532
rect 5404 35474 5460 35486
rect 5404 35422 5406 35474
rect 5458 35422 5460 35474
rect 5292 32564 5348 32574
rect 5292 32470 5348 32508
rect 5180 31826 5236 31836
rect 4620 30882 4676 30894
rect 4620 30830 4622 30882
rect 4674 30830 4676 30882
rect 4620 30772 4676 30830
rect 4620 30716 5012 30772
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4620 30436 4676 30446
rect 4284 30434 4676 30436
rect 4284 30382 4622 30434
rect 4674 30382 4676 30434
rect 4284 30380 4676 30382
rect 4620 30324 4676 30380
rect 4620 30258 4676 30268
rect 4844 30436 4900 30446
rect 4844 30210 4900 30380
rect 4844 30158 4846 30210
rect 4898 30158 4900 30210
rect 4844 30146 4900 30158
rect 4284 29988 4340 29998
rect 4956 29988 5012 30716
rect 5404 30548 5460 35422
rect 5964 35476 6020 35534
rect 5964 35410 6020 35420
rect 6188 35476 6244 38612
rect 6412 38052 6468 38062
rect 6412 37380 6468 37996
rect 6636 38052 6692 38670
rect 6748 38164 6804 38782
rect 6748 38098 6804 38108
rect 7196 38834 7588 38836
rect 7196 38782 7534 38834
rect 7586 38782 7588 38834
rect 7196 38780 7588 38782
rect 6636 37986 6692 37996
rect 6636 37828 6692 37838
rect 6636 37734 6692 37772
rect 6636 37380 6692 37390
rect 6412 37378 6692 37380
rect 6412 37326 6638 37378
rect 6690 37326 6692 37378
rect 6412 37324 6692 37326
rect 6636 37314 6692 37324
rect 7084 37266 7140 37278
rect 7084 37214 7086 37266
rect 7138 37214 7140 37266
rect 7084 36708 7140 37214
rect 7196 36708 7252 38780
rect 7532 38770 7588 38780
rect 7756 38948 7812 38958
rect 7420 38612 7476 38622
rect 7308 38556 7420 38612
rect 7308 38050 7364 38556
rect 7420 38546 7476 38556
rect 7308 37998 7310 38050
rect 7362 37998 7364 38050
rect 7308 37986 7364 37998
rect 7532 37938 7588 37950
rect 7532 37886 7534 37938
rect 7586 37886 7588 37938
rect 7532 37378 7588 37886
rect 7532 37326 7534 37378
rect 7586 37326 7588 37378
rect 7532 37314 7588 37326
rect 7644 37940 7700 37950
rect 7196 36652 7588 36708
rect 7084 36642 7140 36652
rect 7196 36484 7252 36494
rect 7084 36482 7252 36484
rect 7084 36430 7198 36482
rect 7250 36430 7252 36482
rect 7084 36428 7252 36430
rect 6188 35410 6244 35420
rect 6300 36260 6356 36270
rect 6300 34468 6356 36204
rect 6860 34580 6916 34590
rect 6300 34412 6692 34468
rect 5516 33404 5796 33460
rect 5516 32788 5572 33404
rect 5740 33348 5796 33404
rect 5740 33254 5796 33292
rect 6300 33346 6356 33358
rect 6300 33294 6302 33346
rect 6354 33294 6356 33346
rect 5628 33234 5684 33246
rect 5628 33182 5630 33234
rect 5682 33182 5684 33234
rect 5628 32900 5684 33182
rect 6300 33124 6356 33294
rect 6300 33058 6356 33068
rect 5628 32844 6020 32900
rect 5516 32722 5572 32732
rect 5852 32676 5908 32686
rect 5852 32582 5908 32620
rect 5964 32674 6020 32844
rect 5964 32622 5966 32674
rect 6018 32622 6020 32674
rect 5964 32610 6020 32622
rect 5628 32562 5684 32574
rect 5628 32510 5630 32562
rect 5682 32510 5684 32562
rect 5628 32340 5684 32510
rect 6412 32452 6468 32462
rect 6412 32450 6580 32452
rect 6412 32398 6414 32450
rect 6466 32398 6580 32450
rect 6412 32396 6580 32398
rect 6412 32386 6468 32396
rect 5628 32274 5684 32284
rect 6524 32340 6580 32396
rect 5740 31892 5796 31902
rect 5740 31778 5796 31836
rect 5740 31726 5742 31778
rect 5794 31726 5796 31778
rect 5740 31714 5796 31726
rect 6412 31666 6468 31678
rect 6412 31614 6414 31666
rect 6466 31614 6468 31666
rect 6412 31556 6468 31614
rect 6412 31490 6468 31500
rect 5404 30482 5460 30492
rect 6188 30548 6244 30558
rect 5964 30436 6020 30446
rect 5964 30098 6020 30380
rect 5964 30046 5966 30098
rect 6018 30046 6020 30098
rect 5964 30034 6020 30046
rect 5628 29988 5684 29998
rect 4956 29986 5684 29988
rect 4956 29934 5630 29986
rect 5682 29934 5684 29986
rect 4956 29932 5684 29934
rect 4284 29894 4340 29932
rect 4172 29708 4340 29764
rect 3948 28690 4004 28700
rect 3052 28590 3054 28642
rect 3106 28590 3108 28642
rect 3052 28578 3108 28590
rect 4172 28644 4228 28654
rect 4172 28550 4228 28588
rect 2492 27970 2660 27972
rect 2492 27918 2494 27970
rect 2546 27918 2660 27970
rect 2492 27916 2660 27918
rect 2492 27906 2548 27916
rect 2380 27570 2436 27580
rect 2492 26068 2548 26078
rect 2492 25618 2548 26012
rect 2492 25566 2494 25618
rect 2546 25566 2548 25618
rect 2492 25554 2548 25566
rect 1820 25454 1822 25506
rect 1874 25454 1876 25506
rect 1820 25442 1876 25454
rect 4172 24722 4228 24734
rect 4172 24670 4174 24722
rect 4226 24670 4228 24722
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 4172 24500 4228 24670
rect 4284 24724 4340 29708
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4844 28980 4900 28990
rect 4396 28756 4452 28766
rect 4732 28756 4788 28766
rect 4396 28642 4452 28700
rect 4620 28700 4732 28756
rect 4396 28590 4398 28642
rect 4450 28590 4452 28642
rect 4396 28578 4452 28590
rect 4508 28644 4564 28654
rect 4508 27748 4564 28588
rect 4620 28642 4676 28700
rect 4732 28690 4788 28700
rect 4620 28590 4622 28642
rect 4674 28590 4676 28642
rect 4620 28578 4676 28590
rect 4844 28642 4900 28924
rect 5628 28868 5684 29932
rect 5852 29202 5908 29214
rect 5852 29150 5854 29202
rect 5906 29150 5908 29202
rect 5740 28868 5796 28878
rect 5628 28812 5740 28868
rect 5740 28802 5796 28812
rect 5852 28756 5908 29150
rect 5964 29204 6020 29214
rect 5964 29202 6132 29204
rect 5964 29150 5966 29202
rect 6018 29150 6132 29202
rect 5964 29148 6132 29150
rect 5964 29138 6020 29148
rect 6076 29092 6132 29148
rect 5852 28690 5908 28700
rect 5964 28868 6020 28878
rect 4844 28590 4846 28642
rect 4898 28590 4900 28642
rect 4844 28578 4900 28590
rect 5068 28644 5124 28654
rect 5628 28644 5684 28654
rect 5068 28642 5684 28644
rect 5068 28590 5070 28642
rect 5122 28590 5630 28642
rect 5682 28590 5684 28642
rect 5068 28588 5684 28590
rect 5068 28578 5124 28588
rect 4620 27748 4676 27758
rect 4508 27746 4676 27748
rect 4508 27694 4622 27746
rect 4674 27694 4676 27746
rect 4508 27692 4676 27694
rect 4620 27682 4676 27692
rect 5628 27748 5684 28588
rect 5740 28644 5796 28654
rect 5740 28530 5796 28588
rect 5964 28642 6020 28812
rect 5964 28590 5966 28642
rect 6018 28590 6020 28642
rect 5964 28578 6020 28590
rect 5740 28478 5742 28530
rect 5794 28478 5796 28530
rect 5740 28466 5796 28478
rect 5852 27860 5908 27870
rect 5852 27766 5908 27804
rect 5628 27682 5684 27692
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 6076 26908 6132 29036
rect 5964 26852 6132 26908
rect 6188 29202 6244 30492
rect 6300 30324 6356 30334
rect 6356 30268 6468 30324
rect 6300 30258 6356 30268
rect 6188 29150 6190 29202
rect 6242 29150 6244 29202
rect 5068 26460 5684 26516
rect 4844 26292 4900 26302
rect 4844 26198 4900 26236
rect 5068 26290 5124 26460
rect 5068 26238 5070 26290
rect 5122 26238 5124 26290
rect 5068 26226 5124 26238
rect 5292 26292 5348 26302
rect 5292 26290 5572 26292
rect 5292 26238 5294 26290
rect 5346 26238 5572 26290
rect 5292 26236 5572 26238
rect 5292 26226 5348 26236
rect 4732 26068 4788 26106
rect 4732 26002 4788 26012
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 5516 25732 5572 26236
rect 5628 26068 5684 26460
rect 5964 26290 6020 26852
rect 6188 26516 6244 29150
rect 6300 29202 6356 29214
rect 6300 29150 6302 29202
rect 6354 29150 6356 29202
rect 6300 28084 6356 29150
rect 6412 28642 6468 30268
rect 6524 29540 6580 32284
rect 6636 30772 6692 34412
rect 6860 34354 6916 34524
rect 6860 34302 6862 34354
rect 6914 34302 6916 34354
rect 6860 34290 6916 34302
rect 7084 31220 7140 36428
rect 7196 36418 7252 36428
rect 7532 36372 7588 36652
rect 7644 36482 7700 37884
rect 7756 37154 7812 38892
rect 8204 38948 8260 39340
rect 7980 38836 8036 38846
rect 7868 38724 7924 38762
rect 7980 38742 8036 38780
rect 7868 38658 7924 38668
rect 8092 37268 8148 37278
rect 8204 37268 8260 38892
rect 8316 38946 8372 38958
rect 8316 38894 8318 38946
rect 8370 38894 8372 38946
rect 8316 38836 8372 38894
rect 8764 38836 8820 43484
rect 8876 43428 8932 43438
rect 8876 42866 8932 43372
rect 8876 42814 8878 42866
rect 8930 42814 8932 42866
rect 8876 42802 8932 42814
rect 8988 42084 9044 42094
rect 8988 40964 9044 42028
rect 8988 40962 9156 40964
rect 8988 40910 8990 40962
rect 9042 40910 9156 40962
rect 8988 40908 9156 40910
rect 8988 40898 9044 40908
rect 8988 40628 9044 40638
rect 8988 40290 9044 40572
rect 8988 40238 8990 40290
rect 9042 40238 9044 40290
rect 8988 39284 9044 40238
rect 9100 39396 9156 40908
rect 9772 40514 9828 45612
rect 9996 45602 10052 45612
rect 10108 45330 10164 46732
rect 10556 45890 10612 46732
rect 10556 45838 10558 45890
rect 10610 45838 10612 45890
rect 10556 45826 10612 45838
rect 11676 46732 12180 46788
rect 11676 45890 11732 46732
rect 11676 45838 11678 45890
rect 11730 45838 11732 45890
rect 11676 45826 11732 45838
rect 10332 45668 10388 45678
rect 10108 45278 10110 45330
rect 10162 45278 10164 45330
rect 10108 45266 10164 45278
rect 10220 45666 10388 45668
rect 10220 45614 10334 45666
rect 10386 45614 10388 45666
rect 10220 45612 10388 45614
rect 10220 43764 10276 45612
rect 10332 45602 10388 45612
rect 11900 45668 11956 45678
rect 11900 45666 12068 45668
rect 11900 45614 11902 45666
rect 11954 45614 12068 45666
rect 11900 45612 12068 45614
rect 11900 45602 11956 45612
rect 9996 43708 10276 43764
rect 9996 41970 10052 43708
rect 10108 43538 10164 43550
rect 10108 43486 10110 43538
rect 10162 43486 10164 43538
rect 10108 42194 10164 43486
rect 10556 43538 10612 43550
rect 10556 43486 10558 43538
rect 10610 43486 10612 43538
rect 10332 43428 10388 43438
rect 10332 43334 10388 43372
rect 10108 42142 10110 42194
rect 10162 42142 10164 42194
rect 10108 42130 10164 42142
rect 10556 42196 10612 43486
rect 10780 43540 10836 43550
rect 11900 43540 11956 43550
rect 10780 43538 11172 43540
rect 10780 43486 10782 43538
rect 10834 43486 11172 43538
rect 10780 43484 11172 43486
rect 10780 43474 10836 43484
rect 11004 42868 11060 42878
rect 10556 42130 10612 42140
rect 10892 42866 11060 42868
rect 10892 42814 11006 42866
rect 11058 42814 11060 42866
rect 10892 42812 11060 42814
rect 9996 41918 9998 41970
rect 10050 41918 10052 41970
rect 9996 41906 10052 41918
rect 10892 41970 10948 42812
rect 11004 42802 11060 42812
rect 11116 42644 11172 43484
rect 11004 42588 11172 42644
rect 11004 42194 11060 42588
rect 11452 42532 11508 42542
rect 11004 42142 11006 42194
rect 11058 42142 11060 42194
rect 11004 42130 11060 42142
rect 11340 42530 11508 42532
rect 11340 42478 11454 42530
rect 11506 42478 11508 42530
rect 11340 42476 11508 42478
rect 11116 42084 11172 42094
rect 11116 41990 11172 42028
rect 10892 41918 10894 41970
rect 10946 41918 10948 41970
rect 9772 40462 9774 40514
rect 9826 40462 9828 40514
rect 9772 40450 9828 40462
rect 10108 40740 10164 40750
rect 9884 40404 9940 40414
rect 9884 40310 9940 40348
rect 10108 39620 10164 40684
rect 10668 40740 10724 40750
rect 10220 40628 10276 40638
rect 10220 40534 10276 40572
rect 10668 40290 10724 40684
rect 10668 40238 10670 40290
rect 10722 40238 10724 40290
rect 10668 40226 10724 40238
rect 10556 39620 10612 39630
rect 10108 39618 10276 39620
rect 10108 39566 10110 39618
rect 10162 39566 10276 39618
rect 10108 39564 10276 39566
rect 10108 39554 10164 39564
rect 9212 39396 9268 39406
rect 9100 39394 9268 39396
rect 9100 39342 9214 39394
rect 9266 39342 9268 39394
rect 9100 39340 9268 39342
rect 8988 39228 9156 39284
rect 8988 38836 9044 38846
rect 8764 38834 9044 38836
rect 8764 38782 8990 38834
rect 9042 38782 9044 38834
rect 8764 38780 9044 38782
rect 8316 38770 8372 38780
rect 8988 38612 9044 38780
rect 8988 38546 9044 38556
rect 8652 38052 8708 38062
rect 8652 37958 8708 37996
rect 8092 37266 8260 37268
rect 8092 37214 8094 37266
rect 8146 37214 8260 37266
rect 8092 37212 8260 37214
rect 8092 37202 8148 37212
rect 7756 37102 7758 37154
rect 7810 37102 7812 37154
rect 7756 37090 7812 37102
rect 8988 36708 9044 36718
rect 7644 36430 7646 36482
rect 7698 36430 7700 36482
rect 7644 36418 7700 36430
rect 7868 36484 7924 36494
rect 7868 36390 7924 36428
rect 8316 36372 8372 36382
rect 7532 35698 7588 36316
rect 7980 36370 8372 36372
rect 7980 36318 8318 36370
rect 8370 36318 8372 36370
rect 7980 36316 8372 36318
rect 7532 35646 7534 35698
rect 7586 35646 7588 35698
rect 7532 35634 7588 35646
rect 7756 36258 7812 36270
rect 7756 36206 7758 36258
rect 7810 36206 7812 36258
rect 7756 35364 7812 36206
rect 7980 35588 8036 36316
rect 8316 36306 8372 36316
rect 8428 36372 8484 36382
rect 8484 36316 8596 36372
rect 8428 36278 8484 36316
rect 8540 36036 8596 36316
rect 8652 36260 8708 36270
rect 8652 36166 8708 36204
rect 8540 35980 8708 36036
rect 7756 35298 7812 35308
rect 7868 35586 8036 35588
rect 7868 35534 7982 35586
rect 8034 35534 8036 35586
rect 7868 35532 8036 35534
rect 7420 34580 7476 34590
rect 7308 34524 7420 34580
rect 7308 34354 7364 34524
rect 7420 34514 7476 34524
rect 7644 34356 7700 34366
rect 7868 34356 7924 35532
rect 7980 35522 8036 35532
rect 8316 35700 8372 35710
rect 8316 35474 8372 35644
rect 8316 35422 8318 35474
rect 8370 35422 8372 35474
rect 8316 35410 8372 35422
rect 8540 35364 8596 35374
rect 8428 34580 8484 34590
rect 7308 34302 7310 34354
rect 7362 34302 7364 34354
rect 7308 34290 7364 34302
rect 7420 34354 7924 34356
rect 7420 34302 7646 34354
rect 7698 34302 7924 34354
rect 7420 34300 7924 34302
rect 8316 34524 8428 34580
rect 7420 33460 7476 34300
rect 7644 34290 7700 34300
rect 8092 34018 8148 34030
rect 8092 33966 8094 34018
rect 8146 33966 8148 34018
rect 8092 33908 8148 33966
rect 7420 33366 7476 33404
rect 7644 33852 8148 33908
rect 7196 33236 7252 33246
rect 7196 32562 7252 33180
rect 7308 33124 7364 33134
rect 7308 33030 7364 33068
rect 7196 32510 7198 32562
rect 7250 32510 7252 32562
rect 7196 32498 7252 32510
rect 7644 31892 7700 33852
rect 8204 33236 8260 33246
rect 8204 33142 8260 33180
rect 8316 33124 8372 34524
rect 8428 34514 8484 34524
rect 8428 33460 8484 33470
rect 8428 33346 8484 33404
rect 8428 33294 8430 33346
rect 8482 33294 8484 33346
rect 8428 33282 8484 33294
rect 8316 33068 8484 33124
rect 7756 32844 8260 32900
rect 7756 32786 7812 32844
rect 7756 32734 7758 32786
rect 7810 32734 7812 32786
rect 7756 32722 7812 32734
rect 8204 32676 8260 32844
rect 8204 32674 8372 32676
rect 8204 32622 8206 32674
rect 8258 32622 8372 32674
rect 8204 32620 8372 32622
rect 8204 32610 8260 32620
rect 8092 32452 8148 32462
rect 8092 32450 8260 32452
rect 8092 32398 8094 32450
rect 8146 32398 8260 32450
rect 8092 32396 8260 32398
rect 8092 32386 8148 32396
rect 7756 31892 7812 31902
rect 7644 31836 7756 31892
rect 7756 31826 7812 31836
rect 7196 31220 7252 31230
rect 7084 31218 7252 31220
rect 7084 31166 7198 31218
rect 7250 31166 7252 31218
rect 7084 31164 7252 31166
rect 7196 31154 7252 31164
rect 6636 30706 6692 30716
rect 7420 31106 7476 31118
rect 7420 31054 7422 31106
rect 7474 31054 7476 31106
rect 7196 30436 7252 30446
rect 6524 29484 6804 29540
rect 6636 29092 6692 29102
rect 6636 28866 6692 29036
rect 6636 28814 6638 28866
rect 6690 28814 6692 28866
rect 6636 28802 6692 28814
rect 6748 28644 6804 29484
rect 6412 28590 6414 28642
rect 6466 28590 6468 28642
rect 6412 28578 6468 28590
rect 6636 28588 6804 28644
rect 7196 28642 7252 30380
rect 7420 30212 7476 31054
rect 8204 31108 8260 32396
rect 8316 32116 8372 32620
rect 8428 32674 8484 33068
rect 8428 32622 8430 32674
rect 8482 32622 8484 32674
rect 8428 32610 8484 32622
rect 8540 32340 8596 35308
rect 8652 34914 8708 35980
rect 8652 34862 8654 34914
rect 8706 34862 8708 34914
rect 8652 34850 8708 34862
rect 8764 35698 8820 35710
rect 8764 35646 8766 35698
rect 8818 35646 8820 35698
rect 8764 34802 8820 35646
rect 8988 35698 9044 36652
rect 9100 36594 9156 39228
rect 9212 38724 9268 39340
rect 10108 39396 10164 39406
rect 9548 38948 9604 38958
rect 9548 38854 9604 38892
rect 9212 38658 9268 38668
rect 9660 38836 9716 38846
rect 9660 38834 9828 38836
rect 9660 38782 9662 38834
rect 9714 38782 9828 38834
rect 9660 38780 9828 38782
rect 9660 38612 9716 38780
rect 9660 38546 9716 38556
rect 9660 38050 9716 38062
rect 9660 37998 9662 38050
rect 9714 37998 9716 38050
rect 9660 37940 9716 37998
rect 9660 37874 9716 37884
rect 9100 36542 9102 36594
rect 9154 36542 9156 36594
rect 9100 36530 9156 36542
rect 9548 37826 9604 37838
rect 9548 37774 9550 37826
rect 9602 37774 9604 37826
rect 9212 36258 9268 36270
rect 9212 36206 9214 36258
rect 9266 36206 9268 36258
rect 9212 35924 9268 36206
rect 9548 36036 9604 37774
rect 9660 37268 9716 37278
rect 9660 37154 9716 37212
rect 9660 37102 9662 37154
rect 9714 37102 9716 37154
rect 9660 37090 9716 37102
rect 9548 35980 9716 36036
rect 9212 35868 9604 35924
rect 9548 35810 9604 35868
rect 9548 35758 9550 35810
rect 9602 35758 9604 35810
rect 9548 35746 9604 35758
rect 8988 35646 8990 35698
rect 9042 35646 9044 35698
rect 8988 35634 9044 35646
rect 9660 35476 9716 35980
rect 8764 34750 8766 34802
rect 8818 34750 8820 34802
rect 8764 33572 8820 34750
rect 9324 35420 9716 35476
rect 8764 33506 8820 33516
rect 9212 33684 9268 33694
rect 9212 33570 9268 33628
rect 9212 33518 9214 33570
rect 9266 33518 9268 33570
rect 9212 33506 9268 33518
rect 8764 33348 8820 33358
rect 9100 33348 9156 33358
rect 8820 33346 9156 33348
rect 8820 33294 9102 33346
rect 9154 33294 9156 33346
rect 8820 33292 9156 33294
rect 8764 33254 8820 33292
rect 9100 33282 9156 33292
rect 9212 33348 9268 33358
rect 8652 33122 8708 33134
rect 8652 33070 8654 33122
rect 8706 33070 8708 33122
rect 8652 32788 8708 33070
rect 8652 32732 9044 32788
rect 8652 32564 8708 32574
rect 8652 32470 8708 32508
rect 8540 32284 8708 32340
rect 8316 32060 8596 32116
rect 8428 31892 8484 31902
rect 8428 31218 8484 31836
rect 8540 31890 8596 32060
rect 8540 31838 8542 31890
rect 8594 31838 8596 31890
rect 8540 31826 8596 31838
rect 8428 31166 8430 31218
rect 8482 31166 8484 31218
rect 8428 31154 8484 31166
rect 8204 31042 8260 31052
rect 7532 30994 7588 31006
rect 7532 30942 7534 30994
rect 7586 30942 7588 30994
rect 7532 30436 7588 30942
rect 7532 30370 7588 30380
rect 7644 30324 7700 30334
rect 7644 30212 7700 30268
rect 7420 30156 7700 30212
rect 7196 28590 7198 28642
rect 7250 28590 7252 28642
rect 6636 28196 6692 28588
rect 7196 28578 7252 28590
rect 7644 28642 7700 30156
rect 7644 28590 7646 28642
rect 7698 28590 7700 28642
rect 7644 28578 7700 28590
rect 8092 29316 8148 29326
rect 6636 28130 6692 28140
rect 7644 28420 7700 28430
rect 6300 28028 6580 28084
rect 6524 27972 6580 28028
rect 6636 27972 6692 27982
rect 6524 27970 6692 27972
rect 6524 27918 6638 27970
rect 6690 27918 6692 27970
rect 6524 27916 6692 27918
rect 6636 27906 6692 27916
rect 7644 27186 7700 28364
rect 7644 27134 7646 27186
rect 7698 27134 7700 27186
rect 7644 26908 7700 27134
rect 5964 26238 5966 26290
rect 6018 26238 6020 26290
rect 5628 26066 5908 26068
rect 5628 26014 5630 26066
rect 5682 26014 5908 26066
rect 5628 26012 5908 26014
rect 5628 26002 5684 26012
rect 5628 25732 5684 25742
rect 5516 25730 5684 25732
rect 5516 25678 5630 25730
rect 5682 25678 5684 25730
rect 5516 25676 5684 25678
rect 5628 25666 5684 25676
rect 4620 25618 4676 25630
rect 4620 25566 4622 25618
rect 4674 25566 4676 25618
rect 4620 25284 4676 25566
rect 5740 25508 5796 25518
rect 5740 25394 5796 25452
rect 5740 25342 5742 25394
rect 5794 25342 5796 25394
rect 5740 25330 5796 25342
rect 4620 25218 4676 25228
rect 4284 24658 4340 24668
rect 4172 24434 4228 24444
rect 5628 24610 5684 24622
rect 5628 24558 5630 24610
rect 5682 24558 5684 24610
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4620 24050 4676 24062
rect 4620 23998 4622 24050
rect 4674 23998 4676 24050
rect 1820 23940 1876 23950
rect 2044 23940 2100 23950
rect 1820 23938 2044 23940
rect 1820 23886 1822 23938
rect 1874 23886 2044 23938
rect 1820 23884 2044 23886
rect 1708 23154 1764 23166
rect 1708 23102 1710 23154
rect 1762 23102 1764 23154
rect 1708 22932 1764 23102
rect 1708 22866 1764 22876
rect 1820 22370 1876 23884
rect 2044 23874 2100 23884
rect 2492 23828 2548 23838
rect 2492 23826 2884 23828
rect 2492 23774 2494 23826
rect 2546 23774 2884 23826
rect 2492 23772 2884 23774
rect 2492 23762 2548 23772
rect 1820 22318 1822 22370
rect 1874 22318 1876 22370
rect 1708 22260 1764 22270
rect 1708 20802 1764 22204
rect 1708 20750 1710 20802
rect 1762 20750 1764 20802
rect 1708 20738 1764 20750
rect 1820 20018 1876 22318
rect 2044 23266 2100 23278
rect 2044 23214 2046 23266
rect 2098 23214 2100 23266
rect 2044 21700 2100 23214
rect 2492 23042 2548 23054
rect 2492 22990 2494 23042
rect 2546 22990 2548 23042
rect 2492 22932 2548 22990
rect 2828 23042 2884 23772
rect 4620 23604 4676 23998
rect 5068 23940 5124 23950
rect 5068 23846 5124 23884
rect 5516 23714 5572 23726
rect 5516 23662 5518 23714
rect 5570 23662 5572 23714
rect 4620 23538 4676 23548
rect 5292 23604 5348 23614
rect 3612 23380 3668 23390
rect 2940 23266 2996 23278
rect 2940 23214 2942 23266
rect 2994 23214 2996 23266
rect 2940 23156 2996 23214
rect 2940 23090 2996 23100
rect 2828 22990 2830 23042
rect 2882 22990 2884 23042
rect 2828 22978 2884 22990
rect 3164 23044 3220 23054
rect 3164 22950 3220 22988
rect 2492 22866 2548 22876
rect 2044 21634 2100 21644
rect 2380 22260 2436 22270
rect 1932 21476 1988 21486
rect 1932 21382 1988 21420
rect 2044 21028 2100 21038
rect 2044 20690 2100 20972
rect 2380 20916 2436 22204
rect 2492 22258 2548 22270
rect 2492 22206 2494 22258
rect 2546 22206 2548 22258
rect 2492 21924 2548 22206
rect 2492 21858 2548 21868
rect 2492 20916 2548 20926
rect 2380 20914 2548 20916
rect 2380 20862 2494 20914
rect 2546 20862 2548 20914
rect 2380 20860 2548 20862
rect 2492 20850 2548 20860
rect 3276 20916 3332 20926
rect 3276 20802 3332 20860
rect 3276 20750 3278 20802
rect 3330 20750 3332 20802
rect 3276 20738 3332 20750
rect 2044 20638 2046 20690
rect 2098 20638 2100 20690
rect 2044 20626 2100 20638
rect 2828 20690 2884 20702
rect 2828 20638 2830 20690
rect 2882 20638 2884 20690
rect 2828 20188 2884 20638
rect 2828 20132 3108 20188
rect 1820 19966 1822 20018
rect 1874 19966 1876 20018
rect 1820 18452 1876 19966
rect 2492 19908 2548 19918
rect 2492 19906 2772 19908
rect 2492 19854 2494 19906
rect 2546 19854 2772 19906
rect 2492 19852 2772 19854
rect 2492 19842 2548 19852
rect 2716 19458 2772 19852
rect 2716 19406 2718 19458
rect 2770 19406 2772 19458
rect 2716 19394 2772 19406
rect 3052 19458 3108 20132
rect 3052 19406 3054 19458
rect 3106 19406 3108 19458
rect 3052 19394 3108 19406
rect 2828 19348 2884 19358
rect 2828 19122 2884 19292
rect 3500 19348 3556 19358
rect 3612 19348 3668 23324
rect 5292 23154 5348 23548
rect 5292 23102 5294 23154
rect 5346 23102 5348 23154
rect 5292 23090 5348 23102
rect 5516 23154 5572 23662
rect 5516 23102 5518 23154
rect 5570 23102 5572 23154
rect 5516 23090 5572 23102
rect 4620 23044 4676 23054
rect 4620 22950 4676 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4620 22482 4676 22494
rect 4620 22430 4622 22482
rect 4674 22430 4676 22482
rect 4620 22260 4676 22430
rect 4620 22194 4676 22204
rect 5068 22148 5124 22158
rect 4284 21588 4340 21598
rect 4284 21494 4340 21532
rect 4956 21364 5012 21374
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4620 21028 4676 21038
rect 4620 20934 4676 20972
rect 4956 21026 5012 21308
rect 4956 20974 4958 21026
rect 5010 20974 5012 21026
rect 4956 20962 5012 20974
rect 3724 20802 3780 20814
rect 3724 20750 3726 20802
rect 3778 20750 3780 20802
rect 3724 20132 3780 20750
rect 4844 20802 4900 20814
rect 4844 20750 4846 20802
rect 4898 20750 4900 20802
rect 4508 20692 4564 20702
rect 3724 20066 3780 20076
rect 3836 20690 4564 20692
rect 3836 20638 4510 20690
rect 4562 20638 4564 20690
rect 3836 20636 4564 20638
rect 3500 19346 3612 19348
rect 3500 19294 3502 19346
rect 3554 19294 3612 19346
rect 3500 19292 3612 19294
rect 3500 19282 3556 19292
rect 3612 19282 3668 19292
rect 2828 19070 2830 19122
rect 2882 19070 2884 19122
rect 2828 19058 2884 19070
rect 3836 18788 3892 20636
rect 4508 20626 4564 20636
rect 4844 20132 4900 20750
rect 4844 20066 4900 20076
rect 4620 19908 4676 19918
rect 4620 19906 4900 19908
rect 4620 19854 4622 19906
rect 4674 19854 4900 19906
rect 4620 19852 4900 19854
rect 4620 19842 4676 19852
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4844 19236 4900 19852
rect 5068 19906 5124 22092
rect 5628 21588 5684 24558
rect 5852 23940 5908 26012
rect 5964 25730 6020 26238
rect 6076 26460 6244 26516
rect 7420 26852 7700 26908
rect 7756 27860 7812 27870
rect 7756 27076 7812 27804
rect 7420 26514 7476 26852
rect 7420 26462 7422 26514
rect 7474 26462 7476 26514
rect 6076 26292 6132 26460
rect 7420 26450 7476 26462
rect 6076 26226 6132 26236
rect 7084 26402 7140 26414
rect 7084 26350 7086 26402
rect 7138 26350 7140 26402
rect 7084 26292 7140 26350
rect 7084 26226 7140 26236
rect 5964 25678 5966 25730
rect 6018 25678 6020 25730
rect 5964 24834 6020 25678
rect 6188 26178 6244 26190
rect 6188 26126 6190 26178
rect 6242 26126 6244 26178
rect 6188 25508 6244 26126
rect 6636 25508 6692 25518
rect 6188 25452 6636 25508
rect 6636 25394 6692 25452
rect 7756 25506 7812 27020
rect 8092 26402 8148 29260
rect 8652 28642 8708 32284
rect 8988 31778 9044 32732
rect 9100 32340 9156 32350
rect 9100 32246 9156 32284
rect 8988 31726 8990 31778
rect 9042 31726 9044 31778
rect 8988 31714 9044 31726
rect 9212 31890 9268 33292
rect 9212 31838 9214 31890
rect 9266 31838 9268 31890
rect 9100 31556 9156 31566
rect 9100 31462 9156 31500
rect 9212 31332 9268 31838
rect 8988 31276 9268 31332
rect 8764 31108 8820 31118
rect 8764 31014 8820 31052
rect 8988 31106 9044 31276
rect 8988 31054 8990 31106
rect 9042 31054 9044 31106
rect 8988 31042 9044 31054
rect 8876 30882 8932 30894
rect 8876 30830 8878 30882
rect 8930 30830 8932 30882
rect 8876 29428 8932 30830
rect 8876 29362 8932 29372
rect 9324 29204 9380 35420
rect 9772 35364 9828 38780
rect 10108 38834 10164 39340
rect 10108 38782 10110 38834
rect 10162 38782 10164 38834
rect 10108 38770 10164 38782
rect 10220 37940 10276 39564
rect 10556 39526 10612 39564
rect 10668 39060 10724 39070
rect 10892 39060 10948 41918
rect 11228 40516 11284 40526
rect 11228 40422 11284 40460
rect 11004 40404 11060 40414
rect 11004 40310 11060 40348
rect 11228 40068 11284 40078
rect 11228 39506 11284 40012
rect 11228 39454 11230 39506
rect 11282 39454 11284 39506
rect 11228 39442 11284 39454
rect 10668 39058 10948 39060
rect 10668 39006 10670 39058
rect 10722 39006 10948 39058
rect 10668 39004 10948 39006
rect 11004 39396 11060 39406
rect 10668 38994 10724 39004
rect 11004 38946 11060 39340
rect 11004 38894 11006 38946
rect 11058 38894 11060 38946
rect 11004 38668 11060 38894
rect 11116 38836 11172 38846
rect 11116 38742 11172 38780
rect 11340 38724 11396 42476
rect 11452 42466 11508 42476
rect 11900 42308 11956 43484
rect 11452 42196 11508 42206
rect 11452 40514 11508 42140
rect 11900 42194 11956 42252
rect 11900 42142 11902 42194
rect 11954 42142 11956 42194
rect 11900 42130 11956 42142
rect 11564 41972 11620 41982
rect 11564 41970 11732 41972
rect 11564 41918 11566 41970
rect 11618 41918 11732 41970
rect 11564 41916 11732 41918
rect 11564 41906 11620 41916
rect 11452 40462 11454 40514
rect 11506 40462 11508 40514
rect 11452 40450 11508 40462
rect 11564 40402 11620 40414
rect 11564 40350 11566 40402
rect 11618 40350 11620 40402
rect 11564 39730 11620 40350
rect 11676 40068 11732 41916
rect 12012 40516 12068 45612
rect 12124 45330 12180 46732
rect 12796 46004 12852 49200
rect 12348 45948 12852 46004
rect 12348 45890 12404 45948
rect 12348 45838 12350 45890
rect 12402 45838 12404 45890
rect 12348 45826 12404 45838
rect 12572 45668 12628 45678
rect 12572 45574 12628 45612
rect 12124 45278 12126 45330
rect 12178 45278 12180 45330
rect 12124 45266 12180 45278
rect 12796 45330 12852 45948
rect 13468 46004 13524 49200
rect 13468 46002 13748 46004
rect 13468 45950 13470 46002
rect 13522 45950 13748 46002
rect 13468 45948 13748 45950
rect 13468 45938 13524 45948
rect 13692 45890 13748 45948
rect 13692 45838 13694 45890
rect 13746 45838 13748 45890
rect 13692 45826 13748 45838
rect 14812 45890 14868 49200
rect 14812 45838 14814 45890
rect 14866 45838 14868 45890
rect 12796 45278 12798 45330
rect 12850 45278 12852 45330
rect 12796 45266 12852 45278
rect 13468 45668 13524 45678
rect 12124 40516 12180 40526
rect 12012 40514 12180 40516
rect 12012 40462 12126 40514
rect 12178 40462 12180 40514
rect 12012 40460 12180 40462
rect 12124 40450 12180 40460
rect 11676 40002 11732 40012
rect 12236 40178 12292 40190
rect 12236 40126 12238 40178
rect 12290 40126 12292 40178
rect 11564 39678 11566 39730
rect 11618 39678 11620 39730
rect 11564 39666 11620 39678
rect 11676 39620 11732 39630
rect 11452 39396 11508 39406
rect 11452 39302 11508 39340
rect 11676 39060 11732 39564
rect 12236 39618 12292 40126
rect 12236 39566 12238 39618
rect 12290 39566 12292 39618
rect 12236 39554 12292 39566
rect 12684 39506 12740 39518
rect 12684 39454 12686 39506
rect 12738 39454 12740 39506
rect 12460 39394 12516 39406
rect 12460 39342 12462 39394
rect 12514 39342 12516 39394
rect 11676 39004 11844 39060
rect 11004 38612 11172 38668
rect 11340 38658 11396 38668
rect 11452 38836 11508 38846
rect 10556 38164 10612 38174
rect 10220 37874 10276 37884
rect 10444 38050 10500 38062
rect 10444 37998 10446 38050
rect 10498 37998 10500 38050
rect 10108 37268 10164 37278
rect 10164 37212 10276 37268
rect 10108 37202 10164 37212
rect 9660 35308 9828 35364
rect 9996 35698 10052 35710
rect 9996 35646 9998 35698
rect 10050 35646 10052 35698
rect 9660 32900 9716 35308
rect 9772 35140 9828 35150
rect 9772 34914 9828 35084
rect 9772 34862 9774 34914
rect 9826 34862 9828 34914
rect 9772 34850 9828 34862
rect 9996 34356 10052 35646
rect 10108 34356 10164 34366
rect 9996 34300 10108 34356
rect 10108 34290 10164 34300
rect 10108 34132 10164 34142
rect 10220 34132 10276 37212
rect 10444 36484 10500 37998
rect 10444 36418 10500 36428
rect 10556 35698 10612 38108
rect 10780 37268 10836 37278
rect 10780 36482 10836 37212
rect 10892 36708 10948 36718
rect 10892 36614 10948 36652
rect 10780 36430 10782 36482
rect 10834 36430 10836 36482
rect 10780 36418 10836 36430
rect 10556 35646 10558 35698
rect 10610 35646 10612 35698
rect 10556 35140 10612 35646
rect 10556 35074 10612 35084
rect 10668 35922 10724 35934
rect 10668 35870 10670 35922
rect 10722 35870 10724 35922
rect 10108 34130 10276 34132
rect 10108 34078 10110 34130
rect 10162 34078 10276 34130
rect 10108 34076 10276 34078
rect 10332 34916 10388 34926
rect 10108 34066 10164 34076
rect 10220 33908 10276 33918
rect 9996 33906 10276 33908
rect 9996 33854 10222 33906
rect 10274 33854 10276 33906
rect 9996 33852 10276 33854
rect 9996 33684 10052 33852
rect 10220 33842 10276 33852
rect 9884 33628 9996 33684
rect 9884 33570 9940 33628
rect 9996 33590 10052 33628
rect 9884 33518 9886 33570
rect 9938 33518 9940 33570
rect 9884 33506 9940 33518
rect 9884 33348 9940 33358
rect 9884 33122 9940 33292
rect 9884 33070 9886 33122
rect 9938 33070 9940 33122
rect 9884 33058 9940 33070
rect 9996 33346 10052 33358
rect 9996 33294 9998 33346
rect 10050 33294 10052 33346
rect 9996 33124 10052 33294
rect 9660 32844 9940 32900
rect 9884 32788 9940 32844
rect 9884 32694 9940 32732
rect 9996 32676 10052 33068
rect 9996 32610 10052 32620
rect 10220 33348 10276 33358
rect 10332 33348 10388 34860
rect 10556 34244 10612 34254
rect 10556 34150 10612 34188
rect 10668 34132 10724 35870
rect 10892 35924 10948 35934
rect 11116 35924 11172 38612
rect 11452 38050 11508 38780
rect 11676 38834 11732 38846
rect 11676 38782 11678 38834
rect 11730 38782 11732 38834
rect 11676 38724 11732 38782
rect 11676 38658 11732 38668
rect 11788 38668 11844 39004
rect 12348 38948 12404 38958
rect 12460 38948 12516 39342
rect 12348 38946 12516 38948
rect 12348 38894 12350 38946
rect 12402 38894 12516 38946
rect 12348 38892 12516 38894
rect 12348 38882 12404 38892
rect 12460 38724 12516 38734
rect 11788 38612 11956 38668
rect 11452 37998 11454 38050
rect 11506 37998 11508 38050
rect 11452 37986 11508 37998
rect 11788 37380 11844 37390
rect 11788 37286 11844 37324
rect 11564 36260 11620 36270
rect 10892 35922 11060 35924
rect 10892 35870 10894 35922
rect 10946 35870 11060 35922
rect 10892 35868 11060 35870
rect 10892 35858 10948 35868
rect 10780 35140 10836 35150
rect 10780 35046 10836 35084
rect 10892 35028 10948 35038
rect 10668 34066 10724 34076
rect 10780 34356 10836 34366
rect 10780 34130 10836 34300
rect 10892 34244 10948 34972
rect 11004 34916 11060 35868
rect 11116 35858 11172 35868
rect 11452 35924 11508 35934
rect 11340 35700 11396 35710
rect 11340 35606 11396 35644
rect 11452 35140 11508 35868
rect 11564 35922 11620 36204
rect 11564 35870 11566 35922
rect 11618 35870 11620 35922
rect 11564 35858 11620 35870
rect 11788 35924 11844 35934
rect 11900 35924 11956 38612
rect 12012 38164 12068 38174
rect 12012 38070 12068 38108
rect 12460 37826 12516 38668
rect 12684 38668 12740 39454
rect 12908 39508 12964 39518
rect 12908 39414 12964 39452
rect 12684 38612 13188 38668
rect 12460 37774 12462 37826
rect 12514 37774 12516 37826
rect 12460 37268 12516 37774
rect 13132 37492 13188 38612
rect 13132 37398 13188 37436
rect 13020 37380 13076 37390
rect 13020 37286 13076 37324
rect 12572 37268 12628 37278
rect 12460 37266 12628 37268
rect 12460 37214 12574 37266
rect 12626 37214 12628 37266
rect 12460 37212 12628 37214
rect 12572 36596 12628 37212
rect 12908 37266 12964 37278
rect 12908 37214 12910 37266
rect 12962 37214 12964 37266
rect 12908 36708 12964 37214
rect 13356 37268 13412 37278
rect 13356 37174 13412 37212
rect 12908 36642 12964 36652
rect 12796 36596 12852 36606
rect 12572 36594 12852 36596
rect 12572 36542 12798 36594
rect 12850 36542 12852 36594
rect 12572 36540 12852 36542
rect 12796 36530 12852 36540
rect 13468 36482 13524 45612
rect 14028 45668 14084 45678
rect 14028 45666 14532 45668
rect 14028 45614 14030 45666
rect 14082 45614 14532 45666
rect 14028 45612 14532 45614
rect 14028 45602 14084 45612
rect 14252 45108 14308 45118
rect 14252 44322 14308 45052
rect 14252 44270 14254 44322
rect 14306 44270 14308 44322
rect 14252 44258 14308 44270
rect 14476 42866 14532 45612
rect 14812 45330 14868 45838
rect 15484 45892 15540 49200
rect 16044 46786 16100 46798
rect 16044 46734 16046 46786
rect 16098 46734 16100 46786
rect 15596 45892 15652 45902
rect 16044 45892 16100 46734
rect 16156 46116 16212 49200
rect 16156 46050 16212 46060
rect 15484 45890 15652 45892
rect 15484 45838 15598 45890
rect 15650 45838 15652 45890
rect 15484 45836 15652 45838
rect 14812 45278 14814 45330
rect 14866 45278 14868 45330
rect 14812 45266 14868 45278
rect 15036 45666 15092 45678
rect 15372 45668 15428 45678
rect 15036 45614 15038 45666
rect 15090 45614 15092 45666
rect 14924 45108 14980 45118
rect 14924 44436 14980 45052
rect 14476 42814 14478 42866
rect 14530 42814 14532 42866
rect 14476 42802 14532 42814
rect 14812 44380 14980 44436
rect 13580 42754 13636 42766
rect 13580 42702 13582 42754
rect 13634 42702 13636 42754
rect 13580 41972 13636 42702
rect 13804 42754 13860 42766
rect 13804 42702 13806 42754
rect 13858 42702 13860 42754
rect 13804 42196 13860 42702
rect 14140 42756 14196 42766
rect 14364 42756 14420 42766
rect 14140 42754 14420 42756
rect 14140 42702 14142 42754
rect 14194 42702 14366 42754
rect 14418 42702 14420 42754
rect 14140 42700 14420 42702
rect 14140 42690 14196 42700
rect 14364 42690 14420 42700
rect 13916 42532 13972 42542
rect 13916 42530 14196 42532
rect 13916 42478 13918 42530
rect 13970 42478 14196 42530
rect 13916 42476 14196 42478
rect 13916 42466 13972 42476
rect 13804 42130 13860 42140
rect 14140 42082 14196 42476
rect 14140 42030 14142 42082
rect 14194 42030 14196 42082
rect 14140 42018 14196 42030
rect 14700 42196 14756 42206
rect 13580 41906 13636 41916
rect 13580 40068 13636 40078
rect 13580 39732 13636 40012
rect 13580 39506 13636 39676
rect 13580 39454 13582 39506
rect 13634 39454 13636 39506
rect 13580 39442 13636 39454
rect 13916 39508 13972 39518
rect 13916 39414 13972 39452
rect 13804 39396 13860 39406
rect 13804 39302 13860 39340
rect 14028 39394 14084 39406
rect 14028 39342 14030 39394
rect 14082 39342 14084 39394
rect 14028 38668 14084 39342
rect 14476 38722 14532 38734
rect 14476 38670 14478 38722
rect 14530 38670 14532 38722
rect 14476 38668 14532 38670
rect 14028 38612 14532 38668
rect 14028 37828 14084 37838
rect 14028 37826 14196 37828
rect 14028 37774 14030 37826
rect 14082 37774 14196 37826
rect 14028 37772 14196 37774
rect 14028 37762 14084 37772
rect 13580 37266 13636 37278
rect 13580 37214 13582 37266
rect 13634 37214 13636 37266
rect 13580 36706 13636 37214
rect 14140 37268 14196 37772
rect 14252 37380 14308 37390
rect 14252 37286 14308 37324
rect 13580 36654 13582 36706
rect 13634 36654 13636 36706
rect 13580 36642 13636 36654
rect 14028 37156 14084 37166
rect 13468 36430 13470 36482
rect 13522 36430 13524 36482
rect 13468 36418 13524 36430
rect 13692 36596 13748 36606
rect 13580 36372 13636 36382
rect 13692 36372 13748 36540
rect 13580 36370 13860 36372
rect 13580 36318 13582 36370
rect 13634 36318 13860 36370
rect 13580 36316 13860 36318
rect 13580 36306 13636 36316
rect 11900 35868 12068 35924
rect 11788 35830 11844 35868
rect 11900 35700 11956 35710
rect 11788 35698 11956 35700
rect 11788 35646 11902 35698
rect 11954 35646 11956 35698
rect 11788 35644 11956 35646
rect 11676 35586 11732 35598
rect 11676 35534 11678 35586
rect 11730 35534 11732 35586
rect 11564 35140 11620 35150
rect 11452 35138 11620 35140
rect 11452 35086 11566 35138
rect 11618 35086 11620 35138
rect 11452 35084 11620 35086
rect 11564 35074 11620 35084
rect 11116 34916 11172 34926
rect 11004 34914 11172 34916
rect 11004 34862 11118 34914
rect 11170 34862 11172 34914
rect 11004 34860 11172 34862
rect 11004 34580 11060 34860
rect 11116 34850 11172 34860
rect 11676 34692 11732 35534
rect 11788 34916 11844 35644
rect 11900 35634 11956 35644
rect 11788 34822 11844 34860
rect 12012 34916 12068 35868
rect 13804 35922 13860 36316
rect 13804 35870 13806 35922
rect 13858 35870 13860 35922
rect 13804 35858 13860 35870
rect 13244 35700 13300 35710
rect 13020 34916 13076 34926
rect 12012 34914 12852 34916
rect 12012 34862 12014 34914
rect 12066 34862 12852 34914
rect 12012 34860 12852 34862
rect 11676 34636 11956 34692
rect 11004 34514 11060 34524
rect 11004 34244 11060 34254
rect 10892 34242 11060 34244
rect 10892 34190 11006 34242
rect 11058 34190 11060 34242
rect 10892 34188 11060 34190
rect 11004 34178 11060 34188
rect 10780 34078 10782 34130
rect 10834 34078 10836 34130
rect 10220 33346 10388 33348
rect 10220 33294 10222 33346
rect 10274 33294 10388 33346
rect 10220 33292 10388 33294
rect 10220 32450 10276 33292
rect 10444 33236 10500 33246
rect 10780 33236 10836 34078
rect 11116 34020 11172 34030
rect 11116 34018 11508 34020
rect 11116 33966 11118 34018
rect 11170 33966 11508 34018
rect 11116 33964 11508 33966
rect 11116 33954 11172 33964
rect 11452 33570 11508 33964
rect 11452 33518 11454 33570
rect 11506 33518 11508 33570
rect 11452 33506 11508 33518
rect 11900 33572 11956 34636
rect 12012 34130 12068 34860
rect 12796 34802 12852 34860
rect 12796 34750 12798 34802
rect 12850 34750 12852 34802
rect 12796 34738 12852 34750
rect 12908 34802 12964 34814
rect 12908 34750 12910 34802
rect 12962 34750 12964 34802
rect 12012 34078 12014 34130
rect 12066 34078 12068 34130
rect 12012 34066 12068 34078
rect 12124 34690 12180 34702
rect 12124 34638 12126 34690
rect 12178 34638 12180 34690
rect 12124 33684 12180 34638
rect 12236 34692 12292 34702
rect 12236 34598 12292 34636
rect 12572 34690 12628 34702
rect 12572 34638 12574 34690
rect 12626 34638 12628 34690
rect 12572 34244 12628 34638
rect 12908 34692 12964 34750
rect 12908 34626 12964 34636
rect 12124 33628 12404 33684
rect 11900 33516 12180 33572
rect 11228 33460 11284 33470
rect 11228 33366 11284 33404
rect 12124 33346 12180 33516
rect 12124 33294 12126 33346
rect 12178 33294 12180 33346
rect 12124 33282 12180 33294
rect 12348 33460 12404 33628
rect 10500 33180 10836 33236
rect 12348 33234 12404 33404
rect 12348 33182 12350 33234
rect 12402 33182 12404 33234
rect 10444 32674 10500 33180
rect 12348 33170 12404 33182
rect 12460 33234 12516 33246
rect 12460 33182 12462 33234
rect 12514 33182 12516 33234
rect 10892 33124 10948 33134
rect 10444 32622 10446 32674
rect 10498 32622 10500 32674
rect 10444 32610 10500 32622
rect 10556 33068 10892 33124
rect 10220 32398 10222 32450
rect 10274 32398 10276 32450
rect 10220 32386 10276 32398
rect 9436 31778 9492 31790
rect 9436 31726 9438 31778
rect 9490 31726 9492 31778
rect 9436 29986 9492 31726
rect 10556 31780 10612 33068
rect 10892 33030 10948 33068
rect 11788 33122 11844 33134
rect 11788 33070 11790 33122
rect 11842 33070 11844 33122
rect 11004 32788 11060 32798
rect 11004 32694 11060 32732
rect 10780 32676 10836 32686
rect 10780 32582 10836 32620
rect 11788 32674 11844 33070
rect 11788 32622 11790 32674
rect 11842 32622 11844 32674
rect 11788 32610 11844 32622
rect 11116 32452 11172 32462
rect 11116 32358 11172 32396
rect 11228 32340 11284 32350
rect 11116 31892 11172 31902
rect 11116 31798 11172 31836
rect 10556 31686 10612 31724
rect 10108 30882 10164 30894
rect 10108 30830 10110 30882
rect 10162 30830 10164 30882
rect 9884 30212 9940 30222
rect 10108 30212 10164 30830
rect 9884 30210 10164 30212
rect 9884 30158 9886 30210
rect 9938 30158 10164 30210
rect 9884 30156 10164 30158
rect 9884 30146 9940 30156
rect 9436 29934 9438 29986
rect 9490 29934 9492 29986
rect 9436 29316 9492 29934
rect 9436 29250 9492 29260
rect 8652 28590 8654 28642
rect 8706 28590 8708 28642
rect 8652 28578 8708 28590
rect 8876 29148 9380 29204
rect 8876 28642 8932 29148
rect 8876 28590 8878 28642
rect 8930 28590 8932 28642
rect 8876 28578 8932 28590
rect 9660 28980 9716 28990
rect 9660 28644 9716 28924
rect 9884 28866 9940 28878
rect 9884 28814 9886 28866
rect 9938 28814 9940 28866
rect 9772 28756 9828 28766
rect 9772 28662 9828 28700
rect 9660 28550 9716 28588
rect 9884 28308 9940 28814
rect 9884 28242 9940 28252
rect 9996 28644 10052 28654
rect 9996 28082 10052 28588
rect 9996 28030 9998 28082
rect 10050 28030 10052 28082
rect 9996 28018 10052 28030
rect 9772 27972 9828 27982
rect 9660 27916 9772 27972
rect 9548 27858 9604 27870
rect 9548 27806 9550 27858
rect 9602 27806 9604 27858
rect 8764 27748 8820 27758
rect 8764 27654 8820 27692
rect 9548 27748 9604 27806
rect 9100 27188 9156 27198
rect 9100 27094 9156 27132
rect 9436 27188 9492 27198
rect 9548 27188 9604 27692
rect 9660 27298 9716 27916
rect 9772 27878 9828 27916
rect 9884 27860 9940 27870
rect 9884 27766 9940 27804
rect 9660 27246 9662 27298
rect 9714 27246 9716 27298
rect 9660 27234 9716 27246
rect 9436 27186 9604 27188
rect 9436 27134 9438 27186
rect 9490 27134 9604 27186
rect 9436 27132 9604 27134
rect 9436 27122 9492 27132
rect 10108 27076 10164 30156
rect 10556 30100 10612 30110
rect 10332 30098 10612 30100
rect 10332 30046 10558 30098
rect 10610 30046 10612 30098
rect 10332 30044 10612 30046
rect 10332 29650 10388 30044
rect 10556 30034 10612 30044
rect 10332 29598 10334 29650
rect 10386 29598 10388 29650
rect 10332 29586 10388 29598
rect 10220 29428 10276 29438
rect 10220 29334 10276 29372
rect 10444 29428 10500 29438
rect 10444 29334 10500 29372
rect 11228 29426 11284 32284
rect 11900 31780 11956 31790
rect 11900 30996 11956 31724
rect 12460 31444 12516 33182
rect 12572 33234 12628 34188
rect 13020 34130 13076 34860
rect 13020 34078 13022 34130
rect 13074 34078 13076 34130
rect 13020 34066 13076 34078
rect 12572 33182 12574 33234
rect 12626 33182 12628 33234
rect 12572 33170 12628 33182
rect 12908 33458 12964 33470
rect 12908 33406 12910 33458
rect 12962 33406 12964 33458
rect 12908 33236 12964 33406
rect 12908 33170 12964 33180
rect 12908 33012 12964 33022
rect 12460 31378 12516 31388
rect 12684 31668 12740 31678
rect 12684 31108 12740 31612
rect 12908 31218 12964 32956
rect 13244 32562 13300 35644
rect 14028 35698 14084 37100
rect 14140 36708 14196 37212
rect 14476 37044 14532 38612
rect 14588 37266 14644 37278
rect 14588 37214 14590 37266
rect 14642 37214 14644 37266
rect 14588 37156 14644 37214
rect 14588 37090 14644 37100
rect 14476 36978 14532 36988
rect 14140 36642 14196 36652
rect 14028 35646 14030 35698
rect 14082 35646 14084 35698
rect 14028 35634 14084 35646
rect 14476 35924 14532 35934
rect 14700 35924 14756 42140
rect 14812 41970 14868 44380
rect 14924 44210 14980 44222
rect 14924 44158 14926 44210
rect 14978 44158 14980 44210
rect 14924 43652 14980 44158
rect 14924 43586 14980 43596
rect 14812 41918 14814 41970
rect 14866 41918 14868 41970
rect 14812 40404 14868 41918
rect 14924 42308 14980 42318
rect 14924 41298 14980 42252
rect 14924 41246 14926 41298
rect 14978 41246 14980 41298
rect 14924 41234 14980 41246
rect 14812 39618 14868 40348
rect 14812 39566 14814 39618
rect 14866 39566 14868 39618
rect 14812 36484 14868 39566
rect 14924 37380 14980 37390
rect 15036 37380 15092 45614
rect 15148 45666 15428 45668
rect 15148 45614 15374 45666
rect 15426 45614 15428 45666
rect 15148 45612 15428 45614
rect 15148 40514 15204 45612
rect 15372 45602 15428 45612
rect 15372 45332 15428 45342
rect 15484 45332 15540 45836
rect 15596 45826 15652 45836
rect 15820 45890 16100 45892
rect 15820 45838 16046 45890
rect 16098 45838 16100 45890
rect 15820 45836 16100 45838
rect 15372 45330 15540 45332
rect 15372 45278 15374 45330
rect 15426 45278 15540 45330
rect 15372 45276 15540 45278
rect 15820 45330 15876 45836
rect 16044 45826 16100 45836
rect 16380 45666 16436 45678
rect 16380 45614 16382 45666
rect 16434 45614 16436 45666
rect 15820 45278 15822 45330
rect 15874 45278 15876 45330
rect 15372 45266 15428 45276
rect 15820 45266 15876 45278
rect 16268 45332 16324 45342
rect 16268 45238 16324 45276
rect 15260 42308 15316 42318
rect 15260 42194 15316 42252
rect 15260 42142 15262 42194
rect 15314 42142 15316 42194
rect 15260 42130 15316 42142
rect 15484 42084 15540 42094
rect 15372 41972 15428 41982
rect 15372 41878 15428 41916
rect 15484 40964 15540 42028
rect 15932 41970 15988 41982
rect 15932 41918 15934 41970
rect 15986 41918 15988 41970
rect 15932 41860 15988 41918
rect 16268 41860 16324 41870
rect 15932 41804 16268 41860
rect 16268 41766 16324 41804
rect 15148 40462 15150 40514
rect 15202 40462 15204 40514
rect 15148 40450 15204 40462
rect 15372 40908 15540 40964
rect 16044 41186 16100 41198
rect 16044 41134 16046 41186
rect 16098 41134 16100 41186
rect 15260 40178 15316 40190
rect 15260 40126 15262 40178
rect 15314 40126 15316 40178
rect 15260 38834 15316 40126
rect 15260 38782 15262 38834
rect 15314 38782 15316 38834
rect 15260 38770 15316 38782
rect 14924 37378 15092 37380
rect 14924 37326 14926 37378
rect 14978 37326 15092 37378
rect 14924 37324 15092 37326
rect 14924 37314 14980 37324
rect 15260 37268 15316 37278
rect 15036 37266 15316 37268
rect 15036 37214 15262 37266
rect 15314 37214 15316 37266
rect 15036 37212 15316 37214
rect 14812 36390 14868 36428
rect 14924 37156 14980 37166
rect 14476 35922 14756 35924
rect 14476 35870 14478 35922
rect 14530 35870 14756 35922
rect 14476 35868 14756 35870
rect 14812 35924 14868 35934
rect 14924 35924 14980 37100
rect 15036 37154 15092 37212
rect 15260 37202 15316 37212
rect 15036 37102 15038 37154
rect 15090 37102 15092 37154
rect 15036 37090 15092 37102
rect 14812 35922 14980 35924
rect 14812 35870 14814 35922
rect 14866 35870 14980 35922
rect 14812 35868 14980 35870
rect 15372 36484 15428 40908
rect 16044 40404 16100 41134
rect 16380 40628 16436 45614
rect 16828 45332 16884 49200
rect 17500 46786 17556 49200
rect 17500 46734 17502 46786
rect 17554 46734 17556 46786
rect 17500 46722 17556 46734
rect 18172 46450 18228 49200
rect 18172 46398 18174 46450
rect 18226 46398 18228 46450
rect 18172 46386 18228 46398
rect 17948 46116 18004 46126
rect 17948 46022 18004 46060
rect 17388 45892 17444 45902
rect 18844 45892 18900 49200
rect 19068 46562 19124 46574
rect 19068 46510 19070 46562
rect 19122 46510 19124 46562
rect 17388 45890 17892 45892
rect 17388 45838 17390 45890
rect 17442 45838 17892 45890
rect 17388 45836 17892 45838
rect 18844 45836 19012 45892
rect 17388 45826 17444 45836
rect 16492 45218 16548 45230
rect 16492 45166 16494 45218
rect 16546 45166 16548 45218
rect 16492 43538 16548 45166
rect 16828 45218 16884 45276
rect 16828 45166 16830 45218
rect 16882 45166 16884 45218
rect 16828 45154 16884 45166
rect 17388 45108 17444 45118
rect 17388 45014 17444 45052
rect 17052 44436 17108 44446
rect 17052 44342 17108 44380
rect 17500 43652 17556 43662
rect 17500 43558 17556 43596
rect 16492 43486 16494 43538
rect 16546 43486 16548 43538
rect 16492 43474 16548 43486
rect 16716 43540 16772 43550
rect 16716 43446 16772 43484
rect 17388 43538 17444 43550
rect 17388 43486 17390 43538
rect 17442 43486 17444 43538
rect 16828 43428 16884 43438
rect 16828 43334 16884 43372
rect 17388 42868 17444 43486
rect 17612 43540 17668 43550
rect 17612 43446 17668 43484
rect 17388 42802 17444 42812
rect 17724 43428 17780 43438
rect 17388 42082 17444 42094
rect 17388 42030 17390 42082
rect 17442 42030 17444 42082
rect 17388 41748 17444 42030
rect 17612 41970 17668 41982
rect 17612 41918 17614 41970
rect 17666 41918 17668 41970
rect 17388 41682 17444 41692
rect 17500 41858 17556 41870
rect 17500 41806 17502 41858
rect 17554 41806 17556 41858
rect 17500 41524 17556 41806
rect 16828 41468 17556 41524
rect 16828 41298 16884 41468
rect 16828 41246 16830 41298
rect 16882 41246 16884 41298
rect 16828 41234 16884 41246
rect 16380 40562 16436 40572
rect 17388 40628 17444 40638
rect 16044 40338 16100 40348
rect 17388 40402 17444 40572
rect 17388 40350 17390 40402
rect 17442 40350 17444 40402
rect 17388 40338 17444 40350
rect 17612 40290 17668 41918
rect 17612 40238 17614 40290
rect 17666 40238 17668 40290
rect 17612 40226 17668 40238
rect 17724 40292 17780 43372
rect 17724 40198 17780 40236
rect 17836 40068 17892 45836
rect 18844 45668 18900 45678
rect 18172 44996 18228 45006
rect 18172 44994 18452 44996
rect 18172 44942 18174 44994
rect 18226 44942 18452 44994
rect 18172 44940 18452 44942
rect 18172 44930 18228 44940
rect 18396 44434 18452 44940
rect 18396 44382 18398 44434
rect 18450 44382 18452 44434
rect 18396 44370 18452 44382
rect 18508 44324 18564 44334
rect 18508 44322 18676 44324
rect 18508 44270 18510 44322
rect 18562 44270 18676 44322
rect 18508 44268 18676 44270
rect 18508 44258 18564 44268
rect 18620 44212 18676 44268
rect 18732 44212 18788 44222
rect 18620 44156 18732 44212
rect 18732 44146 18788 44156
rect 17612 40012 17892 40068
rect 18060 44098 18116 44110
rect 18060 44046 18062 44098
rect 18114 44046 18116 44098
rect 18060 43538 18116 44046
rect 18284 44100 18340 44110
rect 18508 44100 18564 44110
rect 18284 44098 18452 44100
rect 18284 44046 18286 44098
rect 18338 44046 18452 44098
rect 18284 44044 18452 44046
rect 18284 44034 18340 44044
rect 18396 43762 18452 44044
rect 18396 43710 18398 43762
rect 18450 43710 18452 43762
rect 18396 43698 18452 43710
rect 18508 43650 18564 44044
rect 18508 43598 18510 43650
rect 18562 43598 18564 43650
rect 18508 43586 18564 43598
rect 18060 43486 18062 43538
rect 18114 43486 18116 43538
rect 18060 41970 18116 43486
rect 18284 43428 18340 43438
rect 18284 43334 18340 43372
rect 18060 41918 18062 41970
rect 18114 41918 18116 41970
rect 17612 39732 17668 40012
rect 17500 39730 17668 39732
rect 17500 39678 17614 39730
rect 17666 39678 17668 39730
rect 17500 39676 17668 39678
rect 15484 39506 15540 39518
rect 15484 39454 15486 39506
rect 15538 39454 15540 39506
rect 15484 39058 15540 39454
rect 15484 39006 15486 39058
rect 15538 39006 15540 39058
rect 15484 38994 15540 39006
rect 15932 39396 15988 39406
rect 15932 38946 15988 39340
rect 15932 38894 15934 38946
rect 15986 38894 15988 38946
rect 15932 38882 15988 38894
rect 15708 38834 15764 38846
rect 15708 38782 15710 38834
rect 15762 38782 15764 38834
rect 15596 37490 15652 37502
rect 15596 37438 15598 37490
rect 15650 37438 15652 37490
rect 15596 36594 15652 37438
rect 15708 37380 15764 38782
rect 17500 38834 17556 39676
rect 17612 39666 17668 39676
rect 18060 39620 18116 41918
rect 18844 40628 18900 45612
rect 18956 45332 19012 45836
rect 18956 45266 19012 45276
rect 19068 44434 19124 46510
rect 19516 46562 19572 49200
rect 19516 46510 19518 46562
rect 19570 46510 19572 46562
rect 19516 46498 19572 46510
rect 20076 46562 20132 46574
rect 20076 46510 20078 46562
rect 20130 46510 20132 46562
rect 20076 45890 20132 46510
rect 21644 46450 21700 46462
rect 21644 46398 21646 46450
rect 21698 46398 21700 46450
rect 20076 45838 20078 45890
rect 20130 45838 20132 45890
rect 20076 45826 20132 45838
rect 20972 45890 21028 45902
rect 20972 45838 20974 45890
rect 21026 45838 21028 45890
rect 19852 45668 19908 45706
rect 19852 45602 19908 45612
rect 20748 45666 20804 45678
rect 20748 45614 20750 45666
rect 20802 45614 20804 45666
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20524 45332 20580 45342
rect 20580 45276 20692 45332
rect 20524 45266 20580 45276
rect 19852 45220 19908 45230
rect 19068 44382 19070 44434
rect 19122 44382 19124 44434
rect 19068 44370 19124 44382
rect 19516 44436 19572 44446
rect 19516 44322 19572 44380
rect 19740 44324 19796 44334
rect 19516 44270 19518 44322
rect 19570 44270 19572 44322
rect 19292 44210 19348 44222
rect 19292 44158 19294 44210
rect 19346 44158 19348 44210
rect 19292 43540 19348 44158
rect 19404 44212 19460 44222
rect 19404 44118 19460 44156
rect 19516 43876 19572 44270
rect 19516 43810 19572 43820
rect 19628 44322 19796 44324
rect 19628 44270 19742 44322
rect 19794 44270 19796 44322
rect 19628 44268 19796 44270
rect 19292 42756 19348 43484
rect 19628 43428 19684 44268
rect 19740 44258 19796 44268
rect 19852 44100 19908 45164
rect 20188 45108 20244 45118
rect 20076 44324 20132 44334
rect 20076 44230 20132 44268
rect 19852 44034 19908 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19740 43764 19796 43774
rect 19740 43650 19796 43708
rect 19740 43598 19742 43650
rect 19794 43598 19796 43650
rect 19740 43586 19796 43598
rect 19628 43092 19684 43372
rect 19852 43316 19908 43326
rect 19852 43222 19908 43260
rect 19628 43036 19908 43092
rect 19852 42978 19908 43036
rect 19852 42926 19854 42978
rect 19906 42926 19908 42978
rect 19852 42914 19908 42926
rect 19516 42868 19572 42878
rect 19516 42774 19572 42812
rect 19404 42756 19460 42766
rect 19292 42754 19460 42756
rect 19292 42702 19406 42754
rect 19458 42702 19460 42754
rect 19292 42700 19460 42702
rect 19404 42690 19460 42700
rect 20076 42756 20132 42766
rect 20076 42662 20132 42700
rect 19628 42642 19684 42654
rect 19628 42590 19630 42642
rect 19682 42590 19684 42642
rect 19516 42196 19572 42206
rect 18956 41300 19012 41310
rect 18956 41206 19012 41244
rect 18956 40628 19012 40638
rect 18844 40626 19012 40628
rect 18844 40574 18958 40626
rect 19010 40574 19012 40626
rect 18844 40572 19012 40574
rect 18956 40562 19012 40572
rect 19516 40402 19572 42140
rect 19628 41972 19684 42590
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 20076 42196 20132 42206
rect 19964 42194 20132 42196
rect 19964 42142 20078 42194
rect 20130 42142 20132 42194
rect 19964 42140 20132 42142
rect 19964 42084 20020 42140
rect 20076 42130 20132 42140
rect 20188 42196 20244 45052
rect 20300 44996 20356 45006
rect 20524 44996 20580 45006
rect 20300 44994 20580 44996
rect 20300 44942 20302 44994
rect 20354 44942 20526 44994
rect 20578 44942 20580 44994
rect 20300 44940 20580 44942
rect 20300 44930 20356 44940
rect 20524 44930 20580 44940
rect 20524 44324 20580 44334
rect 20524 44230 20580 44268
rect 20412 44212 20468 44222
rect 20188 42130 20244 42140
rect 20300 44210 20468 44212
rect 20300 44158 20414 44210
rect 20466 44158 20468 44210
rect 20300 44156 20468 44158
rect 19964 42018 20020 42028
rect 20300 42084 20356 44156
rect 20412 44146 20468 44156
rect 20524 43652 20580 43662
rect 20636 43652 20692 45276
rect 20748 45220 20804 45614
rect 20972 45332 21028 45838
rect 21644 45892 21700 46398
rect 22316 46004 22372 46014
rect 22876 46004 22932 49200
rect 23548 46116 23604 49200
rect 23548 46050 23604 46060
rect 23772 46450 23828 46462
rect 23772 46398 23774 46450
rect 23826 46398 23828 46450
rect 22316 46002 22932 46004
rect 22316 45950 22318 46002
rect 22370 45950 22932 46002
rect 22316 45948 22932 45950
rect 22316 45938 22372 45948
rect 22876 45892 22932 45948
rect 22988 45892 23044 45902
rect 21644 45890 21812 45892
rect 21644 45838 21646 45890
rect 21698 45838 21812 45890
rect 21644 45836 21812 45838
rect 22876 45890 23044 45892
rect 22876 45838 22990 45890
rect 23042 45838 23044 45890
rect 22876 45836 23044 45838
rect 21644 45826 21700 45836
rect 21420 45668 21476 45678
rect 21420 45666 21588 45668
rect 21420 45614 21422 45666
rect 21474 45614 21588 45666
rect 21420 45612 21588 45614
rect 21420 45602 21476 45612
rect 20972 45266 21028 45276
rect 20748 45154 20804 45164
rect 20860 45108 20916 45118
rect 21084 45108 21140 45118
rect 20916 45106 21140 45108
rect 20916 45054 21086 45106
rect 21138 45054 21140 45106
rect 20916 45052 21140 45054
rect 20860 45042 20916 45052
rect 21084 45042 21140 45052
rect 20748 44994 20804 45006
rect 20748 44942 20750 44994
rect 20802 44942 20804 44994
rect 20748 44548 20804 44942
rect 20748 44492 21476 44548
rect 21420 44434 21476 44492
rect 21420 44382 21422 44434
rect 21474 44382 21476 44434
rect 20748 44324 20804 44334
rect 21308 44324 21364 44334
rect 20748 44322 21364 44324
rect 20748 44270 20750 44322
rect 20802 44270 21310 44322
rect 21362 44270 21364 44322
rect 20748 44268 21364 44270
rect 20748 44258 20804 44268
rect 21308 44258 21364 44268
rect 20524 43650 20692 43652
rect 20524 43598 20526 43650
rect 20578 43598 20692 43650
rect 20524 43596 20692 43598
rect 21420 43652 21476 44382
rect 20524 43586 20580 43596
rect 21420 43586 21476 43596
rect 19628 41300 19684 41916
rect 20300 41970 20356 42028
rect 20300 41918 20302 41970
rect 20354 41918 20356 41970
rect 20300 41906 20356 41918
rect 20412 42756 20468 42766
rect 20188 41858 20244 41870
rect 20188 41806 20190 41858
rect 20242 41806 20244 41858
rect 20188 41748 20244 41806
rect 20412 41748 20468 42700
rect 21532 42196 21588 45612
rect 21756 45332 21812 45836
rect 22988 45826 23044 45836
rect 23772 45890 23828 46398
rect 23772 45838 23774 45890
rect 23826 45838 23828 45890
rect 22764 45780 22820 45790
rect 22764 45686 22820 45724
rect 23772 45780 23828 45838
rect 23772 45714 23828 45724
rect 23324 45668 23380 45678
rect 22988 45666 23380 45668
rect 22988 45614 23326 45666
rect 23378 45614 23380 45666
rect 22988 45612 23380 45614
rect 21756 45276 21924 45332
rect 21756 44994 21812 45006
rect 21756 44942 21758 44994
rect 21810 44942 21812 44994
rect 21196 42140 21588 42196
rect 21644 43540 21700 43550
rect 21644 42196 21700 43484
rect 21756 43316 21812 44942
rect 21868 44434 21924 45276
rect 21868 44382 21870 44434
rect 21922 44382 21924 44434
rect 21868 44370 21924 44382
rect 22988 43988 23044 45612
rect 23324 45602 23380 45612
rect 23996 45668 24052 45678
rect 24220 45668 24276 49200
rect 24892 46450 24948 49200
rect 24892 46398 24894 46450
rect 24946 46398 24948 46450
rect 24892 46386 24948 46398
rect 26908 46450 26964 49200
rect 27580 46786 27636 49200
rect 27580 46734 27582 46786
rect 27634 46734 27636 46786
rect 27580 46722 27636 46734
rect 26908 46398 26910 46450
rect 26962 46398 26964 46450
rect 26908 46386 26964 46398
rect 27468 46450 27524 46462
rect 27468 46398 27470 46450
rect 27522 46398 27524 46450
rect 25564 46116 25620 46126
rect 25564 46022 25620 46060
rect 25004 45890 25060 45902
rect 27468 45892 27524 46398
rect 25004 45838 25006 45890
rect 25058 45838 25060 45890
rect 23996 45666 24164 45668
rect 23996 45614 23998 45666
rect 24050 45614 24164 45666
rect 23996 45612 24164 45614
rect 24220 45612 24612 45668
rect 23996 45602 24052 45612
rect 24108 45444 24164 45612
rect 24108 45388 24500 45444
rect 24332 45220 24388 45230
rect 24220 45218 24388 45220
rect 24220 45166 24334 45218
rect 24386 45166 24388 45218
rect 24220 45164 24388 45166
rect 23884 44994 23940 45006
rect 23884 44942 23886 44994
rect 23938 44942 23940 44994
rect 23436 44212 23492 44222
rect 23884 44212 23940 44942
rect 24108 44212 24164 44222
rect 23884 44156 24108 44212
rect 23436 44118 23492 44156
rect 23324 44098 23380 44110
rect 23324 44046 23326 44098
rect 23378 44046 23380 44098
rect 22988 43932 23268 43988
rect 22428 43764 22484 43774
rect 22764 43764 22820 43774
rect 22428 43762 22820 43764
rect 22428 43710 22430 43762
rect 22482 43710 22766 43762
rect 22818 43710 22820 43762
rect 22428 43708 22820 43710
rect 22428 43698 22484 43708
rect 22764 43698 22820 43708
rect 21868 43652 21924 43662
rect 21868 43558 21924 43596
rect 22428 43538 22484 43550
rect 22428 43486 22430 43538
rect 22482 43486 22484 43538
rect 22092 43428 22148 43438
rect 21756 43250 21812 43260
rect 21868 43372 22092 43428
rect 20636 41972 20692 41982
rect 20636 41878 20692 41916
rect 20748 41972 20804 41982
rect 21084 41972 21140 41982
rect 20748 41970 21140 41972
rect 20748 41918 20750 41970
rect 20802 41918 21086 41970
rect 21138 41918 21140 41970
rect 20748 41916 21140 41918
rect 20748 41906 20804 41916
rect 21084 41906 21140 41916
rect 20188 41692 20468 41748
rect 19628 41234 19684 41244
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 20188 40404 20244 40414
rect 20412 40404 20468 40414
rect 19516 40350 19518 40402
rect 19570 40350 19572 40402
rect 18732 40292 18788 40302
rect 18788 40236 18900 40292
rect 18732 40198 18788 40236
rect 18060 39554 18116 39564
rect 18396 39732 18452 39742
rect 18172 39508 18228 39518
rect 18396 39508 18452 39676
rect 17500 38782 17502 38834
rect 17554 38782 17556 38834
rect 17500 38770 17556 38782
rect 17948 39394 18004 39406
rect 17948 39342 17950 39394
rect 18002 39342 18004 39394
rect 17948 38834 18004 39342
rect 18060 39396 18116 39406
rect 18060 39302 18116 39340
rect 17948 38782 17950 38834
rect 18002 38782 18004 38834
rect 17948 38668 18004 38782
rect 15708 37286 15764 37324
rect 17612 38612 18004 38668
rect 18172 38668 18228 39452
rect 18284 39506 18452 39508
rect 18284 39454 18398 39506
rect 18450 39454 18452 39506
rect 18284 39452 18452 39454
rect 18284 39058 18340 39452
rect 18396 39442 18452 39452
rect 18844 39506 18900 40236
rect 19068 40180 19124 40190
rect 19068 40178 19460 40180
rect 19068 40126 19070 40178
rect 19122 40126 19460 40178
rect 19068 40124 19460 40126
rect 19068 40114 19124 40124
rect 19404 39730 19460 40124
rect 19404 39678 19406 39730
rect 19458 39678 19460 39730
rect 19404 39666 19460 39678
rect 19180 39620 19236 39630
rect 19180 39526 19236 39564
rect 18844 39454 18846 39506
rect 18898 39454 18900 39506
rect 18844 39442 18900 39454
rect 18284 39006 18286 39058
rect 18338 39006 18340 39058
rect 18284 38994 18340 39006
rect 18620 38834 18676 38846
rect 18620 38782 18622 38834
rect 18674 38782 18676 38834
rect 18620 38668 18676 38782
rect 19068 38722 19124 38734
rect 19068 38670 19070 38722
rect 19122 38670 19124 38722
rect 19068 38668 19124 38670
rect 18172 38612 18564 38668
rect 18620 38612 19124 38668
rect 15932 37266 15988 37278
rect 15932 37214 15934 37266
rect 15986 37214 15988 37266
rect 15596 36542 15598 36594
rect 15650 36542 15652 36594
rect 15596 36530 15652 36542
rect 15820 37044 15876 37054
rect 13468 35588 13524 35598
rect 13580 35588 13636 35598
rect 13468 35586 13580 35588
rect 13468 35534 13470 35586
rect 13522 35534 13580 35586
rect 13468 35532 13580 35534
rect 13468 35522 13524 35532
rect 13468 35140 13524 35150
rect 13468 34130 13524 35084
rect 13468 34078 13470 34130
rect 13522 34078 13524 34130
rect 13468 34066 13524 34078
rect 13580 33348 13636 35532
rect 14476 34914 14532 35868
rect 14812 35858 14868 35868
rect 15260 35586 15316 35598
rect 15260 35534 15262 35586
rect 15314 35534 15316 35586
rect 15148 35476 15204 35486
rect 14476 34862 14478 34914
rect 14530 34862 14532 34914
rect 14476 34850 14532 34862
rect 14812 35474 15204 35476
rect 14812 35422 15150 35474
rect 15202 35422 15204 35474
rect 14812 35420 15204 35422
rect 14812 34914 14868 35420
rect 15148 35410 15204 35420
rect 14812 34862 14814 34914
rect 14866 34862 14868 34914
rect 14812 34850 14868 34862
rect 15036 35252 15092 35262
rect 15036 34914 15092 35196
rect 15036 34862 15038 34914
rect 15090 34862 15092 34914
rect 15036 34850 15092 34862
rect 13804 34802 13860 34814
rect 13804 34750 13806 34802
rect 13858 34750 13860 34802
rect 13692 34692 13748 34702
rect 13692 34598 13748 34636
rect 13692 34132 13748 34142
rect 13692 34038 13748 34076
rect 13692 33348 13748 33358
rect 13580 33292 13692 33348
rect 13692 33254 13748 33292
rect 13244 32510 13246 32562
rect 13298 32510 13300 32562
rect 13244 32498 13300 32510
rect 13692 32562 13748 32574
rect 13692 32510 13694 32562
rect 13746 32510 13748 32562
rect 12908 31166 12910 31218
rect 12962 31166 12964 31218
rect 12908 31154 12964 31166
rect 13468 32450 13524 32462
rect 13468 32398 13470 32450
rect 13522 32398 13524 32450
rect 11900 30994 12628 30996
rect 11900 30942 11902 30994
rect 11954 30942 12628 30994
rect 11900 30940 12628 30942
rect 11900 30930 11956 30940
rect 12572 29652 12628 30940
rect 12684 30436 12740 31052
rect 13356 30996 13412 31006
rect 13468 30996 13524 32398
rect 13692 32452 13748 32510
rect 13692 32386 13748 32396
rect 13692 31780 13748 31818
rect 13692 31714 13748 31724
rect 13804 31668 13860 34750
rect 15260 34804 15316 35534
rect 15372 34914 15428 36428
rect 15820 35698 15876 36988
rect 15932 36596 15988 37214
rect 15932 36530 15988 36540
rect 15820 35646 15822 35698
rect 15874 35646 15876 35698
rect 15820 35634 15876 35646
rect 16828 36372 16884 36382
rect 16268 35588 16324 35598
rect 16156 35586 16324 35588
rect 16156 35534 16270 35586
rect 16322 35534 16324 35586
rect 16156 35532 16324 35534
rect 16156 35364 16212 35532
rect 16268 35522 16324 35532
rect 15484 35252 15540 35262
rect 15484 35026 15540 35196
rect 15484 34974 15486 35026
rect 15538 34974 15540 35026
rect 15484 34962 15540 34974
rect 15372 34862 15374 34914
rect 15426 34862 15428 34914
rect 15372 34850 15428 34862
rect 16044 34916 16100 34926
rect 16044 34822 16100 34860
rect 15260 34738 15316 34748
rect 14700 34690 14756 34702
rect 14700 34638 14702 34690
rect 14754 34638 14756 34690
rect 14700 33460 14756 34638
rect 15148 34692 15204 34702
rect 15148 34242 15204 34636
rect 15148 34190 15150 34242
rect 15202 34190 15204 34242
rect 15148 34178 15204 34190
rect 15596 34690 15652 34702
rect 15596 34638 15598 34690
rect 15650 34638 15652 34690
rect 14924 34020 14980 34030
rect 14924 34018 15204 34020
rect 14924 33966 14926 34018
rect 14978 33966 15204 34018
rect 14924 33964 15204 33966
rect 14924 33954 14980 33964
rect 14700 33394 14756 33404
rect 14364 33348 14420 33358
rect 14812 33348 14868 33358
rect 14364 33346 14644 33348
rect 14364 33294 14366 33346
rect 14418 33294 14644 33346
rect 14364 33292 14644 33294
rect 14364 33282 14420 33292
rect 13916 33236 13972 33246
rect 13916 33142 13972 33180
rect 14028 33122 14084 33134
rect 14028 33070 14030 33122
rect 14082 33070 14084 33122
rect 14028 31892 14084 33070
rect 14028 31826 14084 31836
rect 14364 31780 14420 31790
rect 14364 31686 14420 31724
rect 13804 31602 13860 31612
rect 14476 31666 14532 31678
rect 14476 31614 14478 31666
rect 14530 31614 14532 31666
rect 13692 31554 13748 31566
rect 13692 31502 13694 31554
rect 13746 31502 13748 31554
rect 13692 31332 13748 31502
rect 13916 31556 13972 31566
rect 13692 31266 13748 31276
rect 13804 31444 13860 31454
rect 13356 30994 13524 30996
rect 13356 30942 13358 30994
rect 13410 30942 13524 30994
rect 13356 30940 13524 30942
rect 13580 31106 13636 31118
rect 13580 31054 13582 31106
rect 13634 31054 13636 31106
rect 13580 30996 13636 31054
rect 13804 31106 13860 31388
rect 13804 31054 13806 31106
rect 13858 31054 13860 31106
rect 13804 31042 13860 31054
rect 13580 30940 13748 30996
rect 13356 30930 13412 30940
rect 12684 30322 12740 30380
rect 12684 30270 12686 30322
rect 12738 30270 12740 30322
rect 12684 30258 12740 30270
rect 13468 30436 13524 30446
rect 12684 29652 12740 29662
rect 12572 29650 12740 29652
rect 12572 29598 12686 29650
rect 12738 29598 12740 29650
rect 12572 29596 12740 29598
rect 12684 29586 12740 29596
rect 11228 29374 11230 29426
rect 11282 29374 11284 29426
rect 10668 29316 10724 29326
rect 10668 29222 10724 29260
rect 10220 28756 10276 28766
rect 10220 27970 10276 28700
rect 10220 27918 10222 27970
rect 10274 27918 10276 27970
rect 10220 27906 10276 27918
rect 10780 28308 10836 28318
rect 10444 27860 10500 27870
rect 10444 27766 10500 27804
rect 10780 27858 10836 28252
rect 10780 27806 10782 27858
rect 10834 27806 10836 27858
rect 10780 27794 10836 27806
rect 11004 27858 11060 27870
rect 11004 27806 11006 27858
rect 11058 27806 11060 27858
rect 8092 26350 8094 26402
rect 8146 26350 8148 26402
rect 8092 26180 8148 26350
rect 8988 26962 9044 26974
rect 8988 26910 8990 26962
rect 9042 26910 9044 26962
rect 8092 26114 8148 26124
rect 8652 26180 8708 26190
rect 8652 26086 8708 26124
rect 7756 25454 7758 25506
rect 7810 25454 7812 25506
rect 7756 25442 7812 25454
rect 7868 26066 7924 26078
rect 7868 26014 7870 26066
rect 7922 26014 7924 26066
rect 6636 25342 6638 25394
rect 6690 25342 6692 25394
rect 6636 25330 6692 25342
rect 5964 24782 5966 24834
rect 6018 24782 6020 24834
rect 5964 24770 6020 24782
rect 6300 25284 6356 25294
rect 6300 24722 6356 25228
rect 6748 24836 6804 24846
rect 6300 24670 6302 24722
rect 6354 24670 6356 24722
rect 6300 24658 6356 24670
rect 6412 24834 6804 24836
rect 6412 24782 6750 24834
rect 6802 24782 6804 24834
rect 6412 24780 6804 24782
rect 5852 23846 5908 23884
rect 5740 23828 5796 23838
rect 5740 23734 5796 23772
rect 6412 23604 6468 24780
rect 6748 24770 6804 24780
rect 6860 24722 6916 24734
rect 6860 24670 6862 24722
rect 6914 24670 6916 24722
rect 6748 23828 6804 23838
rect 6860 23828 6916 24670
rect 7868 24050 7924 26014
rect 8204 26068 8260 26078
rect 8204 26066 8484 26068
rect 8204 26014 8206 26066
rect 8258 26014 8484 26066
rect 8204 26012 8484 26014
rect 8204 26002 8260 26012
rect 8428 25618 8484 26012
rect 8428 25566 8430 25618
rect 8482 25566 8484 25618
rect 8428 25554 8484 25566
rect 8988 25508 9044 26910
rect 9212 26964 9268 27002
rect 10108 26982 10164 27020
rect 10668 27746 10724 27758
rect 10668 27694 10670 27746
rect 10722 27694 10724 27746
rect 10668 26908 10724 27694
rect 10780 27636 10836 27646
rect 10780 27186 10836 27580
rect 10780 27134 10782 27186
rect 10834 27134 10836 27186
rect 10780 27122 10836 27134
rect 11004 27188 11060 27806
rect 11228 27860 11284 29374
rect 11452 29538 11508 29550
rect 11452 29486 11454 29538
rect 11506 29486 11508 29538
rect 11452 29428 11508 29486
rect 11452 29362 11508 29372
rect 12572 29428 12628 29438
rect 11900 29316 11956 29326
rect 11956 29260 12180 29316
rect 11900 29222 11956 29260
rect 11676 28530 11732 28542
rect 11676 28478 11678 28530
rect 11730 28478 11732 28530
rect 11676 28420 11732 28478
rect 11676 28364 12068 28420
rect 11676 28196 11732 28206
rect 11676 27972 11732 28140
rect 11900 28196 11956 28206
rect 11788 27972 11844 27982
rect 11676 27970 11844 27972
rect 11676 27918 11790 27970
rect 11842 27918 11844 27970
rect 11676 27916 11844 27918
rect 11228 27794 11284 27804
rect 11788 27748 11844 27916
rect 11788 27682 11844 27692
rect 11676 27636 11732 27646
rect 11676 27542 11732 27580
rect 11004 27122 11060 27132
rect 9212 26898 9268 26908
rect 10444 26852 10724 26908
rect 11116 27076 11172 27086
rect 8988 25442 9044 25452
rect 9548 26180 9604 26190
rect 9548 24946 9604 26124
rect 9548 24894 9550 24946
rect 9602 24894 9604 24946
rect 9548 24882 9604 24894
rect 9884 24722 9940 24734
rect 9884 24670 9886 24722
rect 9938 24670 9940 24722
rect 9884 24612 9940 24670
rect 10332 24612 10388 24622
rect 9884 24610 10388 24612
rect 9884 24558 10334 24610
rect 10386 24558 10388 24610
rect 9884 24556 10388 24558
rect 7868 23998 7870 24050
rect 7922 23998 7924 24050
rect 7868 23986 7924 23998
rect 6972 23940 7028 23950
rect 6972 23846 7028 23884
rect 7196 23938 7252 23950
rect 7196 23886 7198 23938
rect 7250 23886 7252 23938
rect 6804 23772 6916 23828
rect 6748 23762 6804 23772
rect 6412 23266 6468 23548
rect 7196 23492 7252 23886
rect 10332 23940 10388 24556
rect 10332 23874 10388 23884
rect 8316 23828 8372 23838
rect 8316 23734 8372 23772
rect 7196 23426 7252 23436
rect 8204 23714 8260 23726
rect 8204 23662 8206 23714
rect 8258 23662 8260 23714
rect 8204 23492 8260 23662
rect 6412 23214 6414 23266
rect 6466 23214 6468 23266
rect 6412 23202 6468 23214
rect 8204 23156 8260 23436
rect 9324 23268 9380 23278
rect 8204 23100 8708 23156
rect 6524 22932 6580 22942
rect 8540 22932 8596 22942
rect 6524 22838 6580 22876
rect 8316 22876 8540 22932
rect 8204 22370 8260 22382
rect 8204 22318 8206 22370
rect 8258 22318 8260 22370
rect 6188 22260 6244 22270
rect 6188 22166 6244 22204
rect 7196 22260 7252 22270
rect 6300 22146 6356 22158
rect 6300 22094 6302 22146
rect 6354 22094 6356 22146
rect 5852 21644 6132 21700
rect 5740 21588 5796 21598
rect 5852 21588 5908 21644
rect 5628 21586 5908 21588
rect 5628 21534 5742 21586
rect 5794 21534 5908 21586
rect 5628 21532 5908 21534
rect 5740 21522 5796 21532
rect 5404 21364 5460 21374
rect 5404 21270 5460 21308
rect 5068 19854 5070 19906
rect 5122 19854 5124 19906
rect 4956 19236 5012 19246
rect 4844 19180 4956 19236
rect 4956 19170 5012 19180
rect 3500 18732 3892 18788
rect 1820 16882 1876 18396
rect 2828 18452 2884 18462
rect 2828 18358 2884 18396
rect 3500 18450 3556 18732
rect 3500 18398 3502 18450
rect 3554 18398 3556 18450
rect 3500 18386 3556 18398
rect 5068 18452 5124 19854
rect 1932 18228 1988 18238
rect 1932 17890 1988 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17838 1934 17890
rect 1986 17838 1988 17890
rect 1932 17826 1988 17838
rect 4172 17668 4228 17678
rect 4060 17666 4228 17668
rect 4060 17614 4174 17666
rect 4226 17614 4228 17666
rect 4060 17612 4228 17614
rect 1820 16830 1822 16882
rect 1874 16830 1876 16882
rect 1820 16818 1876 16830
rect 1932 17556 1988 17566
rect 1932 16322 1988 17500
rect 2492 16772 2548 16782
rect 2492 16678 2548 16716
rect 1932 16270 1934 16322
rect 1986 16270 1988 16322
rect 1932 16258 1988 16270
rect 3388 16660 3444 16670
rect 2940 15876 2996 15886
rect 2940 15314 2996 15820
rect 2940 15262 2942 15314
rect 2994 15262 2996 15314
rect 2940 15250 2996 15262
rect 3276 15428 3332 15438
rect 3276 15314 3332 15372
rect 3388 15426 3444 16604
rect 4060 16548 4116 17612
rect 4172 17602 4228 17612
rect 4844 17444 4900 17454
rect 5068 17444 5124 18396
rect 5516 20916 5572 20926
rect 5516 19012 5572 20860
rect 5628 20130 5684 20142
rect 5628 20078 5630 20130
rect 5682 20078 5684 20130
rect 5628 20020 5684 20078
rect 5740 20132 5796 20142
rect 5740 20038 5796 20076
rect 5852 20130 5908 21532
rect 5852 20078 5854 20130
rect 5906 20078 5908 20130
rect 5852 20066 5908 20078
rect 5964 21474 6020 21486
rect 5964 21422 5966 21474
rect 6018 21422 6020 21474
rect 5964 20802 6020 21422
rect 5964 20750 5966 20802
rect 6018 20750 6020 20802
rect 5628 19954 5684 19964
rect 5964 20020 6020 20750
rect 6076 20690 6132 21644
rect 6076 20638 6078 20690
rect 6130 20638 6132 20690
rect 6076 20626 6132 20638
rect 6300 20692 6356 22094
rect 6748 21924 6804 21934
rect 6748 21700 6804 21868
rect 6860 21700 6916 21710
rect 6748 21698 6916 21700
rect 6748 21646 6862 21698
rect 6914 21646 6916 21698
rect 6748 21644 6916 21646
rect 6860 21634 6916 21644
rect 7196 21698 7252 22204
rect 8204 22148 8260 22318
rect 8204 22082 8260 22092
rect 8316 21810 8372 22876
rect 8540 22838 8596 22876
rect 8316 21758 8318 21810
rect 8370 21758 8372 21810
rect 8316 21746 8372 21758
rect 8428 22260 8484 22270
rect 7196 21646 7198 21698
rect 7250 21646 7252 21698
rect 7196 21634 7252 21646
rect 7532 21698 7588 21710
rect 7532 21646 7534 21698
rect 7586 21646 7588 21698
rect 6300 20626 6356 20636
rect 6412 21362 6468 21374
rect 6412 21310 6414 21362
rect 6466 21310 6468 21362
rect 6412 20242 6468 21310
rect 6524 21364 6580 21374
rect 6524 20580 6580 21308
rect 6748 21362 6804 21374
rect 6748 21310 6750 21362
rect 6802 21310 6804 21362
rect 6748 21028 6804 21310
rect 6748 20962 6804 20972
rect 6972 20580 7028 20590
rect 6524 20578 7028 20580
rect 6524 20526 6974 20578
rect 7026 20526 7028 20578
rect 6524 20524 7028 20526
rect 6972 20514 7028 20524
rect 6412 20190 6414 20242
rect 6466 20190 6468 20242
rect 6412 20178 6468 20190
rect 6188 20132 6244 20142
rect 6188 20038 6244 20076
rect 6748 20132 6804 20142
rect 6748 20038 6804 20076
rect 7532 20132 7588 21646
rect 8428 21588 8484 22204
rect 8652 21810 8708 23100
rect 8876 23154 8932 23166
rect 8876 23102 8878 23154
rect 8930 23102 8932 23154
rect 8652 21758 8654 21810
rect 8706 21758 8708 21810
rect 8652 21746 8708 21758
rect 8764 23042 8820 23054
rect 8764 22990 8766 23042
rect 8818 22990 8820 23042
rect 8428 21494 8484 21532
rect 8540 21474 8596 21486
rect 8540 21422 8542 21474
rect 8594 21422 8596 21474
rect 7980 20916 8036 20926
rect 8540 20916 8596 21422
rect 7980 20802 8036 20860
rect 7980 20750 7982 20802
rect 8034 20750 8036 20802
rect 7980 20738 8036 20750
rect 8428 20860 8596 20916
rect 5628 19236 5684 19246
rect 5628 19142 5684 19180
rect 5740 19012 5796 19022
rect 5516 19010 5796 19012
rect 5516 18958 5742 19010
rect 5794 18958 5796 19010
rect 5516 18956 5796 18958
rect 5516 18452 5572 18956
rect 5740 18946 5796 18956
rect 5964 18900 6020 19964
rect 5964 18562 6020 18844
rect 5964 18510 5966 18562
rect 6018 18510 6020 18562
rect 5964 18498 6020 18510
rect 6524 20018 6580 20030
rect 6524 19966 6526 20018
rect 6578 19966 6580 20018
rect 6524 19236 6580 19966
rect 7532 19796 7588 20076
rect 7532 19730 7588 19740
rect 8428 19908 8484 20860
rect 8540 20692 8596 20702
rect 8540 20598 8596 20636
rect 8764 20356 8820 22990
rect 8876 22260 8932 23102
rect 8876 22194 8932 22204
rect 8988 22258 9044 22270
rect 8988 22206 8990 22258
rect 9042 22206 9044 22258
rect 8876 21586 8932 21598
rect 8876 21534 8878 21586
rect 8930 21534 8932 21586
rect 8876 20580 8932 21534
rect 8988 21476 9044 22206
rect 8988 21410 9044 21420
rect 9324 20580 9380 23212
rect 10220 22484 10276 22494
rect 10220 20914 10276 22428
rect 10332 21812 10388 21822
rect 10332 21718 10388 21756
rect 10220 20862 10222 20914
rect 10274 20862 10276 20914
rect 10220 20850 10276 20862
rect 8876 20524 9380 20580
rect 8540 20300 8820 20356
rect 8540 20018 8596 20300
rect 8652 20132 8708 20142
rect 8652 20038 8708 20076
rect 8540 19966 8542 20018
rect 8594 19966 8596 20018
rect 8540 19954 8596 19966
rect 8428 19236 8484 19852
rect 8764 19796 8820 20300
rect 8876 20020 8932 20030
rect 8876 19926 8932 19964
rect 9100 20018 9156 20030
rect 9100 19966 9102 20018
rect 9154 19966 9156 20018
rect 9100 19796 9156 19966
rect 8764 19740 9044 19796
rect 8988 19458 9044 19740
rect 9100 19730 9156 19740
rect 9212 19460 9268 19470
rect 8988 19406 8990 19458
rect 9042 19406 9044 19458
rect 8988 19394 9044 19406
rect 9100 19404 9212 19460
rect 8652 19236 8708 19246
rect 8428 19234 8708 19236
rect 8428 19182 8654 19234
rect 8706 19182 8708 19234
rect 8428 19180 8708 19182
rect 5516 18386 5572 18396
rect 6188 18450 6244 18462
rect 6188 18398 6190 18450
rect 6242 18398 6244 18450
rect 5628 18340 5684 18350
rect 5628 18246 5684 18284
rect 6188 18340 6244 18398
rect 4900 17388 5124 17444
rect 5740 17892 5796 17902
rect 4620 16884 4676 16894
rect 4620 16770 4676 16828
rect 4620 16718 4622 16770
rect 4674 16718 4676 16770
rect 4620 16706 4676 16718
rect 4060 16492 4340 16548
rect 4060 16324 4116 16334
rect 4060 16100 4116 16268
rect 3388 15374 3390 15426
rect 3442 15374 3444 15426
rect 3388 15362 3444 15374
rect 3500 16098 4116 16100
rect 3500 16046 4062 16098
rect 4114 16046 4116 16098
rect 3500 16044 4116 16046
rect 3276 15262 3278 15314
rect 3330 15262 3332 15314
rect 3276 15250 3332 15262
rect 2492 14420 2548 14430
rect 2492 13858 2548 14364
rect 2492 13806 2494 13858
rect 2546 13806 2548 13858
rect 2492 13794 2548 13806
rect 1820 13746 1876 13758
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1820 11396 1876 13694
rect 2492 12068 2548 12078
rect 2492 11506 2548 12012
rect 2492 11454 2494 11506
rect 2546 11454 2548 11506
rect 2492 11442 2548 11454
rect 1820 11302 1876 11340
rect 3500 10500 3556 16044
rect 4060 16034 4116 16044
rect 4172 15764 4228 15774
rect 3836 15428 3892 15438
rect 3836 15334 3892 15372
rect 4172 15426 4228 15708
rect 4172 15374 4174 15426
rect 4226 15374 4228 15426
rect 4172 15362 4228 15374
rect 3948 15202 4004 15214
rect 3948 15150 3950 15202
rect 4002 15150 4004 15202
rect 3948 15148 4004 15150
rect 3948 15092 4116 15148
rect 3948 14980 4004 14990
rect 3724 14530 3780 14542
rect 3724 14478 3726 14530
rect 3778 14478 3780 14530
rect 3612 14420 3668 14430
rect 3612 14326 3668 14364
rect 3724 13412 3780 14478
rect 3948 14530 4004 14924
rect 4060 14754 4116 15092
rect 4284 14756 4340 16492
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4844 16212 4900 17388
rect 5740 17108 5796 17836
rect 6188 17668 6244 18284
rect 6188 17602 6244 17612
rect 6412 17780 6468 17790
rect 5852 17444 5908 17454
rect 5852 17350 5908 17388
rect 5292 17106 5796 17108
rect 5292 17054 5742 17106
rect 5794 17054 5796 17106
rect 5292 17052 5796 17054
rect 5180 16884 5236 16894
rect 5068 16772 5124 16782
rect 5068 16678 5124 16716
rect 4956 16660 5012 16670
rect 5180 16660 5236 16828
rect 5292 16882 5348 17052
rect 5740 17042 5796 17052
rect 5292 16830 5294 16882
rect 5346 16830 5348 16882
rect 5292 16818 5348 16830
rect 6412 16994 6468 17724
rect 6524 17666 6580 19180
rect 8652 19170 8708 19180
rect 8316 19010 8372 19022
rect 8316 18958 8318 19010
rect 8370 18958 8372 19010
rect 6972 18900 7028 18910
rect 6972 18674 7028 18844
rect 6972 18622 6974 18674
rect 7026 18622 7028 18674
rect 6972 18610 7028 18622
rect 7084 18676 7140 18686
rect 7084 18582 7140 18620
rect 8092 18562 8148 18574
rect 8092 18510 8094 18562
rect 8146 18510 8148 18562
rect 6748 18452 6804 18462
rect 6748 18450 7140 18452
rect 6748 18398 6750 18450
rect 6802 18398 7140 18450
rect 6748 18396 7140 18398
rect 6748 18386 6804 18396
rect 6972 18228 7028 18238
rect 6860 18172 6972 18228
rect 6860 17778 6916 18172
rect 6972 18162 7028 18172
rect 6860 17726 6862 17778
rect 6914 17726 6916 17778
rect 6860 17714 6916 17726
rect 6524 17614 6526 17666
rect 6578 17614 6580 17666
rect 6524 17602 6580 17614
rect 6972 17668 7028 17678
rect 6972 17574 7028 17612
rect 6412 16942 6414 16994
rect 6466 16942 6468 16994
rect 5180 16604 5348 16660
rect 4956 16566 5012 16604
rect 5180 16436 5236 16446
rect 4956 16212 5012 16222
rect 4844 16210 5012 16212
rect 4844 16158 4958 16210
rect 5010 16158 5012 16210
rect 4844 16156 5012 16158
rect 4956 16146 5012 16156
rect 5180 15428 5236 16380
rect 5180 15334 5236 15372
rect 5292 15764 5348 16604
rect 6412 16324 6468 16942
rect 6412 16258 6468 16268
rect 6748 17442 6804 17454
rect 6748 17390 6750 17442
rect 6802 17390 6804 17442
rect 6748 16994 6804 17390
rect 6748 16942 6750 16994
rect 6802 16942 6804 16994
rect 6412 16100 6468 16110
rect 6300 16098 6468 16100
rect 6300 16046 6414 16098
rect 6466 16046 6468 16098
rect 6300 16044 6468 16046
rect 6188 15988 6244 15998
rect 6188 15894 6244 15932
rect 5292 15426 5348 15708
rect 5292 15374 5294 15426
rect 5346 15374 5348 15426
rect 5292 15362 5348 15374
rect 5964 15876 6020 15886
rect 4396 15316 4452 15326
rect 4396 15222 4452 15260
rect 5516 15316 5572 15326
rect 5964 15316 6020 15820
rect 6188 15764 6244 15774
rect 5572 15260 6020 15316
rect 5516 15222 5572 15260
rect 4396 15092 4452 15102
rect 4732 15092 4788 15102
rect 4452 15090 4788 15092
rect 4452 15038 4734 15090
rect 4786 15038 4788 15090
rect 4452 15036 4788 15038
rect 4396 15026 4452 15036
rect 4732 15026 4788 15036
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4060 14702 4062 14754
rect 4114 14702 4116 14754
rect 4060 14690 4116 14702
rect 4172 14700 4340 14756
rect 3948 14478 3950 14530
rect 4002 14478 4004 14530
rect 3724 13346 3780 13356
rect 3836 13748 3892 13758
rect 3836 12178 3892 13692
rect 3836 12126 3838 12178
rect 3890 12126 3892 12178
rect 3836 12114 3892 12126
rect 3948 12740 4004 14478
rect 3948 12066 4004 12684
rect 3948 12014 3950 12066
rect 4002 12014 4004 12066
rect 3948 12002 4004 12014
rect 3500 10444 4004 10500
rect 3948 9268 4004 10444
rect 1708 8148 1764 8158
rect 1708 8054 1764 8092
rect 2044 8148 2100 8158
rect 2044 8054 2100 8092
rect 2492 8036 2548 8046
rect 2492 7942 2548 7980
rect 3948 7698 4004 9212
rect 3948 7646 3950 7698
rect 4002 7646 4004 7698
rect 3948 7634 4004 7646
rect 4172 7700 4228 14700
rect 5068 14532 5124 14542
rect 5068 14438 5124 14476
rect 4956 14420 5012 14430
rect 4732 14364 4956 14420
rect 4620 14308 4676 14318
rect 4508 14306 4676 14308
rect 4508 14254 4622 14306
rect 4674 14254 4676 14306
rect 4508 14252 4676 14254
rect 4284 13748 4340 13758
rect 4284 13076 4340 13692
rect 4508 13524 4564 14252
rect 4620 14242 4676 14252
rect 4620 13636 4676 13646
rect 4732 13636 4788 14364
rect 4956 14326 5012 14364
rect 5628 14420 5684 14430
rect 5628 14326 5684 14364
rect 5964 14418 6020 15260
rect 6076 15428 6132 15438
rect 6076 15148 6132 15372
rect 6188 15426 6244 15708
rect 6188 15374 6190 15426
rect 6242 15374 6244 15426
rect 6188 15362 6244 15374
rect 6300 15538 6356 16044
rect 6412 16034 6468 16044
rect 6748 16100 6804 16942
rect 7084 16100 7140 18396
rect 7196 18450 7252 18462
rect 7196 18398 7198 18450
rect 7250 18398 7252 18450
rect 7196 17780 7252 18398
rect 7308 18452 7364 18462
rect 7308 18358 7364 18396
rect 7868 18452 7924 18462
rect 7868 18358 7924 18396
rect 7196 17714 7252 17724
rect 7196 17556 7252 17566
rect 7196 17554 7476 17556
rect 7196 17502 7198 17554
rect 7250 17502 7476 17554
rect 7196 17500 7476 17502
rect 7196 17490 7252 17500
rect 7420 16882 7476 17500
rect 7420 16830 7422 16882
rect 7474 16830 7476 16882
rect 7308 16324 7364 16334
rect 7420 16324 7476 16830
rect 7644 16772 7700 16782
rect 7644 16770 7924 16772
rect 7644 16718 7646 16770
rect 7698 16718 7924 16770
rect 7644 16716 7924 16718
rect 7644 16706 7700 16716
rect 7308 16322 7700 16324
rect 7308 16270 7310 16322
rect 7362 16270 7700 16322
rect 7308 16268 7700 16270
rect 7308 16258 7364 16268
rect 7196 16100 7252 16110
rect 6748 16034 6804 16044
rect 6860 16098 7252 16100
rect 6860 16046 7198 16098
rect 7250 16046 7252 16098
rect 6860 16044 7252 16046
rect 6300 15486 6302 15538
rect 6354 15486 6356 15538
rect 6076 15092 6244 15148
rect 5964 14366 5966 14418
rect 6018 14366 6020 14418
rect 5964 14354 6020 14366
rect 4620 13634 4788 13636
rect 4620 13582 4622 13634
rect 4674 13582 4788 13634
rect 4620 13580 4788 13582
rect 5068 13634 5124 13646
rect 5068 13582 5070 13634
rect 5122 13582 5124 13634
rect 4620 13570 4676 13580
rect 4508 13458 4564 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4396 13076 4452 13086
rect 4284 13074 4452 13076
rect 4284 13022 4398 13074
rect 4450 13022 4452 13074
rect 4284 13020 4452 13022
rect 4396 13010 4452 13020
rect 4732 12852 4788 12862
rect 4732 12758 4788 12796
rect 4844 12290 4900 12302
rect 4844 12238 4846 12290
rect 4898 12238 4900 12290
rect 4844 12180 4900 12238
rect 4844 12114 4900 12124
rect 4284 12068 4340 12078
rect 4620 12068 4676 12078
rect 4284 12066 4676 12068
rect 4284 12014 4286 12066
rect 4338 12014 4622 12066
rect 4674 12014 4676 12066
rect 4284 12012 4676 12014
rect 4284 12002 4340 12012
rect 4620 12002 4676 12012
rect 4732 12068 4788 12078
rect 4732 11974 4788 12012
rect 4844 11956 4900 11966
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4732 11620 4788 11630
rect 4620 11564 4732 11620
rect 4620 11506 4676 11564
rect 4732 11554 4788 11564
rect 4620 11454 4622 11506
rect 4674 11454 4676 11506
rect 4620 11442 4676 11454
rect 4844 10724 4900 11900
rect 5068 11396 5124 13582
rect 6188 13076 6244 15092
rect 6300 14420 6356 15486
rect 6300 14354 6356 14364
rect 6748 14530 6804 14542
rect 6748 14478 6750 14530
rect 6802 14478 6804 14530
rect 6748 13748 6804 14478
rect 6860 13860 6916 16044
rect 7196 16034 7252 16044
rect 7644 16098 7700 16268
rect 7644 16046 7646 16098
rect 7698 16046 7700 16098
rect 7084 15428 7140 15438
rect 7084 15426 7252 15428
rect 7084 15374 7086 15426
rect 7138 15374 7252 15426
rect 7084 15372 7252 15374
rect 7084 15362 7140 15372
rect 6972 15314 7028 15326
rect 6972 15262 6974 15314
rect 7026 15262 7028 15314
rect 6972 14084 7028 15262
rect 7084 15090 7140 15102
rect 7084 15038 7086 15090
rect 7138 15038 7140 15090
rect 7084 14756 7140 15038
rect 7196 15092 7252 15372
rect 7644 15314 7700 16046
rect 7868 16098 7924 16716
rect 8092 16660 8148 18510
rect 8204 18340 8260 18350
rect 8316 18340 8372 18958
rect 8428 19010 8484 19022
rect 8428 18958 8430 19010
rect 8482 18958 8484 19010
rect 8428 18452 8484 18958
rect 8540 19010 8596 19022
rect 8540 18958 8542 19010
rect 8594 18958 8596 19010
rect 8540 18676 8596 18958
rect 8652 18676 8708 18686
rect 8540 18620 8652 18676
rect 8652 18582 8708 18620
rect 8876 18676 8932 18686
rect 9100 18676 9156 19404
rect 9212 19366 9268 19404
rect 9324 18788 9380 20524
rect 10108 20580 10164 20590
rect 10108 20578 10276 20580
rect 10108 20526 10110 20578
rect 10162 20526 10276 20578
rect 10108 20524 10276 20526
rect 10108 20514 10164 20524
rect 9884 20132 9940 20142
rect 9660 19796 9716 19806
rect 9716 19740 9828 19796
rect 9660 19702 9716 19740
rect 9772 19234 9828 19740
rect 9772 19182 9774 19234
rect 9826 19182 9828 19234
rect 9772 19170 9828 19182
rect 9884 19010 9940 20076
rect 9884 18958 9886 19010
rect 9938 18958 9940 19010
rect 9660 18788 9716 18798
rect 9324 18732 9660 18788
rect 8876 18674 9156 18676
rect 8876 18622 8878 18674
rect 8930 18622 9156 18674
rect 8876 18620 9156 18622
rect 8876 18610 8932 18620
rect 8428 18386 8484 18396
rect 8540 18450 8596 18462
rect 8540 18398 8542 18450
rect 8594 18398 8596 18450
rect 8204 18338 8372 18340
rect 8204 18286 8206 18338
rect 8258 18286 8372 18338
rect 8204 18284 8372 18286
rect 8204 18274 8260 18284
rect 8540 18228 8596 18398
rect 8540 18162 8596 18172
rect 8876 18340 8932 18350
rect 8428 16882 8484 16894
rect 8428 16830 8430 16882
rect 8482 16830 8484 16882
rect 7868 16046 7870 16098
rect 7922 16046 7924 16098
rect 7868 15876 7924 16046
rect 7868 15810 7924 15820
rect 7980 16604 8148 16660
rect 8204 16660 8260 16670
rect 7756 15428 7812 15438
rect 7756 15334 7812 15372
rect 7644 15262 7646 15314
rect 7698 15262 7700 15314
rect 7644 15250 7700 15262
rect 7196 15026 7252 15036
rect 7084 14690 7140 14700
rect 7868 14420 7924 14430
rect 7756 14418 7924 14420
rect 7756 14366 7870 14418
rect 7922 14366 7924 14418
rect 7756 14364 7924 14366
rect 6972 14028 7476 14084
rect 7420 13972 7476 14028
rect 7420 13878 7476 13916
rect 7084 13860 7140 13870
rect 6860 13858 7140 13860
rect 6860 13806 7086 13858
rect 7138 13806 7140 13858
rect 6860 13804 7140 13806
rect 6748 13682 6804 13692
rect 5852 13020 6244 13076
rect 5292 12852 5348 12862
rect 5292 12402 5348 12796
rect 5292 12350 5294 12402
rect 5346 12350 5348 12402
rect 5292 11844 5348 12350
rect 5292 11778 5348 11788
rect 5740 12180 5796 12190
rect 5068 11170 5124 11340
rect 5068 11118 5070 11170
rect 5122 11118 5124 11170
rect 4956 10724 5012 10734
rect 4844 10722 5012 10724
rect 4844 10670 4958 10722
rect 5010 10670 5012 10722
rect 4844 10668 5012 10670
rect 4956 10658 5012 10668
rect 4284 10610 4340 10622
rect 4284 10558 4286 10610
rect 4338 10558 4340 10610
rect 4284 10500 4340 10558
rect 4284 10434 4340 10444
rect 5068 10500 5124 11118
rect 5068 10434 5124 10444
rect 5740 11170 5796 12124
rect 5852 12178 5908 13020
rect 6188 12964 6244 13020
rect 6636 13412 6692 13422
rect 6300 12964 6356 12974
rect 6188 12962 6356 12964
rect 6188 12910 6302 12962
rect 6354 12910 6356 12962
rect 6188 12908 6356 12910
rect 6300 12898 6356 12908
rect 6524 12962 6580 12974
rect 6524 12910 6526 12962
rect 6578 12910 6580 12962
rect 6076 12850 6132 12862
rect 6076 12798 6078 12850
rect 6130 12798 6132 12850
rect 5964 12740 6020 12750
rect 6076 12740 6132 12798
rect 6020 12684 6132 12740
rect 6188 12738 6244 12750
rect 6188 12686 6190 12738
rect 6242 12686 6244 12738
rect 5964 12674 6020 12684
rect 5852 12126 5854 12178
rect 5906 12126 5908 12178
rect 5852 12114 5908 12126
rect 6188 12178 6244 12686
rect 6188 12126 6190 12178
rect 6242 12126 6244 12178
rect 6188 12114 6244 12126
rect 6412 12292 6468 12302
rect 6412 12178 6468 12236
rect 6412 12126 6414 12178
rect 6466 12126 6468 12178
rect 6412 12114 6468 12126
rect 6524 12068 6580 12910
rect 6636 12404 6692 13356
rect 6636 12178 6692 12348
rect 6636 12126 6638 12178
rect 6690 12126 6692 12178
rect 6636 12114 6692 12126
rect 6524 12002 6580 12012
rect 6748 11956 6804 11966
rect 6748 11862 6804 11900
rect 5740 11118 5742 11170
rect 5794 11118 5796 11170
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 5740 8372 5796 11118
rect 6972 8484 7028 13804
rect 7084 13794 7140 13804
rect 7196 13860 7252 13870
rect 7196 12404 7252 13804
rect 7756 13860 7812 14364
rect 7868 14354 7924 14364
rect 7308 13748 7364 13758
rect 7308 13654 7364 13692
rect 7532 13748 7588 13758
rect 7308 12404 7364 12414
rect 7196 12402 7364 12404
rect 7196 12350 7310 12402
rect 7362 12350 7364 12402
rect 7196 12348 7364 12350
rect 7308 12338 7364 12348
rect 7196 12178 7252 12190
rect 7196 12126 7198 12178
rect 7250 12126 7252 12178
rect 7084 11396 7140 11406
rect 7196 11396 7252 12126
rect 7420 12068 7476 12078
rect 7420 11506 7476 12012
rect 7532 11956 7588 13692
rect 7756 13746 7812 13804
rect 7756 13694 7758 13746
rect 7810 13694 7812 13746
rect 7756 13682 7812 13694
rect 7980 13748 8036 16604
rect 8204 16566 8260 16604
rect 8204 16212 8260 16222
rect 8204 16118 8260 16156
rect 8092 16100 8148 16110
rect 8092 16006 8148 16044
rect 8204 15874 8260 15886
rect 8204 15822 8206 15874
rect 8258 15822 8260 15874
rect 8204 15428 8260 15822
rect 8428 15764 8484 16830
rect 8876 16882 8932 18284
rect 8876 16830 8878 16882
rect 8930 16830 8932 16882
rect 8876 16818 8932 16830
rect 8428 15698 8484 15708
rect 8764 16100 8820 16110
rect 8204 15362 8260 15372
rect 8764 15426 8820 16044
rect 8764 15374 8766 15426
rect 8818 15374 8820 15426
rect 8764 15362 8820 15374
rect 9100 16098 9156 16110
rect 9100 16046 9102 16098
rect 9154 16046 9156 16098
rect 9100 15428 9156 16046
rect 9660 15764 9716 18732
rect 9660 15698 9716 15708
rect 9772 16210 9828 16222
rect 9772 16158 9774 16210
rect 9826 16158 9828 16210
rect 9100 15362 9156 15372
rect 8428 15316 8484 15326
rect 8316 15202 8372 15214
rect 8316 15150 8318 15202
rect 8370 15150 8372 15202
rect 8316 15148 8372 15150
rect 7980 13682 8036 13692
rect 8204 15092 8372 15148
rect 8204 13746 8260 15036
rect 8204 13694 8206 13746
rect 8258 13694 8260 13746
rect 8204 13636 8260 13694
rect 8316 13748 8372 13758
rect 8316 13654 8372 13692
rect 8204 13570 8260 13580
rect 7756 12404 7812 12414
rect 7756 12310 7812 12348
rect 8428 12068 8484 15260
rect 8988 15316 9044 15326
rect 8988 15222 9044 15260
rect 9772 15316 9828 16158
rect 9772 15250 9828 15260
rect 9884 15148 9940 18958
rect 9996 19794 10052 19806
rect 9996 19742 9998 19794
rect 10050 19742 10052 19794
rect 9996 19012 10052 19742
rect 10220 19124 10276 20524
rect 10332 20020 10388 20030
rect 10332 19926 10388 19964
rect 10444 19796 10500 26852
rect 10556 25618 10612 25630
rect 10556 25566 10558 25618
rect 10610 25566 10612 25618
rect 10556 25172 10612 25566
rect 10556 23828 10612 25116
rect 11116 24722 11172 27020
rect 11788 26964 11844 26974
rect 11900 26908 11956 28140
rect 12012 27970 12068 28364
rect 12012 27918 12014 27970
rect 12066 27918 12068 27970
rect 12012 27906 12068 27918
rect 11788 26852 11956 26908
rect 11340 25956 11396 25966
rect 11340 25506 11396 25900
rect 11340 25454 11342 25506
rect 11394 25454 11396 25506
rect 11340 25442 11396 25454
rect 11564 25508 11620 25518
rect 11564 25414 11620 25452
rect 11788 25506 11844 26852
rect 12124 26180 12180 29260
rect 12348 28868 12404 28878
rect 12348 28642 12404 28812
rect 12572 28754 12628 29372
rect 12572 28702 12574 28754
rect 12626 28702 12628 28754
rect 12572 28690 12628 28702
rect 12348 28590 12350 28642
rect 12402 28590 12404 28642
rect 12348 28578 12404 28590
rect 13468 28644 13524 30380
rect 13580 29876 13636 29886
rect 13580 29650 13636 29820
rect 13580 29598 13582 29650
rect 13634 29598 13636 29650
rect 13580 29586 13636 29598
rect 13692 29316 13748 30940
rect 13804 30884 13860 30894
rect 13804 30324 13860 30828
rect 13804 30098 13860 30268
rect 13916 30322 13972 31500
rect 14476 31556 14532 31614
rect 14476 31490 14532 31500
rect 14588 31220 14644 33292
rect 14588 31154 14644 31164
rect 14812 32674 14868 33292
rect 14924 33122 14980 33134
rect 14924 33070 14926 33122
rect 14978 33070 14980 33122
rect 14924 33012 14980 33070
rect 14924 32946 14980 32956
rect 14812 32622 14814 32674
rect 14866 32622 14868 32674
rect 14476 30884 14532 30894
rect 14476 30790 14532 30828
rect 14812 30660 14868 32622
rect 15036 31780 15092 31790
rect 14364 30604 14868 30660
rect 14924 31668 14980 31678
rect 13916 30270 13918 30322
rect 13970 30270 13972 30322
rect 13916 30258 13972 30270
rect 14252 30324 14308 30334
rect 13804 30046 13806 30098
rect 13858 30046 13860 30098
rect 13804 30034 13860 30046
rect 14028 30098 14084 30110
rect 14028 30046 14030 30098
rect 14082 30046 14084 30098
rect 13916 29316 13972 29326
rect 13692 29314 13972 29316
rect 13692 29262 13918 29314
rect 13970 29262 13972 29314
rect 13692 29260 13972 29262
rect 13580 28868 13636 28878
rect 13580 28774 13636 28812
rect 13468 28588 13636 28644
rect 12460 27748 12516 27758
rect 12460 26908 12516 27692
rect 12908 27186 12964 27198
rect 12908 27134 12910 27186
rect 12962 27134 12964 27186
rect 12908 26964 12964 27134
rect 13580 27076 13636 28588
rect 13580 27010 13636 27020
rect 13692 28530 13748 28542
rect 13692 28478 13694 28530
rect 13746 28478 13748 28530
rect 13692 27858 13748 28478
rect 13692 27806 13694 27858
rect 13746 27806 13748 27858
rect 12460 26852 12852 26908
rect 12908 26898 12964 26908
rect 13468 26962 13524 26974
rect 13468 26910 13470 26962
rect 13522 26910 13524 26962
rect 12124 26114 12180 26124
rect 11788 25454 11790 25506
rect 11842 25454 11844 25506
rect 11788 25442 11844 25454
rect 11900 25956 11956 25966
rect 11228 25282 11284 25294
rect 11228 25230 11230 25282
rect 11282 25230 11284 25282
rect 11228 25172 11284 25230
rect 11228 25106 11284 25116
rect 11452 25282 11508 25294
rect 11452 25230 11454 25282
rect 11506 25230 11508 25282
rect 11116 24670 11118 24722
rect 11170 24670 11172 24722
rect 11116 24658 11172 24670
rect 10556 23762 10612 23772
rect 11452 23380 11508 25230
rect 11900 24836 11956 25900
rect 11788 24780 11956 24836
rect 11788 24164 11844 24780
rect 11900 24612 11956 24622
rect 11900 24610 12516 24612
rect 11900 24558 11902 24610
rect 11954 24558 12516 24610
rect 11900 24556 12516 24558
rect 11900 24546 11956 24556
rect 11900 24164 11956 24174
rect 11788 24162 11956 24164
rect 11788 24110 11902 24162
rect 11954 24110 11956 24162
rect 11788 24108 11956 24110
rect 11900 24098 11956 24108
rect 10780 23324 11508 23380
rect 12012 23826 12068 23838
rect 12012 23774 12014 23826
rect 12066 23774 12068 23826
rect 12012 23716 12068 23774
rect 12348 23716 12404 23726
rect 12012 23714 12404 23716
rect 12012 23662 12350 23714
rect 12402 23662 12404 23714
rect 12012 23660 12404 23662
rect 10556 23044 10612 23054
rect 10556 22148 10612 22988
rect 10556 22082 10612 22092
rect 10668 21588 10724 21598
rect 10668 21494 10724 21532
rect 10780 20130 10836 23324
rect 12012 23268 12068 23660
rect 12348 23650 12404 23660
rect 12012 23202 12068 23212
rect 11340 23154 11396 23166
rect 11340 23102 11342 23154
rect 11394 23102 11396 23154
rect 10892 23042 10948 23054
rect 10892 22990 10894 23042
rect 10946 22990 10948 23042
rect 10892 21588 10948 22990
rect 11116 22484 11172 22494
rect 11340 22484 11396 23102
rect 11900 23044 11956 23054
rect 11900 23042 12068 23044
rect 11900 22990 11902 23042
rect 11954 22990 12068 23042
rect 11900 22988 12068 22990
rect 11900 22978 11956 22988
rect 11172 22428 11396 22484
rect 11788 22930 11844 22942
rect 11788 22878 11790 22930
rect 11842 22878 11844 22930
rect 11116 22390 11172 22428
rect 11452 22148 11508 22158
rect 11004 22146 11508 22148
rect 11004 22094 11454 22146
rect 11506 22094 11508 22146
rect 11004 22092 11508 22094
rect 11004 21810 11060 22092
rect 11004 21758 11006 21810
rect 11058 21758 11060 21810
rect 11004 21746 11060 21758
rect 10892 21522 10948 21532
rect 11116 21588 11172 21598
rect 11116 20578 11172 21532
rect 11116 20526 11118 20578
rect 11170 20526 11172 20578
rect 11116 20188 11172 20526
rect 10780 20078 10782 20130
rect 10834 20078 10836 20130
rect 10780 20066 10836 20078
rect 10892 20132 11172 20188
rect 10556 20020 10612 20030
rect 10556 20018 10724 20020
rect 10556 19966 10558 20018
rect 10610 19966 10724 20018
rect 10556 19964 10724 19966
rect 10556 19954 10612 19964
rect 10444 19740 10612 19796
rect 10556 19234 10612 19740
rect 10668 19348 10724 19964
rect 10668 19282 10724 19292
rect 10556 19182 10558 19234
rect 10610 19182 10612 19234
rect 10556 19170 10612 19182
rect 10780 19236 10836 19246
rect 10220 19068 10388 19124
rect 9996 18946 10052 18956
rect 10108 19012 10164 19022
rect 10108 19010 10276 19012
rect 10108 18958 10110 19010
rect 10162 18958 10276 19010
rect 10108 18956 10276 18958
rect 10108 18946 10164 18956
rect 9996 18452 10052 18462
rect 10220 18452 10276 18956
rect 10332 18676 10388 19068
rect 10332 18610 10388 18620
rect 10444 19122 10500 19134
rect 10444 19070 10446 19122
rect 10498 19070 10500 19122
rect 10444 18674 10500 19070
rect 10444 18622 10446 18674
rect 10498 18622 10500 18674
rect 10444 18610 10500 18622
rect 10556 19012 10612 19022
rect 10332 18452 10388 18462
rect 10220 18450 10388 18452
rect 10220 18398 10334 18450
rect 10386 18398 10388 18450
rect 10220 18396 10388 18398
rect 9996 18358 10052 18396
rect 10332 18386 10388 18396
rect 10556 18450 10612 18956
rect 10556 18398 10558 18450
rect 10610 18398 10612 18450
rect 10556 18386 10612 18398
rect 10780 18450 10836 19180
rect 10780 18398 10782 18450
rect 10834 18398 10836 18450
rect 10780 18386 10836 18398
rect 10892 18228 10948 20132
rect 11004 20018 11060 20030
rect 11004 19966 11006 20018
rect 11058 19966 11060 20018
rect 11004 19908 11060 19966
rect 11004 19842 11060 19852
rect 11116 19906 11172 19918
rect 11116 19854 11118 19906
rect 11170 19854 11172 19906
rect 11004 19460 11060 19470
rect 11116 19460 11172 19854
rect 11228 19460 11284 19470
rect 11116 19458 11284 19460
rect 11116 19406 11230 19458
rect 11282 19406 11284 19458
rect 11116 19404 11284 19406
rect 11004 19366 11060 19404
rect 11228 19394 11284 19404
rect 11340 19236 11396 22092
rect 11452 22082 11508 22092
rect 11564 22146 11620 22158
rect 11564 22094 11566 22146
rect 11618 22094 11620 22146
rect 11564 21586 11620 22094
rect 11676 22146 11732 22158
rect 11676 22094 11678 22146
rect 11730 22094 11732 22146
rect 11676 21812 11732 22094
rect 11788 21924 11844 22878
rect 12012 22036 12068 22988
rect 12348 23042 12404 23054
rect 12348 22990 12350 23042
rect 12402 22990 12404 23042
rect 12348 22484 12404 22990
rect 12124 22428 12348 22484
rect 12124 22370 12180 22428
rect 12348 22418 12404 22428
rect 12460 22482 12516 24556
rect 12572 24500 12628 24510
rect 12572 23938 12628 24444
rect 12572 23886 12574 23938
rect 12626 23886 12628 23938
rect 12572 23874 12628 23886
rect 12796 23268 12852 26852
rect 13468 25844 13524 26910
rect 13692 26964 13748 27806
rect 13692 26898 13748 26908
rect 13804 27074 13860 27086
rect 13804 27022 13806 27074
rect 13858 27022 13860 27074
rect 13692 26740 13748 26750
rect 13468 25788 13636 25844
rect 13468 25620 13524 25630
rect 12796 23212 13076 23268
rect 12796 23044 12852 23054
rect 12460 22430 12462 22482
rect 12514 22430 12516 22482
rect 12460 22418 12516 22430
rect 12684 23042 12852 23044
rect 12684 22990 12798 23042
rect 12850 22990 12852 23042
rect 12684 22988 12852 22990
rect 12124 22318 12126 22370
rect 12178 22318 12180 22370
rect 12124 22306 12180 22318
rect 12348 22258 12404 22270
rect 12348 22206 12350 22258
rect 12402 22206 12404 22258
rect 12012 21980 12180 22036
rect 11788 21868 12068 21924
rect 11676 21746 11732 21756
rect 12012 21698 12068 21868
rect 12012 21646 12014 21698
rect 12066 21646 12068 21698
rect 12012 21634 12068 21646
rect 11564 21534 11566 21586
rect 11618 21534 11620 21586
rect 11564 21522 11620 21534
rect 11676 21588 11732 21598
rect 11900 21588 11956 21598
rect 11676 21494 11732 21532
rect 11788 21586 11956 21588
rect 11788 21534 11902 21586
rect 11954 21534 11956 21586
rect 11788 21532 11956 21534
rect 11788 21476 11844 21532
rect 11900 21522 11956 21532
rect 11788 21410 11844 21420
rect 12124 21252 12180 21980
rect 12348 21812 12404 22206
rect 12684 22258 12740 22988
rect 12796 22978 12852 22988
rect 12684 22206 12686 22258
rect 12738 22206 12740 22258
rect 12460 21812 12516 21822
rect 12348 21810 12516 21812
rect 12348 21758 12462 21810
rect 12514 21758 12516 21810
rect 12348 21756 12516 21758
rect 12460 21746 12516 21756
rect 12572 21700 12628 21710
rect 12572 21606 12628 21644
rect 12684 21588 12740 22206
rect 12908 22260 12964 22270
rect 12908 22166 12964 22204
rect 12684 21522 12740 21532
rect 12124 21186 12180 21196
rect 12908 20692 12964 20702
rect 12908 20130 12964 20636
rect 12908 20078 12910 20130
rect 12962 20078 12964 20130
rect 12908 20066 12964 20078
rect 12124 20020 12180 20030
rect 11116 19180 11396 19236
rect 11788 19964 12124 20020
rect 11004 18452 11060 18462
rect 11004 18358 11060 18396
rect 10892 18172 11060 18228
rect 10892 17668 10948 17678
rect 10892 17574 10948 17612
rect 10444 16882 10500 16894
rect 10444 16830 10446 16882
rect 10498 16830 10500 16882
rect 10220 16324 10276 16334
rect 9996 16100 10052 16110
rect 9996 15986 10052 16044
rect 9996 15934 9998 15986
rect 10050 15934 10052 15986
rect 9996 15922 10052 15934
rect 10108 16098 10164 16110
rect 10108 16046 10110 16098
rect 10162 16046 10164 16098
rect 9996 15764 10052 15774
rect 9996 15314 10052 15708
rect 9996 15262 9998 15314
rect 10050 15262 10052 15314
rect 9996 15250 10052 15262
rect 10108 15148 10164 16046
rect 10220 15988 10276 16268
rect 10444 16100 10500 16830
rect 10556 16882 10612 16894
rect 10556 16830 10558 16882
rect 10610 16830 10612 16882
rect 10556 16212 10612 16830
rect 10892 16882 10948 16894
rect 10892 16830 10894 16882
rect 10946 16830 10948 16882
rect 10780 16772 10836 16782
rect 10780 16678 10836 16716
rect 10892 16660 10948 16830
rect 10892 16594 10948 16604
rect 10612 16156 10948 16212
rect 10556 16146 10612 16156
rect 10444 16034 10500 16044
rect 10220 15316 10276 15932
rect 10220 15250 10276 15260
rect 10444 15314 10500 15326
rect 10444 15262 10446 15314
rect 10498 15262 10500 15314
rect 9884 15092 10052 15148
rect 10108 15092 10276 15148
rect 8764 14532 8820 14542
rect 8764 14438 8820 14476
rect 9324 14420 9380 14430
rect 9324 14326 9380 14364
rect 9660 13972 9716 13982
rect 8652 13860 8708 13870
rect 8652 13766 8708 13804
rect 9660 13858 9716 13916
rect 9660 13806 9662 13858
rect 9714 13806 9716 13858
rect 9660 13794 9716 13806
rect 9884 13860 9940 13870
rect 9884 13766 9940 13804
rect 8540 13634 8596 13646
rect 8540 13582 8542 13634
rect 8594 13582 8596 13634
rect 8540 13076 8596 13582
rect 9548 13636 9604 13646
rect 9548 13542 9604 13580
rect 9884 13524 9940 13534
rect 9212 13188 9268 13198
rect 8540 13010 8596 13020
rect 8988 13132 9212 13188
rect 8988 12850 9044 13132
rect 9212 13122 9268 13132
rect 8988 12798 8990 12850
rect 9042 12798 9044 12850
rect 8988 12786 9044 12798
rect 8876 12740 8932 12750
rect 8764 12628 8820 12638
rect 8652 12292 8708 12302
rect 8652 12198 8708 12236
rect 8428 12002 8484 12012
rect 7532 11900 7700 11956
rect 7420 11454 7422 11506
rect 7474 11454 7476 11506
rect 7420 11442 7476 11454
rect 7084 11394 7252 11396
rect 7084 11342 7086 11394
rect 7138 11342 7252 11394
rect 7084 11340 7252 11342
rect 7084 10498 7140 11340
rect 7084 10446 7086 10498
rect 7138 10446 7140 10498
rect 7084 10434 7140 10446
rect 7532 10500 7588 10510
rect 7308 9828 7364 9838
rect 7532 9828 7588 10444
rect 7308 9826 7588 9828
rect 7308 9774 7310 9826
rect 7362 9774 7588 9826
rect 7308 9772 7588 9774
rect 7308 9762 7364 9772
rect 7196 9268 7252 9278
rect 7196 9174 7252 9212
rect 6972 8428 7364 8484
rect 5740 8306 5796 8316
rect 6972 8260 7028 8270
rect 7196 8260 7252 8270
rect 6972 8258 7252 8260
rect 6972 8206 6974 8258
rect 7026 8206 7198 8258
rect 7250 8206 7252 8258
rect 6972 8204 7252 8206
rect 6972 8194 7028 8204
rect 7196 8194 7252 8204
rect 6860 8148 6916 8158
rect 6860 8054 6916 8092
rect 4172 5796 4228 7644
rect 6188 8036 6244 8046
rect 6188 7586 6244 7980
rect 7308 7924 7364 8428
rect 7420 8260 7476 9772
rect 7532 9604 7588 9772
rect 7532 9538 7588 9548
rect 7532 9156 7588 9166
rect 7644 9156 7700 11900
rect 8764 11508 8820 12572
rect 8876 12402 8932 12684
rect 9324 12738 9380 12750
rect 9772 12740 9828 12750
rect 9324 12686 9326 12738
rect 9378 12686 9380 12738
rect 9324 12628 9380 12686
rect 9324 12562 9380 12572
rect 9660 12684 9772 12740
rect 8876 12350 8878 12402
rect 8930 12350 8932 12402
rect 8876 12338 8932 12350
rect 9548 12178 9604 12190
rect 9548 12126 9550 12178
rect 9602 12126 9604 12178
rect 8988 12068 9044 12078
rect 9548 12068 9604 12126
rect 8988 12066 9604 12068
rect 8988 12014 8990 12066
rect 9042 12014 9604 12066
rect 8988 12012 9604 12014
rect 8988 12002 9044 12012
rect 8876 11508 8932 11518
rect 8764 11506 8932 11508
rect 8764 11454 8878 11506
rect 8930 11454 8932 11506
rect 8764 11452 8932 11454
rect 8876 11442 8932 11452
rect 7980 11396 8036 11406
rect 7980 9938 8036 11340
rect 9212 11284 9268 11294
rect 9212 11190 9268 11228
rect 9548 11284 9604 11294
rect 9660 11284 9716 12684
rect 9772 12646 9828 12684
rect 9884 12738 9940 13468
rect 9996 13188 10052 15092
rect 9996 12962 10052 13132
rect 9996 12910 9998 12962
rect 10050 12910 10052 12962
rect 9996 12898 10052 12910
rect 10108 13076 10164 13086
rect 10108 12962 10164 13020
rect 10108 12910 10110 12962
rect 10162 12910 10164 12962
rect 10108 12898 10164 12910
rect 10220 12852 10276 15092
rect 10444 15092 10500 15262
rect 10668 15314 10724 15326
rect 10668 15262 10670 15314
rect 10722 15262 10724 15314
rect 10444 15026 10500 15036
rect 10556 15202 10612 15214
rect 10556 15150 10558 15202
rect 10610 15150 10612 15202
rect 10332 14644 10388 14654
rect 10332 14306 10388 14588
rect 10332 14254 10334 14306
rect 10386 14254 10388 14306
rect 10332 14242 10388 14254
rect 10556 13860 10612 15150
rect 10668 14532 10724 15262
rect 10892 15316 10948 16156
rect 11004 15540 11060 18172
rect 11116 15652 11172 19180
rect 11676 19124 11732 19134
rect 11676 19030 11732 19068
rect 11340 19012 11396 19022
rect 11340 18918 11396 18956
rect 11452 18788 11508 18798
rect 11452 18674 11508 18732
rect 11452 18622 11454 18674
rect 11506 18622 11508 18674
rect 11452 18610 11508 18622
rect 11340 18564 11396 18574
rect 11228 18562 11396 18564
rect 11228 18510 11342 18562
rect 11394 18510 11396 18562
rect 11228 18508 11396 18510
rect 11228 16324 11284 18508
rect 11340 18498 11396 18508
rect 11228 16258 11284 16268
rect 11676 18450 11732 18462
rect 11676 18398 11678 18450
rect 11730 18398 11732 18450
rect 11340 15988 11396 15998
rect 11340 15986 11620 15988
rect 11340 15934 11342 15986
rect 11394 15934 11620 15986
rect 11340 15932 11620 15934
rect 11340 15922 11396 15932
rect 11116 15596 11508 15652
rect 11004 15484 11284 15540
rect 11004 15316 11060 15326
rect 10892 15314 11060 15316
rect 10892 15262 11006 15314
rect 11058 15262 11060 15314
rect 10892 15260 11060 15262
rect 11004 15250 11060 15260
rect 11116 14756 11172 14766
rect 11116 14662 11172 14700
rect 10668 14466 10724 14476
rect 10892 14418 10948 14430
rect 10892 14366 10894 14418
rect 10946 14366 10948 14418
rect 10892 13972 10948 14366
rect 10892 13906 10948 13916
rect 10556 13794 10612 13804
rect 10332 13748 10388 13758
rect 10332 13654 10388 13692
rect 10556 13524 10612 13534
rect 10444 13522 10612 13524
rect 10444 13470 10558 13522
rect 10610 13470 10612 13522
rect 10444 13468 10612 13470
rect 10444 13186 10500 13468
rect 10556 13458 10612 13468
rect 10444 13134 10446 13186
rect 10498 13134 10500 13186
rect 10444 13122 10500 13134
rect 10668 13412 10724 13422
rect 10220 12786 10276 12796
rect 9884 12686 9886 12738
rect 9938 12686 9940 12738
rect 9884 12674 9940 12686
rect 9772 12516 9828 12526
rect 9772 12178 9828 12460
rect 9772 12126 9774 12178
rect 9826 12126 9828 12178
rect 9772 12114 9828 12126
rect 9996 12404 10052 12414
rect 10556 12404 10612 12414
rect 10668 12404 10724 13356
rect 10052 12402 10724 12404
rect 10052 12350 10558 12402
rect 10610 12350 10724 12402
rect 10052 12348 10724 12350
rect 9996 12178 10052 12348
rect 10556 12338 10612 12348
rect 9996 12126 9998 12178
rect 10050 12126 10052 12178
rect 9996 12114 10052 12126
rect 10108 11954 10164 11966
rect 10108 11902 10110 11954
rect 10162 11902 10164 11954
rect 10108 11396 10164 11902
rect 10108 11330 10164 11340
rect 10780 11394 10836 11406
rect 10780 11342 10782 11394
rect 10834 11342 10836 11394
rect 9548 11282 9716 11284
rect 9548 11230 9550 11282
rect 9602 11230 9716 11282
rect 9548 11228 9716 11230
rect 9548 11218 9604 11228
rect 9884 11172 9940 11182
rect 10220 11172 10276 11182
rect 9884 11170 10276 11172
rect 9884 11118 9886 11170
rect 9938 11118 10222 11170
rect 10274 11118 10276 11170
rect 9884 11116 10276 11118
rect 9884 11106 9940 11116
rect 7980 9886 7982 9938
rect 8034 9886 8036 9938
rect 7980 9874 8036 9886
rect 10108 9938 10164 11116
rect 10220 11106 10276 11116
rect 10780 10724 10836 11342
rect 10780 10658 10836 10668
rect 11116 11284 11172 11294
rect 10108 9886 10110 9938
rect 10162 9886 10164 9938
rect 10108 9874 10164 9886
rect 10780 9828 10836 9838
rect 9660 9604 9716 9614
rect 7532 9154 7812 9156
rect 7532 9102 7534 9154
rect 7586 9102 7812 9154
rect 7532 9100 7812 9102
rect 7532 9090 7588 9100
rect 7644 8260 7700 8270
rect 7420 8204 7588 8260
rect 7420 8036 7476 8046
rect 7420 7942 7476 7980
rect 7308 7858 7364 7868
rect 7420 7700 7476 7710
rect 7532 7700 7588 8204
rect 6188 7534 6190 7586
rect 6242 7534 6244 7586
rect 6188 7522 6244 7534
rect 6972 7698 7588 7700
rect 6972 7646 7422 7698
rect 7474 7646 7588 7698
rect 6972 7644 7588 7646
rect 6972 7474 7028 7644
rect 6972 7422 6974 7474
rect 7026 7422 7028 7474
rect 6972 7410 7028 7422
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 6860 6692 6916 6702
rect 7084 6692 7140 6702
rect 6860 6690 7140 6692
rect 6860 6638 6862 6690
rect 6914 6638 7086 6690
rect 7138 6638 7140 6690
rect 6860 6636 7140 6638
rect 6860 6626 6916 6636
rect 7084 6626 7140 6636
rect 6748 6578 6804 6590
rect 6748 6526 6750 6578
rect 6802 6526 6804 6578
rect 6524 6468 6580 6478
rect 6524 6018 6580 6412
rect 6524 5966 6526 6018
rect 6578 5966 6580 6018
rect 6524 5954 6580 5966
rect 4396 5796 4452 5806
rect 4172 5794 4452 5796
rect 4172 5742 4398 5794
rect 4450 5742 4452 5794
rect 4172 5740 4452 5742
rect 4396 5730 4452 5740
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 6748 4564 6804 6526
rect 7196 6132 7252 7644
rect 7420 7634 7476 7644
rect 7532 6578 7588 6590
rect 7532 6526 7534 6578
rect 7586 6526 7588 6578
rect 7308 6468 7364 6478
rect 7308 6374 7364 6412
rect 7532 6468 7588 6526
rect 7532 6402 7588 6412
rect 7196 5906 7252 6076
rect 7196 5854 7198 5906
rect 7250 5854 7252 5906
rect 7196 5124 7252 5854
rect 7308 5124 7364 5134
rect 7196 5122 7364 5124
rect 7196 5070 7310 5122
rect 7362 5070 7364 5122
rect 7196 5068 7364 5070
rect 7308 5058 7364 5068
rect 6860 5010 6916 5022
rect 6860 4958 6862 5010
rect 6914 4958 6916 5010
rect 6860 4676 6916 4958
rect 7644 5012 7700 8204
rect 7756 8036 7812 9100
rect 9660 9042 9716 9548
rect 10556 9604 10612 9614
rect 10556 9510 10612 9548
rect 9660 8990 9662 9042
rect 9714 8990 9716 9042
rect 9660 8978 9716 8990
rect 10332 8932 10388 8942
rect 9996 8930 10388 8932
rect 9996 8878 10334 8930
rect 10386 8878 10388 8930
rect 9996 8876 10388 8878
rect 9996 8370 10052 8876
rect 10332 8866 10388 8876
rect 9996 8318 9998 8370
rect 10050 8318 10052 8370
rect 9996 8306 10052 8318
rect 7868 8260 7924 8270
rect 8316 8260 8372 8270
rect 7868 8258 8372 8260
rect 7868 8206 7870 8258
rect 7922 8206 8318 8258
rect 8370 8206 8372 8258
rect 7868 8204 8372 8206
rect 7868 8194 7924 8204
rect 8316 8194 8372 8204
rect 9548 8260 9604 8270
rect 9772 8260 9828 8270
rect 9548 8258 9828 8260
rect 9548 8206 9550 8258
rect 9602 8206 9774 8258
rect 9826 8206 9828 8258
rect 9548 8204 9828 8206
rect 9548 8194 9604 8204
rect 9772 8194 9828 8204
rect 10220 8260 10276 8270
rect 10220 8166 10276 8204
rect 9436 8148 9492 8158
rect 8764 8146 9492 8148
rect 8764 8094 9438 8146
rect 9490 8094 9492 8146
rect 8764 8092 9492 8094
rect 8204 8036 8260 8046
rect 7756 8034 8260 8036
rect 7756 7982 8206 8034
rect 8258 7982 8260 8034
rect 7756 7980 8260 7982
rect 8204 7970 8260 7980
rect 8428 8036 8484 8046
rect 8652 8036 8708 8046
rect 8428 7942 8484 7980
rect 8540 8034 8708 8036
rect 8540 7982 8654 8034
rect 8706 7982 8708 8034
rect 8540 7980 8708 7982
rect 8316 7924 8372 7934
rect 8316 7700 8372 7868
rect 8092 7698 8372 7700
rect 8092 7646 8318 7698
rect 8370 7646 8372 7698
rect 8092 7644 8372 7646
rect 7756 6580 7812 6590
rect 7756 6486 7812 6524
rect 7980 6468 8036 6478
rect 7980 6132 8036 6412
rect 8092 6466 8148 7644
rect 8316 7634 8372 7644
rect 8540 6804 8596 7980
rect 8652 7970 8708 7980
rect 8652 7700 8708 7710
rect 8652 7606 8708 7644
rect 8652 6804 8708 6814
rect 8540 6748 8652 6804
rect 8316 6692 8372 6702
rect 8316 6690 8484 6692
rect 8316 6638 8318 6690
rect 8370 6638 8484 6690
rect 8316 6636 8484 6638
rect 8316 6626 8372 6636
rect 8204 6580 8260 6590
rect 8204 6486 8260 6524
rect 8092 6414 8094 6466
rect 8146 6414 8148 6466
rect 8092 6402 8148 6414
rect 8428 6356 8484 6636
rect 8652 6690 8708 6748
rect 8652 6638 8654 6690
rect 8706 6638 8708 6690
rect 8652 6626 8708 6638
rect 8428 6290 8484 6300
rect 8092 6132 8148 6142
rect 7980 6130 8148 6132
rect 7980 6078 8094 6130
rect 8146 6078 8148 6130
rect 7980 6076 8148 6078
rect 8092 6066 8148 6076
rect 8428 6132 8484 6142
rect 8428 6038 8484 6076
rect 8652 5796 8708 5806
rect 7644 4956 8036 5012
rect 6972 4900 7028 4910
rect 7980 4900 8036 4956
rect 6972 4898 7924 4900
rect 6972 4846 6974 4898
rect 7026 4846 7924 4898
rect 6972 4844 7924 4846
rect 6972 4834 7028 4844
rect 6860 4620 7700 4676
rect 6748 4508 7140 4564
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 6860 3556 6916 3566
rect 6412 3444 6468 3482
rect 6860 3462 6916 3500
rect 6412 3378 6468 3388
rect 7084 3442 7140 4508
rect 7308 4228 7364 4238
rect 7308 4226 7588 4228
rect 7308 4174 7310 4226
rect 7362 4174 7588 4226
rect 7308 4172 7588 4174
rect 7308 4162 7364 4172
rect 7084 3390 7086 3442
rect 7138 3390 7140 3442
rect 7084 3378 7140 3390
rect 7308 3444 7364 3454
rect 7420 3444 7476 3482
rect 7364 3442 7476 3444
rect 7364 3390 7422 3442
rect 7474 3390 7476 3442
rect 7364 3388 7476 3390
rect 7308 3378 7364 3388
rect 7420 800 7476 3388
rect 7532 3220 7588 4172
rect 7644 3444 7700 4620
rect 7868 4338 7924 4844
rect 7868 4286 7870 4338
rect 7922 4286 7924 4338
rect 7868 4274 7924 4286
rect 7980 4340 8036 4844
rect 8092 5010 8148 5022
rect 8092 4958 8094 5010
rect 8146 4958 8148 5010
rect 8092 4562 8148 4958
rect 8092 4510 8094 4562
rect 8146 4510 8148 4562
rect 8092 4498 8148 4510
rect 8540 4452 8596 4462
rect 8652 4452 8708 5740
rect 8540 4450 8708 4452
rect 8540 4398 8542 4450
rect 8594 4398 8708 4450
rect 8540 4396 8708 4398
rect 8540 4386 8596 4396
rect 8204 4340 8260 4350
rect 7980 4338 8260 4340
rect 7980 4286 8206 4338
rect 8258 4286 8260 4338
rect 7980 4284 8260 4286
rect 8204 4274 8260 4284
rect 7756 4228 7812 4238
rect 7756 4134 7812 4172
rect 8428 3556 8484 3566
rect 8428 3462 8484 3500
rect 7756 3444 7812 3454
rect 7644 3442 7812 3444
rect 7644 3390 7758 3442
rect 7810 3390 7812 3442
rect 7644 3388 7812 3390
rect 7756 3378 7812 3388
rect 8092 3442 8148 3454
rect 8092 3390 8094 3442
rect 8146 3390 8148 3442
rect 8092 3220 8148 3390
rect 8764 3442 8820 8092
rect 9436 8082 9492 8092
rect 10444 8146 10500 8158
rect 10444 8094 10446 8146
rect 10498 8094 10500 8146
rect 9772 8036 9828 8046
rect 9100 6466 9156 6478
rect 9100 6414 9102 6466
rect 9154 6414 9156 6466
rect 9100 6356 9156 6414
rect 9100 6290 9156 6300
rect 9772 6130 9828 7980
rect 10444 7812 10500 8094
rect 10780 8034 10836 9772
rect 10780 7982 10782 8034
rect 10834 7982 10836 8034
rect 10780 7970 10836 7982
rect 10892 8034 10948 8046
rect 10892 7982 10894 8034
rect 10946 7982 10948 8034
rect 10892 7812 10948 7982
rect 11004 8036 11060 8046
rect 11004 7942 11060 7980
rect 10444 7756 10948 7812
rect 10668 7586 10724 7598
rect 10668 7534 10670 7586
rect 10722 7534 10724 7586
rect 10332 7476 10388 7486
rect 10220 7474 10388 7476
rect 10220 7422 10334 7474
rect 10386 7422 10388 7474
rect 10220 7420 10388 7422
rect 10108 6804 10164 6814
rect 9884 6690 9940 6702
rect 9884 6638 9886 6690
rect 9938 6638 9940 6690
rect 9884 6356 9940 6638
rect 9996 6356 10052 6366
rect 9884 6300 9996 6356
rect 9996 6290 10052 6300
rect 9772 6078 9774 6130
rect 9826 6078 9828 6130
rect 9772 6066 9828 6078
rect 9548 6020 9604 6030
rect 9548 5926 9604 5964
rect 10108 5906 10164 6748
rect 10108 5854 10110 5906
rect 10162 5854 10164 5906
rect 10108 5842 10164 5854
rect 9660 5796 9716 5806
rect 9660 5702 9716 5740
rect 10220 5012 10276 7420
rect 10332 7410 10388 7420
rect 10444 6692 10500 6702
rect 10668 6692 10724 7534
rect 10892 6916 10948 6926
rect 10892 6692 10948 6860
rect 11116 6692 11172 11228
rect 11228 7700 11284 15484
rect 11452 15538 11508 15596
rect 11452 15486 11454 15538
rect 11506 15486 11508 15538
rect 11452 15092 11508 15486
rect 11564 15538 11620 15932
rect 11564 15486 11566 15538
rect 11618 15486 11620 15538
rect 11564 15474 11620 15486
rect 11676 15540 11732 18398
rect 11788 17778 11844 19964
rect 12124 19926 12180 19964
rect 12124 19348 12180 19358
rect 12124 19254 12180 19292
rect 12236 19236 12292 19246
rect 12236 19142 12292 19180
rect 11788 17726 11790 17778
rect 11842 17726 11844 17778
rect 11788 17444 11844 17726
rect 11788 17378 11844 17388
rect 11900 19122 11956 19134
rect 11900 19070 11902 19122
rect 11954 19070 11956 19122
rect 11900 18452 11956 19070
rect 11788 16660 11844 16670
rect 11788 16098 11844 16604
rect 11788 16046 11790 16098
rect 11842 16046 11844 16098
rect 11788 16034 11844 16046
rect 11676 15474 11732 15484
rect 11676 15316 11732 15326
rect 11676 15222 11732 15260
rect 11340 14530 11396 14542
rect 11340 14478 11342 14530
rect 11394 14478 11396 14530
rect 11340 13860 11396 14478
rect 11452 14420 11508 15036
rect 11564 14756 11620 14766
rect 11564 14662 11620 14700
rect 11452 14354 11508 14364
rect 11340 13794 11396 13804
rect 11900 13748 11956 18396
rect 13020 17780 13076 23212
rect 13132 21812 13188 21822
rect 13132 21476 13188 21756
rect 13132 21382 13188 21420
rect 13356 18452 13412 18462
rect 13468 18452 13524 25564
rect 13580 23716 13636 25788
rect 13580 23650 13636 23660
rect 13580 23044 13636 23054
rect 13580 22950 13636 22988
rect 13580 22484 13636 22494
rect 13580 22258 13636 22428
rect 13580 22206 13582 22258
rect 13634 22206 13636 22258
rect 13580 22194 13636 22206
rect 13580 18564 13636 18574
rect 13692 18564 13748 26684
rect 13804 25956 13860 27022
rect 13804 25890 13860 25900
rect 13916 25844 13972 29260
rect 14028 28084 14084 30046
rect 14028 27990 14084 28028
rect 14252 27074 14308 30268
rect 14364 29988 14420 30604
rect 14924 30322 14980 31612
rect 15036 31106 15092 31724
rect 15036 31054 15038 31106
rect 15090 31054 15092 31106
rect 15036 30434 15092 31054
rect 15036 30382 15038 30434
rect 15090 30382 15092 30434
rect 15036 30370 15092 30382
rect 14924 30270 14926 30322
rect 14978 30270 14980 30322
rect 14700 30212 14756 30222
rect 14588 30210 14756 30212
rect 14588 30158 14702 30210
rect 14754 30158 14756 30210
rect 14588 30156 14756 30158
rect 14364 29932 14532 29988
rect 14364 29314 14420 29326
rect 14364 29262 14366 29314
rect 14418 29262 14420 29314
rect 14364 28532 14420 29262
rect 14364 28466 14420 28476
rect 14252 27022 14254 27074
rect 14306 27022 14308 27074
rect 14252 27010 14308 27022
rect 14476 26908 14532 29932
rect 14588 28868 14644 30156
rect 14700 30146 14756 30156
rect 14924 29876 14980 30270
rect 14924 29810 14980 29820
rect 14812 29652 14868 29662
rect 14812 29650 14980 29652
rect 14812 29598 14814 29650
rect 14866 29598 14980 29650
rect 14812 29596 14980 29598
rect 14812 29586 14868 29596
rect 14588 28802 14644 28812
rect 14700 29204 14756 29214
rect 13916 25778 13972 25788
rect 14252 26852 14532 26908
rect 14140 25284 14196 25294
rect 14028 24610 14084 24622
rect 14028 24558 14030 24610
rect 14082 24558 14084 24610
rect 14028 24500 14084 24558
rect 14028 24434 14084 24444
rect 13916 23154 13972 23166
rect 13916 23102 13918 23154
rect 13970 23102 13972 23154
rect 13916 23044 13972 23102
rect 13916 22978 13972 22988
rect 14028 22372 14084 22382
rect 14140 22372 14196 25228
rect 14028 22370 14196 22372
rect 14028 22318 14030 22370
rect 14082 22318 14196 22370
rect 14028 22316 14196 22318
rect 14028 22306 14084 22316
rect 13916 22260 13972 22270
rect 13916 22166 13972 22204
rect 13804 22146 13860 22158
rect 13804 22094 13806 22146
rect 13858 22094 13860 22146
rect 13804 21476 13860 22094
rect 13804 21410 13860 21420
rect 14252 20916 14308 26852
rect 14700 25508 14756 29148
rect 14924 28868 14980 29596
rect 14924 28774 14980 28812
rect 15036 29204 15092 29214
rect 15036 28642 15092 29148
rect 15036 28590 15038 28642
rect 15090 28590 15092 28642
rect 15036 28578 15092 28590
rect 15148 28420 15204 33964
rect 15596 32676 15652 34638
rect 16156 34132 16212 35308
rect 16828 35026 16884 36316
rect 17500 35588 17556 35598
rect 17500 35494 17556 35532
rect 16828 34974 16830 35026
rect 16882 34974 16884 35026
rect 16828 34962 16884 34974
rect 16268 34132 16324 34142
rect 16156 34130 16324 34132
rect 16156 34078 16270 34130
rect 16322 34078 16324 34130
rect 16156 34076 16324 34078
rect 16044 32788 16100 32798
rect 15596 32610 15652 32620
rect 15932 32674 15988 32686
rect 15932 32622 15934 32674
rect 15986 32622 15988 32674
rect 15820 32340 15876 32350
rect 15260 32338 15876 32340
rect 15260 32286 15822 32338
rect 15874 32286 15876 32338
rect 15260 32284 15876 32286
rect 15260 31218 15316 32284
rect 15820 32274 15876 32284
rect 15372 31556 15428 31566
rect 15372 31462 15428 31500
rect 15708 31332 15764 31342
rect 15596 31276 15708 31332
rect 15260 31166 15262 31218
rect 15314 31166 15316 31218
rect 15260 31154 15316 31166
rect 15372 31220 15428 31230
rect 15372 31126 15428 31164
rect 15596 31218 15652 31276
rect 15708 31266 15764 31276
rect 15596 31166 15598 31218
rect 15650 31166 15652 31218
rect 15596 31154 15652 31166
rect 15484 31108 15540 31118
rect 15484 31014 15540 31052
rect 15932 31108 15988 32622
rect 15932 31042 15988 31052
rect 16044 30884 16100 32732
rect 16156 32338 16212 32350
rect 16156 32286 16158 32338
rect 16210 32286 16212 32338
rect 16156 31780 16212 32286
rect 16156 31714 16212 31724
rect 15932 30828 16100 30884
rect 16156 30882 16212 30894
rect 16156 30830 16158 30882
rect 16210 30830 16212 30882
rect 15596 30212 15652 30222
rect 15260 30100 15316 30110
rect 15260 29426 15316 30044
rect 15596 29650 15652 30156
rect 15932 30210 15988 30828
rect 16156 30772 16212 30830
rect 15932 30158 15934 30210
rect 15986 30158 15988 30210
rect 15932 30100 15988 30158
rect 15932 30034 15988 30044
rect 16044 30322 16100 30334
rect 16044 30270 16046 30322
rect 16098 30270 16100 30322
rect 16044 29652 16100 30270
rect 16156 30212 16212 30716
rect 16156 30146 16212 30156
rect 16268 29876 16324 34076
rect 17164 33460 17220 33470
rect 17164 33366 17220 33404
rect 17612 32788 17668 38612
rect 18172 37492 18228 37502
rect 18508 37492 18564 38612
rect 17836 37380 17892 37390
rect 17836 37286 17892 37324
rect 18172 37378 18228 37436
rect 18172 37326 18174 37378
rect 18226 37326 18228 37378
rect 18172 37314 18228 37326
rect 18284 37490 18564 37492
rect 18284 37438 18510 37490
rect 18562 37438 18564 37490
rect 18284 37436 18564 37438
rect 17724 36594 17780 36606
rect 17724 36542 17726 36594
rect 17778 36542 17780 36594
rect 17724 36260 17780 36542
rect 18172 36596 18228 36606
rect 18172 36502 18228 36540
rect 18284 36482 18340 37436
rect 18508 37426 18564 37436
rect 18284 36430 18286 36482
rect 18338 36430 18340 36482
rect 18284 36418 18340 36430
rect 18060 36260 18116 36270
rect 17724 36258 18116 36260
rect 17724 36206 18062 36258
rect 18114 36206 18116 36258
rect 17724 36204 18116 36206
rect 17948 35586 18004 35598
rect 17948 35534 17950 35586
rect 18002 35534 18004 35586
rect 17948 35364 18004 35534
rect 17948 35298 18004 35308
rect 18060 33796 18116 36204
rect 18508 36258 18564 36270
rect 18508 36206 18510 36258
rect 18562 36206 18564 36258
rect 18396 35698 18452 35710
rect 18396 35646 18398 35698
rect 18450 35646 18452 35698
rect 18060 33730 18116 33740
rect 18284 34692 18340 34702
rect 18284 34130 18340 34636
rect 18284 34078 18286 34130
rect 18338 34078 18340 34130
rect 17612 32722 17668 32732
rect 17948 33346 18004 33358
rect 17948 33294 17950 33346
rect 18002 33294 18004 33346
rect 16604 32676 16660 32686
rect 16604 32582 16660 32620
rect 17388 32676 17444 32686
rect 16492 32564 16548 32574
rect 16492 30996 16548 32508
rect 16716 32562 16772 32574
rect 16716 32510 16718 32562
rect 16770 32510 16772 32562
rect 16604 32338 16660 32350
rect 16604 32286 16606 32338
rect 16658 32286 16660 32338
rect 16604 31332 16660 32286
rect 16604 31266 16660 31276
rect 16604 30996 16660 31006
rect 16492 30994 16660 30996
rect 16492 30942 16606 30994
rect 16658 30942 16660 30994
rect 16492 30940 16660 30942
rect 16716 30996 16772 32510
rect 16716 30940 17108 30996
rect 16604 30930 16660 30940
rect 16268 29810 16324 29820
rect 16716 30770 16772 30782
rect 16716 30718 16718 30770
rect 16770 30718 16772 30770
rect 15596 29598 15598 29650
rect 15650 29598 15652 29650
rect 15596 29586 15652 29598
rect 15820 29596 16044 29652
rect 15260 29374 15262 29426
rect 15314 29374 15316 29426
rect 15260 29204 15316 29374
rect 15260 29138 15316 29148
rect 15372 29426 15428 29438
rect 15372 29374 15374 29426
rect 15426 29374 15428 29426
rect 15372 28644 15428 29374
rect 15820 29426 15876 29596
rect 16044 29586 16100 29596
rect 16156 29540 16212 29550
rect 16156 29446 16212 29484
rect 15820 29374 15822 29426
rect 15874 29374 15876 29426
rect 15820 29362 15876 29374
rect 16492 29426 16548 29438
rect 16492 29374 16494 29426
rect 16546 29374 16548 29426
rect 15372 28578 15428 28588
rect 15484 29314 15540 29326
rect 15484 29262 15486 29314
rect 15538 29262 15540 29314
rect 15036 28364 15204 28420
rect 15260 28532 15316 28542
rect 14812 27076 14868 27086
rect 14812 26982 14868 27020
rect 14476 25452 14756 25508
rect 14924 25508 14980 25518
rect 14364 24722 14420 24734
rect 14364 24670 14366 24722
rect 14418 24670 14420 24722
rect 14364 24500 14420 24670
rect 14364 24434 14420 24444
rect 14476 22484 14532 25452
rect 14700 25284 14756 25294
rect 14924 25284 14980 25452
rect 14756 25228 14980 25284
rect 14700 24946 14756 25228
rect 14700 24894 14702 24946
rect 14754 24894 14756 24946
rect 14700 24882 14756 24894
rect 15036 24722 15092 28364
rect 15260 27860 15316 28476
rect 15372 27860 15428 27870
rect 15260 27858 15428 27860
rect 15260 27806 15374 27858
rect 15426 27806 15428 27858
rect 15260 27804 15428 27806
rect 15372 27636 15428 27804
rect 15372 27570 15428 27580
rect 15372 26964 15428 27002
rect 15372 26898 15428 26908
rect 15148 26852 15204 26862
rect 15148 26850 15316 26852
rect 15148 26798 15150 26850
rect 15202 26798 15316 26850
rect 15148 26796 15316 26798
rect 15148 26786 15204 26796
rect 15260 26290 15316 26796
rect 15484 26402 15540 29262
rect 16492 29204 16548 29374
rect 16492 29138 16548 29148
rect 16380 28756 16436 28766
rect 16716 28756 16772 30718
rect 16940 30212 16996 30222
rect 16380 28754 16772 28756
rect 16380 28702 16382 28754
rect 16434 28702 16772 28754
rect 16380 28700 16772 28702
rect 16828 30100 16884 30110
rect 16044 28308 16100 28318
rect 15596 28084 15652 28094
rect 15596 27858 15652 28028
rect 16044 28082 16100 28252
rect 16380 28196 16436 28700
rect 16828 28642 16884 30044
rect 16940 29540 16996 30156
rect 17052 29988 17108 30940
rect 17276 29988 17332 29998
rect 17052 29986 17332 29988
rect 17052 29934 17278 29986
rect 17330 29934 17332 29986
rect 17052 29932 17332 29934
rect 17388 29988 17444 32620
rect 17612 32564 17668 32574
rect 17612 32470 17668 32508
rect 17948 32564 18004 33294
rect 18284 33124 18340 34078
rect 18396 34020 18452 35646
rect 18508 34916 18564 36206
rect 18732 35252 18788 38612
rect 18844 37492 18900 37502
rect 18844 37398 18900 37436
rect 18732 35186 18788 35196
rect 18956 37380 19012 37390
rect 18508 34850 18564 34860
rect 18844 34914 18900 34926
rect 18844 34862 18846 34914
rect 18898 34862 18900 34914
rect 18844 34692 18900 34862
rect 18844 34626 18900 34636
rect 18844 34020 18900 34030
rect 18396 34018 18900 34020
rect 18396 33966 18846 34018
rect 18898 33966 18900 34018
rect 18396 33964 18900 33966
rect 18508 33796 18564 33806
rect 18284 33058 18340 33068
rect 18396 33122 18452 33134
rect 18396 33070 18398 33122
rect 18450 33070 18452 33122
rect 17948 32498 18004 32508
rect 18172 32452 18228 32462
rect 18396 32452 18452 33070
rect 18228 32396 18452 32452
rect 18172 32358 18228 32396
rect 18172 31780 18228 31790
rect 18060 31666 18116 31678
rect 18060 31614 18062 31666
rect 18114 31614 18116 31666
rect 18060 31108 18116 31614
rect 17612 30994 17668 31006
rect 17612 30942 17614 30994
rect 17666 30942 17668 30994
rect 17612 30324 17668 30942
rect 18060 30770 18116 31052
rect 18060 30718 18062 30770
rect 18114 30718 18116 30770
rect 18060 30706 18116 30718
rect 17612 30210 17668 30268
rect 17612 30158 17614 30210
rect 17666 30158 17668 30210
rect 17612 30146 17668 30158
rect 18060 30324 18116 30334
rect 18060 30210 18116 30268
rect 18060 30158 18062 30210
rect 18114 30158 18116 30210
rect 18060 30146 18116 30158
rect 17948 30100 18004 30110
rect 17948 30006 18004 30044
rect 17388 29932 17668 29988
rect 16940 29474 16996 29484
rect 16828 28590 16830 28642
rect 16882 28590 16884 28642
rect 16380 28130 16436 28140
rect 16604 28308 16660 28318
rect 16044 28030 16046 28082
rect 16098 28030 16100 28082
rect 16044 28018 16100 28030
rect 15820 27972 15876 27982
rect 15820 27878 15876 27916
rect 16268 27972 16324 27982
rect 15596 27806 15598 27858
rect 15650 27806 15652 27858
rect 15596 27794 15652 27806
rect 15932 27748 15988 27758
rect 15932 27654 15988 27692
rect 15820 27636 15876 27646
rect 15820 27074 15876 27580
rect 15820 27022 15822 27074
rect 15874 27022 15876 27074
rect 15820 27010 15876 27022
rect 16268 27074 16324 27916
rect 16604 27076 16660 28252
rect 16268 27022 16270 27074
rect 16322 27022 16324 27074
rect 16268 27010 16324 27022
rect 16492 27020 16660 27076
rect 16492 26962 16548 27020
rect 16492 26910 16494 26962
rect 16546 26910 16548 26962
rect 16492 26898 16548 26910
rect 16604 26850 16660 26862
rect 16604 26798 16606 26850
rect 16658 26798 16660 26850
rect 16604 26404 16660 26798
rect 15484 26350 15486 26402
rect 15538 26350 15540 26402
rect 15484 26338 15540 26350
rect 15932 26348 16660 26404
rect 15260 26238 15262 26290
rect 15314 26238 15316 26290
rect 15260 26226 15316 26238
rect 15932 26290 15988 26348
rect 15932 26238 15934 26290
rect 15986 26238 15988 26290
rect 15932 26226 15988 26238
rect 15372 26068 15428 26078
rect 15260 25956 15316 25966
rect 15260 25730 15316 25900
rect 15260 25678 15262 25730
rect 15314 25678 15316 25730
rect 15260 25666 15316 25678
rect 15148 25284 15204 25294
rect 15148 25190 15204 25228
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 15036 24658 15092 24670
rect 14924 23716 14980 23726
rect 14980 23660 15092 23716
rect 14924 23650 14980 23660
rect 14476 22390 14532 22428
rect 14700 23042 14756 23054
rect 14700 22990 14702 23042
rect 14754 22990 14756 23042
rect 14700 21252 14756 22990
rect 14924 21474 14980 21486
rect 14924 21422 14926 21474
rect 14978 21422 14980 21474
rect 14812 21364 14868 21374
rect 14812 21270 14868 21308
rect 14476 21196 14756 21252
rect 14364 21028 14420 21038
rect 14364 20934 14420 20972
rect 14140 20860 14308 20916
rect 14028 19348 14084 19358
rect 13804 19236 13860 19246
rect 13804 19142 13860 19180
rect 13916 19236 13972 19246
rect 14028 19236 14084 19292
rect 13916 19234 14084 19236
rect 13916 19182 13918 19234
rect 13970 19182 14084 19234
rect 13916 19180 14084 19182
rect 13916 19170 13972 19180
rect 13580 18562 13748 18564
rect 13580 18510 13582 18562
rect 13634 18510 13748 18562
rect 13580 18508 13748 18510
rect 13580 18498 13636 18508
rect 13356 18450 13468 18452
rect 13356 18398 13358 18450
rect 13410 18398 13468 18450
rect 13356 18396 13468 18398
rect 14140 18452 14196 20860
rect 14252 20692 14308 20702
rect 14252 20598 14308 20636
rect 14140 18396 14308 18452
rect 13356 18386 13412 18396
rect 13468 18358 13524 18396
rect 13692 18338 13748 18350
rect 13692 18286 13694 18338
rect 13746 18286 13748 18338
rect 13692 17892 13748 18286
rect 13692 17826 13748 17836
rect 13916 18226 13972 18238
rect 13916 18174 13918 18226
rect 13970 18174 13972 18226
rect 13020 17714 13076 17724
rect 13580 17668 13636 17678
rect 13580 16882 13636 17612
rect 13580 16830 13582 16882
rect 13634 16830 13636 16882
rect 13580 16818 13636 16830
rect 12572 16770 12628 16782
rect 12572 16718 12574 16770
rect 12626 16718 12628 16770
rect 12236 16100 12292 16110
rect 12236 16006 12292 16044
rect 12236 15314 12292 15326
rect 12236 15262 12238 15314
rect 12290 15262 12292 15314
rect 12236 15148 12292 15262
rect 12124 15092 12292 15148
rect 12460 15314 12516 15326
rect 12460 15262 12462 15314
rect 12514 15262 12516 15314
rect 12012 14868 12068 14878
rect 12012 14754 12068 14812
rect 12012 14702 12014 14754
rect 12066 14702 12068 14754
rect 12012 14690 12068 14702
rect 12012 13748 12068 13758
rect 11900 13746 12068 13748
rect 11900 13694 12014 13746
rect 12066 13694 12068 13746
rect 11900 13692 12068 13694
rect 11676 13076 11732 13086
rect 11676 11506 11732 13020
rect 11676 11454 11678 11506
rect 11730 11454 11732 11506
rect 11676 11442 11732 11454
rect 11788 11844 11844 11854
rect 11788 11394 11844 11788
rect 11788 11342 11790 11394
rect 11842 11342 11844 11394
rect 11788 11330 11844 11342
rect 11340 11172 11396 11182
rect 11340 11078 11396 11116
rect 11564 11170 11620 11182
rect 11564 11118 11566 11170
rect 11618 11118 11620 11170
rect 11564 9826 11620 11118
rect 11788 11172 11844 11182
rect 11788 10834 11844 11116
rect 11788 10782 11790 10834
rect 11842 10782 11844 10834
rect 11788 10770 11844 10782
rect 11900 10724 11956 10734
rect 11900 10630 11956 10668
rect 11564 9774 11566 9826
rect 11618 9774 11620 9826
rect 11564 9716 11620 9774
rect 11900 9940 11956 9950
rect 12012 9940 12068 13692
rect 12124 13076 12180 15092
rect 12348 15090 12404 15102
rect 12348 15038 12350 15090
rect 12402 15038 12404 15090
rect 12348 14756 12404 15038
rect 12348 14690 12404 14700
rect 12348 14308 12404 14318
rect 12460 14308 12516 15262
rect 12572 15148 12628 16718
rect 13468 16772 13524 16782
rect 13468 16322 13524 16716
rect 13468 16270 13470 16322
rect 13522 16270 13524 16322
rect 13468 16258 13524 16270
rect 13804 16212 13860 16222
rect 13804 16118 13860 16156
rect 12796 16100 12852 16110
rect 12796 15874 12852 16044
rect 12908 15988 12964 15992
rect 13020 15988 13076 15998
rect 12908 15980 13020 15988
rect 12908 15928 12910 15980
rect 12962 15932 13020 15980
rect 12962 15928 12964 15932
rect 12908 15916 12964 15928
rect 13020 15922 13076 15932
rect 13580 15988 13636 15998
rect 12796 15822 12798 15874
rect 12850 15822 12852 15874
rect 12796 15810 12852 15822
rect 13468 15876 13524 15886
rect 12684 15540 12740 15550
rect 12684 15446 12740 15484
rect 12908 15314 12964 15326
rect 12908 15262 12910 15314
rect 12962 15262 12964 15314
rect 12908 15148 12964 15262
rect 12572 15092 12852 15148
rect 12908 15092 13076 15148
rect 12572 14420 12628 14430
rect 12572 14326 12628 14364
rect 12684 14418 12740 14430
rect 12684 14366 12686 14418
rect 12738 14366 12740 14418
rect 12348 14306 12516 14308
rect 12348 14254 12350 14306
rect 12402 14254 12516 14306
rect 12348 14252 12516 14254
rect 12684 14308 12740 14366
rect 12236 13858 12292 13870
rect 12236 13806 12238 13858
rect 12290 13806 12292 13858
rect 12236 13188 12292 13806
rect 12348 13748 12404 14252
rect 12684 14242 12740 14252
rect 12348 13682 12404 13692
rect 12684 13188 12740 13198
rect 12236 13122 12292 13132
rect 12572 13132 12684 13188
rect 12124 13010 12180 13020
rect 12572 11844 12628 13132
rect 12684 13122 12740 13132
rect 12684 12852 12740 12862
rect 12684 12290 12740 12796
rect 12684 12238 12686 12290
rect 12738 12238 12740 12290
rect 12684 12226 12740 12238
rect 11900 9938 12068 9940
rect 11900 9886 11902 9938
rect 11954 9886 12068 9938
rect 11900 9884 12068 9886
rect 12236 11394 12292 11406
rect 12236 11342 12238 11394
rect 12290 11342 12292 11394
rect 11900 9828 11956 9884
rect 11900 9762 11956 9772
rect 12124 9828 12180 9838
rect 12236 9828 12292 11342
rect 12572 11396 12628 11788
rect 12684 11396 12740 11406
rect 12572 11394 12740 11396
rect 12572 11342 12686 11394
rect 12738 11342 12740 11394
rect 12572 11340 12740 11342
rect 12684 11330 12740 11340
rect 12460 11284 12516 11294
rect 12460 11190 12516 11228
rect 12348 11172 12404 11182
rect 12348 11078 12404 11116
rect 12572 11170 12628 11182
rect 12572 11118 12574 11170
rect 12626 11118 12628 11170
rect 12572 11060 12628 11118
rect 12572 10994 12628 11004
rect 12572 10498 12628 10510
rect 12572 10446 12574 10498
rect 12626 10446 12628 10498
rect 12348 9828 12404 9838
rect 12236 9826 12404 9828
rect 12236 9774 12350 9826
rect 12402 9774 12404 9826
rect 12236 9772 12404 9774
rect 11564 9650 11620 9660
rect 11452 8258 11508 8270
rect 11452 8206 11454 8258
rect 11506 8206 11508 8258
rect 11284 7644 11396 7700
rect 11228 7634 11284 7644
rect 10444 6690 10948 6692
rect 10444 6638 10446 6690
rect 10498 6638 10894 6690
rect 10946 6638 10948 6690
rect 10444 6636 10948 6638
rect 10444 6626 10500 6636
rect 10892 6626 10948 6636
rect 11004 6636 11172 6692
rect 11228 6916 11284 6926
rect 10668 6132 10724 6142
rect 10668 6038 10724 6076
rect 10332 6020 10388 6030
rect 10332 5234 10388 5964
rect 11004 6020 11060 6636
rect 11116 6468 11172 6478
rect 11116 6374 11172 6412
rect 11228 6244 11284 6860
rect 11340 6468 11396 7644
rect 11452 6804 11508 8206
rect 11452 6578 11508 6748
rect 11788 8036 11844 8046
rect 11788 6692 11844 7980
rect 11900 7700 11956 7710
rect 11900 7606 11956 7644
rect 11788 6636 11956 6692
rect 11452 6526 11454 6578
rect 11506 6526 11508 6578
rect 11452 6514 11508 6526
rect 11340 6402 11396 6412
rect 11788 6468 11844 6478
rect 11788 6374 11844 6412
rect 11004 5906 11060 5964
rect 11004 5854 11006 5906
rect 11058 5854 11060 5906
rect 11004 5842 11060 5854
rect 11116 6188 11284 6244
rect 11004 5684 11060 5694
rect 10332 5182 10334 5234
rect 10386 5182 10388 5234
rect 10332 5170 10388 5182
rect 10892 5628 11004 5684
rect 10220 4564 10276 4956
rect 10780 4900 10836 4910
rect 10780 4806 10836 4844
rect 10332 4564 10388 4574
rect 10220 4562 10388 4564
rect 10220 4510 10334 4562
rect 10386 4510 10388 4562
rect 10220 4508 10388 4510
rect 10332 4498 10388 4508
rect 9100 4452 9156 4462
rect 9100 4358 9156 4396
rect 9996 4452 10052 4462
rect 9660 4340 9716 4350
rect 9660 4246 9716 4284
rect 8764 3390 8766 3442
rect 8818 3390 8820 3442
rect 8764 3378 8820 3390
rect 9324 4228 9380 4238
rect 9324 3554 9380 4172
rect 9548 4226 9604 4238
rect 9548 4174 9550 4226
rect 9602 4174 9604 4226
rect 9324 3502 9326 3554
rect 9378 3502 9380 3554
rect 9324 3444 9380 3502
rect 9324 3378 9380 3388
rect 9436 3556 9492 3566
rect 7532 3164 8148 3220
rect 8092 800 8148 3164
rect 9436 800 9492 3500
rect 9548 3444 9604 4174
rect 9660 3444 9716 3454
rect 9548 3442 9716 3444
rect 9548 3390 9662 3442
rect 9714 3390 9716 3442
rect 9548 3388 9716 3390
rect 9660 3378 9716 3388
rect 9996 3388 10052 4396
rect 10556 4340 10612 4350
rect 10556 4246 10612 4284
rect 10780 4228 10836 4238
rect 10780 4134 10836 4172
rect 10892 3388 10948 5628
rect 11004 5618 11060 5628
rect 11116 5122 11172 6188
rect 11564 6132 11620 6142
rect 11116 5070 11118 5122
rect 11170 5070 11172 5122
rect 11116 5058 11172 5070
rect 11228 5124 11284 5134
rect 11004 4900 11060 4910
rect 11004 4450 11060 4844
rect 11004 4398 11006 4450
rect 11058 4398 11060 4450
rect 11004 4386 11060 4398
rect 11228 4450 11284 5068
rect 11452 5122 11508 5134
rect 11452 5070 11454 5122
rect 11506 5070 11508 5122
rect 11340 5012 11396 5022
rect 11452 5012 11508 5070
rect 11396 4956 11508 5012
rect 11340 4946 11396 4956
rect 11228 4398 11230 4450
rect 11282 4398 11284 4450
rect 11228 4386 11284 4398
rect 11564 4338 11620 6076
rect 11788 5012 11844 5022
rect 11900 5012 11956 6636
rect 12012 5684 12068 5694
rect 12012 5590 12068 5628
rect 11788 5010 11900 5012
rect 11788 4958 11790 5010
rect 11842 4958 11900 5010
rect 11788 4956 11900 4958
rect 11788 4946 11844 4956
rect 11900 4918 11956 4956
rect 11564 4286 11566 4338
rect 11618 4286 11620 4338
rect 11564 4274 11620 4286
rect 11564 3666 11620 3678
rect 11564 3614 11566 3666
rect 11618 3614 11620 3666
rect 11452 3444 11508 3454
rect 9996 3332 10164 3388
rect 10892 3332 11060 3388
rect 10108 800 10164 3332
rect 11004 2884 11060 3332
rect 10780 2828 11060 2884
rect 10780 800 10836 2828
rect 11452 800 11508 3388
rect 11564 3388 11620 3614
rect 12124 3554 12180 9772
rect 12348 8932 12404 9772
rect 12572 9828 12628 10446
rect 12572 9762 12628 9772
rect 12796 9604 12852 15092
rect 13020 14308 13076 15092
rect 13468 14756 13524 15820
rect 12908 13860 12964 13870
rect 12908 13766 12964 13804
rect 13020 13746 13076 14252
rect 13020 13694 13022 13746
rect 13074 13694 13076 13746
rect 13020 13682 13076 13694
rect 13244 14700 13524 14756
rect 13580 15876 13636 15932
rect 13804 15988 13860 15998
rect 13692 15876 13748 15886
rect 13580 15874 13748 15876
rect 13580 15822 13694 15874
rect 13746 15822 13748 15874
rect 13580 15820 13748 15822
rect 13244 13412 13300 14700
rect 13468 14530 13524 14542
rect 13468 14478 13470 14530
rect 13522 14478 13524 14530
rect 13468 13412 13524 14478
rect 13580 13972 13636 15820
rect 13692 15810 13748 15820
rect 13692 15314 13748 15326
rect 13692 15262 13694 15314
rect 13746 15262 13748 15314
rect 13692 14418 13748 15262
rect 13804 15316 13860 15932
rect 13804 15222 13860 15260
rect 13916 15148 13972 18174
rect 14140 18228 14196 18238
rect 14140 18134 14196 18172
rect 14028 17668 14084 17678
rect 14028 17574 14084 17612
rect 14140 16772 14196 16782
rect 14028 16716 14140 16772
rect 14252 16772 14308 18396
rect 14364 16996 14420 17006
rect 14476 16996 14532 21196
rect 14924 21140 14980 21422
rect 14588 21084 14980 21140
rect 14588 21026 14644 21084
rect 14588 20974 14590 21026
rect 14642 20974 14644 21026
rect 14588 20962 14644 20974
rect 14700 20916 14756 20926
rect 14700 20822 14756 20860
rect 15036 20244 15092 23660
rect 14588 20188 15092 20244
rect 15148 21586 15204 21598
rect 15372 21588 15428 26012
rect 15484 26066 15540 26078
rect 15484 26014 15486 26066
rect 15538 26014 15540 26066
rect 15484 24722 15540 26014
rect 16156 25956 16212 25966
rect 16044 25900 16156 25956
rect 15932 25844 15988 25854
rect 15708 25508 15764 25518
rect 15708 25414 15764 25452
rect 15484 24670 15486 24722
rect 15538 24670 15540 24722
rect 15484 24658 15540 24670
rect 15148 21534 15150 21586
rect 15202 21534 15204 21586
rect 15148 20804 15204 21534
rect 14588 19012 14644 20188
rect 14700 19964 15092 20020
rect 14700 19348 14756 19964
rect 15036 19906 15092 19964
rect 15036 19854 15038 19906
rect 15090 19854 15092 19906
rect 15036 19842 15092 19854
rect 14700 19234 14756 19292
rect 15148 19348 15204 20748
rect 15148 19254 15204 19292
rect 15260 21532 15428 21588
rect 15484 24498 15540 24510
rect 15484 24446 15486 24498
rect 15538 24446 15540 24498
rect 14700 19182 14702 19234
rect 14754 19182 14756 19234
rect 14700 19170 14756 19182
rect 14588 18956 15092 19012
rect 14700 18452 14756 18462
rect 14756 18396 14868 18452
rect 14700 18358 14756 18396
rect 14700 17444 14756 17454
rect 14364 16994 14532 16996
rect 14364 16942 14366 16994
rect 14418 16942 14532 16994
rect 14364 16940 14532 16942
rect 14588 17442 14756 17444
rect 14588 17390 14702 17442
rect 14754 17390 14756 17442
rect 14588 17388 14756 17390
rect 14364 16930 14420 16940
rect 14252 16716 14420 16772
rect 14028 15988 14084 16716
rect 14140 16706 14196 16716
rect 14252 15988 14308 15998
rect 14028 15922 14084 15932
rect 14140 15932 14252 15988
rect 14140 15426 14196 15932
rect 14252 15894 14308 15932
rect 14140 15374 14142 15426
rect 14194 15374 14196 15426
rect 14140 15362 14196 15374
rect 14252 15314 14308 15326
rect 14252 15262 14254 15314
rect 14306 15262 14308 15314
rect 13916 15092 14196 15148
rect 13692 14366 13694 14418
rect 13746 14366 13748 14418
rect 13692 14084 13748 14366
rect 13804 14308 13860 14318
rect 13804 14214 13860 14252
rect 13692 14028 14084 14084
rect 13580 13916 13748 13972
rect 13580 13746 13636 13758
rect 13580 13694 13582 13746
rect 13634 13694 13636 13746
rect 13580 13524 13636 13694
rect 13580 13458 13636 13468
rect 13244 13346 13300 13356
rect 13356 13356 13524 13412
rect 13356 12852 13412 13356
rect 13580 13300 13636 13310
rect 13468 13188 13524 13198
rect 13468 13094 13524 13132
rect 13580 12962 13636 13244
rect 13580 12910 13582 12962
rect 13634 12910 13636 12962
rect 13580 12898 13636 12910
rect 13356 12786 13412 12796
rect 13692 12628 13748 13916
rect 13580 12572 13748 12628
rect 13916 13860 13972 13870
rect 13468 12404 13524 12414
rect 12908 12180 12964 12190
rect 12908 10722 12964 12124
rect 13020 12178 13076 12190
rect 13020 12126 13022 12178
rect 13074 12126 13076 12178
rect 13020 12068 13076 12126
rect 13020 12002 13076 12012
rect 13468 11844 13524 12348
rect 12908 10670 12910 10722
rect 12962 10670 12964 10722
rect 12908 10658 12964 10670
rect 13356 11788 13524 11844
rect 13356 10724 13412 11788
rect 13468 11620 13524 11630
rect 13580 11620 13636 12572
rect 13692 12180 13748 12190
rect 13692 12086 13748 12124
rect 13916 12068 13972 13804
rect 14028 12404 14084 14028
rect 14140 13970 14196 15092
rect 14252 14644 14308 15262
rect 14364 14868 14420 16716
rect 14476 16660 14532 16670
rect 14588 16660 14644 17388
rect 14700 17378 14756 17388
rect 14532 16604 14644 16660
rect 14700 16658 14756 16670
rect 14700 16606 14702 16658
rect 14754 16606 14756 16658
rect 14476 15876 14532 16604
rect 14700 16436 14756 16606
rect 14588 15988 14644 15998
rect 14700 15988 14756 16380
rect 14588 15986 14756 15988
rect 14588 15934 14590 15986
rect 14642 15934 14756 15986
rect 14588 15932 14756 15934
rect 14588 15922 14644 15932
rect 14812 15876 14868 18396
rect 14924 17778 14980 17790
rect 14924 17726 14926 17778
rect 14978 17726 14980 17778
rect 14924 16882 14980 17726
rect 14924 16830 14926 16882
rect 14978 16830 14980 16882
rect 14924 16818 14980 16830
rect 15036 17554 15092 18956
rect 15036 17502 15038 17554
rect 15090 17502 15092 17554
rect 15036 16772 15092 17502
rect 15036 16706 15092 16716
rect 15260 17890 15316 21532
rect 15372 21364 15428 21374
rect 15372 20802 15428 21308
rect 15372 20750 15374 20802
rect 15426 20750 15428 20802
rect 15372 20692 15428 20750
rect 15372 20626 15428 20636
rect 15484 20244 15540 24446
rect 15932 23938 15988 25788
rect 16044 25394 16100 25900
rect 16156 25890 16212 25900
rect 16492 25506 16548 26348
rect 16716 26292 16772 26302
rect 16716 26198 16772 26236
rect 16828 25844 16884 28590
rect 17276 28420 17332 29932
rect 17500 29540 17556 29550
rect 17500 29446 17556 29484
rect 17388 29204 17444 29214
rect 17388 28642 17444 29148
rect 17388 28590 17390 28642
rect 17442 28590 17444 28642
rect 17388 28578 17444 28590
rect 17612 28644 17668 29932
rect 18172 29876 18228 31724
rect 18396 31556 18452 32396
rect 18508 31778 18564 33740
rect 18620 32564 18676 32574
rect 18844 32564 18900 33964
rect 18676 32508 18900 32564
rect 18620 32004 18676 32508
rect 18956 32452 19012 37324
rect 19516 37268 19572 40350
rect 20076 40402 20244 40404
rect 20076 40350 20190 40402
rect 20242 40350 20244 40402
rect 20076 40348 20244 40350
rect 19628 39732 19684 39742
rect 19628 39730 20020 39732
rect 19628 39678 19630 39730
rect 19682 39678 20020 39730
rect 19628 39676 20020 39678
rect 19628 39666 19684 39676
rect 19964 39618 20020 39676
rect 20076 39730 20132 40348
rect 20188 40338 20244 40348
rect 20300 40348 20412 40404
rect 20076 39678 20078 39730
rect 20130 39678 20132 39730
rect 20076 39666 20132 39678
rect 19964 39566 19966 39618
rect 20018 39566 20020 39618
rect 19964 39554 20020 39566
rect 20188 39620 20244 39630
rect 20300 39620 20356 40348
rect 20412 40338 20468 40348
rect 20188 39618 20356 39620
rect 20188 39566 20190 39618
rect 20242 39566 20356 39618
rect 20188 39564 20356 39566
rect 20188 39554 20244 39564
rect 19628 39508 19684 39518
rect 19628 39396 19684 39452
rect 19740 39396 19796 39406
rect 19628 39394 19796 39396
rect 19628 39342 19742 39394
rect 19794 39342 19796 39394
rect 19628 39340 19796 39342
rect 19628 39060 19684 39340
rect 19740 39330 19796 39340
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19964 39060 20020 39070
rect 19628 39058 20020 39060
rect 19628 39006 19966 39058
rect 20018 39006 20020 39058
rect 19628 39004 20020 39006
rect 19964 38994 20020 39004
rect 20300 38836 20356 38846
rect 20300 38742 20356 38780
rect 20188 38050 20244 38062
rect 20188 37998 20190 38050
rect 20242 37998 20244 38050
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19740 37268 19796 37278
rect 19516 37266 19796 37268
rect 19516 37214 19742 37266
rect 19794 37214 19796 37266
rect 19516 37212 19796 37214
rect 19740 37202 19796 37212
rect 19964 36820 20020 36830
rect 19740 36708 19796 36718
rect 19740 36594 19796 36652
rect 19964 36706 20020 36764
rect 19964 36654 19966 36706
rect 20018 36654 20020 36706
rect 19964 36642 20020 36654
rect 20188 36708 20244 37998
rect 20412 37826 20468 37838
rect 20412 37774 20414 37826
rect 20466 37774 20468 37826
rect 20412 37380 20468 37774
rect 21196 37492 21252 42140
rect 21644 42130 21700 42140
rect 21420 41972 21476 41982
rect 21420 41878 21476 41916
rect 21308 41858 21364 41870
rect 21308 41806 21310 41858
rect 21362 41806 21364 41858
rect 21308 41188 21364 41806
rect 21868 41412 21924 43372
rect 22092 43334 22148 43372
rect 22428 42868 22484 43486
rect 22988 43538 23044 43550
rect 22988 43486 22990 43538
rect 23042 43486 23044 43538
rect 22876 43426 22932 43438
rect 22876 43374 22878 43426
rect 22930 43374 22932 43426
rect 22876 43316 22932 43374
rect 22876 43250 22932 43260
rect 22764 43204 22820 43214
rect 22652 43148 22764 43204
rect 22540 42868 22596 42878
rect 22428 42866 22596 42868
rect 22428 42814 22542 42866
rect 22594 42814 22596 42866
rect 22428 42812 22596 42814
rect 22540 42802 22596 42812
rect 22428 42642 22484 42654
rect 22428 42590 22430 42642
rect 22482 42590 22484 42642
rect 22428 42084 22484 42590
rect 22652 42642 22708 43148
rect 22764 43138 22820 43148
rect 22652 42590 22654 42642
rect 22706 42590 22708 42642
rect 22652 42578 22708 42590
rect 22988 42532 23044 43486
rect 23212 42754 23268 43932
rect 23324 43204 23380 44046
rect 23996 43988 24052 43998
rect 23324 43138 23380 43148
rect 23436 43538 23492 43550
rect 23436 43486 23438 43538
rect 23490 43486 23492 43538
rect 23436 43428 23492 43486
rect 23436 42980 23492 43372
rect 23884 43538 23940 43550
rect 23884 43486 23886 43538
rect 23938 43486 23940 43538
rect 23436 42924 23828 42980
rect 23660 42756 23716 42766
rect 23212 42702 23214 42754
rect 23266 42702 23268 42754
rect 23212 42690 23268 42702
rect 23548 42700 23660 42756
rect 23548 42642 23604 42700
rect 23660 42690 23716 42700
rect 23548 42590 23550 42642
rect 23602 42590 23604 42642
rect 23548 42578 23604 42590
rect 23436 42532 23492 42542
rect 22988 42530 23492 42532
rect 22988 42478 23438 42530
rect 23490 42478 23492 42530
rect 22988 42476 23492 42478
rect 23436 42466 23492 42476
rect 23212 42196 23268 42206
rect 23212 42102 23268 42140
rect 22484 42028 22708 42084
rect 22428 42018 22484 42028
rect 21868 41318 21924 41356
rect 22204 41748 22260 41758
rect 22204 41298 22260 41692
rect 22204 41246 22206 41298
rect 22258 41246 22260 41298
rect 22204 41234 22260 41246
rect 21532 41188 21588 41198
rect 21308 41186 21588 41188
rect 21308 41134 21534 41186
rect 21586 41134 21588 41186
rect 21308 41132 21588 41134
rect 21532 41122 21588 41132
rect 22316 41188 22372 41198
rect 22316 41094 22372 41132
rect 22092 41076 22148 41086
rect 22092 41074 22260 41076
rect 22092 41022 22094 41074
rect 22146 41022 22260 41074
rect 22092 41020 22260 41022
rect 22092 41010 22148 41020
rect 22204 40292 22260 41020
rect 22652 40626 22708 42028
rect 23436 41970 23492 41982
rect 23436 41918 23438 41970
rect 23490 41918 23492 41970
rect 23212 41412 23268 41422
rect 23212 41074 23268 41356
rect 23212 41022 23214 41074
rect 23266 41022 23268 41074
rect 23212 41010 23268 41022
rect 23436 40964 23492 41918
rect 23548 41076 23604 41086
rect 23548 40982 23604 41020
rect 22652 40574 22654 40626
rect 22706 40574 22708 40626
rect 22652 40562 22708 40574
rect 22988 40628 23044 40638
rect 22316 40292 22372 40302
rect 22204 40236 22316 40292
rect 22316 40198 22372 40236
rect 22988 38052 23044 40572
rect 23212 38052 23268 38062
rect 22988 38050 23268 38052
rect 22988 37998 23214 38050
rect 23266 37998 23268 38050
rect 22988 37996 23268 37998
rect 21196 37426 21252 37436
rect 22316 37828 22372 37838
rect 20524 37380 20580 37390
rect 20412 37378 20580 37380
rect 20412 37326 20526 37378
rect 20578 37326 20580 37378
rect 20412 37324 20580 37326
rect 20524 37314 20580 37324
rect 20300 36708 20356 36718
rect 20188 36706 20356 36708
rect 20188 36654 20302 36706
rect 20354 36654 20356 36706
rect 20188 36652 20356 36654
rect 20300 36642 20356 36652
rect 20748 36708 20804 36718
rect 20748 36596 20804 36652
rect 19740 36542 19742 36594
rect 19794 36542 19796 36594
rect 19740 36530 19796 36542
rect 20524 36594 20804 36596
rect 20524 36542 20750 36594
rect 20802 36542 20804 36594
rect 20524 36540 20804 36542
rect 19292 36372 19348 36382
rect 19292 36370 19684 36372
rect 19292 36318 19294 36370
rect 19346 36318 19684 36370
rect 19292 36316 19684 36318
rect 19292 36306 19348 36316
rect 19180 36260 19236 36270
rect 19068 36258 19236 36260
rect 19068 36206 19182 36258
rect 19234 36206 19236 36258
rect 19068 36204 19236 36206
rect 19068 35810 19124 36204
rect 19180 36194 19236 36204
rect 19068 35758 19070 35810
rect 19122 35758 19124 35810
rect 19068 35746 19124 35758
rect 19628 35028 19684 36316
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19852 35476 19908 35486
rect 19740 35028 19796 35038
rect 19628 35026 19796 35028
rect 19628 34974 19742 35026
rect 19794 34974 19796 35026
rect 19628 34972 19796 34974
rect 19740 34962 19796 34972
rect 19852 34914 19908 35420
rect 20524 35364 20580 36540
rect 20748 36530 20804 36540
rect 21196 35812 21252 35822
rect 21196 35586 21252 35756
rect 22316 35810 22372 37772
rect 22652 37156 22708 37166
rect 22652 37154 22932 37156
rect 22652 37102 22654 37154
rect 22706 37102 22932 37154
rect 22652 37100 22932 37102
rect 22652 37090 22708 37100
rect 22428 36260 22484 36270
rect 22428 36258 22596 36260
rect 22428 36206 22430 36258
rect 22482 36206 22596 36258
rect 22428 36204 22596 36206
rect 22428 36194 22484 36204
rect 22316 35758 22318 35810
rect 22370 35758 22372 35810
rect 22316 35746 22372 35758
rect 22540 35812 22596 36204
rect 21196 35534 21198 35586
rect 21250 35534 21252 35586
rect 21196 35522 21252 35534
rect 21644 35476 21700 35486
rect 21644 35382 21700 35420
rect 21980 35476 22036 35486
rect 21980 35382 22036 35420
rect 19852 34862 19854 34914
rect 19906 34862 19908 34914
rect 19852 34850 19908 34862
rect 20300 34916 20356 34926
rect 19404 34690 19460 34702
rect 19404 34638 19406 34690
rect 19458 34638 19460 34690
rect 19404 33684 19460 34638
rect 19404 33618 19460 33628
rect 19628 34690 19684 34702
rect 19628 34638 19630 34690
rect 19682 34638 19684 34690
rect 19516 33348 19572 33358
rect 19292 33346 19572 33348
rect 19292 33294 19518 33346
rect 19570 33294 19572 33346
rect 19292 33292 19572 33294
rect 19180 33122 19236 33134
rect 19180 33070 19182 33122
rect 19234 33070 19236 33122
rect 19180 32676 19236 33070
rect 19180 32610 19236 32620
rect 19292 32674 19348 33292
rect 19516 33282 19572 33292
rect 19628 33236 19684 34638
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20188 33684 20244 33694
rect 20076 33460 20132 33470
rect 20076 33346 20132 33404
rect 20076 33294 20078 33346
rect 20130 33294 20132 33346
rect 20076 33282 20132 33294
rect 19628 33142 19684 33180
rect 19292 32622 19294 32674
rect 19346 32622 19348 32674
rect 19292 32610 19348 32622
rect 19404 33122 19460 33134
rect 19404 33070 19406 33122
rect 19458 33070 19460 33122
rect 18956 32396 19236 32452
rect 18620 31938 18676 31948
rect 18508 31726 18510 31778
rect 18562 31726 18564 31778
rect 18508 31714 18564 31726
rect 19180 31780 19236 32396
rect 19404 32002 19460 33070
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19404 31950 19406 32002
rect 19458 31950 19460 32002
rect 19404 31938 19460 31950
rect 19628 32676 19684 32686
rect 19516 31780 19572 31790
rect 19180 31778 19572 31780
rect 19180 31726 19518 31778
rect 19570 31726 19572 31778
rect 19180 31724 19572 31726
rect 19516 31714 19572 31724
rect 19068 31668 19124 31678
rect 18396 31500 18788 31556
rect 18732 30994 18788 31500
rect 18732 30942 18734 30994
rect 18786 30942 18788 30994
rect 18732 30930 18788 30942
rect 19068 30324 19124 31612
rect 19628 31556 19684 32620
rect 19740 32340 19796 32350
rect 19740 32002 19796 32284
rect 19740 31950 19742 32002
rect 19794 31950 19796 32002
rect 19740 31938 19796 31950
rect 19852 31778 19908 31790
rect 19852 31726 19854 31778
rect 19906 31726 19908 31778
rect 19852 31556 19908 31726
rect 19068 30258 19124 30268
rect 19292 31500 19908 31556
rect 20188 31556 20244 33628
rect 20300 31892 20356 34860
rect 20412 34690 20468 34702
rect 20412 34638 20414 34690
rect 20466 34638 20468 34690
rect 20412 33684 20468 34638
rect 20412 33618 20468 33628
rect 20412 33460 20468 33470
rect 20524 33460 20580 35308
rect 22428 35028 22484 35038
rect 22540 35028 22596 35756
rect 22652 36258 22708 36270
rect 22652 36206 22654 36258
rect 22706 36206 22708 36258
rect 22652 35924 22708 36206
rect 22764 36258 22820 36270
rect 22764 36206 22766 36258
rect 22818 36206 22820 36258
rect 22764 36148 22820 36206
rect 22876 36258 22932 37100
rect 23212 36484 23268 37996
rect 23436 37828 23492 40908
rect 23772 40852 23828 42924
rect 23884 42196 23940 43486
rect 23884 42130 23940 42140
rect 23884 40964 23940 40974
rect 23884 40870 23940 40908
rect 23548 40796 23828 40852
rect 23548 39060 23604 40796
rect 23996 40516 24052 43932
rect 24108 43650 24164 44156
rect 24108 43598 24110 43650
rect 24162 43598 24164 43650
rect 24108 43586 24164 43598
rect 24220 41972 24276 45164
rect 24332 45154 24388 45164
rect 24332 43316 24388 43326
rect 24444 43316 24500 45388
rect 24556 45108 24612 45612
rect 24556 45106 24948 45108
rect 24556 45054 24558 45106
rect 24610 45054 24948 45106
rect 24556 45052 24948 45054
rect 24556 45042 24612 45052
rect 24892 44434 24948 45052
rect 24892 44382 24894 44434
rect 24946 44382 24948 44434
rect 24892 44370 24948 44382
rect 25004 43988 25060 45838
rect 27244 45890 27524 45892
rect 27244 45838 27470 45890
rect 27522 45838 27524 45890
rect 27244 45836 27524 45838
rect 25340 45108 25396 45118
rect 25340 45014 25396 45052
rect 26012 44996 26068 45006
rect 25004 43922 25060 43932
rect 25452 44994 26068 44996
rect 25452 44942 26014 44994
rect 26066 44942 26068 44994
rect 25452 44940 26068 44942
rect 24668 43764 24724 43774
rect 25340 43764 25396 43774
rect 25452 43764 25508 44940
rect 26012 44930 26068 44940
rect 26796 44996 26852 45006
rect 24668 43762 25172 43764
rect 24668 43710 24670 43762
rect 24722 43710 25172 43762
rect 24668 43708 25172 43710
rect 24668 43698 24724 43708
rect 25116 43652 25172 43708
rect 25340 43762 25508 43764
rect 25340 43710 25342 43762
rect 25394 43710 25508 43762
rect 25340 43708 25508 43710
rect 26796 43708 26852 44940
rect 27244 44434 27300 45836
rect 27468 45826 27524 45836
rect 28252 46228 28308 49200
rect 28588 46786 28644 46798
rect 28588 46734 28590 46786
rect 28642 46734 28644 46786
rect 28252 46172 28532 46228
rect 27804 45668 27860 45678
rect 27804 45666 28084 45668
rect 27804 45614 27806 45666
rect 27858 45614 28084 45666
rect 27804 45612 28084 45614
rect 27804 45602 27860 45612
rect 27244 44382 27246 44434
rect 27298 44382 27300 44434
rect 27244 44370 27300 44382
rect 25340 43698 25396 43708
rect 25228 43652 25284 43662
rect 25116 43650 25284 43652
rect 25116 43598 25230 43650
rect 25282 43598 25284 43650
rect 25116 43596 25284 43598
rect 25228 43586 25284 43596
rect 25676 43650 25732 43662
rect 25676 43598 25678 43650
rect 25730 43598 25732 43650
rect 24668 43540 24724 43550
rect 25452 43540 25508 43550
rect 24668 43446 24724 43484
rect 25340 43538 25508 43540
rect 25340 43486 25454 43538
rect 25506 43486 25508 43538
rect 25340 43484 25508 43486
rect 24444 43260 24836 43316
rect 24332 43222 24388 43260
rect 24780 42754 24836 43260
rect 25340 43092 25396 43484
rect 25452 43474 25508 43484
rect 25564 43540 25620 43550
rect 25004 43036 25396 43092
rect 25004 42866 25060 43036
rect 25004 42814 25006 42866
rect 25058 42814 25060 42866
rect 25004 42802 25060 42814
rect 25564 42866 25620 43484
rect 25676 43428 25732 43598
rect 26236 43652 26852 43708
rect 27356 43764 27412 43774
rect 27804 43764 27860 43774
rect 27356 43762 27860 43764
rect 27356 43710 27358 43762
rect 27410 43710 27806 43762
rect 27858 43710 27860 43762
rect 27356 43708 27860 43710
rect 27356 43698 27412 43708
rect 27804 43698 27860 43708
rect 28028 43708 28084 45612
rect 28140 44996 28196 45006
rect 28140 44902 28196 44940
rect 28252 44434 28308 46172
rect 28252 44382 28254 44434
rect 28306 44382 28308 44434
rect 28252 44370 28308 44382
rect 28364 45666 28420 45678
rect 28364 45614 28366 45666
rect 28418 45614 28420 45666
rect 28364 43708 28420 45614
rect 28476 45218 28532 46172
rect 28588 45890 28644 46734
rect 28924 46116 28980 49200
rect 28924 46050 28980 46060
rect 30044 46116 30100 46126
rect 30044 46022 30100 46060
rect 28588 45838 28590 45890
rect 28642 45838 28644 45890
rect 28588 45332 28644 45838
rect 28588 45266 28644 45276
rect 29260 45890 29316 45902
rect 29260 45838 29262 45890
rect 29314 45838 29316 45890
rect 28476 45166 28478 45218
rect 28530 45166 28532 45218
rect 28476 45154 28532 45166
rect 28812 45218 28868 45230
rect 28812 45166 28814 45218
rect 28866 45166 28868 45218
rect 28812 43764 28868 45166
rect 28924 43764 28980 43774
rect 28812 43762 28980 43764
rect 28812 43710 28926 43762
rect 28978 43710 28980 43762
rect 28812 43708 28980 43710
rect 28028 43652 28196 43708
rect 26236 43650 26292 43652
rect 26236 43598 26238 43650
rect 26290 43598 26292 43650
rect 26236 43586 26292 43598
rect 26796 43650 26852 43652
rect 26796 43598 26798 43650
rect 26850 43598 26852 43650
rect 26796 43586 26852 43598
rect 25676 43362 25732 43372
rect 26572 43538 26628 43550
rect 26572 43486 26574 43538
rect 26626 43486 26628 43538
rect 26124 43316 26180 43326
rect 25564 42814 25566 42866
rect 25618 42814 25620 42866
rect 25564 42802 25620 42814
rect 25788 43314 26180 43316
rect 25788 43262 26126 43314
rect 26178 43262 26180 43314
rect 25788 43260 26180 43262
rect 24780 42702 24782 42754
rect 24834 42702 24836 42754
rect 24780 42690 24836 42702
rect 25116 42756 25172 42766
rect 25116 42662 25172 42700
rect 25788 42754 25844 43260
rect 26124 43250 26180 43260
rect 25788 42702 25790 42754
rect 25842 42702 25844 42754
rect 25788 42690 25844 42702
rect 25452 42642 25508 42654
rect 25452 42590 25454 42642
rect 25506 42590 25508 42642
rect 25452 41972 25508 42590
rect 24220 41916 24724 41972
rect 24556 41076 24612 41086
rect 24220 40964 24276 40974
rect 24276 40908 24388 40964
rect 24220 40870 24276 40908
rect 23884 40460 24052 40516
rect 23660 40404 23716 40414
rect 23660 40310 23716 40348
rect 23772 40292 23828 40302
rect 23772 40198 23828 40236
rect 23884 39620 23940 40460
rect 24220 40404 24276 40442
rect 24220 40338 24276 40348
rect 23996 40180 24052 40190
rect 24332 40180 24388 40908
rect 23996 40178 24388 40180
rect 23996 40126 23998 40178
rect 24050 40126 24388 40178
rect 23996 40124 24388 40126
rect 23996 40114 24052 40124
rect 24556 39956 24612 41020
rect 23772 39564 23940 39620
rect 24108 39900 24612 39956
rect 23660 39060 23716 39070
rect 23548 39058 23716 39060
rect 23548 39006 23662 39058
rect 23714 39006 23716 39058
rect 23548 39004 23716 39006
rect 23660 38994 23716 39004
rect 23772 38668 23828 39564
rect 23884 39396 23940 39406
rect 23884 39302 23940 39340
rect 23660 38612 23828 38668
rect 23996 38834 24052 38846
rect 23996 38782 23998 38834
rect 24050 38782 24052 38834
rect 23996 38612 24052 38782
rect 23436 37734 23492 37772
rect 23548 38276 23604 38286
rect 23212 36418 23268 36428
rect 23324 36370 23380 36382
rect 23324 36318 23326 36370
rect 23378 36318 23380 36370
rect 23324 36260 23380 36318
rect 22876 36206 22878 36258
rect 22930 36206 22932 36258
rect 22876 36148 22932 36206
rect 23100 36204 23380 36260
rect 23436 36258 23492 36270
rect 23436 36206 23438 36258
rect 23490 36206 23492 36258
rect 23100 36148 23156 36204
rect 22876 36092 23156 36148
rect 22764 36082 22820 36092
rect 22652 35138 22708 35868
rect 23100 35308 23156 36092
rect 23212 36036 23268 36046
rect 23212 35810 23268 35980
rect 23436 36036 23492 36206
rect 23436 35970 23492 35980
rect 23212 35758 23214 35810
rect 23266 35758 23268 35810
rect 23212 35746 23268 35758
rect 23324 35812 23380 35822
rect 23324 35810 23492 35812
rect 23324 35758 23326 35810
rect 23378 35758 23492 35810
rect 23324 35756 23492 35758
rect 23324 35746 23380 35756
rect 23324 35476 23380 35486
rect 23324 35382 23380 35420
rect 22652 35086 22654 35138
rect 22706 35086 22708 35138
rect 22652 35074 22708 35086
rect 22876 35252 23156 35308
rect 22876 35138 22932 35252
rect 22876 35086 22878 35138
rect 22930 35086 22932 35138
rect 22876 35074 22932 35086
rect 23324 35140 23380 35150
rect 23436 35140 23492 35756
rect 23324 35138 23492 35140
rect 23324 35086 23326 35138
rect 23378 35086 23492 35138
rect 23324 35084 23492 35086
rect 22428 35026 22596 35028
rect 22428 34974 22430 35026
rect 22482 34974 22596 35026
rect 22428 34972 22596 34974
rect 22428 34962 22484 34972
rect 23100 34804 23156 34814
rect 20748 34692 20804 34702
rect 20748 34354 20804 34636
rect 20748 34302 20750 34354
rect 20802 34302 20804 34354
rect 20748 34290 20804 34302
rect 22428 34580 22484 34590
rect 20468 33404 20580 33460
rect 20412 33366 20468 33404
rect 22204 33236 22260 33246
rect 22204 32786 22260 33180
rect 22204 32734 22206 32786
rect 22258 32734 22260 32786
rect 22204 32722 22260 32734
rect 22428 32786 22484 34524
rect 23100 33458 23156 34748
rect 23100 33406 23102 33458
rect 23154 33406 23156 33458
rect 23100 33394 23156 33406
rect 23212 33234 23268 33246
rect 23212 33182 23214 33234
rect 23266 33182 23268 33234
rect 22428 32734 22430 32786
rect 22482 32734 22484 32786
rect 22428 32722 22484 32734
rect 22988 33124 23044 33134
rect 22876 32562 22932 32574
rect 22876 32510 22878 32562
rect 22930 32510 22932 32562
rect 21420 32450 21476 32462
rect 21420 32398 21422 32450
rect 21474 32398 21476 32450
rect 21420 32340 21476 32398
rect 21420 32274 21476 32284
rect 22316 32450 22372 32462
rect 22316 32398 22318 32450
rect 22370 32398 22372 32450
rect 21420 32004 21476 32014
rect 20300 31836 21364 31892
rect 20300 31778 20356 31836
rect 20300 31726 20302 31778
rect 20354 31726 20356 31778
rect 20300 31714 20356 31726
rect 20972 31668 21028 31678
rect 20636 31556 20692 31566
rect 20188 31554 20692 31556
rect 20188 31502 20638 31554
rect 20690 31502 20692 31554
rect 20188 31500 20692 31502
rect 18396 30100 18452 30110
rect 17836 29820 18228 29876
rect 18284 30098 18452 30100
rect 18284 30046 18398 30098
rect 18450 30046 18452 30098
rect 18284 30044 18452 30046
rect 17836 28866 17892 29820
rect 17948 29652 18004 29662
rect 17948 29558 18004 29596
rect 18060 29428 18116 29438
rect 18284 29428 18340 30044
rect 18396 30034 18452 30044
rect 18732 30100 18788 30110
rect 19068 30100 19124 30110
rect 18732 30098 19124 30100
rect 18732 30046 18734 30098
rect 18786 30046 19070 30098
rect 19122 30046 19124 30098
rect 18732 30044 19124 30046
rect 18732 30034 18788 30044
rect 19068 30034 19124 30044
rect 18508 29988 18564 29998
rect 18508 29986 18676 29988
rect 18508 29934 18510 29986
rect 18562 29934 18676 29986
rect 18508 29932 18676 29934
rect 18508 29922 18564 29932
rect 18060 29426 18228 29428
rect 18060 29374 18062 29426
rect 18114 29374 18228 29426
rect 18060 29372 18228 29374
rect 18060 29362 18116 29372
rect 17836 28814 17838 28866
rect 17890 28814 17892 28866
rect 17836 28802 17892 28814
rect 17612 28588 17892 28644
rect 17276 28364 17444 28420
rect 17276 28196 17332 28206
rect 16828 25778 16884 25788
rect 16940 27748 16996 27758
rect 16492 25454 16494 25506
rect 16546 25454 16548 25506
rect 16492 25442 16548 25454
rect 16940 25506 16996 27692
rect 17276 26962 17332 28140
rect 17276 26910 17278 26962
rect 17330 26910 17332 26962
rect 17276 26898 17332 26910
rect 17388 26290 17444 28364
rect 17724 27634 17780 27646
rect 17724 27582 17726 27634
rect 17778 27582 17780 27634
rect 17612 27076 17668 27114
rect 17612 27010 17668 27020
rect 17724 26908 17780 27582
rect 17836 27636 17892 28588
rect 18172 28196 18228 29372
rect 18284 29334 18340 29372
rect 18620 29426 18676 29932
rect 19180 29986 19236 29998
rect 19180 29934 19182 29986
rect 19234 29934 19236 29986
rect 19180 29652 19236 29934
rect 19292 29764 19348 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19404 29988 19460 29998
rect 19740 29988 19796 30026
rect 19404 29986 19684 29988
rect 19404 29934 19406 29986
rect 19458 29934 19684 29986
rect 19404 29932 19684 29934
rect 19404 29922 19460 29932
rect 19292 29708 19460 29764
rect 19180 29586 19236 29596
rect 18844 29540 18900 29550
rect 18844 29538 19012 29540
rect 18844 29486 18846 29538
rect 18898 29486 19012 29538
rect 18844 29484 19012 29486
rect 18844 29474 18900 29484
rect 18620 29374 18622 29426
rect 18674 29374 18676 29426
rect 18620 28196 18676 29374
rect 18844 29314 18900 29326
rect 18844 29262 18846 29314
rect 18898 29262 18900 29314
rect 18844 29092 18900 29262
rect 18172 28140 18564 28196
rect 18508 28084 18564 28140
rect 18620 28130 18676 28140
rect 18732 28642 18788 28654
rect 18732 28590 18734 28642
rect 18786 28590 18788 28642
rect 18284 27970 18340 27982
rect 18284 27918 18286 27970
rect 18338 27918 18340 27970
rect 17948 27860 18004 27870
rect 17948 27766 18004 27804
rect 17836 27580 18004 27636
rect 17388 26238 17390 26290
rect 17442 26238 17444 26290
rect 17388 25956 17444 26238
rect 17500 26852 17780 26908
rect 17836 26852 17892 26862
rect 17500 26068 17556 26852
rect 17836 26514 17892 26796
rect 17836 26462 17838 26514
rect 17890 26462 17892 26514
rect 17500 26002 17556 26012
rect 17612 26290 17668 26302
rect 17612 26238 17614 26290
rect 17666 26238 17668 26290
rect 17388 25890 17444 25900
rect 16940 25454 16942 25506
rect 16994 25454 16996 25506
rect 16940 25442 16996 25454
rect 17612 25508 17668 26238
rect 17724 26292 17780 26302
rect 17724 26198 17780 26236
rect 17612 25442 17668 25452
rect 17724 25508 17780 25518
rect 17836 25508 17892 26462
rect 17724 25506 17892 25508
rect 17724 25454 17726 25506
rect 17778 25454 17892 25506
rect 17724 25452 17892 25454
rect 17948 26290 18004 27580
rect 18284 26964 18340 27918
rect 18508 27970 18564 28028
rect 18508 27918 18510 27970
rect 18562 27918 18564 27970
rect 18508 27906 18564 27918
rect 18732 27858 18788 28590
rect 18732 27806 18734 27858
rect 18786 27806 18788 27858
rect 18396 27076 18452 27114
rect 18732 27076 18788 27806
rect 18452 27020 18788 27076
rect 18396 27010 18452 27020
rect 18284 26898 18340 26908
rect 18396 26852 18452 26862
rect 18396 26758 18452 26796
rect 17948 26238 17950 26290
rect 18002 26238 18004 26290
rect 17724 25442 17780 25452
rect 16044 25342 16046 25394
rect 16098 25342 16100 25394
rect 16044 25330 16100 25342
rect 17948 25394 18004 26238
rect 17948 25342 17950 25394
rect 18002 25342 18004 25394
rect 17948 25330 18004 25342
rect 16156 25284 16212 25294
rect 16156 24722 16212 25228
rect 16156 24670 16158 24722
rect 16210 24670 16212 24722
rect 16156 24658 16212 24670
rect 16380 25282 16436 25294
rect 16380 25230 16382 25282
rect 16434 25230 16436 25282
rect 16380 24610 16436 25230
rect 18508 24948 18564 27020
rect 18620 26852 18676 26862
rect 18620 26290 18676 26796
rect 18620 26238 18622 26290
rect 18674 26238 18676 26290
rect 18620 26226 18676 26238
rect 18844 26290 18900 29036
rect 18956 28644 19012 29484
rect 19292 29316 19348 29326
rect 19292 29222 19348 29260
rect 19404 29092 19460 29708
rect 19628 29652 19684 29932
rect 19740 29922 19796 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19628 29596 19908 29652
rect 19516 29426 19572 29438
rect 19516 29374 19518 29426
rect 19570 29374 19572 29426
rect 19516 29204 19572 29374
rect 19516 29138 19572 29148
rect 19628 29426 19684 29438
rect 19628 29374 19630 29426
rect 19682 29374 19684 29426
rect 19292 29036 19460 29092
rect 19628 29092 19684 29374
rect 19852 29426 19908 29596
rect 19852 29374 19854 29426
rect 19906 29374 19908 29426
rect 19852 29362 19908 29374
rect 20300 29428 20356 29438
rect 20524 29428 20580 29438
rect 20300 29426 20580 29428
rect 20300 29374 20302 29426
rect 20354 29374 20526 29426
rect 20578 29374 20580 29426
rect 20300 29372 20580 29374
rect 20300 29362 20356 29372
rect 20524 29362 20580 29372
rect 20636 29316 20692 31500
rect 20636 29250 20692 29260
rect 20748 30994 20804 31006
rect 20748 30942 20750 30994
rect 20802 30942 20804 30994
rect 19180 28980 19236 28990
rect 19068 28644 19124 28654
rect 18956 28642 19124 28644
rect 18956 28590 19070 28642
rect 19122 28590 19124 28642
rect 18956 28588 19124 28590
rect 19068 28308 19124 28588
rect 19068 27858 19124 28252
rect 19068 27806 19070 27858
rect 19122 27806 19124 27858
rect 19068 27794 19124 27806
rect 19180 26852 19236 28924
rect 19180 26786 19236 26796
rect 19292 26516 19348 29036
rect 19628 29026 19684 29036
rect 20748 28980 20804 30942
rect 20972 30996 21028 31612
rect 21308 31666 21364 31836
rect 21308 31614 21310 31666
rect 21362 31614 21364 31666
rect 21308 31332 21364 31614
rect 21308 31266 21364 31276
rect 21420 31220 21476 31948
rect 22204 31892 22260 31902
rect 21644 31556 21700 31566
rect 22092 31556 22148 31566
rect 21644 31554 22148 31556
rect 21644 31502 21646 31554
rect 21698 31502 22094 31554
rect 22146 31502 22148 31554
rect 21644 31500 22148 31502
rect 21644 31490 21700 31500
rect 22092 31444 22148 31500
rect 21756 31332 21812 31342
rect 21420 31164 21588 31220
rect 21420 30996 21476 31006
rect 20972 30994 21476 30996
rect 20972 30942 20974 30994
rect 21026 30942 21422 30994
rect 21474 30942 21476 30994
rect 20972 30940 21476 30942
rect 20972 30930 21028 30940
rect 21420 30930 21476 30940
rect 21532 30212 21588 31164
rect 21756 31106 21812 31276
rect 21756 31054 21758 31106
rect 21810 31054 21812 31106
rect 21756 31042 21812 31054
rect 21980 31220 22036 31230
rect 21980 31106 22036 31164
rect 21980 31054 21982 31106
rect 22034 31054 22036 31106
rect 21980 31042 22036 31054
rect 21644 30212 21700 30222
rect 21532 30210 21700 30212
rect 21532 30158 21646 30210
rect 21698 30158 21700 30210
rect 21532 30156 21700 30158
rect 20748 28914 20804 28924
rect 20860 29538 20916 29550
rect 20860 29486 20862 29538
rect 20914 29486 20916 29538
rect 19404 28644 19460 28654
rect 19404 28550 19460 28588
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 28084 19572 28094
rect 19516 27858 19572 28028
rect 19516 27806 19518 27858
rect 19570 27806 19572 27858
rect 19516 27794 19572 27806
rect 20076 28084 20132 28094
rect 20076 27746 20132 28028
rect 20860 27972 20916 29486
rect 21308 29316 21364 29326
rect 21308 29222 21364 29260
rect 21420 29204 21476 29214
rect 21420 28530 21476 29148
rect 21420 28478 21422 28530
rect 21474 28478 21476 28530
rect 21420 28466 21476 28478
rect 21532 28756 21588 28766
rect 21532 28530 21588 28700
rect 21532 28478 21534 28530
rect 21586 28478 21588 28530
rect 21532 28466 21588 28478
rect 20860 27906 20916 27916
rect 20076 27694 20078 27746
rect 20130 27694 20132 27746
rect 20076 27682 20132 27694
rect 21644 27860 21700 30156
rect 22092 28756 22148 31388
rect 22204 30996 22260 31836
rect 22316 31668 22372 32398
rect 22876 32228 22932 32510
rect 22988 32452 23044 33068
rect 23212 33012 23268 33182
rect 23212 32946 23268 32956
rect 23100 32676 23156 32686
rect 23324 32676 23380 35084
rect 23548 33348 23604 38220
rect 23660 35476 23716 38612
rect 23996 38276 24052 38556
rect 23884 38220 24052 38276
rect 23772 37938 23828 37950
rect 23772 37886 23774 37938
rect 23826 37886 23828 37938
rect 23772 37828 23828 37886
rect 23884 37828 23940 38220
rect 23996 38052 24052 38062
rect 24108 38052 24164 39900
rect 24668 39844 24724 41916
rect 25004 41188 25060 41198
rect 25004 41074 25060 41132
rect 25452 41188 25508 41916
rect 25452 41122 25508 41132
rect 25564 41412 25620 41422
rect 25004 41022 25006 41074
rect 25058 41022 25060 41074
rect 25004 41010 25060 41022
rect 25228 41076 25284 41086
rect 25228 40626 25284 41020
rect 25228 40574 25230 40626
rect 25282 40574 25284 40626
rect 25228 40562 25284 40574
rect 25340 41074 25396 41086
rect 25340 41022 25342 41074
rect 25394 41022 25396 41074
rect 25340 40628 25396 41022
rect 25340 40562 25396 40572
rect 25564 40626 25620 41356
rect 26124 41298 26180 41310
rect 26124 41246 26126 41298
rect 26178 41246 26180 41298
rect 25788 41188 25844 41198
rect 26124 41188 26180 41246
rect 26460 41188 26516 41198
rect 26124 41186 26516 41188
rect 26124 41134 26462 41186
rect 26514 41134 26516 41186
rect 26124 41132 26516 41134
rect 25788 41094 25844 41132
rect 26460 41122 26516 41132
rect 25564 40574 25566 40626
rect 25618 40574 25620 40626
rect 25564 40404 25620 40574
rect 25564 40338 25620 40348
rect 26012 40962 26068 40974
rect 26012 40910 26014 40962
rect 26066 40910 26068 40962
rect 24332 39788 24724 39844
rect 26012 39844 26068 40910
rect 26572 40964 26628 43486
rect 27132 43538 27188 43550
rect 27132 43486 27134 43538
rect 27186 43486 27188 43538
rect 26908 43316 26964 43326
rect 27020 43316 27076 43326
rect 26964 43314 27076 43316
rect 26964 43262 27022 43314
rect 27074 43262 27076 43314
rect 26964 43260 27076 43262
rect 26796 42642 26852 42654
rect 26796 42590 26798 42642
rect 26850 42590 26852 42642
rect 26796 41972 26852 42590
rect 26796 41906 26852 41916
rect 26796 41412 26852 41422
rect 26908 41412 26964 43260
rect 27020 43250 27076 43260
rect 27132 42978 27188 43486
rect 28028 43540 28084 43550
rect 28028 43446 28084 43484
rect 27132 42926 27134 42978
rect 27186 42926 27188 42978
rect 27132 42914 27188 42926
rect 27916 43426 27972 43438
rect 27916 43374 27918 43426
rect 27970 43374 27972 43426
rect 27916 42868 27972 43374
rect 27916 42802 27972 42812
rect 28028 43316 28084 43326
rect 27132 42756 27188 42766
rect 27468 42756 27524 42766
rect 27132 42754 27524 42756
rect 27132 42702 27134 42754
rect 27186 42702 27470 42754
rect 27522 42702 27524 42754
rect 27132 42700 27524 42702
rect 27132 42690 27188 42700
rect 27468 42690 27524 42700
rect 27580 42644 27636 42654
rect 27580 42196 27636 42588
rect 26852 41356 26964 41412
rect 27020 42140 27636 42196
rect 26796 41318 26852 41356
rect 27020 41186 27076 42140
rect 27132 41300 27188 41310
rect 27132 41298 27636 41300
rect 27132 41246 27134 41298
rect 27186 41246 27636 41298
rect 27132 41244 27636 41246
rect 27132 41234 27188 41244
rect 27020 41134 27022 41186
rect 27074 41134 27076 41186
rect 27020 41122 27076 41134
rect 27580 41186 27636 41244
rect 27580 41134 27582 41186
rect 27634 41134 27636 41186
rect 27580 41122 27636 41134
rect 27244 41074 27300 41086
rect 27244 41022 27246 41074
rect 27298 41022 27300 41074
rect 27244 40964 27300 41022
rect 26628 40908 27300 40964
rect 27356 41076 27412 41086
rect 26460 40516 26516 40526
rect 24220 39620 24276 39630
rect 24220 39526 24276 39564
rect 24332 38612 24388 39788
rect 26012 39778 26068 39788
rect 26348 40514 26516 40516
rect 26348 40462 26462 40514
rect 26514 40462 26516 40514
rect 26348 40460 26516 40462
rect 26348 39732 26404 40460
rect 26460 40450 26516 40460
rect 26572 40514 26628 40908
rect 27356 40852 27412 41020
rect 28028 41074 28084 43260
rect 28028 41022 28030 41074
rect 28082 41022 28084 41074
rect 28028 41010 28084 41022
rect 27692 40964 27748 40974
rect 27692 40870 27748 40908
rect 27804 40962 27860 40974
rect 27804 40910 27806 40962
rect 27858 40910 27860 40962
rect 27244 40796 27412 40852
rect 27244 40626 27300 40796
rect 27804 40740 27860 40910
rect 27244 40574 27246 40626
rect 27298 40574 27300 40626
rect 27244 40562 27300 40574
rect 27356 40684 27860 40740
rect 26572 40462 26574 40514
rect 26626 40462 26628 40514
rect 26572 40450 26628 40462
rect 27020 40292 27076 40302
rect 26348 39666 26404 39676
rect 26460 40178 26516 40190
rect 26460 40126 26462 40178
rect 26514 40126 26516 40178
rect 24220 38556 24388 38612
rect 24444 38834 24500 38846
rect 24444 38782 24446 38834
rect 24498 38782 24500 38834
rect 24444 38612 24500 38782
rect 24220 38276 24276 38556
rect 24444 38546 24500 38556
rect 24668 38836 24724 38846
rect 24444 38388 24500 38398
rect 24500 38332 24612 38388
rect 24444 38322 24500 38332
rect 24220 38210 24276 38220
rect 23996 38050 24276 38052
rect 23996 37998 23998 38050
rect 24050 37998 24276 38050
rect 23996 37996 24276 37998
rect 23996 37986 24052 37996
rect 23884 37772 24052 37828
rect 23772 37762 23828 37772
rect 23772 36482 23828 36494
rect 23772 36430 23774 36482
rect 23826 36430 23828 36482
rect 23772 36372 23828 36430
rect 23772 36316 23940 36372
rect 23772 36036 23828 36046
rect 23772 35810 23828 35980
rect 23772 35758 23774 35810
rect 23826 35758 23828 35810
rect 23772 35746 23828 35758
rect 23660 35420 23828 35476
rect 23772 33348 23828 35420
rect 23884 34804 23940 36316
rect 23996 36148 24052 37772
rect 24220 36596 24276 37996
rect 24332 37828 24388 37838
rect 24332 37826 24500 37828
rect 24332 37774 24334 37826
rect 24386 37774 24500 37826
rect 24332 37772 24500 37774
rect 24332 37762 24388 37772
rect 24444 37268 24500 37772
rect 24220 36530 24276 36540
rect 24332 36820 24388 36830
rect 24108 36484 24164 36494
rect 24108 36390 24164 36428
rect 24332 36482 24388 36764
rect 24332 36430 24334 36482
rect 24386 36430 24388 36482
rect 24332 36418 24388 36430
rect 24220 36260 24276 36270
rect 24444 36260 24500 37212
rect 24220 36166 24276 36204
rect 24332 36258 24500 36260
rect 24332 36206 24446 36258
rect 24498 36206 24500 36258
rect 24332 36204 24500 36206
rect 23996 36092 24164 36148
rect 23996 35812 24052 35822
rect 23996 35718 24052 35756
rect 24108 35588 24164 36092
rect 24332 35924 24388 36204
rect 24444 36194 24500 36204
rect 24556 35924 24612 38332
rect 24668 38052 24724 38780
rect 25004 38612 25060 38622
rect 24780 38052 24836 38062
rect 24668 38050 24836 38052
rect 24668 37998 24782 38050
rect 24834 37998 24836 38050
rect 24668 37996 24836 37998
rect 23884 34738 23940 34748
rect 23996 35532 24164 35588
rect 24220 35868 24388 35924
rect 24444 35868 24612 35924
rect 24668 36484 24724 36494
rect 24668 35922 24724 36428
rect 24668 35870 24670 35922
rect 24722 35870 24724 35922
rect 23772 33292 23940 33348
rect 23548 33282 23604 33292
rect 23100 32674 23380 32676
rect 23100 32622 23102 32674
rect 23154 32622 23380 32674
rect 23100 32620 23380 32622
rect 23100 32610 23156 32620
rect 22988 32386 23044 32396
rect 23212 32338 23268 32350
rect 23212 32286 23214 32338
rect 23266 32286 23268 32338
rect 23212 32228 23268 32286
rect 22876 32172 23268 32228
rect 23212 31778 23268 32172
rect 23324 31892 23380 32620
rect 23324 31826 23380 31836
rect 23548 33122 23604 33134
rect 23548 33070 23550 33122
rect 23602 33070 23604 33122
rect 23548 33012 23604 33070
rect 23212 31726 23214 31778
rect 23266 31726 23268 31778
rect 23212 31714 23268 31726
rect 22316 31612 22932 31668
rect 22652 31218 22708 31230
rect 22652 31166 22654 31218
rect 22706 31166 22708 31218
rect 22316 30996 22372 31006
rect 22204 30994 22372 30996
rect 22204 30942 22318 30994
rect 22370 30942 22372 30994
rect 22204 30940 22372 30942
rect 22316 30930 22372 30940
rect 22652 30996 22708 31166
rect 22652 30930 22708 30940
rect 22876 30994 22932 31612
rect 23324 31666 23380 31678
rect 23324 31614 23326 31666
rect 23378 31614 23380 31666
rect 23324 31220 23380 31614
rect 23548 31556 23604 32956
rect 23660 33122 23716 33134
rect 23660 33070 23662 33122
rect 23714 33070 23716 33122
rect 23660 32674 23716 33070
rect 23772 33124 23828 33134
rect 23772 33030 23828 33068
rect 23772 32788 23828 32798
rect 23884 32788 23940 33292
rect 23772 32786 23940 32788
rect 23772 32734 23774 32786
rect 23826 32734 23940 32786
rect 23772 32732 23940 32734
rect 23772 32722 23828 32732
rect 23660 32622 23662 32674
rect 23714 32622 23716 32674
rect 23660 32610 23716 32622
rect 23884 31892 23940 31902
rect 23660 31556 23716 31566
rect 23548 31554 23716 31556
rect 23548 31502 23662 31554
rect 23714 31502 23716 31554
rect 23548 31500 23716 31502
rect 23324 31106 23380 31164
rect 23324 31054 23326 31106
rect 23378 31054 23380 31106
rect 23324 31042 23380 31054
rect 22876 30942 22878 30994
rect 22930 30942 22932 30994
rect 22876 30930 22932 30942
rect 23436 30996 23492 31006
rect 23436 30902 23492 30940
rect 23100 30884 23156 30894
rect 22988 30882 23156 30884
rect 22988 30830 23102 30882
rect 23154 30830 23156 30882
rect 22988 30828 23156 30830
rect 22540 30772 22596 30782
rect 22428 30770 22596 30772
rect 22428 30718 22542 30770
rect 22594 30718 22596 30770
rect 22428 30716 22596 30718
rect 22428 30548 22484 30716
rect 22540 30706 22596 30716
rect 22204 30492 22484 30548
rect 22204 30212 22260 30492
rect 22988 30436 23044 30828
rect 23100 30818 23156 30828
rect 22316 30380 23044 30436
rect 22316 30322 22372 30380
rect 22316 30270 22318 30322
rect 22370 30270 22372 30322
rect 22316 30258 22372 30270
rect 22204 30146 22260 30156
rect 23660 29652 23716 31500
rect 23884 31106 23940 31836
rect 23884 31054 23886 31106
rect 23938 31054 23940 31106
rect 23884 31042 23940 31054
rect 23660 29586 23716 29596
rect 23996 29428 24052 35532
rect 24220 34580 24276 35868
rect 24332 35700 24388 35710
rect 24332 35474 24388 35644
rect 24332 35422 24334 35474
rect 24386 35422 24388 35474
rect 24332 34804 24388 35422
rect 24444 35252 24500 35868
rect 24668 35700 24724 35870
rect 24668 35634 24724 35644
rect 24780 35588 24836 37996
rect 25004 37940 25060 38556
rect 25564 38052 25620 38062
rect 25564 37958 25620 37996
rect 26236 37940 26292 37950
rect 25004 37938 25396 37940
rect 25004 37886 25006 37938
rect 25058 37886 25396 37938
rect 25004 37884 25396 37886
rect 25004 37874 25060 37884
rect 25340 37492 25396 37884
rect 26124 37938 26292 37940
rect 26124 37886 26238 37938
rect 26290 37886 26292 37938
rect 26124 37884 26292 37886
rect 25340 37398 25396 37436
rect 26012 37492 26068 37502
rect 25900 37380 25956 37390
rect 25900 37286 25956 37324
rect 26012 37378 26068 37436
rect 26012 37326 26014 37378
rect 26066 37326 26068 37378
rect 26012 37314 26068 37326
rect 25676 37268 25732 37278
rect 25676 37174 25732 37212
rect 26012 37156 26068 37166
rect 26124 37156 26180 37884
rect 26236 37874 26292 37884
rect 26460 37266 26516 40126
rect 26572 39844 26628 39854
rect 26796 39844 26852 39854
rect 26628 39842 26852 39844
rect 26628 39790 26798 39842
rect 26850 39790 26852 39842
rect 26628 39788 26852 39790
rect 26572 39778 26628 39788
rect 26796 39778 26852 39788
rect 26908 39732 26964 39742
rect 26908 39638 26964 39676
rect 27020 39396 27076 40236
rect 27356 40290 27412 40684
rect 27356 40238 27358 40290
rect 27410 40238 27412 40290
rect 27356 40226 27412 40238
rect 27692 40290 27748 40302
rect 27692 40238 27694 40290
rect 27746 40238 27748 40290
rect 27692 39732 27748 40238
rect 27692 39666 27748 39676
rect 27020 39330 27076 39340
rect 28140 38668 28196 43652
rect 28252 43652 28420 43708
rect 28924 43698 28980 43708
rect 28252 41076 28308 43652
rect 28364 43538 28420 43550
rect 28364 43486 28366 43538
rect 28418 43486 28420 43538
rect 28364 43428 28420 43486
rect 28812 43540 28868 43550
rect 28812 43446 28868 43484
rect 28364 43362 28420 43372
rect 28252 41010 28308 41020
rect 28700 43314 28756 43326
rect 28700 43262 28702 43314
rect 28754 43262 28756 43314
rect 28700 42756 28756 43262
rect 28700 40292 28756 42700
rect 29148 42866 29204 42878
rect 29148 42814 29150 42866
rect 29202 42814 29204 42866
rect 29148 42644 29204 42814
rect 29148 42578 29204 42588
rect 29260 42308 29316 45838
rect 32284 45890 32340 45902
rect 32284 45838 32286 45890
rect 32338 45838 32340 45890
rect 29708 45332 29764 45342
rect 29708 45238 29764 45276
rect 30492 45220 30548 45230
rect 30828 45220 30884 45230
rect 30492 45218 30772 45220
rect 30492 45166 30494 45218
rect 30546 45166 30772 45218
rect 30492 45164 30772 45166
rect 30492 45154 30548 45164
rect 29372 45108 29428 45118
rect 29372 45014 29428 45052
rect 30268 45108 30324 45118
rect 30268 45106 30436 45108
rect 30268 45054 30270 45106
rect 30322 45054 30436 45106
rect 30268 45052 30436 45054
rect 30268 45042 30324 45052
rect 29596 44100 29652 44110
rect 29932 44100 29988 44110
rect 29596 44098 29988 44100
rect 29596 44046 29598 44098
rect 29650 44046 29934 44098
rect 29986 44046 29988 44098
rect 29596 44044 29988 44046
rect 29596 44034 29652 44044
rect 29932 43764 29988 44044
rect 30380 44100 30436 45052
rect 30604 44996 30660 45006
rect 30380 44006 30436 44044
rect 30492 44940 30604 44996
rect 29932 43698 29988 43708
rect 30380 43652 30436 43662
rect 30492 43652 30548 44940
rect 30604 44930 30660 44940
rect 30380 43650 30548 43652
rect 30380 43598 30382 43650
rect 30434 43598 30548 43650
rect 30380 43596 30548 43598
rect 30380 43586 30436 43596
rect 28700 40226 28756 40236
rect 29036 42252 29316 42308
rect 27916 38612 28196 38668
rect 27804 38164 27860 38174
rect 27692 37380 27748 37390
rect 27692 37286 27748 37324
rect 27804 37378 27860 38108
rect 27804 37326 27806 37378
rect 27858 37326 27860 37378
rect 27804 37314 27860 37326
rect 26460 37214 26462 37266
rect 26514 37214 26516 37266
rect 26460 37202 26516 37214
rect 26012 37154 26180 37156
rect 26012 37102 26014 37154
rect 26066 37102 26180 37154
rect 26012 37100 26180 37102
rect 26012 37090 26068 37100
rect 25676 36596 25732 36606
rect 25676 36594 25844 36596
rect 25676 36542 25678 36594
rect 25730 36542 25844 36594
rect 25676 36540 25844 36542
rect 25676 36530 25732 36540
rect 24892 36372 24948 36382
rect 24892 35812 24948 36316
rect 24892 35746 24948 35756
rect 25788 35924 25844 36540
rect 27804 36372 27860 36382
rect 27132 36370 27860 36372
rect 27132 36318 27806 36370
rect 27858 36318 27860 36370
rect 27132 36316 27860 36318
rect 25564 35700 25620 35710
rect 25564 35606 25620 35644
rect 25788 35698 25844 35868
rect 27020 35924 27076 35934
rect 25788 35646 25790 35698
rect 25842 35646 25844 35698
rect 25788 35634 25844 35646
rect 26124 35812 26180 35822
rect 24780 35532 25172 35588
rect 24556 35476 24612 35486
rect 24556 35474 25060 35476
rect 24556 35422 24558 35474
rect 24610 35422 25060 35474
rect 24556 35420 25060 35422
rect 24556 35410 24612 35420
rect 24444 35196 24836 35252
rect 24668 34804 24724 34814
rect 24332 34802 24724 34804
rect 24332 34750 24670 34802
rect 24722 34750 24724 34802
rect 24332 34748 24724 34750
rect 24668 34738 24724 34748
rect 24780 34580 24836 35196
rect 24220 34514 24276 34524
rect 24556 34524 24836 34580
rect 24892 34914 24948 34926
rect 24892 34862 24894 34914
rect 24946 34862 24948 34914
rect 24556 33570 24612 34524
rect 24556 33518 24558 33570
rect 24610 33518 24612 33570
rect 24556 33506 24612 33518
rect 24108 33348 24164 33358
rect 24164 33292 24612 33348
rect 24108 32562 24164 33292
rect 24556 33234 24612 33292
rect 24556 33182 24558 33234
rect 24610 33182 24612 33234
rect 24556 33170 24612 33182
rect 24668 33234 24724 33246
rect 24668 33182 24670 33234
rect 24722 33182 24724 33234
rect 24668 32564 24724 33182
rect 24108 32510 24110 32562
rect 24162 32510 24164 32562
rect 24108 32498 24164 32510
rect 24556 32508 24724 32564
rect 24332 32452 24388 32462
rect 24556 32452 24612 32508
rect 24388 32396 24612 32452
rect 24332 32340 24388 32396
rect 24108 32338 24388 32340
rect 24108 32286 24334 32338
rect 24386 32286 24388 32338
rect 24108 32284 24388 32286
rect 24108 30882 24164 32284
rect 24332 32274 24388 32284
rect 24668 32340 24724 32350
rect 24892 32340 24948 34862
rect 25004 33236 25060 35420
rect 25116 33460 25172 35532
rect 25900 35252 25956 35262
rect 25900 34914 25956 35196
rect 25900 34862 25902 34914
rect 25954 34862 25956 34914
rect 25900 34850 25956 34862
rect 25116 33394 25172 33404
rect 25900 33460 25956 33470
rect 25004 33142 25060 33180
rect 25340 33236 25396 33246
rect 25676 33236 25732 33246
rect 25340 33234 25732 33236
rect 25340 33182 25342 33234
rect 25394 33182 25678 33234
rect 25730 33182 25732 33234
rect 25340 33180 25732 33182
rect 25340 33170 25396 33180
rect 25228 33124 25284 33134
rect 25228 32562 25284 33068
rect 25676 32788 25732 33180
rect 25788 32788 25844 32798
rect 25676 32786 25844 32788
rect 25676 32734 25790 32786
rect 25842 32734 25844 32786
rect 25676 32732 25844 32734
rect 25788 32722 25844 32732
rect 25228 32510 25230 32562
rect 25282 32510 25284 32562
rect 25228 32498 25284 32510
rect 25452 32452 25508 32462
rect 25452 32358 25508 32396
rect 24724 32284 24948 32340
rect 25340 32340 25396 32350
rect 24668 32246 24724 32284
rect 24780 32116 24836 32126
rect 24556 31220 24612 31230
rect 24556 31126 24612 31164
rect 24220 30996 24276 31006
rect 24668 30996 24724 31006
rect 24220 30994 24724 30996
rect 24220 30942 24222 30994
rect 24274 30942 24670 30994
rect 24722 30942 24724 30994
rect 24220 30940 24724 30942
rect 24220 30930 24276 30940
rect 24108 30830 24110 30882
rect 24162 30830 24164 30882
rect 24108 30818 24164 30830
rect 24444 30322 24500 30940
rect 24668 30930 24724 30940
rect 24444 30270 24446 30322
rect 24498 30270 24500 30322
rect 24444 30258 24500 30270
rect 22092 28662 22148 28700
rect 23548 29372 24052 29428
rect 24220 30212 24276 30222
rect 20636 27076 20692 27086
rect 20412 26964 20468 26974
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 18844 26238 18846 26290
rect 18898 26238 18900 26290
rect 18844 26226 18900 26238
rect 18956 26460 19348 26516
rect 18620 24948 18676 24958
rect 18508 24946 18676 24948
rect 18508 24894 18622 24946
rect 18674 24894 18676 24946
rect 18508 24892 18676 24894
rect 18620 24882 18676 24892
rect 16380 24558 16382 24610
rect 16434 24558 16436 24610
rect 16380 24546 16436 24558
rect 15932 23886 15934 23938
rect 15986 23886 15988 23938
rect 15596 23716 15652 23726
rect 15596 23622 15652 23660
rect 15932 23548 15988 23886
rect 15820 23492 15988 23548
rect 18396 23716 18452 23726
rect 15820 23044 15876 23492
rect 17388 23436 17780 23492
rect 15820 22978 15876 22988
rect 16828 23044 16884 23054
rect 16828 22950 16884 22988
rect 17388 21698 17444 23436
rect 17612 23268 17668 23278
rect 17724 23268 17780 23436
rect 18060 23380 18116 23390
rect 18396 23380 18452 23660
rect 18116 23324 18452 23380
rect 18844 23380 18900 23390
rect 18060 23286 18116 23324
rect 18844 23286 18900 23324
rect 17836 23268 17892 23278
rect 17724 23266 17892 23268
rect 17724 23214 17838 23266
rect 17890 23214 17892 23266
rect 17724 23212 17892 23214
rect 17612 22372 17668 23212
rect 17836 23202 17892 23212
rect 18508 23266 18564 23278
rect 18508 23214 18510 23266
rect 18562 23214 18564 23266
rect 18172 22932 18228 22942
rect 18172 22930 18340 22932
rect 18172 22878 18174 22930
rect 18226 22878 18340 22930
rect 18172 22876 18340 22878
rect 18172 22866 18228 22876
rect 18284 22482 18340 22876
rect 18284 22430 18286 22482
rect 18338 22430 18340 22482
rect 18284 22418 18340 22430
rect 17612 22370 18116 22372
rect 17612 22318 17614 22370
rect 17666 22318 18116 22370
rect 17612 22316 18116 22318
rect 17612 22306 17668 22316
rect 17388 21646 17390 21698
rect 17442 21646 17444 21698
rect 17388 21634 17444 21646
rect 17836 21588 17892 21598
rect 17500 21586 17892 21588
rect 17500 21534 17838 21586
rect 17890 21534 17892 21586
rect 17500 21532 17892 21534
rect 15708 20916 15764 20926
rect 15708 20822 15764 20860
rect 16156 20804 16212 20814
rect 16156 20710 16212 20748
rect 16604 20804 16660 20814
rect 15260 17838 15262 17890
rect 15314 17838 15316 17890
rect 15260 16772 15316 17838
rect 15260 15988 15316 16716
rect 15372 20188 15540 20244
rect 15372 16548 15428 20188
rect 15484 20020 15540 20030
rect 15484 19926 15540 19964
rect 16604 19908 16660 20748
rect 16716 20692 16772 20702
rect 16716 20598 16772 20636
rect 17500 20356 17556 21532
rect 17836 21522 17892 21532
rect 17836 20804 17892 20814
rect 17836 20710 17892 20748
rect 16828 20300 17556 20356
rect 17724 20690 17780 20702
rect 17724 20638 17726 20690
rect 17778 20638 17780 20690
rect 16828 20242 16884 20300
rect 16828 20190 16830 20242
rect 16882 20190 16884 20242
rect 16828 20178 16884 20190
rect 16716 19908 16772 19918
rect 16604 19906 16772 19908
rect 16604 19854 16718 19906
rect 16770 19854 16772 19906
rect 16604 19852 16772 19854
rect 15820 19348 15876 19358
rect 15820 17666 15876 19292
rect 16268 17780 16324 17790
rect 16604 17780 16660 19852
rect 16716 19842 16772 19852
rect 16828 18452 16884 18462
rect 16828 17780 16884 18396
rect 16268 17778 16660 17780
rect 16268 17726 16270 17778
rect 16322 17726 16660 17778
rect 16268 17724 16660 17726
rect 16716 17724 16884 17780
rect 16268 17714 16324 17724
rect 15820 17614 15822 17666
rect 15874 17614 15876 17666
rect 15820 17602 15876 17614
rect 16044 17668 16100 17678
rect 16044 17666 16212 17668
rect 16044 17614 16046 17666
rect 16098 17614 16212 17666
rect 16044 17612 16212 17614
rect 16044 17602 16100 17612
rect 15596 17554 15652 17566
rect 15596 17502 15598 17554
rect 15650 17502 15652 17554
rect 15484 16772 15540 16782
rect 15484 16678 15540 16716
rect 15372 16492 15540 16548
rect 15372 16100 15428 16110
rect 15372 16006 15428 16044
rect 14476 15810 14532 15820
rect 14700 15820 14868 15876
rect 14924 15876 14980 15886
rect 14924 15874 15204 15876
rect 14924 15822 14926 15874
rect 14978 15822 15204 15874
rect 14924 15820 15204 15822
rect 14700 15428 14756 15820
rect 14924 15810 14980 15820
rect 14476 15372 14756 15428
rect 14812 15652 14868 15662
rect 14476 15148 14532 15372
rect 14700 15202 14756 15214
rect 14700 15150 14702 15202
rect 14754 15150 14756 15202
rect 14476 15092 14644 15148
rect 14364 14802 14420 14812
rect 14476 14644 14532 14654
rect 14252 14578 14308 14588
rect 14364 14588 14476 14644
rect 14140 13918 14142 13970
rect 14194 13918 14196 13970
rect 14140 13906 14196 13918
rect 14364 12516 14420 14588
rect 14476 14578 14532 14588
rect 14476 14418 14532 14430
rect 14476 14366 14478 14418
rect 14530 14366 14532 14418
rect 14476 13636 14532 14366
rect 14588 13860 14644 15092
rect 14700 14980 14756 15150
rect 14700 14914 14756 14924
rect 14812 14756 14868 15596
rect 15148 15538 15204 15820
rect 15260 15764 15316 15932
rect 15484 15986 15540 16492
rect 15484 15934 15486 15986
rect 15538 15934 15540 15986
rect 15484 15922 15540 15934
rect 15260 15708 15540 15764
rect 15148 15486 15150 15538
rect 15202 15486 15204 15538
rect 15148 15148 15204 15486
rect 15484 15316 15540 15708
rect 15596 15652 15652 17502
rect 15932 17442 15988 17454
rect 15932 17390 15934 17442
rect 15986 17390 15988 17442
rect 15932 17220 15988 17390
rect 15820 17164 15988 17220
rect 15820 16772 15876 17164
rect 16044 17108 16100 17118
rect 16156 17108 16212 17612
rect 16492 17556 16548 17566
rect 16492 17554 16660 17556
rect 16492 17502 16494 17554
rect 16546 17502 16660 17554
rect 16492 17500 16660 17502
rect 16492 17490 16548 17500
rect 16044 17106 16548 17108
rect 16044 17054 16046 17106
rect 16098 17054 16548 17106
rect 16044 17052 16548 17054
rect 16044 17042 16100 17052
rect 15820 16706 15876 16716
rect 15932 16996 15988 17006
rect 15596 15586 15652 15596
rect 15932 15428 15988 16940
rect 16492 16994 16548 17052
rect 16492 16942 16494 16994
rect 16546 16942 16548 16994
rect 16492 16930 16548 16942
rect 16156 16884 16212 16894
rect 16156 16790 16212 16828
rect 16156 16212 16212 16222
rect 16604 16212 16660 17500
rect 16716 16770 16772 17724
rect 16940 17668 16996 20300
rect 17724 20132 17780 20638
rect 17164 19348 17220 19358
rect 17724 19348 17780 20076
rect 17164 19346 17780 19348
rect 17164 19294 17166 19346
rect 17218 19294 17780 19346
rect 17164 19292 17780 19294
rect 18060 20018 18116 22316
rect 18284 21474 18340 21486
rect 18284 21422 18286 21474
rect 18338 21422 18340 21474
rect 18284 20804 18340 21422
rect 18508 21252 18564 23214
rect 18508 21186 18564 21196
rect 18732 21362 18788 21374
rect 18732 21310 18734 21362
rect 18786 21310 18788 21362
rect 18284 20738 18340 20748
rect 18732 20132 18788 21310
rect 18844 21362 18900 21374
rect 18844 21310 18846 21362
rect 18898 21310 18900 21362
rect 18844 21252 18900 21310
rect 18844 21186 18900 21196
rect 18844 20132 18900 20142
rect 18732 20130 18900 20132
rect 18732 20078 18846 20130
rect 18898 20078 18900 20130
rect 18732 20076 18900 20078
rect 18844 20066 18900 20076
rect 18060 19966 18062 20018
rect 18114 19966 18116 20018
rect 17164 19282 17220 19292
rect 17052 19012 17108 19022
rect 17612 19012 17668 19022
rect 17052 19010 17332 19012
rect 17052 18958 17054 19010
rect 17106 18958 17332 19010
rect 17052 18956 17332 18958
rect 17052 18946 17108 18956
rect 17276 17780 17332 18956
rect 17612 18562 17668 18956
rect 17612 18510 17614 18562
rect 17666 18510 17668 18562
rect 17612 18498 17668 18510
rect 17388 18452 17444 18462
rect 17388 18358 17444 18396
rect 17948 18450 18004 18462
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17836 18340 17892 18350
rect 17836 18246 17892 18284
rect 17276 17724 17444 17780
rect 17052 17668 17108 17678
rect 16940 17666 17108 17668
rect 16940 17614 17054 17666
rect 17106 17614 17108 17666
rect 16940 17612 17108 17614
rect 17052 17602 17108 17612
rect 17388 17668 17444 17724
rect 17388 17666 17668 17668
rect 17388 17614 17390 17666
rect 17442 17614 17668 17666
rect 17388 17612 17668 17614
rect 17388 17602 17444 17612
rect 16828 17556 16884 17566
rect 16828 17554 16996 17556
rect 16828 17502 16830 17554
rect 16882 17502 16996 17554
rect 16828 17500 16996 17502
rect 16828 17490 16884 17500
rect 16828 17108 16884 17118
rect 16828 16882 16884 17052
rect 16940 16996 16996 17500
rect 17164 17442 17220 17454
rect 17164 17390 17166 17442
rect 17218 17390 17220 17442
rect 17164 17108 17220 17390
rect 16940 16940 17108 16996
rect 16828 16830 16830 16882
rect 16882 16830 16884 16882
rect 16828 16818 16884 16830
rect 16716 16718 16718 16770
rect 16770 16718 16772 16770
rect 16716 16706 16772 16718
rect 17052 16324 17108 16940
rect 17164 16772 17220 17052
rect 17276 17442 17332 17454
rect 17276 17390 17278 17442
rect 17330 17390 17332 17442
rect 17276 16996 17332 17390
rect 17276 16930 17332 16940
rect 17500 16884 17556 16894
rect 17388 16882 17556 16884
rect 17388 16830 17502 16882
rect 17554 16830 17556 16882
rect 17388 16828 17556 16830
rect 17388 16772 17444 16828
rect 17500 16818 17556 16828
rect 17612 16884 17668 17612
rect 17948 17108 18004 18398
rect 18060 18452 18116 19966
rect 18060 18386 18116 18396
rect 18060 17108 18116 17118
rect 17948 17106 18116 17108
rect 17948 17054 18062 17106
rect 18114 17054 18116 17106
rect 17948 17052 18116 17054
rect 18060 17042 18116 17052
rect 17612 16818 17668 16828
rect 17164 16716 17444 16772
rect 17724 16772 17780 16782
rect 17724 16678 17780 16716
rect 17500 16660 17556 16670
rect 17556 16604 17668 16660
rect 17500 16594 17556 16604
rect 16828 16268 17108 16324
rect 16604 16156 16772 16212
rect 16156 16118 16212 16156
rect 16380 16098 16436 16110
rect 16380 16046 16382 16098
rect 16434 16046 16436 16098
rect 16156 15986 16212 15998
rect 16156 15934 16158 15986
rect 16210 15934 16212 15986
rect 16156 15540 16212 15934
rect 16156 15474 16212 15484
rect 15932 15362 15988 15372
rect 15484 15222 15540 15260
rect 16156 15316 16212 15326
rect 15708 15204 15764 15242
rect 16156 15222 16212 15260
rect 16380 15148 16436 16046
rect 15148 15092 15316 15148
rect 15708 15138 15764 15148
rect 14588 13794 14644 13804
rect 14700 14700 14868 14756
rect 14700 13636 14756 14700
rect 15260 14642 15316 15092
rect 15260 14590 15262 14642
rect 15314 14590 15316 14642
rect 15260 14578 15316 14590
rect 16156 15092 16436 15148
rect 16604 15428 16660 15438
rect 14476 13580 14756 13636
rect 14812 14532 14868 14542
rect 14476 12962 14532 13580
rect 14812 13524 14868 14476
rect 15484 14530 15540 14542
rect 15484 14478 15486 14530
rect 15538 14478 15540 14530
rect 15484 14196 15540 14478
rect 15820 14308 15876 14318
rect 15820 14306 15988 14308
rect 15820 14254 15822 14306
rect 15874 14254 15988 14306
rect 15820 14252 15988 14254
rect 15820 14242 15876 14252
rect 15484 14130 15540 14140
rect 14476 12910 14478 12962
rect 14530 12910 14532 12962
rect 14476 12740 14532 12910
rect 14700 12964 14756 12974
rect 14700 12870 14756 12908
rect 14476 12684 14756 12740
rect 14364 12450 14420 12460
rect 14028 12178 14084 12348
rect 14588 12292 14644 12302
rect 14028 12126 14030 12178
rect 14082 12126 14084 12178
rect 14028 12114 14084 12126
rect 14476 12290 14644 12292
rect 14476 12238 14590 12290
rect 14642 12238 14644 12290
rect 14476 12236 14644 12238
rect 14364 12068 14420 12078
rect 13916 12002 13972 12012
rect 14140 12066 14420 12068
rect 14140 12014 14366 12066
rect 14418 12014 14420 12066
rect 14140 12012 14420 12014
rect 14140 11844 14196 12012
rect 14364 12002 14420 12012
rect 13468 11618 13636 11620
rect 13468 11566 13470 11618
rect 13522 11566 13636 11618
rect 13468 11564 13636 11566
rect 13692 11788 14196 11844
rect 13468 11554 13524 11564
rect 13692 11394 13748 11788
rect 13692 11342 13694 11394
rect 13746 11342 13748 11394
rect 13692 11330 13748 11342
rect 14252 11396 14308 11406
rect 14252 11302 14308 11340
rect 13804 11284 13860 11294
rect 13804 11190 13860 11228
rect 13356 10658 13412 10668
rect 13916 11060 13972 11070
rect 12908 9828 12964 9838
rect 12908 9734 12964 9772
rect 13916 9826 13972 11004
rect 14476 10948 14532 12236
rect 14588 12226 14644 12236
rect 14700 12180 14756 12684
rect 14700 12114 14756 12124
rect 13916 9774 13918 9826
rect 13970 9774 13972 9826
rect 12796 9268 12852 9548
rect 12908 9268 12964 9278
rect 12796 9266 12964 9268
rect 12796 9214 12910 9266
rect 12962 9214 12964 9266
rect 12796 9212 12964 9214
rect 12460 8932 12516 8942
rect 12348 8930 12516 8932
rect 12348 8878 12462 8930
rect 12514 8878 12516 8930
rect 12348 8876 12516 8878
rect 12460 8866 12516 8876
rect 12348 7700 12404 7710
rect 12348 7606 12404 7644
rect 12796 7588 12852 9212
rect 12908 9202 12964 9212
rect 13580 8372 13636 8382
rect 13020 7700 13076 7710
rect 13580 7700 13636 8316
rect 12796 7532 12964 7588
rect 12684 7476 12740 7486
rect 12684 7382 12740 7420
rect 12236 7364 12292 7374
rect 12236 7362 12628 7364
rect 12236 7310 12238 7362
rect 12290 7310 12628 7362
rect 12236 7308 12628 7310
rect 12236 7298 12292 7308
rect 12236 6468 12292 6478
rect 12236 6374 12292 6412
rect 12572 5460 12628 7308
rect 12796 7362 12852 7374
rect 12796 7310 12798 7362
rect 12850 7310 12852 7362
rect 12796 6580 12852 7310
rect 12908 6692 12964 7532
rect 13020 7586 13076 7644
rect 13020 7534 13022 7586
rect 13074 7534 13076 7586
rect 13020 7522 13076 7534
rect 13468 7698 13636 7700
rect 13468 7646 13582 7698
rect 13634 7646 13636 7698
rect 13468 7644 13636 7646
rect 13132 7476 13188 7486
rect 13132 7382 13188 7420
rect 12908 6598 12964 6636
rect 13244 6804 13300 6814
rect 12796 6514 12852 6524
rect 12572 5404 12964 5460
rect 12460 5124 12516 5134
rect 12460 5030 12516 5068
rect 12572 5012 12628 5022
rect 12572 4918 12628 4956
rect 12348 4898 12404 4910
rect 12348 4846 12350 4898
rect 12402 4846 12404 4898
rect 12348 4788 12404 4846
rect 12908 4900 12964 5404
rect 13020 5124 13076 5134
rect 13244 5124 13300 6748
rect 13468 6356 13524 7644
rect 13580 7634 13636 7644
rect 13804 7700 13860 7710
rect 13804 7606 13860 7644
rect 13692 7476 13748 7486
rect 13692 7382 13748 7420
rect 13580 6692 13636 6702
rect 13580 6598 13636 6636
rect 13468 6290 13524 6300
rect 13020 5122 13300 5124
rect 13020 5070 13022 5122
rect 13074 5070 13300 5122
rect 13020 5068 13300 5070
rect 13020 5058 13076 5068
rect 13692 4900 13748 4910
rect 12908 4844 13188 4900
rect 12348 4722 12404 4732
rect 12348 4228 12404 4238
rect 12348 4134 12404 4172
rect 12124 3502 12126 3554
rect 12178 3502 12180 3554
rect 12124 3490 12180 3502
rect 13132 3442 13188 4844
rect 13468 4898 13748 4900
rect 13468 4846 13694 4898
rect 13746 4846 13748 4898
rect 13468 4844 13748 4846
rect 13356 3556 13412 3566
rect 13468 3556 13524 4844
rect 13692 4834 13748 4844
rect 13804 4788 13860 4798
rect 13916 4788 13972 9774
rect 14252 10892 14532 10948
rect 14588 12068 14644 12078
rect 14252 9828 14308 10892
rect 14588 10836 14644 12012
rect 14812 11732 14868 13468
rect 14924 13076 14980 13086
rect 14924 12962 14980 13020
rect 15596 13076 15652 13086
rect 15260 12964 15316 12974
rect 14924 12910 14926 12962
rect 14978 12910 14980 12962
rect 14924 12898 14980 12910
rect 15148 12908 15260 12964
rect 15148 12850 15204 12908
rect 15260 12898 15316 12908
rect 15148 12798 15150 12850
rect 15202 12798 15204 12850
rect 15148 12786 15204 12798
rect 15036 12740 15092 12750
rect 14924 12738 15092 12740
rect 14924 12686 15038 12738
rect 15090 12686 15092 12738
rect 14924 12684 15092 12686
rect 15596 12740 15652 13020
rect 15708 12964 15764 12974
rect 15708 12870 15764 12908
rect 15932 12962 15988 14252
rect 15932 12910 15934 12962
rect 15986 12910 15988 12962
rect 15820 12852 15876 12862
rect 15820 12758 15876 12796
rect 15596 12684 15764 12740
rect 14924 11732 14980 12684
rect 15036 12674 15092 12684
rect 15036 12180 15092 12190
rect 15036 12086 15092 12124
rect 14924 11676 15540 11732
rect 14812 11666 14868 11676
rect 15036 11396 15092 11406
rect 15036 11302 15092 11340
rect 15484 11394 15540 11676
rect 15484 11342 15486 11394
rect 15538 11342 15540 11394
rect 15484 11330 15540 11342
rect 15596 11172 15652 11182
rect 14700 10836 14756 10846
rect 14588 10834 14756 10836
rect 14588 10782 14702 10834
rect 14754 10782 14756 10834
rect 14588 10780 14756 10782
rect 14700 10770 14756 10780
rect 15596 10834 15652 11116
rect 15708 10948 15764 12684
rect 15932 12292 15988 12910
rect 16156 12402 16212 15092
rect 16380 12740 16436 12750
rect 16380 12646 16436 12684
rect 16156 12350 16158 12402
rect 16210 12350 16212 12402
rect 16156 12338 16212 12350
rect 16268 12404 16324 12414
rect 15932 12226 15988 12236
rect 15820 12178 15876 12190
rect 15820 12126 15822 12178
rect 15874 12126 15876 12178
rect 15820 11394 15876 12126
rect 15820 11342 15822 11394
rect 15874 11342 15876 11394
rect 15820 11330 15876 11342
rect 16044 12178 16100 12190
rect 16044 12126 16046 12178
rect 16098 12126 16100 12178
rect 16044 11396 16100 12126
rect 16156 11508 16212 11518
rect 16268 11508 16324 12348
rect 16492 12178 16548 12190
rect 16492 12126 16494 12178
rect 16546 12126 16548 12178
rect 16156 11506 16324 11508
rect 16156 11454 16158 11506
rect 16210 11454 16324 11506
rect 16156 11452 16324 11454
rect 16380 11732 16436 11742
rect 16156 11442 16212 11452
rect 16044 10948 16100 11340
rect 15708 10892 15876 10948
rect 16044 10892 16212 10948
rect 15596 10782 15598 10834
rect 15650 10782 15652 10834
rect 15596 10770 15652 10782
rect 14476 10722 14532 10734
rect 14476 10670 14478 10722
rect 14530 10670 14532 10722
rect 14364 10610 14420 10622
rect 14364 10558 14366 10610
rect 14418 10558 14420 10610
rect 14364 9938 14420 10558
rect 14476 10052 14532 10670
rect 15148 10722 15204 10734
rect 15148 10670 15150 10722
rect 15202 10670 15204 10722
rect 14476 9996 14980 10052
rect 14364 9886 14366 9938
rect 14418 9886 14420 9938
rect 14364 9874 14420 9886
rect 14252 9762 14308 9772
rect 14476 9828 14532 9838
rect 14028 9604 14084 9614
rect 14028 9510 14084 9548
rect 14252 9602 14308 9614
rect 14252 9550 14254 9602
rect 14306 9550 14308 9602
rect 14252 9268 14308 9550
rect 14252 9202 14308 9212
rect 14364 9492 14420 9502
rect 14364 9266 14420 9436
rect 14364 9214 14366 9266
rect 14418 9214 14420 9266
rect 14364 9202 14420 9214
rect 14252 9044 14308 9054
rect 14476 9044 14532 9772
rect 14812 9154 14868 9996
rect 14924 9938 14980 9996
rect 15148 9940 15204 10670
rect 15708 10724 15764 10734
rect 15708 10610 15764 10668
rect 15708 10558 15710 10610
rect 15762 10558 15764 10610
rect 14924 9886 14926 9938
rect 14978 9886 14980 9938
rect 14924 9874 14980 9886
rect 15036 9884 15428 9940
rect 15036 9826 15092 9884
rect 15036 9774 15038 9826
rect 15090 9774 15092 9826
rect 15036 9762 15092 9774
rect 14924 9716 14980 9726
rect 14924 9622 14980 9660
rect 15260 9602 15316 9614
rect 15260 9550 15262 9602
rect 15314 9550 15316 9602
rect 15260 9492 15316 9550
rect 15260 9426 15316 9436
rect 15372 9266 15428 9884
rect 15484 9716 15540 9726
rect 15484 9714 15652 9716
rect 15484 9662 15486 9714
rect 15538 9662 15652 9714
rect 15484 9660 15652 9662
rect 15484 9650 15540 9660
rect 15372 9214 15374 9266
rect 15426 9214 15428 9266
rect 15372 9202 15428 9214
rect 15484 9268 15540 9278
rect 14812 9102 14814 9154
rect 14866 9102 14868 9154
rect 14812 9090 14868 9102
rect 14252 9042 14532 9044
rect 14252 8990 14254 9042
rect 14306 8990 14532 9042
rect 14252 8988 14532 8990
rect 14588 9042 14644 9054
rect 14588 8990 14590 9042
rect 14642 8990 14644 9042
rect 14252 8978 14308 8988
rect 14588 8372 14644 8990
rect 15484 8930 15540 9212
rect 15484 8878 15486 8930
rect 15538 8878 15540 8930
rect 14588 7700 14644 8316
rect 14588 7634 14644 7644
rect 15148 8372 15204 8382
rect 15148 7698 15204 8316
rect 15148 7646 15150 7698
rect 15202 7646 15204 7698
rect 15148 7634 15204 7646
rect 14028 7586 14084 7598
rect 14028 7534 14030 7586
rect 14082 7534 14084 7586
rect 14028 7476 14084 7534
rect 14028 6804 14084 7420
rect 15484 7474 15540 8878
rect 15596 8708 15652 9660
rect 15708 9492 15764 10558
rect 15820 10612 15876 10892
rect 16044 10612 16100 10622
rect 15820 10610 16100 10612
rect 15820 10558 16046 10610
rect 16098 10558 16100 10610
rect 15820 10556 16100 10558
rect 15708 8820 15764 9436
rect 15820 9604 15876 9614
rect 15932 9604 15988 9614
rect 15876 9602 15988 9604
rect 15876 9550 15934 9602
rect 15986 9550 15988 9602
rect 15876 9548 15988 9550
rect 15820 9044 15876 9548
rect 15932 9538 15988 9548
rect 15820 8950 15876 8988
rect 15932 9042 15988 9054
rect 15932 8990 15934 9042
rect 15986 8990 15988 9042
rect 15932 8820 15988 8990
rect 15708 8764 15988 8820
rect 16044 8708 16100 10556
rect 16156 9602 16212 10892
rect 16380 10834 16436 11676
rect 16492 11508 16548 12126
rect 16492 11442 16548 11452
rect 16380 10782 16382 10834
rect 16434 10782 16436 10834
rect 16380 10770 16436 10782
rect 16156 9550 16158 9602
rect 16210 9550 16212 9602
rect 16156 9538 16212 9550
rect 16380 9826 16436 9838
rect 16380 9774 16382 9826
rect 16434 9774 16436 9826
rect 15596 8652 16100 8708
rect 15484 7422 15486 7474
rect 15538 7422 15540 7474
rect 15484 7364 15540 7422
rect 15932 7364 15988 7374
rect 15484 7362 15988 7364
rect 15484 7310 15934 7362
rect 15986 7310 15988 7362
rect 15484 7308 15988 7310
rect 14028 6738 14084 6748
rect 14924 6692 14980 6702
rect 14252 6580 14308 6590
rect 14252 6486 14308 6524
rect 14812 4900 14868 4910
rect 13860 4732 13972 4788
rect 14476 4844 14812 4900
rect 13804 4722 13860 4732
rect 14476 4226 14532 4844
rect 14812 4806 14868 4844
rect 14924 4562 14980 6636
rect 15932 6692 15988 7308
rect 15932 6626 15988 6636
rect 15820 5236 15876 5246
rect 16044 5236 16100 8652
rect 16380 7698 16436 9774
rect 16604 8372 16660 15372
rect 16716 13076 16772 16156
rect 16716 13010 16772 13020
rect 16828 11060 16884 16268
rect 17388 15988 17444 15998
rect 17052 15932 17388 15988
rect 17612 15988 17668 16604
rect 18508 16098 18564 16110
rect 18508 16046 18510 16098
rect 18562 16046 18564 16098
rect 17724 15988 17780 15998
rect 17612 15986 17780 15988
rect 17612 15934 17726 15986
rect 17778 15934 17780 15986
rect 17612 15932 17780 15934
rect 16940 15540 16996 15550
rect 17052 15540 17108 15932
rect 17388 15894 17444 15932
rect 17724 15922 17780 15932
rect 18060 15988 18116 15998
rect 18060 15894 18116 15932
rect 18508 15988 18564 16046
rect 18508 15922 18564 15932
rect 18732 16100 18788 16110
rect 18732 15986 18788 16044
rect 18732 15934 18734 15986
rect 18786 15934 18788 15986
rect 18732 15922 18788 15934
rect 16940 15538 17108 15540
rect 16940 15486 16942 15538
rect 16994 15486 17108 15538
rect 16940 15484 17108 15486
rect 16940 15474 16996 15484
rect 17388 15202 17444 15214
rect 17388 15150 17390 15202
rect 17442 15150 17444 15202
rect 17388 14532 17444 15150
rect 18956 15148 19012 26460
rect 19180 26292 19236 26302
rect 19516 26292 19572 26302
rect 19180 26290 19572 26292
rect 19180 26238 19182 26290
rect 19234 26238 19518 26290
rect 19570 26238 19572 26290
rect 19180 26236 19572 26238
rect 19180 26226 19236 26236
rect 19516 26226 19572 26236
rect 19180 26068 19236 26078
rect 19740 26068 19796 26078
rect 19236 26066 19796 26068
rect 19236 26014 19742 26066
rect 19794 26014 19796 26066
rect 19236 26012 19796 26014
rect 19180 25618 19236 26012
rect 19740 26002 19796 26012
rect 19964 26068 20020 26078
rect 19964 25974 20020 26012
rect 20076 26066 20132 26078
rect 20076 26014 20078 26066
rect 20130 26014 20132 26066
rect 19180 25566 19182 25618
rect 19234 25566 19236 25618
rect 19180 25554 19236 25566
rect 20076 25284 20132 26014
rect 20076 25228 20244 25284
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24836 20244 25228
rect 20188 24770 20244 24780
rect 19852 23940 19908 23950
rect 19852 23846 19908 23884
rect 20412 23940 20468 26908
rect 20412 23846 20468 23884
rect 20524 26178 20580 26190
rect 20524 26126 20526 26178
rect 20578 26126 20580 26178
rect 20524 26068 20580 26126
rect 19292 23716 19348 23726
rect 19180 23660 19292 23716
rect 19068 21362 19124 21374
rect 19068 21310 19070 21362
rect 19122 21310 19124 21362
rect 19068 20916 19124 21310
rect 19068 20850 19124 20860
rect 19180 20468 19236 23660
rect 19292 23650 19348 23660
rect 19628 23716 19684 23726
rect 19628 23622 19684 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20524 23492 20580 26012
rect 19836 23482 20100 23492
rect 20300 23436 20580 23492
rect 19292 23380 19348 23390
rect 19292 23286 19348 23324
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19292 21586 19348 21598
rect 19292 21534 19294 21586
rect 19346 21534 19348 21586
rect 19292 21364 19348 21534
rect 19292 21298 19348 21308
rect 19740 20916 19796 20926
rect 19796 20860 19908 20916
rect 19740 20850 19796 20860
rect 19628 20804 19684 20814
rect 19628 20710 19684 20748
rect 19852 20802 19908 20860
rect 19852 20750 19854 20802
rect 19906 20750 19908 20802
rect 19852 20738 19908 20750
rect 19964 20802 20020 20814
rect 19964 20750 19966 20802
rect 20018 20750 20020 20802
rect 19516 20692 19572 20702
rect 19516 20598 19572 20636
rect 19964 20580 20020 20750
rect 19964 20514 20020 20524
rect 20188 20802 20244 20814
rect 20188 20750 20190 20802
rect 20242 20750 20244 20802
rect 19180 20412 19684 20468
rect 19628 19348 19684 20412
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20132 20244 20750
rect 20188 20066 20244 20076
rect 20300 19908 20356 23436
rect 20524 23268 20580 23278
rect 20524 23154 20580 23212
rect 20524 23102 20526 23154
rect 20578 23102 20580 23154
rect 20524 23090 20580 23102
rect 20524 22146 20580 22158
rect 20524 22094 20526 22146
rect 20578 22094 20580 22146
rect 20412 20580 20468 20590
rect 20524 20580 20580 22094
rect 20468 20524 20580 20580
rect 20412 20514 20468 20524
rect 20524 19908 20580 19918
rect 20188 19852 20356 19908
rect 20412 19852 20524 19908
rect 19628 19346 20020 19348
rect 19628 19294 19630 19346
rect 19682 19294 20020 19346
rect 19628 19292 20020 19294
rect 19628 19282 19684 19292
rect 19964 19234 20020 19292
rect 19964 19182 19966 19234
rect 20018 19182 20020 19234
rect 19964 19170 20020 19182
rect 20188 19236 20244 19852
rect 20300 19460 20356 19470
rect 20412 19460 20468 19852
rect 20524 19842 20580 19852
rect 20300 19458 20468 19460
rect 20300 19406 20302 19458
rect 20354 19406 20468 19458
rect 20300 19404 20468 19406
rect 20300 19394 20356 19404
rect 20188 19180 20468 19236
rect 20188 19010 20244 19022
rect 20188 18958 20190 19010
rect 20242 18958 20244 19010
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20188 18676 20244 18958
rect 20076 18620 20244 18676
rect 20076 18562 20132 18620
rect 20076 18510 20078 18562
rect 20130 18510 20132 18562
rect 20076 18498 20132 18510
rect 19292 18452 19348 18462
rect 19068 17780 19124 17790
rect 19068 16210 19124 17724
rect 19292 17778 19348 18396
rect 19292 17726 19294 17778
rect 19346 17726 19348 17778
rect 19292 17714 19348 17726
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19068 16158 19070 16210
rect 19122 16158 19124 16210
rect 19068 16146 19124 16158
rect 19180 16772 19236 16782
rect 19180 15988 19236 16716
rect 19852 16772 19908 16782
rect 19852 16770 20244 16772
rect 19852 16718 19854 16770
rect 19906 16718 20244 16770
rect 19852 16716 20244 16718
rect 19852 16706 19908 16716
rect 20076 16212 20132 16222
rect 19628 16100 19684 16110
rect 20076 16100 20132 16156
rect 19684 16098 20132 16100
rect 19684 16046 20078 16098
rect 20130 16046 20132 16098
rect 19684 16044 20132 16046
rect 19628 16006 19684 16044
rect 20076 16034 20132 16044
rect 18844 15092 18900 15102
rect 18956 15092 19124 15148
rect 18508 15036 18844 15092
rect 17612 14756 17668 14766
rect 18172 14756 18228 14766
rect 17612 14754 18228 14756
rect 17612 14702 17614 14754
rect 17666 14702 18174 14754
rect 18226 14702 18228 14754
rect 17612 14700 18228 14702
rect 17612 14690 17668 14700
rect 18172 14690 18228 14700
rect 18508 14754 18564 15036
rect 18844 15026 18900 15036
rect 18508 14702 18510 14754
rect 18562 14702 18564 14754
rect 18508 14690 18564 14702
rect 17276 14420 17332 14430
rect 17276 14326 17332 14364
rect 17388 13972 17444 14476
rect 17612 14530 17668 14542
rect 17612 14478 17614 14530
rect 17666 14478 17668 14530
rect 17612 14196 17668 14478
rect 18060 14532 18116 14542
rect 18060 14530 18340 14532
rect 18060 14478 18062 14530
rect 18114 14478 18340 14530
rect 18060 14476 18340 14478
rect 18060 14466 18116 14476
rect 17612 14140 17892 14196
rect 17724 13972 17780 13982
rect 17388 13970 17780 13972
rect 17388 13918 17726 13970
rect 17778 13918 17780 13970
rect 17388 13916 17780 13918
rect 17724 13906 17780 13916
rect 17836 13636 17892 14140
rect 18172 13636 18228 13646
rect 17836 13634 18228 13636
rect 17836 13582 18174 13634
rect 18226 13582 18228 13634
rect 17836 13580 18228 13582
rect 17612 13412 17668 13422
rect 17500 13300 17556 13310
rect 17500 12404 17556 13244
rect 17500 12310 17556 12348
rect 17612 11620 17668 13356
rect 17836 12962 17892 12974
rect 17836 12910 17838 12962
rect 17890 12910 17892 12962
rect 17836 12740 17892 12910
rect 18172 12964 18228 13580
rect 17836 12674 17892 12684
rect 18060 12738 18116 12750
rect 18060 12686 18062 12738
rect 18114 12686 18116 12738
rect 18060 12628 18116 12686
rect 16828 10994 16884 11004
rect 17500 11564 17668 11620
rect 17836 12404 17892 12414
rect 17500 10948 17556 11564
rect 16604 8306 16660 8316
rect 17164 10892 17556 10948
rect 17164 9714 17220 10892
rect 17500 10834 17556 10892
rect 17500 10782 17502 10834
rect 17554 10782 17556 10834
rect 17500 10770 17556 10782
rect 17612 11394 17668 11406
rect 17612 11342 17614 11394
rect 17666 11342 17668 11394
rect 17388 10724 17444 10734
rect 17276 9828 17332 9838
rect 17276 9734 17332 9772
rect 17164 9662 17166 9714
rect 17218 9662 17220 9714
rect 16380 7646 16382 7698
rect 16434 7646 16436 7698
rect 16380 6802 16436 7646
rect 16380 6750 16382 6802
rect 16434 6750 16436 6802
rect 16380 6738 16436 6750
rect 17052 7476 17108 7486
rect 16828 6690 16884 6702
rect 16828 6638 16830 6690
rect 16882 6638 16884 6690
rect 16828 6468 16884 6638
rect 16828 6402 16884 6412
rect 16940 6692 16996 6702
rect 15820 5234 16100 5236
rect 15820 5182 15822 5234
rect 15874 5182 16100 5234
rect 15820 5180 16100 5182
rect 16268 5348 16324 5358
rect 16268 5234 16324 5292
rect 16268 5182 16270 5234
rect 16322 5182 16324 5234
rect 15820 5170 15876 5180
rect 16268 5170 16324 5182
rect 15596 5124 15652 5134
rect 15596 5122 15764 5124
rect 15596 5070 15598 5122
rect 15650 5070 15764 5122
rect 15596 5068 15764 5070
rect 15596 5058 15652 5068
rect 15148 4900 15204 4910
rect 15036 4898 15204 4900
rect 15036 4846 15150 4898
rect 15202 4846 15204 4898
rect 15036 4844 15204 4846
rect 15036 4788 15092 4844
rect 15148 4834 15204 4844
rect 15708 4900 15764 5068
rect 15036 4722 15092 4732
rect 14924 4510 14926 4562
rect 14978 4510 14980 4562
rect 14924 4498 14980 4510
rect 14476 4174 14478 4226
rect 14530 4174 14532 4226
rect 14476 4162 14532 4174
rect 13356 3554 13524 3556
rect 13356 3502 13358 3554
rect 13410 3502 13524 3554
rect 13356 3500 13524 3502
rect 15708 3556 15764 4844
rect 15932 3556 15988 3566
rect 15708 3554 15988 3556
rect 15708 3502 15934 3554
rect 15986 3502 15988 3554
rect 15708 3500 15988 3502
rect 13356 3490 13412 3500
rect 13132 3390 13134 3442
rect 13186 3390 13188 3442
rect 11564 3332 11956 3388
rect 13132 3378 13188 3390
rect 11900 980 11956 3332
rect 11900 924 12180 980
rect 12124 800 12180 924
rect 13468 800 13524 3500
rect 15932 3490 15988 3500
rect 16940 3554 16996 6636
rect 17052 6580 17108 7420
rect 17052 6486 17108 6524
rect 17164 6132 17220 9662
rect 17388 9380 17444 10668
rect 17612 10612 17668 11342
rect 17836 10836 17892 12348
rect 18060 11732 18116 12572
rect 18172 12178 18228 12908
rect 18284 12628 18340 14476
rect 18396 14530 18452 14542
rect 18396 14478 18398 14530
rect 18450 14478 18452 14530
rect 18396 14308 18452 14478
rect 18396 14242 18452 14252
rect 18620 14420 18676 14430
rect 18284 12562 18340 12572
rect 18508 12740 18564 12750
rect 18172 12126 18174 12178
rect 18226 12126 18228 12178
rect 18172 12114 18228 12126
rect 18060 11676 18452 11732
rect 17948 11508 18004 11518
rect 17948 11414 18004 11452
rect 17836 10780 18116 10836
rect 17836 10612 17892 10622
rect 17612 10610 17892 10612
rect 17612 10558 17838 10610
rect 17890 10558 17892 10610
rect 17612 10556 17892 10558
rect 17836 9938 17892 10556
rect 17836 9886 17838 9938
rect 17890 9886 17892 9938
rect 17836 9716 17892 9886
rect 17836 9650 17892 9660
rect 17948 10386 18004 10398
rect 17948 10334 17950 10386
rect 18002 10334 18004 10386
rect 17948 9828 18004 10334
rect 17276 9324 17444 9380
rect 17276 7364 17332 9324
rect 17948 9156 18004 9772
rect 17948 9090 18004 9100
rect 17836 9044 17892 9054
rect 17836 8950 17892 8988
rect 17388 8932 17444 8942
rect 17388 8930 17780 8932
rect 17388 8878 17390 8930
rect 17442 8878 17780 8930
rect 17388 8876 17780 8878
rect 17388 8866 17444 8876
rect 17724 8482 17780 8876
rect 17724 8430 17726 8482
rect 17778 8430 17780 8482
rect 17724 8418 17780 8430
rect 17500 8372 17556 8382
rect 17500 8146 17556 8316
rect 17500 8094 17502 8146
rect 17554 8094 17556 8146
rect 17500 8082 17556 8094
rect 17612 8036 17668 8046
rect 17612 7942 17668 7980
rect 17388 7364 17444 7374
rect 17276 7362 17444 7364
rect 17276 7310 17390 7362
rect 17442 7310 17444 7362
rect 17276 7308 17444 7310
rect 17388 7298 17444 7308
rect 17500 6692 17556 6702
rect 17500 6468 17556 6636
rect 17500 6402 17556 6412
rect 17164 6066 17220 6076
rect 18060 6020 18116 10780
rect 18284 10724 18340 10734
rect 18284 10630 18340 10668
rect 18396 10612 18452 11676
rect 18508 11394 18564 12684
rect 18620 12290 18676 14364
rect 18844 14308 18900 14318
rect 18732 13636 18788 13646
rect 18844 13636 18900 14252
rect 18788 13580 18900 13636
rect 18732 13542 18788 13580
rect 18732 12852 18788 12862
rect 18732 12758 18788 12796
rect 18844 12850 18900 12862
rect 18844 12798 18846 12850
rect 18898 12798 18900 12850
rect 18620 12238 18622 12290
rect 18674 12238 18676 12290
rect 18620 12226 18676 12238
rect 18844 12180 18900 12798
rect 18956 12850 19012 12862
rect 18956 12798 18958 12850
rect 19010 12798 19012 12850
rect 18956 12628 19012 12798
rect 18956 12562 19012 12572
rect 18508 11342 18510 11394
rect 18562 11342 18564 11394
rect 18508 11330 18564 11342
rect 18732 12124 18844 12180
rect 18732 11282 18788 12124
rect 18844 12114 18900 12124
rect 19068 11508 19124 15092
rect 19180 14532 19236 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15316 20244 16716
rect 20412 16100 20468 19180
rect 20636 16772 20692 27020
rect 20860 24836 20916 24846
rect 20860 24742 20916 24780
rect 21644 24722 21700 27804
rect 21756 28418 21812 28430
rect 21756 28366 21758 28418
rect 21810 28366 21812 28418
rect 21756 27076 21812 28366
rect 22988 28084 23044 28094
rect 22204 27972 22260 27982
rect 22204 27878 22260 27916
rect 22876 27860 22932 27870
rect 22876 27766 22932 27804
rect 21868 27076 21924 27086
rect 21756 27020 21868 27076
rect 21868 26982 21924 27020
rect 22540 27076 22596 27086
rect 22540 26982 22596 27020
rect 22092 26850 22148 26862
rect 22092 26798 22094 26850
rect 22146 26798 22148 26850
rect 22092 26516 22148 26798
rect 22428 26516 22484 26526
rect 22988 26516 23044 28028
rect 23436 27970 23492 27982
rect 23436 27918 23438 27970
rect 23490 27918 23492 27970
rect 22092 26514 23044 26516
rect 22092 26462 22430 26514
rect 22482 26462 22990 26514
rect 23042 26462 23044 26514
rect 22092 26460 23044 26462
rect 22428 26450 22484 26460
rect 22988 26450 23044 26460
rect 23212 27074 23268 27086
rect 23212 27022 23214 27074
rect 23266 27022 23268 27074
rect 21644 24670 21646 24722
rect 21698 24670 21700 24722
rect 21644 24658 21700 24670
rect 21868 26178 21924 26190
rect 21868 26126 21870 26178
rect 21922 26126 21924 26178
rect 21196 23042 21252 23054
rect 21196 22990 21198 23042
rect 21250 22990 21252 23042
rect 21196 22484 21252 22990
rect 21196 22418 21252 22428
rect 21308 21364 21364 21374
rect 21308 21028 21364 21308
rect 21308 20934 21364 20972
rect 21420 20692 21476 20702
rect 21420 20598 21476 20636
rect 20972 20132 21028 20142
rect 20972 19906 21028 20076
rect 20972 19854 20974 19906
rect 21026 19854 21028 19906
rect 20972 19842 21028 19854
rect 21644 19908 21700 19918
rect 21644 19814 21700 19852
rect 20748 17668 20804 17678
rect 21868 17668 21924 26126
rect 22764 25396 22820 25406
rect 22092 25394 22820 25396
rect 22092 25342 22766 25394
rect 22818 25342 22820 25394
rect 22092 25340 22820 25342
rect 22092 24946 22148 25340
rect 22764 25330 22820 25340
rect 23100 25284 23156 25294
rect 22988 25282 23156 25284
rect 22988 25230 23102 25282
rect 23154 25230 23156 25282
rect 22988 25228 23156 25230
rect 22092 24894 22094 24946
rect 22146 24894 22148 24946
rect 22092 24882 22148 24894
rect 22204 24892 22484 24948
rect 22092 23938 22148 23950
rect 22092 23886 22094 23938
rect 22146 23886 22148 23938
rect 22092 23268 22148 23886
rect 22092 23202 22148 23212
rect 21980 22258 22036 22270
rect 21980 22206 21982 22258
rect 22034 22206 22036 22258
rect 21980 21028 22036 22206
rect 22092 22146 22148 22158
rect 22092 22094 22094 22146
rect 22146 22094 22148 22146
rect 22092 21924 22148 22094
rect 22092 21858 22148 21868
rect 21980 20962 22036 20972
rect 22204 21026 22260 24892
rect 22428 24836 22484 24892
rect 22652 24836 22708 24846
rect 22428 24834 22708 24836
rect 22428 24782 22654 24834
rect 22706 24782 22708 24834
rect 22428 24780 22708 24782
rect 22652 24770 22708 24780
rect 22316 24722 22372 24734
rect 22316 24670 22318 24722
rect 22370 24670 22372 24722
rect 22316 22372 22372 24670
rect 22876 24722 22932 24734
rect 22876 24670 22878 24722
rect 22930 24670 22932 24722
rect 22876 24612 22932 24670
rect 22876 24546 22932 24556
rect 22876 24052 22932 24062
rect 22988 24052 23044 25228
rect 23100 25218 23156 25228
rect 22876 24050 23044 24052
rect 22876 23998 22878 24050
rect 22930 23998 23044 24050
rect 22876 23996 23044 23998
rect 23100 24610 23156 24622
rect 23100 24558 23102 24610
rect 23154 24558 23156 24610
rect 22876 23986 22932 23996
rect 23100 23940 23156 24558
rect 23100 23874 23156 23884
rect 22652 22484 22708 22494
rect 22652 22390 22708 22428
rect 23100 22484 23156 22494
rect 22540 22372 22596 22382
rect 22316 22370 22596 22372
rect 22316 22318 22318 22370
rect 22370 22318 22542 22370
rect 22594 22318 22596 22370
rect 22316 22316 22596 22318
rect 22316 22306 22372 22316
rect 22540 22306 22596 22316
rect 22876 22370 22932 22382
rect 22876 22318 22878 22370
rect 22930 22318 22932 22370
rect 22876 22148 22932 22318
rect 22876 22082 22932 22092
rect 22988 22370 23044 22382
rect 22988 22318 22990 22370
rect 23042 22318 23044 22370
rect 22988 21028 23044 22318
rect 23100 22370 23156 22428
rect 23100 22318 23102 22370
rect 23154 22318 23156 22370
rect 23100 22036 23156 22318
rect 23100 21970 23156 21980
rect 22204 20974 22206 21026
rect 22258 20974 22260 21026
rect 22204 20962 22260 20974
rect 22876 20972 23044 21028
rect 22092 20692 22148 20702
rect 22092 20598 22148 20636
rect 22204 20580 22260 20590
rect 22204 20578 22708 20580
rect 22204 20526 22206 20578
rect 22258 20526 22708 20578
rect 22204 20524 22708 20526
rect 22204 20514 22260 20524
rect 22540 20356 22596 20366
rect 22316 20020 22372 20030
rect 22316 19926 22372 19964
rect 22540 20018 22596 20300
rect 22540 19966 22542 20018
rect 22594 19966 22596 20018
rect 22540 19954 22596 19966
rect 22204 18338 22260 18350
rect 22204 18286 22206 18338
rect 22258 18286 22260 18338
rect 22204 18116 22260 18286
rect 22204 18050 22260 18060
rect 22652 17890 22708 20524
rect 22876 20356 22932 20972
rect 22876 20290 22932 20300
rect 22988 20802 23044 20814
rect 22988 20750 22990 20802
rect 23042 20750 23044 20802
rect 22988 20692 23044 20750
rect 22988 20018 23044 20636
rect 23100 20804 23156 20814
rect 23100 20130 23156 20748
rect 23100 20078 23102 20130
rect 23154 20078 23156 20130
rect 23100 20066 23156 20078
rect 22988 19966 22990 20018
rect 23042 19966 23044 20018
rect 22988 19954 23044 19966
rect 22876 18450 22932 18462
rect 22876 18398 22878 18450
rect 22930 18398 22932 18450
rect 22876 18116 22932 18398
rect 22876 18050 22932 18060
rect 23100 18338 23156 18350
rect 23100 18286 23102 18338
rect 23154 18286 23156 18338
rect 23100 18004 23156 18286
rect 23100 17938 23156 17948
rect 22652 17838 22654 17890
rect 22706 17838 22708 17890
rect 21868 17612 22036 17668
rect 20748 16996 20804 17612
rect 21420 17444 21476 17454
rect 21868 17444 21924 17454
rect 21420 17442 21924 17444
rect 21420 17390 21422 17442
rect 21474 17390 21870 17442
rect 21922 17390 21924 17442
rect 21420 17388 21924 17390
rect 21420 17378 21476 17388
rect 20972 16996 21028 17006
rect 20748 16940 20972 16996
rect 20972 16882 21028 16940
rect 21868 16996 21924 17388
rect 21868 16930 21924 16940
rect 20972 16830 20974 16882
rect 21026 16830 21028 16882
rect 20972 16818 21028 16830
rect 21420 16882 21476 16894
rect 21420 16830 21422 16882
rect 21474 16830 21476 16882
rect 20636 16706 20692 16716
rect 21420 16212 21476 16830
rect 21756 16770 21812 16782
rect 21756 16718 21758 16770
rect 21810 16718 21812 16770
rect 21756 16436 21812 16718
rect 21756 16370 21812 16380
rect 21420 16146 21476 16156
rect 21756 16210 21812 16222
rect 21756 16158 21758 16210
rect 21810 16158 21812 16210
rect 20524 16100 20580 16110
rect 20412 16098 20580 16100
rect 20412 16046 20526 16098
rect 20578 16046 20580 16098
rect 20412 16044 20580 16046
rect 20524 15988 20580 16044
rect 21644 16100 21700 16110
rect 20524 15922 20580 15932
rect 21420 15986 21476 15998
rect 21420 15934 21422 15986
rect 21474 15934 21476 15986
rect 19516 15202 19572 15214
rect 19516 15150 19518 15202
rect 19570 15150 19572 15202
rect 19516 15092 19572 15150
rect 19516 15026 19572 15036
rect 19628 14532 19684 14542
rect 19180 14530 19684 14532
rect 19180 14478 19182 14530
rect 19234 14478 19630 14530
rect 19682 14478 19684 14530
rect 19180 14476 19684 14478
rect 19180 14466 19236 14476
rect 19628 14466 19684 14476
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13748 20244 15260
rect 20972 15316 21028 15326
rect 20972 15222 21028 15260
rect 21420 15148 21476 15934
rect 21644 15986 21700 16044
rect 21644 15934 21646 15986
rect 21698 15934 21700 15986
rect 21644 15922 21700 15934
rect 21756 15426 21812 16158
rect 21980 16100 22036 17612
rect 22540 17556 22596 17566
rect 22540 17462 22596 17500
rect 22652 17108 22708 17838
rect 22764 17108 22820 17118
rect 22652 17106 22820 17108
rect 22652 17054 22766 17106
rect 22818 17054 22820 17106
rect 22652 17052 22820 17054
rect 22764 17042 22820 17052
rect 22428 16882 22484 16894
rect 22428 16830 22430 16882
rect 22482 16830 22484 16882
rect 22428 16324 22484 16830
rect 22428 16258 22484 16268
rect 23100 16882 23156 16894
rect 23100 16830 23102 16882
rect 23154 16830 23156 16882
rect 23100 16324 23156 16830
rect 23100 16258 23156 16268
rect 21980 16034 22036 16044
rect 22092 16212 22148 16222
rect 22092 16098 22148 16156
rect 22092 16046 22094 16098
rect 22146 16046 22148 16098
rect 22092 16034 22148 16046
rect 22876 16100 22932 16110
rect 21756 15374 21758 15426
rect 21810 15374 21812 15426
rect 21756 15362 21812 15374
rect 22428 15874 22484 15886
rect 22428 15822 22430 15874
rect 22482 15822 22484 15874
rect 21308 15092 21476 15148
rect 22428 15148 22484 15822
rect 22876 15148 22932 16044
rect 22428 15092 22596 15148
rect 21308 14642 21364 15092
rect 21308 14590 21310 14642
rect 21362 14590 21364 14642
rect 21308 14578 21364 14590
rect 21756 14868 21812 14878
rect 21756 14532 21812 14812
rect 22204 14532 22260 14542
rect 21756 14530 22036 14532
rect 21756 14478 21758 14530
rect 21810 14478 22036 14530
rect 21756 14476 22036 14478
rect 21756 14466 21812 14476
rect 20188 13746 20692 13748
rect 20188 13694 20190 13746
rect 20242 13694 20692 13746
rect 20188 13692 20692 13694
rect 20188 13682 20244 13692
rect 19628 12852 19684 12862
rect 19404 12738 19460 12750
rect 19404 12686 19406 12738
rect 19458 12686 19460 12738
rect 19404 12292 19460 12686
rect 18732 11230 18734 11282
rect 18786 11230 18788 11282
rect 18732 11218 18788 11230
rect 18844 11452 19124 11508
rect 19292 12180 19348 12190
rect 18844 10724 18900 11452
rect 18956 11284 19012 11294
rect 18956 11190 19012 11228
rect 19292 10836 19348 12124
rect 18284 9044 18340 9054
rect 18396 9044 18452 10556
rect 18284 9042 18452 9044
rect 18284 8990 18286 9042
rect 18338 8990 18452 9042
rect 18284 8988 18452 8990
rect 18732 10668 18900 10724
rect 18956 10834 19348 10836
rect 18956 10782 19294 10834
rect 19346 10782 19348 10834
rect 18956 10780 19348 10782
rect 18284 8978 18340 8988
rect 18732 8932 18788 10668
rect 18844 10500 18900 10510
rect 18956 10500 19012 10780
rect 19292 10770 19348 10780
rect 19180 10666 19236 10678
rect 19068 10612 19124 10622
rect 19180 10614 19182 10666
rect 19234 10614 19236 10666
rect 19180 10612 19236 10614
rect 19124 10556 19236 10612
rect 19068 10546 19124 10556
rect 18844 10498 19012 10500
rect 18844 10446 18846 10498
rect 18898 10446 19012 10498
rect 18844 10444 19012 10446
rect 18844 10434 18900 10444
rect 19292 10388 19348 10398
rect 18956 10386 19348 10388
rect 18956 10334 19294 10386
rect 19346 10334 19348 10386
rect 18956 10332 19348 10334
rect 18956 9154 19012 10332
rect 19292 10322 19348 10332
rect 18956 9102 18958 9154
rect 19010 9102 19012 9154
rect 18956 9090 19012 9102
rect 19180 9156 19236 9166
rect 19180 9062 19236 9100
rect 19404 9042 19460 12236
rect 19628 12290 19684 12796
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19628 12238 19630 12290
rect 19682 12238 19684 12290
rect 19516 11508 19572 11518
rect 19628 11508 19684 12238
rect 19740 12180 19796 12190
rect 19740 12086 19796 12124
rect 19572 11452 19684 11508
rect 19516 11442 19572 11452
rect 19628 11282 19684 11294
rect 19628 11230 19630 11282
rect 19682 11230 19684 11282
rect 19628 11172 19684 11230
rect 19628 11106 19684 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20636 9826 20692 13692
rect 20860 13634 20916 13646
rect 20860 13582 20862 13634
rect 20914 13582 20916 13634
rect 20860 11620 20916 13582
rect 21420 13636 21476 13646
rect 21420 12516 21476 13580
rect 21196 12068 21252 12078
rect 21196 11974 21252 12012
rect 21308 11620 21364 11630
rect 20860 11618 21364 11620
rect 20860 11566 21310 11618
rect 21362 11566 21364 11618
rect 20860 11564 21364 11566
rect 21308 11554 21364 11564
rect 21420 11618 21476 12460
rect 21980 12404 22036 14476
rect 22204 14530 22372 14532
rect 22204 14478 22206 14530
rect 22258 14478 22372 14530
rect 22204 14476 22372 14478
rect 22204 14466 22260 14476
rect 22092 13300 22148 13310
rect 22092 13074 22148 13244
rect 22092 13022 22094 13074
rect 22146 13022 22148 13074
rect 22092 13010 22148 13022
rect 21532 12292 21588 12302
rect 21532 12178 21588 12236
rect 21980 12290 22036 12348
rect 21980 12238 21982 12290
rect 22034 12238 22036 12290
rect 21980 12226 22036 12238
rect 22204 12740 22260 12750
rect 22204 12290 22260 12684
rect 22204 12238 22206 12290
rect 22258 12238 22260 12290
rect 22204 12226 22260 12238
rect 22316 12292 22372 14476
rect 22428 12852 22484 12862
rect 22428 12758 22484 12796
rect 22316 12226 22372 12236
rect 21532 12126 21534 12178
rect 21586 12126 21588 12178
rect 21532 12114 21588 12126
rect 21756 12066 21812 12078
rect 21756 12014 21758 12066
rect 21810 12014 21812 12066
rect 21420 11566 21422 11618
rect 21474 11566 21476 11618
rect 20860 11396 20916 11406
rect 21420 11396 21476 11566
rect 21644 11620 21700 11630
rect 21756 11620 21812 12014
rect 22540 11956 22596 15092
rect 21644 11618 21812 11620
rect 21644 11566 21646 11618
rect 21698 11566 21812 11618
rect 21644 11564 21812 11566
rect 22428 11900 22596 11956
rect 22652 15092 22932 15148
rect 21644 11554 21700 11564
rect 21756 11396 21812 11406
rect 20860 11394 21476 11396
rect 20860 11342 20862 11394
rect 20914 11342 21476 11394
rect 20860 11340 21476 11342
rect 21644 11340 21756 11396
rect 20860 11330 20916 11340
rect 21644 9938 21700 11340
rect 21756 11302 21812 11340
rect 21644 9886 21646 9938
rect 21698 9886 21700 9938
rect 21644 9874 21700 9886
rect 22428 9940 22484 11900
rect 22540 11506 22596 11518
rect 22540 11454 22542 11506
rect 22594 11454 22596 11506
rect 22540 11396 22596 11454
rect 22652 11396 22708 15092
rect 22988 13634 23044 13646
rect 22988 13582 22990 13634
rect 23042 13582 23044 13634
rect 22764 12740 22820 12750
rect 22988 12740 23044 13582
rect 23212 13076 23268 27022
rect 23436 27076 23492 27918
rect 23436 27010 23492 27020
rect 23548 24612 23604 29372
rect 23660 28756 23716 28766
rect 23660 27074 23716 28700
rect 24220 28530 24276 30156
rect 24332 28644 24388 28654
rect 24780 28644 24836 32060
rect 25340 30322 25396 32284
rect 25788 32116 25844 32126
rect 25900 32116 25956 33404
rect 26012 33346 26068 33358
rect 26012 33294 26014 33346
rect 26066 33294 26068 33346
rect 26012 33124 26068 33294
rect 26012 33058 26068 33068
rect 25844 32060 25956 32116
rect 25788 32050 25844 32060
rect 26124 30660 26180 35756
rect 26460 35588 26516 35598
rect 26796 35588 26852 35598
rect 26460 35586 26852 35588
rect 26460 35534 26462 35586
rect 26514 35534 26798 35586
rect 26850 35534 26852 35586
rect 26460 35532 26852 35534
rect 26460 35522 26516 35532
rect 26796 35522 26852 35532
rect 26236 35364 26292 35374
rect 26236 34802 26292 35308
rect 26684 35252 26740 35262
rect 26684 35026 26740 35196
rect 26684 34974 26686 35026
rect 26738 34974 26740 35026
rect 26684 34962 26740 34974
rect 26236 34750 26238 34802
rect 26290 34750 26292 34802
rect 26236 31220 26292 34750
rect 26460 33460 26516 33470
rect 26460 33366 26516 33404
rect 27020 33236 27076 35868
rect 27132 35586 27188 36316
rect 27804 36306 27860 36316
rect 27132 35534 27134 35586
rect 27186 35534 27188 35586
rect 27132 35522 27188 35534
rect 27468 35252 27524 35262
rect 27132 33236 27188 33246
rect 27020 33234 27188 33236
rect 27020 33182 27134 33234
rect 27186 33182 27188 33234
rect 27020 33180 27188 33182
rect 27132 33170 27188 33180
rect 27468 33234 27524 35196
rect 27916 33460 27972 38612
rect 28364 38164 28420 38174
rect 28364 38070 28420 38108
rect 29036 38164 29092 42252
rect 30716 41972 30772 45164
rect 30828 45126 30884 45164
rect 31164 45220 31220 45230
rect 31836 45220 31892 45230
rect 31164 45218 31444 45220
rect 31164 45166 31166 45218
rect 31218 45166 31444 45218
rect 31164 45164 31444 45166
rect 31164 45154 31220 45164
rect 30940 44436 30996 44446
rect 30940 44342 30996 44380
rect 31164 44100 31220 44110
rect 31164 44006 31220 44044
rect 30828 43540 30884 43550
rect 30828 43446 30884 43484
rect 31276 43428 31332 43438
rect 31276 43334 31332 43372
rect 31276 42868 31332 42878
rect 31276 42774 31332 42812
rect 30828 41972 30884 41982
rect 30716 41916 30828 41972
rect 31388 41972 31444 45164
rect 31612 45106 31668 45118
rect 31612 45054 31614 45106
rect 31666 45054 31668 45106
rect 31500 44098 31556 44110
rect 31500 44046 31502 44098
rect 31554 44046 31556 44098
rect 31500 43876 31556 44046
rect 31500 43810 31556 43820
rect 31612 43764 31668 45054
rect 31836 44324 31892 45164
rect 32172 45220 32228 45230
rect 32284 45220 32340 45838
rect 32844 45890 32900 45902
rect 32844 45838 32846 45890
rect 32898 45838 32900 45890
rect 32508 45668 32564 45678
rect 32508 45574 32564 45612
rect 32508 45220 32564 45230
rect 32284 45218 32564 45220
rect 32284 45166 32510 45218
rect 32562 45166 32564 45218
rect 32284 45164 32564 45166
rect 32172 45126 32228 45164
rect 31836 44230 31892 44268
rect 31948 45108 32004 45118
rect 31612 43698 31668 43708
rect 31500 43650 31556 43662
rect 31500 43598 31502 43650
rect 31554 43598 31556 43650
rect 31500 43428 31556 43598
rect 31724 43540 31780 43550
rect 31724 43446 31780 43484
rect 31500 43362 31556 43372
rect 31948 42754 32004 45052
rect 32508 44996 32564 45164
rect 32508 44940 32788 44996
rect 32172 44548 32228 44558
rect 32172 44210 32228 44492
rect 32620 44324 32676 44334
rect 32620 44230 32676 44268
rect 32172 44158 32174 44210
rect 32226 44158 32228 44210
rect 32172 44146 32228 44158
rect 32396 44100 32452 44110
rect 32284 43538 32340 43550
rect 32284 43486 32286 43538
rect 32338 43486 32340 43538
rect 32284 43428 32340 43486
rect 32284 43362 32340 43372
rect 31948 42702 31950 42754
rect 32002 42702 32004 42754
rect 31388 41916 31780 41972
rect 30828 41906 30884 41916
rect 30940 41860 30996 41870
rect 30828 41188 30884 41198
rect 30604 41132 30828 41188
rect 29820 40964 29876 40974
rect 29820 40514 29876 40908
rect 29820 40462 29822 40514
rect 29874 40462 29876 40514
rect 29820 40450 29876 40462
rect 30604 40404 30660 41132
rect 30828 41094 30884 41132
rect 30604 40310 30660 40348
rect 30940 40964 30996 41804
rect 30940 40402 30996 40908
rect 30940 40350 30942 40402
rect 30994 40350 30996 40402
rect 30940 40338 30996 40350
rect 31388 40402 31444 40414
rect 31388 40350 31390 40402
rect 31442 40350 31444 40402
rect 29260 40292 29316 40302
rect 29148 38836 29204 38846
rect 29260 38836 29316 40236
rect 30604 39396 30660 39406
rect 31276 39396 31332 39406
rect 31388 39396 31444 40350
rect 31612 39396 31668 39406
rect 29148 38834 29316 38836
rect 29148 38782 29150 38834
rect 29202 38782 29316 38834
rect 29148 38780 29316 38782
rect 29148 38770 29204 38780
rect 29036 38098 29092 38108
rect 29260 38052 29316 38780
rect 30492 39394 31668 39396
rect 30492 39342 30606 39394
rect 30658 39342 31278 39394
rect 31330 39342 31614 39394
rect 31666 39342 31668 39394
rect 30492 39340 31668 39342
rect 29820 38722 29876 38734
rect 29820 38670 29822 38722
rect 29874 38670 29876 38722
rect 29820 38668 29876 38670
rect 30268 38724 30324 38734
rect 29820 38612 29988 38668
rect 29932 38274 29988 38612
rect 29932 38222 29934 38274
rect 29986 38222 29988 38274
rect 29932 38210 29988 38222
rect 30268 38274 30324 38668
rect 30268 38222 30270 38274
rect 30322 38222 30324 38274
rect 30268 38210 30324 38222
rect 29260 36594 29316 37996
rect 30044 37828 30100 37838
rect 30044 37826 30212 37828
rect 30044 37774 30046 37826
rect 30098 37774 30212 37826
rect 30044 37772 30212 37774
rect 30044 37762 30100 37772
rect 29260 36542 29262 36594
rect 29314 36542 29316 36594
rect 28588 36484 28644 36494
rect 28588 36390 28644 36428
rect 29260 36484 29316 36542
rect 29260 36418 29316 36428
rect 29820 36484 29876 36494
rect 29820 36390 29876 36428
rect 30156 36036 30212 37772
rect 30156 35980 30436 36036
rect 29148 35924 29204 35934
rect 27468 33182 27470 33234
rect 27522 33182 27524 33234
rect 27468 33170 27524 33182
rect 27804 33348 27860 33358
rect 27916 33348 27972 33404
rect 27804 33346 27972 33348
rect 27804 33294 27806 33346
rect 27858 33294 27972 33346
rect 27804 33292 27972 33294
rect 28476 34692 28532 34702
rect 26348 33124 26404 33134
rect 26796 33124 26852 33134
rect 26404 33122 26852 33124
rect 26404 33070 26798 33122
rect 26850 33070 26852 33122
rect 26404 33068 26852 33070
rect 26348 33030 26404 33068
rect 26796 33058 26852 33068
rect 27132 32788 27188 32798
rect 27132 32694 27188 32732
rect 27804 32788 27860 33292
rect 27804 32722 27860 32732
rect 26796 32674 26852 32686
rect 26796 32622 26798 32674
rect 26850 32622 26852 32674
rect 26796 31444 26852 32622
rect 28476 32564 28532 34636
rect 29148 33346 29204 35868
rect 30156 35924 30212 35980
rect 30156 35858 30212 35868
rect 30380 35698 30436 35980
rect 30380 35646 30382 35698
rect 30434 35646 30436 35698
rect 30380 35634 30436 35646
rect 30492 35252 30548 39340
rect 30604 39330 30660 39340
rect 31276 39330 31332 39340
rect 31612 39330 31668 39340
rect 31724 38052 31780 41916
rect 31948 41860 32004 42702
rect 32396 42644 32452 44044
rect 32508 43988 32564 43998
rect 32732 43988 32788 44940
rect 32844 44210 32900 45838
rect 32956 45220 33012 49200
rect 33628 46228 33684 49200
rect 33628 46172 34132 46228
rect 33180 45220 33236 45230
rect 33516 45220 33572 45230
rect 32956 45218 33236 45220
rect 32956 45166 33182 45218
rect 33234 45166 33236 45218
rect 32956 45164 33236 45166
rect 32956 44996 33012 45164
rect 33180 45154 33236 45164
rect 33404 45218 33572 45220
rect 33404 45166 33518 45218
rect 33570 45166 33572 45218
rect 33404 45164 33572 45166
rect 32956 44930 33012 44940
rect 32844 44158 32846 44210
rect 32898 44158 32900 44210
rect 32844 44146 32900 44158
rect 33180 44098 33236 44110
rect 33180 44046 33182 44098
rect 33234 44046 33236 44098
rect 33180 43988 33236 44046
rect 32732 43932 33236 43988
rect 32508 43650 32564 43932
rect 32508 43598 32510 43650
rect 32562 43598 32564 43650
rect 32508 43586 32564 43598
rect 33180 43428 33236 43438
rect 33236 43372 33348 43428
rect 33180 43334 33236 43372
rect 32844 42756 32900 42766
rect 32508 42644 32564 42654
rect 32396 42642 32564 42644
rect 32396 42590 32510 42642
rect 32562 42590 32564 42642
rect 32396 42588 32564 42590
rect 31836 41188 31892 41198
rect 31948 41188 32004 41804
rect 31892 41132 32004 41188
rect 32172 41860 32228 41870
rect 32508 41860 32564 42588
rect 32844 42642 32900 42700
rect 32844 42590 32846 42642
rect 32898 42590 32900 42642
rect 32844 42578 32900 42590
rect 33292 42754 33348 43372
rect 33292 42702 33294 42754
rect 33346 42702 33348 42754
rect 33292 42308 33348 42702
rect 33292 42242 33348 42252
rect 32172 41858 32564 41860
rect 32172 41806 32174 41858
rect 32226 41806 32564 41858
rect 32172 41804 32564 41806
rect 33180 41860 33236 41870
rect 33236 41804 33348 41860
rect 31836 41094 31892 41132
rect 31948 39394 32004 39406
rect 31948 39342 31950 39394
rect 32002 39342 32004 39394
rect 31948 39060 32004 39342
rect 32172 39172 32228 41804
rect 33180 41766 33236 41804
rect 32508 41074 32564 41086
rect 32508 41022 32510 41074
rect 32562 41022 32564 41074
rect 32508 40404 32564 41022
rect 32508 40338 32564 40348
rect 32396 39172 32452 39182
rect 32172 39116 32396 39172
rect 32396 39106 32452 39116
rect 31948 38994 32004 39004
rect 32508 39060 32564 39070
rect 32508 38966 32564 39004
rect 33180 38948 33236 38958
rect 33180 38854 33236 38892
rect 32396 38836 32452 38846
rect 31948 38834 32452 38836
rect 31948 38782 32398 38834
rect 32450 38782 32452 38834
rect 31948 38780 32452 38782
rect 31948 38722 32004 38780
rect 32396 38770 32452 38780
rect 31948 38670 31950 38722
rect 32002 38670 32004 38722
rect 31948 38658 32004 38670
rect 33068 38724 33124 38762
rect 33292 38668 33348 41804
rect 33404 39956 33460 45164
rect 33516 45154 33572 45164
rect 33852 45220 33908 45230
rect 33852 45218 34020 45220
rect 33852 45166 33854 45218
rect 33906 45166 34020 45218
rect 33852 45164 34020 45166
rect 33852 45154 33908 45164
rect 33852 44322 33908 44334
rect 33852 44270 33854 44322
rect 33906 44270 33908 44322
rect 33516 44100 33572 44110
rect 33516 44006 33572 44044
rect 33852 43988 33908 44270
rect 33852 43922 33908 43932
rect 33628 43764 33684 43774
rect 33628 43538 33684 43708
rect 33852 43650 33908 43662
rect 33852 43598 33854 43650
rect 33906 43598 33908 43650
rect 33628 43486 33630 43538
rect 33682 43486 33684 43538
rect 33628 43316 33684 43486
rect 33628 43250 33684 43260
rect 33740 43540 33796 43550
rect 33516 42644 33572 42654
rect 33516 42550 33572 42588
rect 33740 42084 33796 43484
rect 33852 43428 33908 43598
rect 33852 43362 33908 43372
rect 33852 42756 33908 42766
rect 33852 42662 33908 42700
rect 33740 41970 33796 42028
rect 33740 41918 33742 41970
rect 33794 41918 33796 41970
rect 33740 41906 33796 41918
rect 33516 41860 33572 41870
rect 33572 41804 33684 41860
rect 33516 41794 33572 41804
rect 33628 40628 33684 41804
rect 33740 40628 33796 40638
rect 33628 40626 33796 40628
rect 33628 40574 33742 40626
rect 33794 40574 33796 40626
rect 33628 40572 33796 40574
rect 33740 40562 33796 40572
rect 33964 40180 34020 45164
rect 34076 45106 34132 46172
rect 34972 46116 35028 49200
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 34972 46050 35028 46060
rect 36988 46116 37044 46126
rect 36988 46022 37044 46060
rect 40348 46116 40404 49200
rect 40348 46050 40404 46060
rect 35196 46002 35252 46014
rect 35196 45950 35198 46002
rect 35250 45950 35252 46002
rect 34076 45054 34078 45106
rect 34130 45054 34132 45106
rect 34076 44436 34132 45054
rect 34076 44370 34132 44380
rect 34300 45668 34356 45678
rect 34300 43538 34356 45612
rect 35196 45444 35252 45950
rect 35196 45378 35252 45388
rect 35980 45890 36036 45902
rect 35980 45838 35982 45890
rect 36034 45838 36036 45890
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34524 43652 34580 43662
rect 34524 43558 34580 43596
rect 34300 43486 34302 43538
rect 34354 43486 34356 43538
rect 34076 42082 34132 42094
rect 34076 42030 34078 42082
rect 34130 42030 34132 42082
rect 34076 40852 34132 42030
rect 34300 41748 34356 43486
rect 35084 43538 35140 43550
rect 35084 43486 35086 43538
rect 35138 43486 35140 43538
rect 34412 43428 34468 43438
rect 34468 43372 34692 43428
rect 34412 43362 34468 43372
rect 34524 42084 34580 42094
rect 34300 41682 34356 41692
rect 34412 41970 34468 41982
rect 34412 41918 34414 41970
rect 34466 41918 34468 41970
rect 34412 41076 34468 41918
rect 34076 40786 34132 40796
rect 34188 41020 34468 41076
rect 34076 40628 34132 40638
rect 34188 40628 34244 41020
rect 34076 40626 34244 40628
rect 34076 40574 34078 40626
rect 34130 40574 34244 40626
rect 34076 40572 34244 40574
rect 34076 40562 34132 40572
rect 33404 39890 33460 39900
rect 33628 40124 34020 40180
rect 34412 40178 34468 40190
rect 34412 40126 34414 40178
rect 34466 40126 34468 40178
rect 33404 39396 33460 39406
rect 33404 38946 33460 39340
rect 33404 38894 33406 38946
rect 33458 38894 33460 38946
rect 33404 38882 33460 38894
rect 33516 39172 33572 39182
rect 33068 38658 33124 38668
rect 31724 37986 31780 37996
rect 33180 38612 33348 38668
rect 33180 38050 33236 38612
rect 33180 37998 33182 38050
rect 33234 37998 33236 38050
rect 32172 37828 32228 37838
rect 32844 37828 32900 37838
rect 33180 37828 33236 37998
rect 32172 37826 33236 37828
rect 32172 37774 32174 37826
rect 32226 37774 32846 37826
rect 32898 37774 33236 37826
rect 32172 37772 33236 37774
rect 32172 37762 32228 37772
rect 32844 37762 32900 37772
rect 32732 36594 32788 36606
rect 32732 36542 32734 36594
rect 32786 36542 32788 36594
rect 30604 36370 30660 36382
rect 30604 36318 30606 36370
rect 30658 36318 30660 36370
rect 30604 35922 30660 36318
rect 30604 35870 30606 35922
rect 30658 35870 30660 35922
rect 30604 35858 30660 35870
rect 31164 35698 31220 35710
rect 31164 35646 31166 35698
rect 31218 35646 31220 35698
rect 30716 35588 30772 35598
rect 31052 35588 31108 35598
rect 30716 35586 31108 35588
rect 30716 35534 30718 35586
rect 30770 35534 31054 35586
rect 31106 35534 31108 35586
rect 30716 35532 31108 35534
rect 30716 35522 30772 35532
rect 31052 35522 31108 35532
rect 30492 35186 30548 35196
rect 29148 33294 29150 33346
rect 29202 33294 29204 33346
rect 29148 33282 29204 33294
rect 29260 34914 29316 34926
rect 29260 34862 29262 34914
rect 29314 34862 29316 34914
rect 29260 32676 29316 34862
rect 29932 34804 29988 34814
rect 29596 34802 29988 34804
rect 29596 34750 29934 34802
rect 29986 34750 29988 34802
rect 29596 34748 29988 34750
rect 29596 33458 29652 34748
rect 29932 34738 29988 34748
rect 31164 34468 31220 35646
rect 31724 35698 31780 35710
rect 31724 35646 31726 35698
rect 31778 35646 31780 35698
rect 31724 34804 31780 35646
rect 32508 35588 32564 35598
rect 31724 34738 31780 34748
rect 32060 35026 32116 35038
rect 32060 34974 32062 35026
rect 32114 34974 32116 35026
rect 29596 33406 29598 33458
rect 29650 33406 29652 33458
rect 29596 33394 29652 33406
rect 30940 34412 31220 34468
rect 30940 33458 30996 34412
rect 30940 33406 30942 33458
rect 30994 33406 30996 33458
rect 30940 33394 30996 33406
rect 31052 34242 31108 34254
rect 31052 34190 31054 34242
rect 31106 34190 31108 34242
rect 31052 33460 31108 34190
rect 31724 34242 31780 34254
rect 31724 34190 31726 34242
rect 31778 34190 31780 34242
rect 31388 34132 31444 34142
rect 31724 34132 31780 34190
rect 31388 34130 31780 34132
rect 31388 34078 31390 34130
rect 31442 34078 31780 34130
rect 31388 34076 31780 34078
rect 32060 34132 32116 34974
rect 31052 33404 31332 33460
rect 28476 32470 28532 32508
rect 29148 32620 29260 32676
rect 28812 32450 28868 32462
rect 28812 32398 28814 32450
rect 28866 32398 28868 32450
rect 28812 32004 28868 32398
rect 28812 31938 28868 31948
rect 29036 32338 29092 32350
rect 29036 32286 29038 32338
rect 29090 32286 29092 32338
rect 29036 31666 29092 32286
rect 29036 31614 29038 31666
rect 29090 31614 29092 31666
rect 29036 31602 29092 31614
rect 26796 31378 26852 31388
rect 27356 31276 27748 31332
rect 27132 31220 27188 31230
rect 27356 31220 27412 31276
rect 26236 31218 26628 31220
rect 26236 31166 26238 31218
rect 26290 31166 26628 31218
rect 26236 31164 26628 31166
rect 26236 31154 26292 31164
rect 26572 30994 26628 31164
rect 27132 31218 27412 31220
rect 27132 31166 27134 31218
rect 27186 31166 27412 31218
rect 27132 31164 27412 31166
rect 27132 31154 27188 31164
rect 26572 30942 26574 30994
rect 26626 30942 26628 30994
rect 26572 30930 26628 30942
rect 27468 31106 27524 31118
rect 27468 31054 27470 31106
rect 27522 31054 27524 31106
rect 26796 30884 26852 30894
rect 26796 30790 26852 30828
rect 26124 30604 26292 30660
rect 25340 30270 25342 30322
rect 25394 30270 25396 30322
rect 25340 30258 25396 30270
rect 25116 30212 25172 30222
rect 25116 30118 25172 30156
rect 25676 30210 25732 30222
rect 25676 30158 25678 30210
rect 25730 30158 25732 30210
rect 25676 29764 25732 30158
rect 26236 29986 26292 30604
rect 26236 29934 26238 29986
rect 26290 29934 26292 29986
rect 26236 29922 26292 29934
rect 26572 29986 26628 29998
rect 26572 29934 26574 29986
rect 26626 29934 26628 29986
rect 26572 29764 26628 29934
rect 25676 29708 26628 29764
rect 24332 28642 24836 28644
rect 24332 28590 24334 28642
rect 24386 28590 24836 28642
rect 24332 28588 24836 28590
rect 24892 28756 24948 28766
rect 24332 28578 24388 28588
rect 24220 28478 24222 28530
rect 24274 28478 24276 28530
rect 23996 28418 24052 28430
rect 23996 28366 23998 28418
rect 24050 28366 24052 28418
rect 23772 28084 23828 28094
rect 23996 28084 24052 28366
rect 24108 28084 24164 28094
rect 23772 28082 24164 28084
rect 23772 28030 23774 28082
rect 23826 28030 24110 28082
rect 24162 28030 24164 28082
rect 23772 28028 24164 28030
rect 23772 28018 23828 28028
rect 23660 27022 23662 27074
rect 23714 27022 23716 27074
rect 23660 27010 23716 27022
rect 24108 27074 24164 28028
rect 24108 27022 24110 27074
rect 24162 27022 24164 27074
rect 24108 27010 24164 27022
rect 23548 24052 23604 24556
rect 23548 23986 23604 23996
rect 24220 23940 24276 28478
rect 24556 27746 24612 27758
rect 24556 27694 24558 27746
rect 24610 27694 24612 27746
rect 24220 23874 24276 23884
rect 24332 27524 24388 27534
rect 24556 27524 24612 27694
rect 24388 27468 24612 27524
rect 23324 23042 23380 23054
rect 23324 22990 23326 23042
rect 23378 22990 23380 23042
rect 23324 22372 23380 22990
rect 24332 22484 24388 27468
rect 24668 27188 24724 27198
rect 24444 26964 24500 26974
rect 24668 26964 24724 27132
rect 24892 27186 24948 28700
rect 25340 28644 25396 28654
rect 25340 27860 25396 28588
rect 25340 27858 25732 27860
rect 25340 27806 25342 27858
rect 25394 27806 25732 27858
rect 25340 27804 25732 27806
rect 25340 27794 25396 27804
rect 24892 27134 24894 27186
rect 24946 27134 24948 27186
rect 24892 27122 24948 27134
rect 25340 27524 25396 27534
rect 25340 27186 25396 27468
rect 25340 27134 25342 27186
rect 25394 27134 25396 27186
rect 25340 27122 25396 27134
rect 24444 26962 24724 26964
rect 24444 26910 24446 26962
rect 24498 26910 24724 26962
rect 24444 26908 24724 26910
rect 24444 26898 24500 26908
rect 24668 25620 24724 26908
rect 24668 25618 25060 25620
rect 24668 25566 24670 25618
rect 24722 25566 25060 25618
rect 24668 25564 25060 25566
rect 24668 25554 24724 25564
rect 24668 24724 24724 24734
rect 24668 24630 24724 24668
rect 24444 22484 24500 22494
rect 24388 22482 24500 22484
rect 24388 22430 24446 22482
rect 24498 22430 24500 22482
rect 24388 22428 24500 22430
rect 24332 22390 24388 22428
rect 24444 22418 24500 22428
rect 24780 22372 24836 25564
rect 25004 25506 25060 25564
rect 25004 25454 25006 25506
rect 25058 25454 25060 25506
rect 25004 25442 25060 25454
rect 25676 25506 25732 27804
rect 26012 27748 26068 27758
rect 25900 27746 26068 27748
rect 25900 27694 26014 27746
rect 26066 27694 26068 27746
rect 25900 27692 26068 27694
rect 25788 27524 25844 27534
rect 25788 26962 25844 27468
rect 25900 27186 25956 27692
rect 26012 27682 26068 27692
rect 26012 27300 26068 27310
rect 26012 27206 26068 27244
rect 25900 27134 25902 27186
rect 25954 27134 25956 27186
rect 25900 27122 25956 27134
rect 25788 26910 25790 26962
rect 25842 26910 25844 26962
rect 25788 26898 25844 26910
rect 26572 26516 26628 29708
rect 27468 29538 27524 31054
rect 27692 30994 27748 31276
rect 27692 30942 27694 30994
rect 27746 30942 27748 30994
rect 27692 30930 27748 30942
rect 27468 29486 27470 29538
rect 27522 29486 27524 29538
rect 27468 29474 27524 29486
rect 26796 29426 26852 29438
rect 26796 29374 26798 29426
rect 26850 29374 26852 29426
rect 26796 28644 26852 29374
rect 26796 28578 26852 28588
rect 29148 28644 29204 32620
rect 29260 32610 29316 32620
rect 29484 33346 29540 33358
rect 29484 33294 29486 33346
rect 29538 33294 29540 33346
rect 29260 32340 29316 32350
rect 29260 32338 29428 32340
rect 29260 32286 29262 32338
rect 29314 32286 29428 32338
rect 29260 32284 29428 32286
rect 29260 32274 29316 32284
rect 29260 31666 29316 31678
rect 29260 31614 29262 31666
rect 29314 31614 29316 31666
rect 29260 31220 29316 31614
rect 29372 31332 29428 32284
rect 29484 31892 29540 33294
rect 29708 33234 29764 33246
rect 29708 33182 29710 33234
rect 29762 33182 29764 33234
rect 29708 32786 29764 33182
rect 30604 33236 30660 33246
rect 30828 33236 30884 33246
rect 30604 33234 30772 33236
rect 30604 33182 30606 33234
rect 30658 33182 30772 33234
rect 30604 33180 30772 33182
rect 30604 33170 30660 33180
rect 29708 32734 29710 32786
rect 29762 32734 29764 32786
rect 29708 32722 29764 32734
rect 30268 33124 30324 33134
rect 29484 31826 29540 31836
rect 29820 32564 29876 32574
rect 29932 32564 29988 32574
rect 30268 32564 30324 33068
rect 29876 32562 30324 32564
rect 29876 32510 29934 32562
rect 29986 32510 30324 32562
rect 29876 32508 30324 32510
rect 29708 31780 29764 31790
rect 29708 31686 29764 31724
rect 29484 31554 29540 31566
rect 29484 31502 29486 31554
rect 29538 31502 29540 31554
rect 29484 31444 29540 31502
rect 29596 31556 29652 31566
rect 29596 31462 29652 31500
rect 29484 31378 29540 31388
rect 29372 31266 29428 31276
rect 29260 31126 29316 31164
rect 29372 30996 29428 31006
rect 29372 30902 29428 30940
rect 29260 30772 29316 30782
rect 29708 30772 29764 30782
rect 29260 30770 29764 30772
rect 29260 30718 29262 30770
rect 29314 30718 29710 30770
rect 29762 30718 29764 30770
rect 29260 30716 29764 30718
rect 29260 30706 29316 30716
rect 29708 30706 29764 30716
rect 29596 29316 29652 29326
rect 29596 29222 29652 29260
rect 29204 28588 29316 28644
rect 29148 28550 29204 28588
rect 28924 28420 28980 28430
rect 28924 27858 28980 28364
rect 28924 27806 28926 27858
rect 28978 27806 28980 27858
rect 28140 27748 28196 27758
rect 28140 27654 28196 27692
rect 28924 27748 28980 27806
rect 29260 27860 29316 28588
rect 28924 27682 28980 27692
rect 29148 27748 29204 27758
rect 29148 27654 29204 27692
rect 28588 27634 28644 27646
rect 28588 27582 28590 27634
rect 28642 27582 28644 27634
rect 28588 27300 28644 27582
rect 28588 27234 28644 27244
rect 26572 26450 26628 26460
rect 26460 26402 26516 26414
rect 26460 26350 26462 26402
rect 26514 26350 26516 26402
rect 25676 25454 25678 25506
rect 25730 25454 25732 25506
rect 25676 25442 25732 25454
rect 26236 26290 26292 26302
rect 26236 26238 26238 26290
rect 26290 26238 26292 26290
rect 25340 25282 25396 25294
rect 25340 25230 25342 25282
rect 25394 25230 25396 25282
rect 25340 24836 25396 25230
rect 25340 24770 25396 24780
rect 25228 24724 25284 24734
rect 25228 24630 25284 24668
rect 26236 24162 26292 26238
rect 26460 25618 26516 26350
rect 26460 25566 26462 25618
rect 26514 25566 26516 25618
rect 26460 25554 26516 25566
rect 28588 25618 28644 25630
rect 28588 25566 28590 25618
rect 28642 25566 28644 25618
rect 28588 25172 28644 25566
rect 29260 25506 29316 27804
rect 29596 27076 29652 27086
rect 29596 26982 29652 27020
rect 29260 25454 29262 25506
rect 29314 25454 29316 25506
rect 29260 25442 29316 25454
rect 26236 24110 26238 24162
rect 26290 24110 26292 24162
rect 26236 24098 26292 24110
rect 28364 25116 28588 25172
rect 23324 22316 23828 22372
rect 23772 22260 23828 22316
rect 24556 22370 24836 22372
rect 24556 22318 24782 22370
rect 24834 22318 24836 22370
rect 24556 22316 24836 22318
rect 23772 22258 23940 22260
rect 23772 22206 23774 22258
rect 23826 22206 23940 22258
rect 23772 22204 23940 22206
rect 23772 22194 23828 22204
rect 23660 22148 23716 22158
rect 23548 22036 23604 22046
rect 23548 21476 23604 21980
rect 23660 21700 23716 22092
rect 23660 21644 23828 21700
rect 23660 21476 23716 21486
rect 23548 21474 23716 21476
rect 23548 21422 23662 21474
rect 23714 21422 23716 21474
rect 23548 21420 23716 21422
rect 23660 21410 23716 21420
rect 23436 20804 23492 20814
rect 23660 20804 23716 20814
rect 23492 20802 23716 20804
rect 23492 20750 23662 20802
rect 23714 20750 23716 20802
rect 23492 20748 23716 20750
rect 23436 20710 23492 20748
rect 23660 20738 23716 20748
rect 23324 20578 23380 20590
rect 23324 20526 23326 20578
rect 23378 20526 23380 20578
rect 23324 20356 23380 20526
rect 23324 20290 23380 20300
rect 23436 20468 23492 20478
rect 23436 17556 23492 20412
rect 23772 18340 23828 21644
rect 23884 20580 23940 22204
rect 23884 20486 23940 20524
rect 23996 21924 24052 21934
rect 23996 20690 24052 21868
rect 24556 21810 24612 22316
rect 24780 22306 24836 22316
rect 25004 24050 25060 24062
rect 25004 23998 25006 24050
rect 25058 23998 25060 24050
rect 25004 21924 25060 23998
rect 25452 23940 25508 23950
rect 25452 23846 25508 23884
rect 25676 23940 25732 23950
rect 25676 23846 25732 23884
rect 26684 23940 26740 23950
rect 26684 23846 26740 23884
rect 28364 23938 28420 25116
rect 28588 25106 28644 25116
rect 29820 24834 29876 32508
rect 29932 32498 29988 32508
rect 30604 32004 30660 32014
rect 30156 31892 30212 31902
rect 30156 31798 30212 31836
rect 30604 31778 30660 31948
rect 30604 31726 30606 31778
rect 30658 31726 30660 31778
rect 30044 31556 30100 31566
rect 30044 31462 30100 31500
rect 30268 31556 30324 31566
rect 29932 31332 29988 31342
rect 29932 30994 29988 31276
rect 30268 31332 30324 31500
rect 30604 31332 30660 31726
rect 30716 31668 30772 33180
rect 30828 33142 30884 33180
rect 31164 33236 31220 33246
rect 31052 33122 31108 33134
rect 31052 33070 31054 33122
rect 31106 33070 31108 33122
rect 31052 33012 31108 33070
rect 31052 32946 31108 32956
rect 31052 32676 31108 32686
rect 31052 32450 31108 32620
rect 31052 32398 31054 32450
rect 31106 32398 31108 32450
rect 31052 32386 31108 32398
rect 31164 31778 31220 33180
rect 31164 31726 31166 31778
rect 31218 31726 31220 31778
rect 30940 31668 30996 31678
rect 30716 31666 30996 31668
rect 30716 31614 30942 31666
rect 30994 31614 30996 31666
rect 30716 31612 30996 31614
rect 30828 31444 30884 31454
rect 30604 31276 30772 31332
rect 30268 31266 30324 31276
rect 30156 31220 30212 31230
rect 30156 31126 30212 31164
rect 29932 30942 29934 30994
rect 29986 30942 29988 30994
rect 29932 30930 29988 30942
rect 30380 30994 30436 31006
rect 30380 30942 30382 30994
rect 30434 30942 30436 30994
rect 30268 30884 30324 30894
rect 30268 30790 30324 30828
rect 30380 30660 30436 30942
rect 30268 30604 30436 30660
rect 30492 30996 30548 31006
rect 30268 30100 30324 30604
rect 30380 30436 30436 30446
rect 30492 30436 30548 30940
rect 30380 30434 30548 30436
rect 30380 30382 30382 30434
rect 30434 30382 30548 30434
rect 30380 30380 30548 30382
rect 30604 30884 30660 30894
rect 30380 30370 30436 30380
rect 30492 30212 30548 30222
rect 30604 30212 30660 30828
rect 30492 30210 30660 30212
rect 30492 30158 30494 30210
rect 30546 30158 30660 30210
rect 30492 30156 30660 30158
rect 30492 30146 30548 30156
rect 30268 30034 30324 30044
rect 30380 29988 30436 29998
rect 30716 29988 30772 31276
rect 30828 31218 30884 31388
rect 30828 31166 30830 31218
rect 30882 31166 30884 31218
rect 30828 31154 30884 31166
rect 30940 30100 30996 31612
rect 31164 31444 31220 31726
rect 31276 32004 31332 33404
rect 31388 33012 31444 34076
rect 32060 34038 32116 34076
rect 32508 33458 32564 35532
rect 32732 34916 32788 36542
rect 33180 36258 33236 37772
rect 33180 36206 33182 36258
rect 33234 36206 33236 36258
rect 33180 35700 33236 36206
rect 33404 35700 33460 35710
rect 33180 35698 33460 35700
rect 33180 35646 33406 35698
rect 33458 35646 33460 35698
rect 33180 35644 33460 35646
rect 33404 35588 33460 35644
rect 33404 35522 33460 35532
rect 32844 34916 32900 34926
rect 32732 34914 33460 34916
rect 32732 34862 32846 34914
rect 32898 34862 33460 34914
rect 32732 34860 33460 34862
rect 32844 34850 32900 34860
rect 32620 34804 32676 34814
rect 32620 34710 32676 34748
rect 33180 34692 33236 34702
rect 33236 34636 33348 34692
rect 33180 34626 33236 34636
rect 32508 33406 32510 33458
rect 32562 33406 32564 33458
rect 32508 33394 32564 33406
rect 33180 34018 33236 34030
rect 33180 33966 33182 34018
rect 33234 33966 33236 34018
rect 33180 33348 33236 33966
rect 33180 33282 33236 33292
rect 33292 33460 33348 34636
rect 33404 34130 33460 34860
rect 33404 34078 33406 34130
rect 33458 34078 33460 34130
rect 33404 34066 33460 34078
rect 31388 32946 31444 32956
rect 32844 33012 32900 33022
rect 31612 32564 31668 32574
rect 31276 31780 31332 31948
rect 31500 32004 31556 32014
rect 31500 31910 31556 31948
rect 31388 31780 31444 31790
rect 31276 31778 31444 31780
rect 31276 31726 31390 31778
rect 31442 31726 31444 31778
rect 31276 31724 31444 31726
rect 31388 31714 31444 31724
rect 31500 31780 31556 31790
rect 31164 31378 31220 31388
rect 30940 30034 30996 30044
rect 31052 30994 31108 31006
rect 31052 30942 31054 30994
rect 31106 30942 31108 30994
rect 30380 29986 30772 29988
rect 30380 29934 30382 29986
rect 30434 29934 30772 29986
rect 30380 29932 30772 29934
rect 30380 29922 30436 29932
rect 31052 29316 31108 30942
rect 31500 30884 31556 31724
rect 31612 31778 31668 32508
rect 31612 31726 31614 31778
rect 31666 31726 31668 31778
rect 31612 31714 31668 31726
rect 32060 31666 32116 31678
rect 32060 31614 32062 31666
rect 32114 31614 32116 31666
rect 32060 31220 32116 31614
rect 32844 31666 32900 32956
rect 33292 32564 33348 33404
rect 33516 32900 33572 39116
rect 33628 35028 33684 40124
rect 33740 39956 33796 39966
rect 33740 38946 33796 39900
rect 34412 39732 34468 40126
rect 34188 39676 34412 39732
rect 34188 39060 34244 39676
rect 34412 39666 34468 39676
rect 33740 38894 33742 38946
rect 33794 38894 33796 38946
rect 33740 38882 33796 38894
rect 33852 38948 33908 38958
rect 33852 38854 33908 38892
rect 33964 38948 34020 38958
rect 34188 38948 34244 39004
rect 33964 38946 34244 38948
rect 33964 38894 33966 38946
rect 34018 38894 34244 38946
rect 33964 38892 34244 38894
rect 34300 39508 34356 39518
rect 34524 39508 34580 42028
rect 34636 41524 34692 43372
rect 34748 42196 34804 42206
rect 34748 42102 34804 42140
rect 35084 42194 35140 43486
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35084 42142 35086 42194
rect 35138 42142 35140 42194
rect 35084 42130 35140 42142
rect 35420 42308 35476 42318
rect 35420 41972 35476 42252
rect 35980 42196 36036 45838
rect 39228 45892 39284 45902
rect 40460 45892 40516 45902
rect 38220 45780 38276 45790
rect 36988 45108 37044 45118
rect 36876 45106 37044 45108
rect 36876 45054 36990 45106
rect 37042 45054 37044 45106
rect 36876 45052 37044 45054
rect 36428 44884 36484 44894
rect 36428 44790 36484 44828
rect 36764 44772 36820 44782
rect 36540 44716 36764 44772
rect 36540 44660 36596 44716
rect 36764 44706 36820 44716
rect 36204 44604 36596 44660
rect 36204 44546 36260 44604
rect 36204 44494 36206 44546
rect 36258 44494 36260 44546
rect 36204 44482 36260 44494
rect 36204 42980 36260 42990
rect 36204 42886 36260 42924
rect 35980 42130 36036 42140
rect 35868 41972 35924 41982
rect 35420 41970 35588 41972
rect 35420 41918 35422 41970
rect 35474 41918 35588 41970
rect 35420 41916 35588 41918
rect 35420 41906 35476 41916
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 34636 41468 34804 41524
rect 35196 41514 35460 41524
rect 34636 41298 34692 41310
rect 34636 41246 34638 41298
rect 34690 41246 34692 41298
rect 34636 41188 34692 41246
rect 34636 40514 34692 41132
rect 34636 40462 34638 40514
rect 34690 40462 34692 40514
rect 34636 40450 34692 40462
rect 34300 39506 34580 39508
rect 34300 39454 34302 39506
rect 34354 39454 34580 39506
rect 34300 39452 34580 39454
rect 33964 38882 34020 38892
rect 34300 38668 34356 39452
rect 34636 39396 34692 39406
rect 34524 39340 34636 39396
rect 34524 39058 34580 39340
rect 34636 39330 34692 39340
rect 34524 39006 34526 39058
rect 34578 39006 34580 39058
rect 34524 38994 34580 39006
rect 34300 38612 34692 38668
rect 33964 37940 34020 37950
rect 33964 37846 34020 37884
rect 34188 35588 34244 35598
rect 34188 35586 34580 35588
rect 34188 35534 34190 35586
rect 34242 35534 34580 35586
rect 34188 35532 34580 35534
rect 34188 35522 34244 35532
rect 33740 35028 33796 35038
rect 33628 35026 33796 35028
rect 33628 34974 33742 35026
rect 33794 34974 33796 35026
rect 33628 34972 33796 34974
rect 33740 34962 33796 34972
rect 34524 35026 34580 35532
rect 34636 35476 34692 38612
rect 34748 35700 34804 41468
rect 35532 41412 35588 41916
rect 35868 41970 36036 41972
rect 35868 41918 35870 41970
rect 35922 41918 36036 41970
rect 35868 41916 36036 41918
rect 35868 41906 35924 41916
rect 35420 41356 35588 41412
rect 35084 41186 35140 41198
rect 35084 41134 35086 41186
rect 35138 41134 35140 41186
rect 35084 40964 35140 41134
rect 34860 40908 35084 40964
rect 35420 40964 35476 41356
rect 35532 41188 35588 41198
rect 35532 41094 35588 41132
rect 35420 40908 35588 40964
rect 34860 39844 34916 40908
rect 35084 40898 35140 40908
rect 35084 40628 35140 40638
rect 35084 40402 35140 40572
rect 35084 40350 35086 40402
rect 35138 40350 35140 40402
rect 35084 40338 35140 40350
rect 35308 40402 35364 40414
rect 35308 40350 35310 40402
rect 35362 40350 35364 40402
rect 35308 40180 35364 40350
rect 35420 40404 35476 40414
rect 35420 40310 35476 40348
rect 34860 39730 34916 39788
rect 34860 39678 34862 39730
rect 34914 39678 34916 39730
rect 34860 39666 34916 39678
rect 35084 40124 35364 40180
rect 34860 37940 34916 37950
rect 34916 37884 35028 37940
rect 34860 37874 34916 37884
rect 34972 37490 35028 37884
rect 34972 37438 34974 37490
rect 35026 37438 35028 37490
rect 34972 37426 35028 37438
rect 34748 35634 34804 35644
rect 34860 37266 34916 37278
rect 34860 37214 34862 37266
rect 34914 37214 34916 37266
rect 34636 35420 34804 35476
rect 34524 34974 34526 35026
rect 34578 34974 34580 35026
rect 34524 34962 34580 34974
rect 34636 34914 34692 34926
rect 34636 34862 34638 34914
rect 34690 34862 34692 34914
rect 34412 34804 34468 34814
rect 34412 34710 34468 34748
rect 33852 34690 33908 34702
rect 33852 34638 33854 34690
rect 33906 34638 33908 34690
rect 33852 34580 33908 34638
rect 34636 34580 34692 34862
rect 33852 34524 34692 34580
rect 33628 34132 33684 34142
rect 33628 34038 33684 34076
rect 34076 33908 34132 33918
rect 33964 33906 34132 33908
rect 33964 33854 34078 33906
rect 34130 33854 34132 33906
rect 33964 33852 34132 33854
rect 33628 33572 33684 33582
rect 33628 33346 33684 33516
rect 33628 33294 33630 33346
rect 33682 33294 33684 33346
rect 33628 33124 33684 33294
rect 33628 33058 33684 33068
rect 33516 32834 33572 32844
rect 33292 32470 33348 32508
rect 33516 32564 33572 32574
rect 33516 32470 33572 32508
rect 33068 32450 33124 32462
rect 33068 32398 33070 32450
rect 33122 32398 33124 32450
rect 33068 31780 33124 32398
rect 33964 31892 34020 33852
rect 34076 33842 34132 33852
rect 34412 33572 34468 33582
rect 33964 31826 34020 31836
rect 34076 33570 34468 33572
rect 34076 33518 34414 33570
rect 34466 33518 34468 33570
rect 34076 33516 34468 33518
rect 33068 31686 33124 31724
rect 33740 31778 33796 31790
rect 33740 31726 33742 31778
rect 33794 31726 33796 31778
rect 32844 31614 32846 31666
rect 32898 31614 32900 31666
rect 32844 31602 32900 31614
rect 32508 31556 32564 31566
rect 32396 31554 32564 31556
rect 32396 31502 32510 31554
rect 32562 31502 32564 31554
rect 32396 31500 32564 31502
rect 32396 31444 32452 31500
rect 32508 31490 32564 31500
rect 33292 31556 33348 31566
rect 32116 31164 32228 31220
rect 32060 31154 32116 31164
rect 31500 30818 31556 30828
rect 31500 30100 31556 30110
rect 31500 30006 31556 30044
rect 32172 30098 32228 31164
rect 32172 30046 32174 30098
rect 32226 30046 32228 30098
rect 32172 30034 32228 30046
rect 31836 29986 31892 29998
rect 31836 29934 31838 29986
rect 31890 29934 31892 29986
rect 31836 29764 31892 29934
rect 31836 29698 31892 29708
rect 32172 29652 32228 29662
rect 32396 29652 32452 31388
rect 33292 30322 33348 31500
rect 33740 31444 33796 31726
rect 34076 31778 34132 33516
rect 34412 33506 34468 33516
rect 34636 33348 34692 34524
rect 34748 34468 34804 35420
rect 34860 34804 34916 37214
rect 35084 37266 35140 40124
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35308 39396 35364 39406
rect 35532 39396 35588 40908
rect 35644 40962 35700 40974
rect 35644 40910 35646 40962
rect 35698 40910 35700 40962
rect 35644 40628 35700 40910
rect 35644 40562 35700 40572
rect 35756 40962 35812 40974
rect 35756 40910 35758 40962
rect 35810 40910 35812 40962
rect 35308 39394 35588 39396
rect 35308 39342 35310 39394
rect 35362 39342 35588 39394
rect 35308 39340 35588 39342
rect 35644 40404 35700 40414
rect 35308 38668 35364 39340
rect 35644 39284 35700 40348
rect 35756 40292 35812 40910
rect 35756 40226 35812 40236
rect 35980 39842 36036 41916
rect 36540 41860 36596 41870
rect 36540 41766 36596 41804
rect 36876 41412 36932 45052
rect 36988 45042 37044 45052
rect 37772 45106 37828 45118
rect 37772 45054 37774 45106
rect 37826 45054 37828 45106
rect 37772 44548 37828 45054
rect 38220 44548 38276 45724
rect 38892 45778 38948 45790
rect 38892 45726 38894 45778
rect 38946 45726 38948 45778
rect 37772 44482 37828 44492
rect 37884 44492 38276 44548
rect 37548 44322 37604 44334
rect 37548 44270 37550 44322
rect 37602 44270 37604 44322
rect 37100 44098 37156 44110
rect 37100 44046 37102 44098
rect 37154 44046 37156 44098
rect 36988 43876 37044 43886
rect 36988 42530 37044 43820
rect 37100 43204 37156 44046
rect 37548 43988 37604 44270
rect 37772 44212 37828 44222
rect 37772 44118 37828 44156
rect 37884 43988 37940 44492
rect 37548 43932 37940 43988
rect 37996 44324 38052 44334
rect 37436 43428 37492 43438
rect 37212 43316 37268 43326
rect 37212 43222 37268 43260
rect 37100 43138 37156 43148
rect 37436 43204 37492 43372
rect 36988 42478 36990 42530
rect 37042 42478 37044 42530
rect 36988 42084 37044 42478
rect 37324 42530 37380 42542
rect 37324 42478 37326 42530
rect 37378 42478 37380 42530
rect 37324 42420 37380 42478
rect 37436 42420 37492 43148
rect 37660 42754 37716 43932
rect 37660 42702 37662 42754
rect 37714 42702 37716 42754
rect 37660 42690 37716 42702
rect 37772 43538 37828 43550
rect 37772 43486 37774 43538
rect 37826 43486 37828 43538
rect 37772 42644 37828 43486
rect 37772 42578 37828 42588
rect 37996 42642 38052 44268
rect 37996 42590 37998 42642
rect 38050 42590 38052 42642
rect 37996 42578 38052 42590
rect 38220 44322 38276 44492
rect 38220 44270 38222 44322
rect 38274 44270 38276 44322
rect 38220 42532 38276 44270
rect 38444 45108 38500 45118
rect 38444 44210 38500 45052
rect 38444 44158 38446 44210
rect 38498 44158 38500 44210
rect 38444 44146 38500 44158
rect 38780 44322 38836 44334
rect 38780 44270 38782 44322
rect 38834 44270 38836 44322
rect 38780 44100 38836 44270
rect 38780 44034 38836 44044
rect 38332 43652 38388 43662
rect 38332 42754 38388 43596
rect 38892 43652 38948 45726
rect 39228 45778 39284 45836
rect 40124 45890 40516 45892
rect 40124 45838 40462 45890
rect 40514 45838 40516 45890
rect 40124 45836 40516 45838
rect 39228 45726 39230 45778
rect 39282 45726 39284 45778
rect 39228 45714 39284 45726
rect 39788 45780 39844 45790
rect 39788 45686 39844 45724
rect 40124 45778 40180 45836
rect 40460 45826 40516 45836
rect 40124 45726 40126 45778
rect 40178 45726 40180 45778
rect 40124 45714 40180 45726
rect 41020 45332 41076 49200
rect 41468 46116 41524 46126
rect 41468 46022 41524 46060
rect 41692 46116 41748 49200
rect 41692 46050 41748 46060
rect 41020 45266 41076 45276
rect 42252 45332 42308 45342
rect 42252 45238 42308 45276
rect 41132 45220 41188 45230
rect 40124 44884 40180 44894
rect 40124 44790 40180 44828
rect 41132 44546 41188 45164
rect 41132 44494 41134 44546
rect 41186 44494 41188 44546
rect 41132 44482 41188 44494
rect 41244 45106 41300 45118
rect 41244 45054 41246 45106
rect 41298 45054 41300 45106
rect 41244 44212 41300 45054
rect 42364 44996 42420 49200
rect 42364 44930 42420 44940
rect 43036 44548 43092 49200
rect 43708 46900 43764 49200
rect 44044 47796 44100 47806
rect 43708 46844 43876 46900
rect 43708 45892 43764 45902
rect 43708 45798 43764 45836
rect 43036 44482 43092 44492
rect 43820 44434 43876 46844
rect 43820 44382 43822 44434
rect 43874 44382 43876 44434
rect 43820 44370 43876 44382
rect 43932 44436 43988 44446
rect 41692 44324 41748 44334
rect 41692 44230 41748 44268
rect 41244 44146 41300 44156
rect 42812 44212 42868 44222
rect 38892 43586 38948 43596
rect 41244 43652 41300 43662
rect 38332 42702 38334 42754
rect 38386 42702 38388 42754
rect 38332 42690 38388 42702
rect 38668 43540 38724 43550
rect 38668 42642 38724 43484
rect 41244 43538 41300 43596
rect 41244 43486 41246 43538
rect 41298 43486 41300 43538
rect 41244 43428 41300 43486
rect 41244 43362 41300 43372
rect 41468 43650 41524 43662
rect 41468 43598 41470 43650
rect 41522 43598 41524 43650
rect 40124 43314 40180 43326
rect 40124 43262 40126 43314
rect 40178 43262 40180 43314
rect 40124 43092 40180 43262
rect 40124 43026 40180 43036
rect 39004 42756 39060 42766
rect 38668 42590 38670 42642
rect 38722 42590 38724 42642
rect 38668 42578 38724 42590
rect 38892 42754 39060 42756
rect 38892 42702 39006 42754
rect 39058 42702 39060 42754
rect 38892 42700 39060 42702
rect 38220 42476 38500 42532
rect 37324 42364 37940 42420
rect 36988 42028 37492 42084
rect 37100 41860 37156 41870
rect 36876 41356 37044 41412
rect 36204 41188 36260 41198
rect 36428 41188 36484 41198
rect 36204 41186 36372 41188
rect 36204 41134 36206 41186
rect 36258 41134 36372 41186
rect 36204 41132 36372 41134
rect 36204 41122 36260 41132
rect 36204 40402 36260 40414
rect 36204 40350 36206 40402
rect 36258 40350 36260 40402
rect 36204 40292 36260 40350
rect 36204 40226 36260 40236
rect 35980 39790 35982 39842
rect 36034 39790 36036 39842
rect 35980 39730 36036 39790
rect 35980 39678 35982 39730
rect 36034 39678 36036 39730
rect 35980 39666 36036 39678
rect 36316 39732 36372 41132
rect 36428 41074 36484 41132
rect 36428 41022 36430 41074
rect 36482 41022 36484 41074
rect 36428 41010 36484 41022
rect 36876 41186 36932 41198
rect 36876 41134 36878 41186
rect 36930 41134 36932 41186
rect 36540 40516 36596 40526
rect 36876 40516 36932 41134
rect 36988 40628 37044 41356
rect 37100 41298 37156 41804
rect 37100 41246 37102 41298
rect 37154 41246 37156 41298
rect 37100 41234 37156 41246
rect 37324 41074 37380 41086
rect 37324 41022 37326 41074
rect 37378 41022 37380 41074
rect 37100 40628 37156 40638
rect 36988 40626 37156 40628
rect 36988 40574 37102 40626
rect 37154 40574 37156 40626
rect 36988 40572 37156 40574
rect 37100 40562 37156 40572
rect 36540 40514 36932 40516
rect 36540 40462 36542 40514
rect 36594 40462 36932 40514
rect 36540 40460 36932 40462
rect 36540 40404 36596 40460
rect 36540 40338 36596 40348
rect 36988 40292 37044 40302
rect 36540 39842 36596 39854
rect 36540 39790 36542 39842
rect 36594 39790 36596 39842
rect 36428 39732 36484 39742
rect 36316 39730 36484 39732
rect 36316 39678 36430 39730
rect 36482 39678 36484 39730
rect 36316 39676 36484 39678
rect 35644 39218 35700 39228
rect 36428 38668 36484 39676
rect 36540 39060 36596 39790
rect 36988 39618 37044 40236
rect 37324 39956 37380 41022
rect 37436 40404 37492 42028
rect 37772 41972 37828 41982
rect 37548 41860 37604 41870
rect 37548 41186 37604 41804
rect 37548 41134 37550 41186
rect 37602 41134 37604 41186
rect 37548 41122 37604 41134
rect 37436 40310 37492 40348
rect 37772 40402 37828 41916
rect 37772 40350 37774 40402
rect 37826 40350 37828 40402
rect 37772 40338 37828 40350
rect 36988 39566 36990 39618
rect 37042 39566 37044 39618
rect 36652 39060 36708 39070
rect 36540 39004 36652 39060
rect 36652 38966 36708 39004
rect 36988 38946 37044 39566
rect 36988 38894 36990 38946
rect 37042 38894 37044 38946
rect 36988 38836 37044 38894
rect 36988 38770 37044 38780
rect 37100 39900 37380 39956
rect 35308 38612 35588 38668
rect 36428 38612 36596 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35532 38276 35588 38612
rect 35084 37214 35086 37266
rect 35138 37214 35140 37266
rect 35084 37156 35140 37214
rect 35084 37090 35140 37100
rect 35308 38220 35588 38276
rect 35308 37044 35364 38220
rect 36092 38164 36148 38174
rect 36148 38108 36260 38164
rect 36092 38070 36148 38108
rect 36092 37492 36148 37502
rect 36092 37398 36148 37436
rect 36204 37490 36260 38108
rect 36204 37438 36206 37490
rect 36258 37438 36260 37490
rect 36204 37426 36260 37438
rect 35420 37380 35476 37390
rect 35420 37286 35476 37324
rect 35980 37268 36036 37278
rect 35980 37174 36036 37212
rect 35644 37156 35700 37166
rect 35308 36988 35588 37044
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 34972 35588 35028 35598
rect 34972 34914 35028 35532
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34972 34862 34974 34914
rect 35026 34862 35028 34914
rect 34972 34850 35028 34862
rect 35532 34916 35588 36988
rect 35644 36594 35700 37100
rect 35644 36542 35646 36594
rect 35698 36542 35700 36594
rect 35644 36530 35700 36542
rect 35756 36370 35812 36382
rect 35756 36318 35758 36370
rect 35810 36318 35812 36370
rect 35756 35924 35812 36318
rect 36540 36148 36596 38612
rect 36988 38164 37044 38174
rect 36988 38070 37044 38108
rect 37100 37826 37156 39900
rect 37772 39844 37828 39854
rect 37772 39730 37828 39788
rect 37772 39678 37774 39730
rect 37826 39678 37828 39730
rect 37324 39396 37380 39406
rect 37324 39302 37380 39340
rect 37100 37774 37102 37826
rect 37154 37774 37156 37826
rect 36652 37268 36708 37278
rect 36652 37266 36932 37268
rect 36652 37214 36654 37266
rect 36706 37214 36932 37266
rect 36652 37212 36932 37214
rect 36652 37202 36708 37212
rect 36876 36484 36932 37212
rect 37100 36932 37156 37774
rect 37212 39060 37268 39070
rect 37212 37266 37268 39004
rect 37772 39060 37828 39678
rect 37772 38994 37828 39004
rect 37324 38834 37380 38846
rect 37324 38782 37326 38834
rect 37378 38782 37380 38834
rect 37324 38668 37380 38782
rect 37660 38834 37716 38846
rect 37660 38782 37662 38834
rect 37714 38782 37716 38834
rect 37660 38668 37716 38782
rect 37324 38612 37716 38668
rect 37884 38668 37940 42364
rect 38108 41748 38164 41758
rect 38108 41186 38164 41692
rect 38108 41134 38110 41186
rect 38162 41134 38164 41186
rect 38108 41122 38164 41134
rect 38444 41074 38500 42476
rect 38668 42196 38724 42206
rect 38668 41858 38724 42140
rect 38668 41806 38670 41858
rect 38722 41806 38724 41858
rect 38668 41794 38724 41806
rect 38892 41636 38948 42700
rect 39004 42690 39060 42700
rect 39228 42644 39284 42654
rect 39228 42196 39284 42588
rect 39228 42102 39284 42140
rect 39788 42642 39844 42654
rect 39788 42590 39790 42642
rect 39842 42590 39844 42642
rect 39004 42084 39060 42094
rect 39004 41990 39060 42028
rect 39676 41970 39732 41982
rect 39676 41918 39678 41970
rect 39730 41918 39732 41970
rect 39116 41860 39172 41870
rect 39116 41766 39172 41804
rect 38444 41022 38446 41074
rect 38498 41022 38500 41074
rect 38444 41010 38500 41022
rect 38668 41580 38948 41636
rect 39676 41748 39732 41918
rect 39788 41972 39844 42590
rect 39788 41906 39844 41916
rect 40124 42532 40180 42542
rect 40124 41970 40180 42476
rect 41132 42308 41188 42318
rect 40124 41918 40126 41970
rect 40178 41918 40180 41970
rect 40124 41906 40180 41918
rect 40348 42082 40404 42094
rect 40348 42030 40350 42082
rect 40402 42030 40404 42082
rect 40348 41860 40404 42030
rect 40348 41794 40404 41804
rect 40796 42084 40852 42094
rect 38108 39620 38164 39630
rect 38668 39620 38724 41580
rect 39452 41524 39508 41534
rect 38780 41188 38836 41198
rect 38780 41094 38836 41132
rect 39452 40514 39508 41468
rect 39452 40462 39454 40514
rect 39506 40462 39508 40514
rect 39452 40450 39508 40462
rect 39676 40180 39732 41692
rect 40684 40628 40740 40638
rect 40460 40572 40684 40628
rect 39676 40114 39732 40124
rect 40236 40404 40292 40414
rect 40012 39844 40068 39854
rect 38108 39618 38836 39620
rect 38108 39566 38110 39618
rect 38162 39566 38836 39618
rect 38108 39564 38836 39566
rect 38108 39172 38164 39564
rect 38108 39106 38164 39116
rect 38444 39060 38500 39070
rect 37996 38948 38052 38958
rect 37996 38854 38052 38892
rect 38332 38836 38388 38846
rect 38332 38742 38388 38780
rect 38444 38668 38500 39004
rect 38668 39060 38724 39070
rect 38668 38966 38724 39004
rect 38780 38668 38836 39564
rect 38892 39508 38948 39518
rect 38892 39506 39508 39508
rect 38892 39454 38894 39506
rect 38946 39454 39508 39506
rect 38892 39452 39508 39454
rect 38892 39442 38948 39452
rect 39340 39284 39396 39294
rect 39340 38946 39396 39228
rect 39452 39058 39508 39452
rect 39452 39006 39454 39058
rect 39506 39006 39508 39058
rect 39452 38994 39508 39006
rect 39340 38894 39342 38946
rect 39394 38894 39396 38946
rect 39340 38882 39396 38894
rect 39676 38834 39732 38846
rect 39676 38782 39678 38834
rect 39730 38782 39732 38834
rect 37884 38612 38164 38668
rect 38444 38612 38612 38668
rect 38780 38612 38948 38668
rect 37212 37214 37214 37266
rect 37266 37214 37268 37266
rect 37212 37202 37268 37214
rect 37324 36932 37380 36942
rect 37100 36876 37324 36932
rect 37324 36866 37380 36876
rect 36876 36428 37156 36484
rect 37100 36260 37156 36428
rect 36540 36092 37044 36148
rect 36316 35924 36372 35934
rect 35756 35868 36316 35924
rect 36316 35586 36372 35868
rect 36876 35924 36932 35934
rect 36876 35830 36932 35868
rect 36316 35534 36318 35586
rect 36370 35534 36372 35586
rect 36316 35522 36372 35534
rect 36652 35812 36708 35822
rect 35644 34916 35700 34926
rect 35532 34860 35644 34916
rect 35644 34850 35700 34860
rect 34860 34738 34916 34748
rect 34748 34402 34804 34412
rect 36652 34356 36708 35756
rect 36988 35700 37044 36092
rect 37100 35922 37156 36204
rect 37100 35870 37102 35922
rect 37154 35870 37156 35922
rect 37100 35858 37156 35870
rect 36876 35644 37044 35700
rect 36764 35588 36820 35598
rect 36764 35494 36820 35532
rect 36652 34290 36708 34300
rect 36764 34018 36820 34030
rect 36764 33966 36766 34018
rect 36818 33966 36820 34018
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 36764 33684 36820 33966
rect 36876 33796 36932 35644
rect 37212 34914 37268 34926
rect 37212 34862 37214 34914
rect 37266 34862 37268 34914
rect 36988 34692 37044 34702
rect 36988 34598 37044 34636
rect 36876 33730 36932 33740
rect 37212 34130 37268 34862
rect 37436 34356 37492 34366
rect 37436 34262 37492 34300
rect 37212 34078 37214 34130
rect 37266 34078 37268 34130
rect 36764 33618 36820 33628
rect 34412 33292 34692 33348
rect 34748 33460 34804 33470
rect 34748 33346 34804 33404
rect 34972 33348 35028 33358
rect 34748 33294 34750 33346
rect 34802 33294 34804 33346
rect 34300 33236 34356 33246
rect 34300 33142 34356 33180
rect 34076 31726 34078 31778
rect 34130 31726 34132 31778
rect 34076 31714 34132 31726
rect 33740 30884 33796 31388
rect 33740 30818 33796 30828
rect 33964 31666 34020 31678
rect 33964 31614 33966 31666
rect 34018 31614 34020 31666
rect 33964 30548 34020 31614
rect 33964 30492 34244 30548
rect 34188 30436 34244 30492
rect 34188 30434 34356 30436
rect 34188 30382 34190 30434
rect 34242 30382 34356 30434
rect 34188 30380 34356 30382
rect 34188 30370 34244 30380
rect 33292 30270 33294 30322
rect 33346 30270 33348 30322
rect 33292 30258 33348 30270
rect 32508 30212 32564 30222
rect 32508 30118 32564 30156
rect 32844 30210 32900 30222
rect 32844 30158 32846 30210
rect 32898 30158 32900 30210
rect 32844 30100 32900 30158
rect 32844 30034 32900 30044
rect 33068 30212 33124 30222
rect 32172 29650 32452 29652
rect 32172 29598 32174 29650
rect 32226 29598 32452 29650
rect 32172 29596 32452 29598
rect 32508 29764 32564 29774
rect 32172 29586 32228 29596
rect 32284 29428 32340 29438
rect 32508 29428 32564 29708
rect 33068 29650 33124 30156
rect 33068 29598 33070 29650
rect 33122 29598 33124 29650
rect 33068 29586 33124 29598
rect 33740 30210 33796 30222
rect 33740 30158 33742 30210
rect 33794 30158 33796 30210
rect 32284 29426 32564 29428
rect 32284 29374 32286 29426
rect 32338 29374 32564 29426
rect 32284 29372 32564 29374
rect 32284 29362 32340 29372
rect 31052 29250 31108 29260
rect 33180 29316 33236 29326
rect 33180 29222 33236 29260
rect 33740 29316 33796 30158
rect 34300 29876 34356 30380
rect 34412 30100 34468 33292
rect 34748 33282 34804 33294
rect 34860 33292 34972 33348
rect 34524 33122 34580 33134
rect 34524 33070 34526 33122
rect 34578 33070 34580 33122
rect 34524 33012 34580 33070
rect 34524 32946 34580 32956
rect 34860 32450 34916 33292
rect 34972 33254 35028 33292
rect 36316 33348 36372 33358
rect 36316 33254 36372 33292
rect 35308 33236 35364 33246
rect 34860 32398 34862 32450
rect 34914 32398 34916 32450
rect 34860 32386 34916 32398
rect 35084 33234 35364 33236
rect 35084 33182 35310 33234
rect 35362 33182 35364 33234
rect 35084 33180 35364 33182
rect 34972 31892 35028 31902
rect 35084 31892 35140 33180
rect 35308 33170 35364 33180
rect 35532 33236 35588 33246
rect 35532 32564 35588 33180
rect 35868 33234 35924 33246
rect 35868 33182 35870 33234
rect 35922 33182 35924 33234
rect 35756 33124 35812 33134
rect 35756 33030 35812 33068
rect 35532 32498 35588 32508
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35868 32004 35924 33182
rect 36204 33236 36260 33246
rect 36204 33142 36260 33180
rect 36988 33124 37044 33134
rect 36988 32674 37044 33068
rect 37212 32788 37268 34078
rect 37268 32732 37492 32788
rect 37212 32722 37268 32732
rect 36988 32622 36990 32674
rect 37042 32622 37044 32674
rect 36988 32610 37044 32622
rect 35868 31938 35924 31948
rect 34972 31890 35140 31892
rect 34972 31838 34974 31890
rect 35026 31838 35140 31890
rect 34972 31836 35140 31838
rect 35532 31892 35588 31902
rect 34972 31826 35028 31836
rect 35532 31778 35588 31836
rect 37100 31892 37156 31902
rect 37100 31798 37156 31836
rect 35532 31726 35534 31778
rect 35586 31726 35588 31778
rect 35532 31714 35588 31726
rect 35644 31780 35700 31790
rect 34524 31556 34580 31566
rect 34860 31556 34916 31566
rect 34524 31554 34916 31556
rect 34524 31502 34526 31554
rect 34578 31502 34862 31554
rect 34914 31502 34916 31554
rect 34524 31500 34916 31502
rect 34524 31490 34580 31500
rect 34860 31490 34916 31500
rect 35084 31556 35140 31566
rect 35084 31462 35140 31500
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34860 30436 34916 30446
rect 34636 30100 34692 30110
rect 34412 30098 34692 30100
rect 34412 30046 34638 30098
rect 34690 30046 34692 30098
rect 34412 30044 34692 30046
rect 34636 30034 34692 30044
rect 34300 29652 34356 29820
rect 34524 29652 34580 29662
rect 34300 29650 34580 29652
rect 34300 29598 34526 29650
rect 34578 29598 34580 29650
rect 34300 29596 34580 29598
rect 34524 29586 34580 29596
rect 34860 29650 34916 30380
rect 35644 30436 35700 31724
rect 36316 31554 36372 31566
rect 36316 31502 36318 31554
rect 36370 31502 36372 31554
rect 36316 31332 36372 31502
rect 35980 31276 36932 31332
rect 35756 31108 35812 31118
rect 35980 31108 36036 31276
rect 35812 31106 36036 31108
rect 35812 31054 35982 31106
rect 36034 31054 36036 31106
rect 35812 31052 36036 31054
rect 35756 31014 35812 31052
rect 35980 31042 36036 31052
rect 36092 31108 36148 31118
rect 36652 31108 36708 31118
rect 36092 31106 36708 31108
rect 36092 31054 36094 31106
rect 36146 31054 36654 31106
rect 36706 31054 36708 31106
rect 36092 31052 36708 31054
rect 36092 31042 36148 31052
rect 36092 30772 36148 30782
rect 36092 30678 36148 30716
rect 35644 30342 35700 30380
rect 35308 30212 35364 30222
rect 35308 30118 35364 30156
rect 34860 29598 34862 29650
rect 34914 29598 34916 29650
rect 34860 29586 34916 29598
rect 35868 30098 35924 30110
rect 35868 30046 35870 30098
rect 35922 30046 35924 30098
rect 35644 29540 35700 29550
rect 35644 29446 35700 29484
rect 35868 29540 35924 30046
rect 36092 30100 36148 30110
rect 36092 30006 36148 30044
rect 35980 29988 36036 29998
rect 35980 29894 36036 29932
rect 35868 29474 35924 29484
rect 36092 29428 36148 29438
rect 36092 29334 36148 29372
rect 33740 29250 33796 29260
rect 32172 29204 32228 29214
rect 32172 29110 32228 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 32060 28756 32116 28766
rect 32060 28754 32228 28756
rect 32060 28702 32062 28754
rect 32114 28702 32228 28754
rect 32060 28700 32228 28702
rect 32060 28690 32116 28700
rect 29932 28530 29988 28542
rect 29932 28478 29934 28530
rect 29986 28478 29988 28530
rect 29932 27970 29988 28478
rect 29932 27918 29934 27970
rect 29986 27918 29988 27970
rect 29932 27906 29988 27918
rect 30380 27748 30436 27758
rect 30380 27654 30436 27692
rect 30828 27748 30884 27758
rect 30828 27654 30884 27692
rect 31388 27748 31444 27758
rect 30044 27634 30100 27646
rect 30044 27582 30046 27634
rect 30098 27582 30100 27634
rect 30044 27076 30100 27582
rect 30268 27634 30324 27646
rect 30268 27582 30270 27634
rect 30322 27582 30324 27634
rect 30044 27010 30100 27020
rect 30156 27524 30212 27534
rect 30156 27074 30212 27468
rect 30268 27186 30324 27582
rect 30492 27636 30548 27646
rect 30492 27298 30548 27580
rect 31164 27636 31220 27646
rect 31164 27542 31220 27580
rect 31388 27524 31444 27692
rect 32172 27748 32228 28700
rect 32396 28082 32452 28094
rect 32396 28030 32398 28082
rect 32450 28030 32452 28082
rect 32396 27972 32452 28030
rect 32396 27906 32452 27916
rect 33852 27972 33908 27982
rect 33852 27878 33908 27916
rect 32172 27682 32228 27692
rect 32508 27858 32564 27870
rect 32508 27806 32510 27858
rect 32562 27806 32564 27858
rect 31388 27458 31444 27468
rect 32060 27634 32116 27646
rect 32060 27582 32062 27634
rect 32114 27582 32116 27634
rect 30492 27246 30494 27298
rect 30546 27246 30548 27298
rect 30492 27234 30548 27246
rect 30268 27134 30270 27186
rect 30322 27134 30324 27186
rect 30268 27122 30324 27134
rect 30156 27022 30158 27074
rect 30210 27022 30212 27074
rect 30156 27010 30212 27022
rect 31612 27076 31668 27086
rect 32060 27076 32116 27582
rect 32284 27634 32340 27646
rect 32284 27582 32286 27634
rect 32338 27582 32340 27634
rect 32284 27412 32340 27582
rect 32508 27636 32564 27806
rect 33068 27860 33124 27870
rect 33124 27804 33460 27860
rect 33068 27766 33124 27804
rect 32508 27570 32564 27580
rect 33180 27636 33236 27646
rect 32284 27356 32788 27412
rect 32732 27298 32788 27356
rect 32732 27246 32734 27298
rect 32786 27246 32788 27298
rect 32732 27234 32788 27246
rect 31668 27020 32116 27076
rect 32844 27076 32900 27086
rect 31612 26982 31668 27020
rect 32844 26962 32900 27020
rect 32844 26910 32846 26962
rect 32898 26910 32900 26962
rect 32844 26898 32900 26910
rect 33068 26962 33124 26974
rect 33068 26910 33070 26962
rect 33122 26910 33124 26962
rect 33068 26908 33124 26910
rect 32956 26852 33124 26908
rect 32508 26404 32564 26414
rect 32172 26292 32228 26302
rect 32508 26292 32564 26348
rect 32172 26198 32228 26236
rect 32396 26290 32564 26292
rect 32396 26238 32510 26290
rect 32562 26238 32564 26290
rect 32396 26236 32564 26238
rect 32060 25620 32116 25630
rect 31836 25618 32116 25620
rect 31836 25566 32062 25618
rect 32114 25566 32116 25618
rect 31836 25564 32116 25566
rect 31500 25508 31556 25518
rect 29932 25394 29988 25406
rect 29932 25342 29934 25394
rect 29986 25342 29988 25394
rect 29932 24948 29988 25342
rect 29932 24882 29988 24892
rect 30940 24948 30996 24958
rect 29820 24782 29822 24834
rect 29874 24782 29876 24834
rect 28364 23886 28366 23938
rect 28418 23886 28420 23938
rect 28364 23874 28420 23886
rect 28588 23940 28644 23950
rect 25788 23828 25844 23838
rect 25788 23734 25844 23772
rect 28588 23826 28644 23884
rect 29708 23940 29764 23950
rect 29708 23846 29764 23884
rect 28588 23774 28590 23826
rect 28642 23774 28644 23826
rect 28588 23762 28644 23774
rect 29148 23828 29204 23838
rect 29148 23734 29204 23772
rect 25340 23154 25396 23166
rect 25340 23102 25342 23154
rect 25394 23102 25396 23154
rect 25004 21858 25060 21868
rect 25116 22146 25172 22158
rect 25116 22094 25118 22146
rect 25170 22094 25172 22146
rect 24556 21758 24558 21810
rect 24610 21758 24612 21810
rect 24556 21746 24612 21758
rect 23996 20638 23998 20690
rect 24050 20638 24052 20690
rect 23996 20468 24052 20638
rect 23996 20402 24052 20412
rect 24556 20802 24612 20814
rect 24892 20804 24948 20814
rect 24556 20750 24558 20802
rect 24610 20750 24612 20802
rect 24556 20356 24612 20750
rect 24556 20290 24612 20300
rect 24780 20802 24948 20804
rect 24780 20750 24894 20802
rect 24946 20750 24948 20802
rect 24780 20748 24948 20750
rect 24668 20130 24724 20142
rect 24668 20078 24670 20130
rect 24722 20078 24724 20130
rect 24108 20020 24164 20030
rect 24164 19964 24276 20020
rect 24108 19926 24164 19964
rect 24220 18564 24276 19964
rect 24332 19908 24388 19918
rect 24332 19814 24388 19852
rect 24332 18564 24388 18574
rect 24220 18562 24388 18564
rect 24220 18510 24334 18562
rect 24386 18510 24388 18562
rect 24220 18508 24388 18510
rect 24108 18452 24164 18462
rect 24108 18358 24164 18396
rect 23884 18340 23940 18350
rect 23772 18338 23940 18340
rect 23772 18286 23886 18338
rect 23938 18286 23940 18338
rect 23772 18284 23940 18286
rect 23660 18228 23716 18238
rect 23436 17490 23492 17500
rect 23548 18226 23716 18228
rect 23548 18174 23662 18226
rect 23714 18174 23716 18226
rect 23548 18172 23716 18174
rect 23548 17108 23604 18172
rect 23660 18162 23716 18172
rect 23884 18228 23940 18284
rect 23884 18162 23940 18172
rect 24220 18338 24276 18350
rect 24220 18286 24222 18338
rect 24274 18286 24276 18338
rect 23772 18116 23828 18126
rect 23660 17668 23716 17678
rect 23772 17668 23828 18060
rect 23996 17780 24052 17790
rect 24220 17780 24276 18286
rect 24332 18004 24388 18508
rect 24668 18228 24724 20078
rect 24668 18162 24724 18172
rect 24780 18116 24836 20748
rect 24892 20738 24948 20748
rect 24892 20578 24948 20590
rect 24892 20526 24894 20578
rect 24946 20526 24948 20578
rect 24892 19460 24948 20526
rect 25116 20132 25172 22094
rect 25340 20804 25396 23102
rect 26012 23044 26068 23054
rect 25676 23042 26068 23044
rect 25676 22990 26014 23042
rect 26066 22990 26068 23042
rect 25676 22988 26068 22990
rect 25452 22484 25508 22494
rect 25452 22370 25508 22428
rect 25676 22482 25732 22988
rect 26012 22978 26068 22988
rect 28140 23042 28196 23054
rect 28140 22990 28142 23042
rect 28194 22990 28196 23042
rect 25676 22430 25678 22482
rect 25730 22430 25732 22482
rect 25676 22418 25732 22430
rect 26908 22482 26964 22494
rect 26908 22430 26910 22482
rect 26962 22430 26964 22482
rect 25452 22318 25454 22370
rect 25506 22318 25508 22370
rect 25452 22306 25508 22318
rect 25788 22260 25844 22270
rect 26572 22260 26628 22270
rect 25788 22258 26628 22260
rect 25788 22206 25790 22258
rect 25842 22206 26574 22258
rect 26626 22206 26628 22258
rect 25788 22204 26628 22206
rect 25788 22194 25844 22204
rect 26572 22194 26628 22204
rect 25340 20748 25732 20804
rect 25228 20690 25284 20702
rect 25228 20638 25230 20690
rect 25282 20638 25284 20690
rect 25228 20244 25284 20638
rect 25228 20188 25396 20244
rect 25116 20066 25172 20076
rect 24892 19394 24948 19404
rect 25228 20020 25284 20030
rect 25228 18452 25284 19964
rect 25228 18386 25284 18396
rect 25340 18676 25396 20188
rect 25452 20132 25508 20142
rect 25452 19458 25508 20076
rect 25676 20020 25732 20748
rect 25676 19954 25732 19964
rect 26908 20020 26964 22430
rect 27244 22372 27300 22382
rect 28028 22372 28084 22382
rect 28140 22372 28196 22990
rect 27244 22370 27860 22372
rect 27244 22318 27246 22370
rect 27298 22318 27860 22370
rect 27244 22316 27860 22318
rect 27244 22306 27300 22316
rect 26012 19906 26068 19918
rect 26012 19854 26014 19906
rect 26066 19854 26068 19906
rect 25452 19406 25454 19458
rect 25506 19406 25508 19458
rect 25452 19348 25508 19406
rect 25676 19460 25732 19470
rect 25676 19366 25732 19404
rect 25452 19282 25508 19292
rect 25900 19236 25956 19246
rect 25900 19142 25956 19180
rect 25788 19012 25844 19022
rect 26012 19012 26068 19854
rect 26908 19236 26964 19964
rect 27804 21810 27860 22316
rect 27804 21758 27806 21810
rect 27858 21758 27860 21810
rect 26908 19122 26964 19180
rect 27132 19908 27188 19918
rect 27132 19234 27188 19852
rect 27132 19182 27134 19234
rect 27186 19182 27188 19234
rect 27132 19170 27188 19182
rect 26908 19070 26910 19122
rect 26962 19070 26964 19122
rect 26908 19058 26964 19070
rect 25788 19010 26068 19012
rect 25788 18958 25790 19010
rect 25842 18958 26068 19010
rect 25788 18956 26068 18958
rect 25788 18946 25844 18956
rect 25340 18450 25396 18620
rect 27132 18676 27188 18686
rect 27132 18582 27188 18620
rect 27356 18674 27412 18686
rect 27356 18622 27358 18674
rect 27410 18622 27412 18674
rect 25340 18398 25342 18450
rect 25394 18398 25396 18450
rect 25340 18386 25396 18398
rect 25228 18228 25284 18238
rect 25228 18134 25284 18172
rect 26124 18228 26180 18238
rect 24780 18050 24836 18060
rect 24332 17938 24388 17948
rect 25676 18004 25732 18014
rect 24220 17724 25172 17780
rect 23660 17666 23828 17668
rect 23660 17614 23662 17666
rect 23714 17614 23828 17666
rect 23660 17612 23828 17614
rect 23884 17668 23940 17678
rect 23660 17602 23716 17612
rect 23884 17574 23940 17612
rect 23996 17666 24052 17724
rect 23996 17614 23998 17666
rect 24050 17614 24052 17666
rect 23996 17602 24052 17614
rect 24220 17554 24276 17566
rect 24220 17502 24222 17554
rect 24274 17502 24276 17554
rect 23772 17442 23828 17454
rect 23772 17390 23774 17442
rect 23826 17390 23828 17442
rect 23548 17052 23716 17108
rect 23660 16994 23716 17052
rect 23660 16942 23662 16994
rect 23714 16942 23716 16994
rect 23548 16324 23604 16334
rect 22764 12738 23044 12740
rect 22764 12686 22766 12738
rect 22818 12686 23044 12738
rect 22764 12684 23044 12686
rect 23100 13020 23268 13076
rect 23324 14308 23380 14318
rect 22764 12292 22820 12684
rect 22764 12226 22820 12236
rect 22876 12404 22932 12414
rect 23100 12404 23156 13020
rect 23324 12850 23380 14252
rect 23548 13412 23604 16268
rect 23660 15428 23716 16942
rect 23660 15362 23716 15372
rect 23772 14532 23828 17390
rect 23884 17444 23940 17454
rect 23884 16882 23940 17388
rect 23884 16830 23886 16882
rect 23938 16830 23940 16882
rect 23884 16818 23940 16830
rect 23996 16884 24052 16894
rect 23996 16770 24052 16828
rect 23996 16718 23998 16770
rect 24050 16718 24052 16770
rect 23996 16706 24052 16718
rect 24220 15316 24276 17502
rect 25116 16098 25172 17724
rect 25340 17668 25396 17678
rect 25340 17574 25396 17612
rect 25564 17554 25620 17566
rect 25564 17502 25566 17554
rect 25618 17502 25620 17554
rect 25564 17444 25620 17502
rect 25340 17388 25620 17444
rect 25340 16884 25396 17388
rect 25676 17332 25732 17948
rect 25452 17276 25732 17332
rect 25900 17666 25956 17678
rect 25900 17614 25902 17666
rect 25954 17614 25956 17666
rect 25452 16994 25508 17276
rect 25452 16942 25454 16994
rect 25506 16942 25508 16994
rect 25452 16930 25508 16942
rect 25564 17108 25620 17118
rect 25900 17108 25956 17614
rect 25564 17106 25956 17108
rect 25564 17054 25566 17106
rect 25618 17054 25956 17106
rect 25564 17052 25956 17054
rect 25228 16212 25284 16222
rect 25228 16118 25284 16156
rect 25116 16046 25118 16098
rect 25170 16046 25172 16098
rect 25116 16034 25172 16046
rect 25340 16098 25396 16828
rect 25340 16046 25342 16098
rect 25394 16046 25396 16098
rect 25340 16034 25396 16046
rect 25564 15986 25620 17052
rect 25564 15934 25566 15986
rect 25618 15934 25620 15986
rect 25564 15922 25620 15934
rect 25676 16882 25732 16894
rect 25676 16830 25678 16882
rect 25730 16830 25732 16882
rect 25676 16772 25732 16830
rect 26124 16882 26180 18172
rect 26572 17890 26628 17902
rect 26572 17838 26574 17890
rect 26626 17838 26628 17890
rect 26572 17668 26628 17838
rect 27356 17780 27412 18622
rect 27804 18564 27860 21758
rect 27916 22370 28196 22372
rect 27916 22318 28030 22370
rect 28082 22318 28196 22370
rect 27916 22316 28196 22318
rect 27916 21698 27972 22316
rect 28028 22306 28084 22316
rect 27916 21646 27918 21698
rect 27970 21646 27972 21698
rect 27916 21634 27972 21646
rect 28252 22146 28308 22158
rect 28252 22094 28254 22146
rect 28306 22094 28308 22146
rect 28252 20132 28308 22094
rect 29260 20860 29652 20916
rect 29260 20690 29316 20860
rect 29260 20638 29262 20690
rect 29314 20638 29316 20690
rect 29260 20626 29316 20638
rect 29372 20690 29428 20702
rect 29372 20638 29374 20690
rect 29426 20638 29428 20690
rect 29372 20468 29428 20638
rect 28140 19906 28196 19918
rect 28140 19854 28142 19906
rect 28194 19854 28196 19906
rect 28140 18676 28196 19854
rect 28140 18610 28196 18620
rect 27804 18498 27860 18508
rect 27580 18452 27636 18462
rect 27580 18450 27748 18452
rect 27580 18398 27582 18450
rect 27634 18398 27748 18450
rect 27580 18396 27748 18398
rect 27580 18386 27636 18396
rect 26572 17602 26628 17612
rect 26796 17724 27412 17780
rect 26796 17666 26852 17724
rect 26796 17614 26798 17666
rect 26850 17614 26852 17666
rect 26796 17602 26852 17614
rect 27132 17106 27188 17724
rect 27132 17054 27134 17106
rect 27186 17054 27188 17106
rect 27132 17042 27188 17054
rect 26124 16830 26126 16882
rect 26178 16830 26180 16882
rect 26124 16818 26180 16830
rect 26572 16994 26628 17006
rect 26572 16942 26574 16994
rect 26626 16942 26628 16994
rect 25676 15540 25732 16716
rect 25676 15538 26068 15540
rect 25676 15486 25678 15538
rect 25730 15486 26068 15538
rect 25676 15484 26068 15486
rect 25676 15474 25732 15484
rect 23772 14466 23828 14476
rect 23884 15202 23940 15214
rect 23884 15150 23886 15202
rect 23938 15150 23940 15202
rect 23884 14308 23940 15150
rect 24220 15148 24276 15260
rect 25228 15428 25284 15438
rect 25228 15148 25284 15372
rect 24220 15092 24388 15148
rect 23884 14242 23940 14252
rect 24220 14308 24276 14318
rect 24220 14214 24276 14252
rect 23548 13346 23604 13356
rect 23436 13300 23492 13310
rect 23436 12962 23492 13244
rect 23436 12910 23438 12962
rect 23490 12910 23492 12962
rect 23436 12898 23492 12910
rect 23996 12964 24052 12974
rect 23324 12798 23326 12850
rect 23378 12798 23380 12850
rect 23324 12786 23380 12798
rect 22876 12178 22932 12348
rect 22876 12126 22878 12178
rect 22930 12126 22932 12178
rect 22876 12114 22932 12126
rect 22988 12348 23156 12404
rect 23436 12740 23492 12750
rect 22652 11340 22820 11396
rect 22540 11330 22596 11340
rect 22652 11172 22708 11182
rect 22652 10612 22708 11116
rect 22652 10546 22708 10556
rect 22428 9884 22596 9940
rect 20636 9774 20638 9826
rect 20690 9774 20692 9826
rect 19964 9714 20020 9726
rect 19964 9662 19966 9714
rect 20018 9662 20020 9714
rect 19964 9604 20020 9662
rect 19628 9548 20020 9604
rect 19628 9268 19684 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19740 9268 19796 9278
rect 19628 9266 19796 9268
rect 19628 9214 19742 9266
rect 19794 9214 19796 9266
rect 19628 9212 19796 9214
rect 19740 9202 19796 9212
rect 19404 8990 19406 9042
rect 19458 8990 19460 9042
rect 19404 8978 19460 8990
rect 19516 9042 19572 9054
rect 19516 8990 19518 9042
rect 19570 8990 19572 9042
rect 18732 8876 19012 8932
rect 18172 8372 18228 8382
rect 18172 8278 18228 8316
rect 18956 6690 19012 8876
rect 19516 8820 19572 8990
rect 19516 8754 19572 8764
rect 20188 8930 20244 8942
rect 20188 8878 20190 8930
rect 20242 8878 20244 8930
rect 20188 8820 20244 8878
rect 20188 8754 20244 8764
rect 19516 8036 19572 8046
rect 19516 7586 19572 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19516 7534 19518 7586
rect 19570 7534 19572 7586
rect 19516 7522 19572 7534
rect 20300 7476 20356 7486
rect 20636 7476 20692 9774
rect 21980 9828 22036 9838
rect 21980 9734 22036 9772
rect 22428 9716 22484 9726
rect 22316 9714 22484 9716
rect 22316 9662 22430 9714
rect 22482 9662 22484 9714
rect 22316 9660 22484 9662
rect 22316 8932 22372 9660
rect 22428 9650 22484 9660
rect 21868 8876 22372 8932
rect 21868 8482 21924 8876
rect 22428 8820 22484 8830
rect 22540 8820 22596 9884
rect 22484 8764 22596 8820
rect 22428 8754 22484 8764
rect 22764 8596 22820 11340
rect 22876 11284 22932 11294
rect 22876 11190 22932 11228
rect 21868 8430 21870 8482
rect 21922 8430 21924 8482
rect 21868 8418 21924 8430
rect 22316 8540 22820 8596
rect 21532 8372 21588 8382
rect 21420 8370 21588 8372
rect 21420 8318 21534 8370
rect 21586 8318 21588 8370
rect 21420 8316 21588 8318
rect 21420 7586 21476 8316
rect 21532 8306 21588 8316
rect 21644 8372 21700 8382
rect 21644 8146 21700 8316
rect 22316 8372 22372 8540
rect 22316 8278 22372 8316
rect 21644 8094 21646 8146
rect 21698 8094 21700 8146
rect 21644 8082 21700 8094
rect 21420 7534 21422 7586
rect 21474 7534 21476 7586
rect 21420 7522 21476 7534
rect 20300 7474 20636 7476
rect 20300 7422 20302 7474
rect 20354 7422 20636 7474
rect 20300 7420 20636 7422
rect 20300 7410 20356 7420
rect 20636 7382 20692 7420
rect 21532 7476 21588 7486
rect 19404 6916 19460 6926
rect 19404 6822 19460 6860
rect 18956 6638 18958 6690
rect 19010 6638 19012 6690
rect 18956 6626 19012 6638
rect 19628 6690 19684 6702
rect 19628 6638 19630 6690
rect 19682 6638 19684 6690
rect 18956 6132 19012 6142
rect 18172 6020 18228 6030
rect 18060 6018 18228 6020
rect 18060 5966 18174 6018
rect 18226 5966 18228 6018
rect 18060 5964 18228 5966
rect 18172 5954 18228 5964
rect 18508 5794 18564 5806
rect 18508 5742 18510 5794
rect 18562 5742 18564 5794
rect 18508 5348 18564 5742
rect 18956 5794 19012 6076
rect 19628 6020 19684 6638
rect 19852 6690 19908 6702
rect 19852 6638 19854 6690
rect 19906 6638 19908 6690
rect 19852 6468 19908 6638
rect 20636 6580 20692 6590
rect 20412 6468 20468 6478
rect 19852 6466 20468 6468
rect 19852 6414 20414 6466
rect 20466 6414 20468 6466
rect 19852 6412 20468 6414
rect 20412 6356 20468 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20412 6290 20468 6300
rect 19836 6234 20100 6244
rect 20188 6132 20244 6142
rect 20076 6020 20132 6030
rect 19628 5964 20076 6020
rect 18956 5742 18958 5794
rect 19010 5742 19012 5794
rect 18956 5730 19012 5742
rect 19404 5906 19460 5918
rect 19404 5854 19406 5906
rect 19458 5854 19460 5906
rect 18508 5282 18564 5292
rect 19404 5348 19460 5854
rect 20076 5906 20132 5964
rect 20076 5854 20078 5906
rect 20130 5854 20132 5906
rect 20076 5842 20132 5854
rect 19404 5282 19460 5292
rect 19180 5124 19236 5134
rect 19628 5124 19684 5134
rect 19180 5030 19236 5068
rect 19292 5122 19684 5124
rect 19292 5070 19630 5122
rect 19682 5070 19684 5122
rect 19292 5068 19684 5070
rect 18396 5010 18452 5022
rect 18396 4958 18398 5010
rect 18450 4958 18452 5010
rect 18396 4564 18452 4958
rect 18396 4498 18452 4508
rect 19180 4564 19236 4574
rect 19292 4564 19348 5068
rect 19628 5058 19684 5068
rect 20188 5122 20244 6076
rect 20300 6018 20356 6030
rect 20300 5966 20302 6018
rect 20354 5966 20356 6018
rect 20300 5908 20356 5966
rect 20300 5842 20356 5852
rect 20636 5460 20692 6524
rect 21308 6468 21364 6478
rect 21196 6466 21364 6468
rect 21196 6414 21310 6466
rect 21362 6414 21364 6466
rect 21196 6412 21364 6414
rect 20748 6132 20804 6142
rect 20748 6038 20804 6076
rect 20524 5236 20580 5246
rect 20188 5070 20190 5122
rect 20242 5070 20244 5122
rect 20188 5058 20244 5070
rect 20300 5122 20356 5134
rect 20300 5070 20302 5122
rect 20354 5070 20356 5122
rect 19180 4562 19348 4564
rect 19180 4510 19182 4562
rect 19234 4510 19348 4562
rect 19180 4508 19348 4510
rect 19516 4898 19572 4910
rect 19516 4846 19518 4898
rect 19570 4846 19572 4898
rect 19180 4498 19236 4508
rect 19516 4450 19572 4846
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4564 19684 4574
rect 20300 4564 20356 5070
rect 20412 5012 20468 5022
rect 20412 4918 20468 4956
rect 19628 4470 19684 4508
rect 20076 4508 20356 4564
rect 19516 4398 19518 4450
rect 19570 4398 19572 4450
rect 19516 4386 19572 4398
rect 19852 4452 19908 4462
rect 19852 4358 19908 4396
rect 20076 4450 20132 4508
rect 20076 4398 20078 4450
rect 20130 4398 20132 4450
rect 20076 4386 20132 4398
rect 18844 4338 18900 4350
rect 18844 4286 18846 4338
rect 18898 4286 18900 4338
rect 18172 4226 18228 4238
rect 18172 4174 18174 4226
rect 18226 4174 18228 4226
rect 18172 4004 18228 4174
rect 18172 3938 18228 3948
rect 18620 4226 18676 4238
rect 18620 4174 18622 4226
rect 18674 4174 18676 4226
rect 16940 3502 16942 3554
rect 16994 3502 16996 3554
rect 16940 3490 16996 3502
rect 18620 3556 18676 4174
rect 18844 4004 18900 4286
rect 20524 4338 20580 5180
rect 20636 5010 20692 5404
rect 20860 5908 20916 5918
rect 20636 4958 20638 5010
rect 20690 4958 20692 5010
rect 20636 4946 20692 4958
rect 20748 5348 20804 5358
rect 20636 4452 20692 4462
rect 20636 4358 20692 4396
rect 20524 4286 20526 4338
rect 20578 4286 20580 4338
rect 20524 4274 20580 4286
rect 18844 3938 18900 3948
rect 19516 4004 19572 4014
rect 18620 3490 18676 3500
rect 18844 3668 18900 3678
rect 14812 3442 14868 3454
rect 14812 3390 14814 3442
rect 14866 3390 14868 3442
rect 14812 800 14868 3390
rect 15484 3444 15540 3454
rect 15484 800 15540 3388
rect 18508 3444 18564 3482
rect 18508 3378 18564 3388
rect 18844 800 18900 3612
rect 19516 800 19572 3948
rect 19852 3556 19908 3566
rect 19852 3462 19908 3500
rect 20748 3554 20804 5292
rect 20860 4452 20916 5852
rect 20972 5012 21028 5022
rect 21196 5012 21252 6412
rect 21308 6402 21364 6412
rect 21532 5124 21588 7420
rect 22876 7476 22932 7486
rect 22876 6690 22932 7420
rect 22876 6638 22878 6690
rect 22930 6638 22932 6690
rect 22876 6626 22932 6638
rect 22988 6692 23044 12348
rect 23436 12290 23492 12684
rect 23996 12402 24052 12908
rect 24108 12962 24164 12974
rect 24108 12910 24110 12962
rect 24162 12910 24164 12962
rect 24108 12740 24164 12910
rect 24332 12852 24388 15092
rect 25004 15092 25284 15148
rect 25452 15314 25508 15326
rect 25452 15262 25454 15314
rect 25506 15262 25508 15314
rect 24780 14868 24836 14878
rect 24780 14642 24836 14812
rect 24780 14590 24782 14642
rect 24834 14590 24836 14642
rect 24780 14578 24836 14590
rect 24556 13634 24612 13646
rect 24556 13582 24558 13634
rect 24610 13582 24612 13634
rect 24556 13412 24612 13582
rect 24612 13356 24948 13412
rect 24556 13346 24612 13356
rect 24332 12850 24612 12852
rect 24332 12798 24334 12850
rect 24386 12798 24612 12850
rect 24332 12796 24612 12798
rect 24332 12786 24388 12796
rect 24108 12674 24164 12684
rect 24220 12738 24276 12750
rect 24220 12686 24222 12738
rect 24274 12686 24276 12738
rect 24220 12628 24276 12686
rect 24220 12562 24276 12572
rect 23996 12350 23998 12402
rect 24050 12350 24052 12402
rect 23996 12338 24052 12350
rect 24556 12404 24612 12796
rect 24892 12850 24948 13356
rect 24892 12798 24894 12850
rect 24946 12798 24948 12850
rect 24892 12786 24948 12798
rect 24556 12310 24612 12348
rect 23436 12238 23438 12290
rect 23490 12238 23492 12290
rect 23436 12226 23492 12238
rect 23884 12292 23940 12302
rect 23884 12198 23940 12236
rect 24668 12292 24724 12302
rect 23212 12068 23268 12078
rect 23212 11394 23268 12012
rect 23212 11342 23214 11394
rect 23266 11342 23268 11394
rect 23212 11330 23268 11342
rect 23324 11954 23380 11966
rect 23324 11902 23326 11954
rect 23378 11902 23380 11954
rect 23324 11284 23380 11902
rect 23324 11218 23380 11228
rect 23436 11396 23492 11406
rect 23436 10722 23492 11340
rect 24332 11284 24388 11294
rect 23436 10670 23438 10722
rect 23490 10670 23492 10722
rect 23436 10658 23492 10670
rect 23548 10724 23604 10734
rect 23548 10722 23716 10724
rect 23548 10670 23550 10722
rect 23602 10670 23716 10722
rect 23548 10668 23716 10670
rect 23548 10658 23604 10668
rect 23212 10612 23268 10622
rect 23212 9826 23268 10556
rect 23212 9774 23214 9826
rect 23266 9774 23268 9826
rect 23212 9762 23268 9774
rect 23660 9716 23716 10668
rect 23772 10612 23828 10622
rect 23772 10610 23940 10612
rect 23772 10558 23774 10610
rect 23826 10558 23940 10610
rect 23772 10556 23940 10558
rect 23772 10546 23828 10556
rect 23548 8930 23604 8942
rect 23548 8878 23550 8930
rect 23602 8878 23604 8930
rect 23548 8820 23604 8878
rect 23548 8754 23604 8764
rect 23548 7364 23604 7374
rect 23660 7364 23716 9660
rect 23884 9154 23940 10556
rect 24332 9714 24388 11228
rect 24332 9662 24334 9714
rect 24386 9662 24388 9714
rect 24332 9650 24388 9662
rect 24444 9604 24500 9614
rect 24444 9380 24500 9548
rect 24668 9492 24724 12236
rect 24332 9324 24500 9380
rect 24556 9436 24724 9492
rect 23884 9102 23886 9154
rect 23938 9102 23940 9154
rect 23884 9090 23940 9102
rect 24108 9156 24164 9166
rect 24108 9062 24164 9100
rect 24332 9042 24388 9324
rect 24332 8990 24334 9042
rect 24386 8990 24388 9042
rect 24332 8978 24388 8990
rect 24220 8258 24276 8270
rect 24220 8206 24222 8258
rect 24274 8206 24276 8258
rect 24220 7476 24276 8206
rect 24220 7410 24276 7420
rect 23548 7362 23716 7364
rect 23548 7310 23550 7362
rect 23602 7310 23716 7362
rect 23548 7308 23716 7310
rect 24108 7362 24164 7374
rect 24108 7310 24110 7362
rect 24162 7310 24164 7362
rect 23548 7298 23604 7308
rect 24108 7252 24164 7310
rect 24220 7252 24276 7262
rect 24108 7196 24220 7252
rect 24220 7186 24276 7196
rect 21644 6466 21700 6478
rect 21644 6414 21646 6466
rect 21698 6414 21700 6466
rect 21644 6020 21700 6414
rect 22988 6132 23044 6636
rect 24332 6804 24388 6814
rect 23660 6580 23716 6590
rect 23660 6578 23940 6580
rect 23660 6526 23662 6578
rect 23714 6526 23940 6578
rect 23660 6524 23940 6526
rect 23660 6514 23716 6524
rect 22988 6066 23044 6076
rect 23884 6130 23940 6524
rect 23884 6078 23886 6130
rect 23938 6078 23940 6130
rect 23884 6066 23940 6078
rect 21644 5954 21700 5964
rect 24332 6018 24388 6748
rect 24332 5966 24334 6018
rect 24386 5966 24388 6018
rect 24332 5954 24388 5966
rect 23436 5908 23492 5918
rect 23660 5908 23716 5918
rect 23436 5906 23716 5908
rect 23436 5854 23438 5906
rect 23490 5854 23662 5906
rect 23714 5854 23716 5906
rect 23436 5852 23716 5854
rect 23436 5842 23492 5852
rect 23660 5842 23716 5852
rect 24108 5908 24164 5918
rect 24108 5814 24164 5852
rect 23324 5794 23380 5806
rect 23324 5742 23326 5794
rect 23378 5742 23380 5794
rect 21028 4956 21252 5012
rect 21420 5010 21476 5022
rect 21420 4958 21422 5010
rect 21474 4958 21476 5010
rect 20972 4946 21028 4956
rect 21308 4900 21364 4910
rect 20860 4386 20916 4396
rect 21084 4898 21364 4900
rect 21084 4846 21310 4898
rect 21362 4846 21364 4898
rect 21084 4844 21364 4846
rect 21084 4338 21140 4844
rect 21308 4834 21364 4844
rect 21420 4564 21476 4958
rect 21084 4286 21086 4338
rect 21138 4286 21140 4338
rect 21084 4274 21140 4286
rect 21196 4508 21476 4564
rect 20860 4228 20916 4238
rect 20860 4134 20916 4172
rect 20748 3502 20750 3554
rect 20802 3502 20804 3554
rect 20748 3490 20804 3502
rect 20188 3442 20244 3454
rect 20188 3390 20190 3442
rect 20242 3390 20244 3442
rect 20188 3388 20244 3390
rect 21196 3388 21252 4508
rect 21420 4340 21476 4350
rect 21532 4340 21588 5068
rect 21756 5460 21812 5470
rect 21756 5122 21812 5404
rect 22316 5236 22372 5246
rect 22316 5142 22372 5180
rect 21756 5070 21758 5122
rect 21810 5070 21812 5122
rect 21756 5058 21812 5070
rect 23324 5124 23380 5742
rect 24556 5460 24612 9436
rect 24668 9268 24724 9278
rect 24668 9266 24948 9268
rect 24668 9214 24670 9266
rect 24722 9214 24948 9266
rect 24668 9212 24948 9214
rect 24668 9202 24724 9212
rect 24668 9042 24724 9054
rect 24668 8990 24670 9042
rect 24722 8990 24724 9042
rect 24668 8820 24724 8990
rect 24668 8754 24724 8764
rect 24892 8370 24948 9212
rect 24892 8318 24894 8370
rect 24946 8318 24948 8370
rect 24892 8306 24948 8318
rect 24668 7476 24724 7486
rect 24668 7382 24724 7420
rect 25004 5908 25060 15092
rect 25116 14418 25172 14430
rect 25116 14366 25118 14418
rect 25170 14366 25172 14418
rect 25116 14308 25172 14366
rect 25116 14242 25172 14252
rect 25228 14308 25284 14318
rect 25452 14308 25508 15262
rect 25788 15314 25844 15326
rect 25788 15262 25790 15314
rect 25842 15262 25844 15314
rect 25564 15202 25620 15214
rect 25564 15150 25566 15202
rect 25618 15150 25620 15202
rect 25564 15092 25620 15150
rect 25788 15204 25844 15262
rect 25788 15138 25844 15148
rect 25564 15026 25620 15036
rect 25900 14756 25956 14766
rect 25900 14662 25956 14700
rect 25228 14306 25508 14308
rect 25228 14254 25230 14306
rect 25282 14254 25508 14306
rect 25228 14252 25508 14254
rect 25564 14420 25620 14430
rect 25228 12962 25284 14252
rect 25228 12910 25230 12962
rect 25282 12910 25284 12962
rect 25228 12898 25284 12910
rect 25564 12964 25620 14364
rect 25788 14306 25844 14318
rect 25788 14254 25790 14306
rect 25842 14254 25844 14306
rect 25564 12898 25620 12908
rect 25676 12962 25732 12974
rect 25676 12910 25678 12962
rect 25730 12910 25732 12962
rect 25228 12740 25284 12750
rect 25228 12290 25284 12684
rect 25452 12404 25508 12414
rect 25452 12310 25508 12348
rect 25228 12238 25230 12290
rect 25282 12238 25284 12290
rect 25228 12226 25284 12238
rect 25676 12292 25732 12910
rect 25676 12226 25732 12236
rect 25564 12068 25620 12078
rect 25564 11974 25620 12012
rect 25788 11508 25844 14254
rect 26012 12180 26068 15484
rect 26124 15314 26180 15326
rect 26124 15262 26126 15314
rect 26178 15262 26180 15314
rect 26124 14868 26180 15262
rect 26460 15316 26516 15326
rect 26460 15222 26516 15260
rect 26348 15202 26404 15214
rect 26348 15150 26350 15202
rect 26402 15150 26404 15202
rect 26348 14980 26404 15150
rect 26348 14914 26404 14924
rect 26124 14802 26180 14812
rect 26236 14532 26292 14542
rect 26236 13636 26292 14476
rect 26348 14420 26404 14430
rect 26572 14420 26628 16942
rect 27692 16996 27748 18396
rect 28252 18450 28308 20076
rect 29260 20412 29428 20468
rect 29484 20690 29540 20702
rect 29484 20638 29486 20690
rect 29538 20638 29540 20690
rect 29260 20132 29316 20412
rect 29484 20188 29540 20638
rect 29036 20018 29092 20030
rect 29036 19966 29038 20018
rect 29090 19966 29092 20018
rect 29036 19908 29092 19966
rect 29036 19842 29092 19852
rect 28812 19796 28868 19806
rect 29260 19796 29316 20076
rect 29372 20132 29540 20188
rect 29372 20020 29428 20132
rect 29372 19954 29428 19964
rect 29484 20018 29540 20030
rect 29484 19966 29486 20018
rect 29538 19966 29540 20018
rect 29484 19796 29540 19966
rect 29260 19740 29540 19796
rect 28812 19702 28868 19740
rect 29484 19460 29540 19740
rect 29596 20018 29652 20860
rect 29820 20188 29876 24782
rect 30940 24834 30996 24892
rect 30940 24782 30942 24834
rect 30994 24782 30996 24834
rect 30940 24770 30996 24782
rect 31052 24836 31108 24846
rect 31052 24722 31108 24780
rect 31388 24724 31444 24734
rect 31500 24724 31556 25452
rect 31836 24724 31892 25564
rect 32060 25554 32116 25564
rect 32396 25618 32452 26236
rect 32508 26226 32564 26236
rect 32620 26292 32676 26302
rect 32396 25566 32398 25618
rect 32450 25566 32452 25618
rect 32396 25554 32452 25566
rect 32508 26066 32564 26078
rect 32508 26014 32510 26066
rect 32562 26014 32564 26066
rect 32508 24948 32564 26014
rect 32620 25732 32676 26236
rect 32620 25638 32676 25676
rect 32956 25732 33012 26852
rect 33068 26516 33124 26526
rect 33180 26516 33236 27580
rect 33068 26514 33236 26516
rect 33068 26462 33070 26514
rect 33122 26462 33236 26514
rect 33068 26460 33236 26462
rect 33068 26450 33124 26460
rect 33404 26068 33460 27804
rect 35980 27746 36036 27758
rect 35980 27694 35982 27746
rect 36034 27694 36036 27746
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 33852 27076 33908 27086
rect 33628 26404 33684 26414
rect 33628 26310 33684 26348
rect 33516 26292 33572 26302
rect 33516 26198 33572 26236
rect 33852 26290 33908 27020
rect 35868 27076 35924 27086
rect 35868 26982 35924 27020
rect 35980 26852 36036 27694
rect 35980 26786 36036 26796
rect 35420 26516 35476 26526
rect 35420 26422 35476 26460
rect 33852 26238 33854 26290
rect 33906 26238 33908 26290
rect 33852 26226 33908 26238
rect 35868 26402 35924 26414
rect 35868 26350 35870 26402
rect 35922 26350 35924 26402
rect 33404 26012 33684 26068
rect 32956 25730 33348 25732
rect 32956 25678 32958 25730
rect 33010 25678 33348 25730
rect 32956 25676 33348 25678
rect 32956 25666 33012 25676
rect 32508 24892 33236 24948
rect 31052 24670 31054 24722
rect 31106 24670 31108 24722
rect 31052 24658 31108 24670
rect 31164 24722 31556 24724
rect 31164 24670 31390 24722
rect 31442 24670 31556 24722
rect 31164 24668 31556 24670
rect 31724 24722 31892 24724
rect 31724 24670 31838 24722
rect 31890 24670 31892 24722
rect 31724 24668 31892 24670
rect 31164 24276 31220 24668
rect 31388 24658 31444 24668
rect 31724 24612 31780 24668
rect 31836 24658 31892 24668
rect 31500 24556 31780 24612
rect 31276 24500 31332 24510
rect 31276 24406 31332 24444
rect 30716 24220 31220 24276
rect 29932 24050 29988 24062
rect 29932 23998 29934 24050
rect 29986 23998 29988 24050
rect 29932 23380 29988 23998
rect 29932 23378 30212 23380
rect 29932 23326 29934 23378
rect 29986 23326 30212 23378
rect 29932 23324 30212 23326
rect 29932 23314 29988 23324
rect 30156 22370 30212 23324
rect 30716 23378 30772 24220
rect 30716 23326 30718 23378
rect 30770 23326 30772 23378
rect 30716 23314 30772 23326
rect 30156 22318 30158 22370
rect 30210 22318 30212 22370
rect 30156 22306 30212 22318
rect 30268 23156 30324 23166
rect 30268 22930 30324 23100
rect 31164 23156 31220 23166
rect 31388 23156 31444 23166
rect 31164 23154 31332 23156
rect 31164 23102 31166 23154
rect 31218 23102 31332 23154
rect 31164 23100 31332 23102
rect 31164 23090 31220 23100
rect 30492 23044 30548 23054
rect 30492 23042 30660 23044
rect 30492 22990 30494 23042
rect 30546 22990 30660 23042
rect 30492 22988 30660 22990
rect 30492 22978 30548 22988
rect 30268 22878 30270 22930
rect 30322 22878 30324 22930
rect 29932 20804 29988 20814
rect 29932 20710 29988 20748
rect 29820 20132 29988 20188
rect 29596 19966 29598 20018
rect 29650 19966 29652 20018
rect 29596 19684 29652 19966
rect 29596 19618 29652 19628
rect 29708 20018 29764 20030
rect 29708 19966 29710 20018
rect 29762 19966 29764 20018
rect 29708 19572 29764 19966
rect 29932 19684 29988 20132
rect 30044 20020 30100 20030
rect 30044 19926 30100 19964
rect 30268 19796 30324 22878
rect 30492 22484 30548 22494
rect 30492 22258 30548 22428
rect 30492 22206 30494 22258
rect 30546 22206 30548 22258
rect 30492 22194 30548 22206
rect 30604 21700 30660 22988
rect 31276 22820 31332 23100
rect 31388 23062 31444 23100
rect 31500 23044 31556 24556
rect 31836 24500 31892 24510
rect 32172 24500 32228 24510
rect 31836 24406 31892 24444
rect 31948 24498 32228 24500
rect 31948 24446 32174 24498
rect 32226 24446 32228 24498
rect 31948 24444 32228 24446
rect 33180 24500 33236 24892
rect 33292 24722 33348 25676
rect 33628 25506 33684 26012
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 33628 25454 33630 25506
rect 33682 25454 33684 25506
rect 33628 25442 33684 25454
rect 34300 25396 34356 25406
rect 33852 25394 34356 25396
rect 33852 25342 34302 25394
rect 34354 25342 34356 25394
rect 33852 25340 34356 25342
rect 33292 24670 33294 24722
rect 33346 24670 33348 24722
rect 33292 24658 33348 24670
rect 33740 24836 33796 24846
rect 33740 24722 33796 24780
rect 33852 24834 33908 25340
rect 34300 25330 34356 25340
rect 33852 24782 33854 24834
rect 33906 24782 33908 24834
rect 33852 24770 33908 24782
rect 34636 24836 34692 24846
rect 33740 24670 33742 24722
rect 33794 24670 33796 24722
rect 33740 24658 33796 24670
rect 33516 24500 33572 24510
rect 33180 24498 33572 24500
rect 33180 24446 33518 24498
rect 33570 24446 33572 24498
rect 33180 24444 33572 24446
rect 31612 23268 31668 23278
rect 31612 23266 31892 23268
rect 31612 23214 31614 23266
rect 31666 23214 31892 23266
rect 31612 23212 31892 23214
rect 31612 23202 31668 23212
rect 31724 23044 31780 23054
rect 31500 23042 31780 23044
rect 31500 22990 31726 23042
rect 31778 22990 31780 23042
rect 31500 22988 31780 22990
rect 31612 22820 31668 22830
rect 31276 22764 31612 22820
rect 31612 22594 31668 22764
rect 31612 22542 31614 22594
rect 31666 22542 31668 22594
rect 31612 22530 31668 22542
rect 30604 21634 30660 21644
rect 31388 22484 31444 22494
rect 31388 21586 31444 22428
rect 31724 22372 31780 22988
rect 31388 21534 31390 21586
rect 31442 21534 31444 21586
rect 31388 21522 31444 21534
rect 31612 22316 31780 22372
rect 31164 21476 31220 21486
rect 31164 21382 31220 21420
rect 30828 21364 30884 21374
rect 30604 21362 30884 21364
rect 30604 21310 30830 21362
rect 30882 21310 30884 21362
rect 30604 21308 30884 21310
rect 30380 20804 30436 20814
rect 30380 20710 30436 20748
rect 30492 20802 30548 20814
rect 30492 20750 30494 20802
rect 30546 20750 30548 20802
rect 30380 20244 30436 20254
rect 30492 20244 30548 20750
rect 30380 20242 30548 20244
rect 30380 20190 30382 20242
rect 30434 20190 30548 20242
rect 30380 20188 30548 20190
rect 30380 20178 30436 20188
rect 30268 19730 30324 19740
rect 30380 20018 30436 20030
rect 30380 19966 30382 20018
rect 30434 19966 30436 20018
rect 29708 19506 29764 19516
rect 29820 19628 29988 19684
rect 29484 19394 29540 19404
rect 28252 18398 28254 18450
rect 28306 18398 28308 18450
rect 28252 18386 28308 18398
rect 28364 18562 28420 18574
rect 28364 18510 28366 18562
rect 28418 18510 28420 18562
rect 27916 18004 27972 18014
rect 27692 16940 27860 16996
rect 27020 16882 27076 16894
rect 27020 16830 27022 16882
rect 27074 16830 27076 16882
rect 27020 16212 27076 16830
rect 27356 16884 27412 16894
rect 27356 16882 27636 16884
rect 27356 16830 27358 16882
rect 27410 16830 27636 16882
rect 27356 16828 27636 16830
rect 27356 16818 27412 16828
rect 27020 16146 27076 16156
rect 27580 16098 27636 16828
rect 27692 16770 27748 16782
rect 27692 16718 27694 16770
rect 27746 16718 27748 16770
rect 27692 16660 27748 16718
rect 27692 16594 27748 16604
rect 27580 16046 27582 16098
rect 27634 16046 27636 16098
rect 27580 16034 27636 16046
rect 27692 15876 27748 15886
rect 27692 15782 27748 15820
rect 27356 15426 27412 15438
rect 27356 15374 27358 15426
rect 27410 15374 27412 15426
rect 26684 15314 26740 15326
rect 27356 15316 27412 15374
rect 26684 15262 26686 15314
rect 26738 15262 26740 15314
rect 26684 14756 26740 15262
rect 27132 15260 27412 15316
rect 27468 15314 27524 15326
rect 27468 15262 27470 15314
rect 27522 15262 27524 15314
rect 27020 15092 27076 15102
rect 26796 14756 26852 14766
rect 26684 14700 26796 14756
rect 26796 14642 26852 14700
rect 26796 14590 26798 14642
rect 26850 14590 26852 14642
rect 26796 14578 26852 14590
rect 27020 14754 27076 15036
rect 27020 14702 27022 14754
rect 27074 14702 27076 14754
rect 26348 14418 26516 14420
rect 26348 14366 26350 14418
rect 26402 14366 26516 14418
rect 26348 14364 26516 14366
rect 26572 14364 26852 14420
rect 26348 14354 26404 14364
rect 26236 13570 26292 13580
rect 26348 13076 26404 13086
rect 26236 12964 26292 12974
rect 26236 12870 26292 12908
rect 26236 12404 26292 12414
rect 26348 12404 26404 13020
rect 26460 12852 26516 14364
rect 26572 13524 26628 13534
rect 26572 13074 26628 13468
rect 26572 13022 26574 13074
rect 26626 13022 26628 13074
rect 26572 13010 26628 13022
rect 26684 12852 26740 12862
rect 26460 12796 26628 12852
rect 26236 12402 26404 12404
rect 26236 12350 26238 12402
rect 26290 12350 26404 12402
rect 26236 12348 26404 12350
rect 26460 12404 26516 12414
rect 26236 12338 26292 12348
rect 26012 12124 26292 12180
rect 25676 11452 25844 11508
rect 26124 11954 26180 11966
rect 26124 11902 26126 11954
rect 26178 11902 26180 11954
rect 25228 11394 25284 11406
rect 25228 11342 25230 11394
rect 25282 11342 25284 11394
rect 25228 10612 25284 11342
rect 25228 9828 25284 10556
rect 25228 9734 25284 9772
rect 25676 7474 25732 11452
rect 25788 11284 25844 11294
rect 26124 11284 26180 11902
rect 25788 11282 26180 11284
rect 25788 11230 25790 11282
rect 25842 11230 26180 11282
rect 25788 11228 26180 11230
rect 25788 9940 25844 11228
rect 25788 9714 25844 9884
rect 25788 9662 25790 9714
rect 25842 9662 25844 9714
rect 25788 9156 25844 9662
rect 25788 9090 25844 9100
rect 26124 10164 26180 10174
rect 25676 7422 25678 7474
rect 25730 7422 25732 7474
rect 25676 6804 25732 7422
rect 26124 7476 26180 10108
rect 26124 7382 26180 7420
rect 26124 7252 26180 7262
rect 26236 7252 26292 12124
rect 26460 12178 26516 12348
rect 26460 12126 26462 12178
rect 26514 12126 26516 12178
rect 26460 12114 26516 12126
rect 26460 10612 26516 10622
rect 26460 9154 26516 10556
rect 26572 10612 26628 12796
rect 26684 12404 26740 12796
rect 26684 12338 26740 12348
rect 26796 11396 26852 14364
rect 27020 13860 27076 14702
rect 27020 13794 27076 13804
rect 27132 14532 27188 15260
rect 27468 15148 27524 15262
rect 27132 13634 27188 14476
rect 27356 15090 27412 15102
rect 27468 15092 27748 15148
rect 27356 15038 27358 15090
rect 27410 15038 27412 15090
rect 27356 14530 27412 15038
rect 27692 14868 27748 15092
rect 27692 14802 27748 14812
rect 27356 14478 27358 14530
rect 27410 14478 27412 14530
rect 27356 14466 27412 14478
rect 27692 14532 27748 14542
rect 27692 14438 27748 14476
rect 27468 14306 27524 14318
rect 27468 14254 27470 14306
rect 27522 14254 27524 14306
rect 27468 14196 27524 14254
rect 27580 14308 27636 14318
rect 27580 14214 27636 14252
rect 27132 13582 27134 13634
rect 27186 13582 27188 13634
rect 26796 11330 26852 11340
rect 27020 12850 27076 12862
rect 27020 12798 27022 12850
rect 27074 12798 27076 12850
rect 26796 11170 26852 11182
rect 26796 11118 26798 11170
rect 26850 11118 26852 11170
rect 26796 10836 26852 11118
rect 26796 10770 26852 10780
rect 26684 10612 26740 10622
rect 26572 10610 26740 10612
rect 26572 10558 26686 10610
rect 26738 10558 26740 10610
rect 26572 10556 26740 10558
rect 26572 10164 26628 10556
rect 26684 10546 26740 10556
rect 26908 10612 26964 10622
rect 26908 10518 26964 10556
rect 26572 10098 26628 10108
rect 26908 10388 26964 10398
rect 26796 9604 26852 9614
rect 26796 9510 26852 9548
rect 26460 9102 26462 9154
rect 26514 9102 26516 9154
rect 26460 9090 26516 9102
rect 26908 7588 26964 10332
rect 27020 9828 27076 12798
rect 27020 9762 27076 9772
rect 27132 9492 27188 13582
rect 27244 14140 27524 14196
rect 27244 13076 27300 14140
rect 27468 13860 27524 13870
rect 27468 13766 27524 13804
rect 27356 13748 27412 13758
rect 27356 13654 27412 13692
rect 27244 13010 27300 13020
rect 27468 13636 27524 13646
rect 27244 12740 27300 12750
rect 27300 12684 27412 12740
rect 27244 12646 27300 12684
rect 27244 12180 27300 12190
rect 27244 9716 27300 12124
rect 27356 10388 27412 12684
rect 27468 12178 27524 13580
rect 27804 12964 27860 16940
rect 27916 16098 27972 17948
rect 28028 17556 28084 17566
rect 28028 16994 28084 17500
rect 28028 16942 28030 16994
rect 28082 16942 28084 16994
rect 28028 16930 28084 16942
rect 28252 16882 28308 16894
rect 28252 16830 28254 16882
rect 28306 16830 28308 16882
rect 28140 16772 28196 16782
rect 28140 16678 28196 16716
rect 27916 16046 27918 16098
rect 27970 16046 27972 16098
rect 27916 16034 27972 16046
rect 28252 16660 28308 16830
rect 28252 15148 28308 16604
rect 28028 15092 28308 15148
rect 27916 14980 27972 14990
rect 27916 13746 27972 14924
rect 27916 13694 27918 13746
rect 27970 13694 27972 13746
rect 27916 13682 27972 13694
rect 28028 13300 28084 15092
rect 28252 14868 28308 14878
rect 28140 14084 28196 14094
rect 28140 13970 28196 14028
rect 28140 13918 28142 13970
rect 28194 13918 28196 13970
rect 28140 13906 28196 13918
rect 28028 13234 28084 13244
rect 28252 13748 28308 14812
rect 28252 13074 28308 13692
rect 28252 13022 28254 13074
rect 28306 13022 28308 13074
rect 28252 13010 28308 13022
rect 27916 12964 27972 12974
rect 27804 12962 27972 12964
rect 27804 12910 27918 12962
rect 27970 12910 27972 12962
rect 27804 12908 27972 12910
rect 27468 12126 27470 12178
rect 27522 12126 27524 12178
rect 27468 12114 27524 12126
rect 27916 12178 27972 12908
rect 28364 12964 28420 18510
rect 29260 18564 29316 18574
rect 28812 17780 28868 17790
rect 28700 17220 28756 17230
rect 28588 16660 28644 16670
rect 28700 16660 28756 17164
rect 28812 16882 28868 17724
rect 28812 16830 28814 16882
rect 28866 16830 28868 16882
rect 28812 16818 28868 16830
rect 28588 16658 28756 16660
rect 28588 16606 28590 16658
rect 28642 16606 28756 16658
rect 28588 16604 28756 16606
rect 28588 16594 28644 16604
rect 28476 15986 28532 15998
rect 28476 15934 28478 15986
rect 28530 15934 28532 15986
rect 28476 15316 28532 15934
rect 28588 15988 28644 15998
rect 28588 15894 28644 15932
rect 28924 15316 28980 15326
rect 28476 15260 28924 15316
rect 28924 15202 28980 15260
rect 28924 15150 28926 15202
rect 28978 15150 28980 15202
rect 28924 15138 28980 15150
rect 29260 15148 29316 18508
rect 29708 18452 29764 18462
rect 29708 18358 29764 18396
rect 29596 18340 29652 18350
rect 29372 17668 29428 17678
rect 29372 17574 29428 17612
rect 29596 17666 29652 18284
rect 29596 17614 29598 17666
rect 29650 17614 29652 17666
rect 29596 17602 29652 17614
rect 29596 16996 29652 17006
rect 29820 16996 29876 19628
rect 30380 19460 30436 19966
rect 30380 19394 30436 19404
rect 30492 20020 30548 20030
rect 30492 19348 30548 19964
rect 30492 19282 30548 19292
rect 30156 19236 30212 19246
rect 30380 19236 30436 19246
rect 30044 19234 30212 19236
rect 30044 19182 30158 19234
rect 30210 19182 30212 19234
rect 30044 19180 30212 19182
rect 29932 19122 29988 19134
rect 29932 19070 29934 19122
rect 29986 19070 29988 19122
rect 29932 18004 29988 19070
rect 29932 17938 29988 17948
rect 29652 16940 29876 16996
rect 29932 17778 29988 17790
rect 29932 17726 29934 17778
rect 29986 17726 29988 17778
rect 29596 16210 29652 16940
rect 29596 16158 29598 16210
rect 29650 16158 29652 16210
rect 29596 16146 29652 16158
rect 29708 16772 29764 16782
rect 29708 16098 29764 16716
rect 29708 16046 29710 16098
rect 29762 16046 29764 16098
rect 29708 16034 29764 16046
rect 29820 16436 29876 16446
rect 29484 15988 29540 15998
rect 29540 15932 29652 15988
rect 29484 15922 29540 15932
rect 29484 15652 29540 15662
rect 29260 15092 29428 15148
rect 29372 14530 29428 15092
rect 29484 14642 29540 15596
rect 29484 14590 29486 14642
rect 29538 14590 29540 14642
rect 29484 14578 29540 14590
rect 29372 14478 29374 14530
rect 29426 14478 29428 14530
rect 29372 14466 29428 14478
rect 29596 14532 29652 15932
rect 29820 15148 29876 16380
rect 29932 16322 29988 17726
rect 30044 16884 30100 19180
rect 30156 19170 30212 19180
rect 30268 19234 30436 19236
rect 30268 19182 30382 19234
rect 30434 19182 30436 19234
rect 30268 19180 30436 19182
rect 30156 19010 30212 19022
rect 30156 18958 30158 19010
rect 30210 18958 30212 19010
rect 30156 17668 30212 18958
rect 30268 18004 30324 19180
rect 30380 19170 30436 19180
rect 30604 18564 30660 21308
rect 30828 21298 30884 21308
rect 30940 21362 30996 21374
rect 30940 21310 30942 21362
rect 30994 21310 30996 21362
rect 30940 20916 30996 21310
rect 30716 20860 30996 20916
rect 30716 20802 30772 20860
rect 30716 20750 30718 20802
rect 30770 20750 30772 20802
rect 30716 20244 30772 20750
rect 31164 20804 31220 20814
rect 31164 20710 31220 20748
rect 30716 20178 30772 20188
rect 30828 20690 30884 20702
rect 30828 20638 30830 20690
rect 30882 20638 30884 20690
rect 30380 18508 30660 18564
rect 30716 20018 30772 20030
rect 30716 19966 30718 20018
rect 30770 19966 30772 20018
rect 30716 19684 30772 19966
rect 30716 18564 30772 19628
rect 30380 18450 30436 18508
rect 30716 18498 30772 18508
rect 30380 18398 30382 18450
rect 30434 18398 30436 18450
rect 30380 18386 30436 18398
rect 30268 17780 30324 17948
rect 30268 17714 30324 17724
rect 30156 17602 30212 17612
rect 30492 17666 30548 17678
rect 30492 17614 30494 17666
rect 30546 17614 30548 17666
rect 30492 17220 30548 17614
rect 30716 17668 30772 17678
rect 30716 17574 30772 17612
rect 30828 17332 30884 20638
rect 31612 20692 31668 22316
rect 31836 21700 31892 23212
rect 31948 22594 32004 24444
rect 32172 24434 32228 24444
rect 33516 24434 33572 24444
rect 33516 23940 33572 23978
rect 33740 23940 33796 23950
rect 33404 23884 33516 23940
rect 33292 23826 33348 23838
rect 33292 23774 33294 23826
rect 33346 23774 33348 23826
rect 33068 22932 33124 22942
rect 33068 22838 33124 22876
rect 31948 22542 31950 22594
rect 32002 22542 32004 22594
rect 31948 21812 32004 22542
rect 33292 22484 33348 23774
rect 33404 23268 33460 23884
rect 33516 23874 33572 23884
rect 33628 23938 33796 23940
rect 33628 23886 33742 23938
rect 33794 23886 33796 23938
rect 33628 23884 33796 23886
rect 33516 23714 33572 23726
rect 33516 23662 33518 23714
rect 33570 23662 33572 23714
rect 33516 23492 33572 23662
rect 33516 23426 33572 23436
rect 33516 23268 33572 23278
rect 33404 23266 33572 23268
rect 33404 23214 33518 23266
rect 33570 23214 33572 23266
rect 33404 23212 33572 23214
rect 33404 22484 33460 22494
rect 33292 22428 33404 22484
rect 33404 22370 33460 22428
rect 33404 22318 33406 22370
rect 33458 22318 33460 22370
rect 33404 22306 33460 22318
rect 33180 22260 33236 22270
rect 33180 22166 33236 22204
rect 33292 22258 33348 22270
rect 33292 22206 33294 22258
rect 33346 22206 33348 22258
rect 33292 22148 33348 22206
rect 33516 22148 33572 23212
rect 33628 23154 33684 23884
rect 33740 23874 33796 23884
rect 34188 23492 34244 23502
rect 34244 23436 34356 23492
rect 34188 23426 34244 23436
rect 33628 23102 33630 23154
rect 33682 23102 33684 23154
rect 33628 22260 33684 23102
rect 33852 23154 33908 23166
rect 33852 23102 33854 23154
rect 33906 23102 33908 23154
rect 33852 22596 33908 23102
rect 33852 22530 33908 22540
rect 34300 22594 34356 23436
rect 34300 22542 34302 22594
rect 34354 22542 34356 22594
rect 34300 22530 34356 22542
rect 34636 22594 34692 24780
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 34972 23156 35028 23166
rect 34972 23062 35028 23100
rect 35644 23042 35700 23054
rect 35644 22990 35646 23042
rect 35698 22990 35700 23042
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34636 22542 34638 22594
rect 34690 22542 34692 22594
rect 34412 22484 34468 22494
rect 33852 22372 33908 22382
rect 34412 22372 34468 22428
rect 33852 22370 34468 22372
rect 33852 22318 33854 22370
rect 33906 22318 34468 22370
rect 33852 22316 34468 22318
rect 33852 22306 33908 22316
rect 33628 22194 33684 22204
rect 33292 22092 33572 22148
rect 34188 22148 34244 22158
rect 31948 21746 32004 21756
rect 33964 21812 34020 21822
rect 31836 21634 31892 21644
rect 32060 21588 32116 21598
rect 31836 21476 31892 21486
rect 31836 21382 31892 21420
rect 31612 20626 31668 20636
rect 31724 21362 31780 21374
rect 31724 21310 31726 21362
rect 31778 21310 31780 21362
rect 31276 20578 31332 20590
rect 31276 20526 31278 20578
rect 31330 20526 31332 20578
rect 31164 20020 31220 20030
rect 31276 20020 31332 20526
rect 31388 20580 31444 20590
rect 31388 20578 31556 20580
rect 31388 20526 31390 20578
rect 31442 20526 31556 20578
rect 31388 20524 31556 20526
rect 31388 20514 31444 20524
rect 31388 20020 31444 20030
rect 31276 20018 31444 20020
rect 31276 19966 31390 20018
rect 31442 19966 31444 20018
rect 31276 19964 31444 19966
rect 31164 19926 31220 19964
rect 31388 19954 31444 19964
rect 31052 19796 31108 19806
rect 31500 19796 31556 20524
rect 31612 20020 31668 20030
rect 31724 20020 31780 21310
rect 31612 20018 31780 20020
rect 31612 19966 31614 20018
rect 31666 19966 31780 20018
rect 31612 19964 31780 19966
rect 31612 19954 31668 19964
rect 31724 19908 31780 19964
rect 31724 19842 31780 19852
rect 31052 19702 31108 19740
rect 31388 19740 31556 19796
rect 31948 19796 32004 19806
rect 31388 19572 31444 19740
rect 31164 19236 31220 19246
rect 31164 18452 31220 19180
rect 30940 17890 30996 17902
rect 30940 17838 30942 17890
rect 30994 17838 30996 17890
rect 30940 17556 30996 17838
rect 30940 17490 30996 17500
rect 30828 17276 31108 17332
rect 30492 17154 30548 17164
rect 30492 16996 30548 17006
rect 30044 16828 30324 16884
rect 29932 16270 29934 16322
rect 29986 16270 29988 16322
rect 29932 16258 29988 16270
rect 30268 15988 30324 16828
rect 30492 16882 30548 16940
rect 30492 16830 30494 16882
rect 30546 16830 30548 16882
rect 30492 16818 30548 16830
rect 30268 15986 30996 15988
rect 30268 15934 30270 15986
rect 30322 15934 30996 15986
rect 30268 15932 30996 15934
rect 30268 15922 30324 15932
rect 30044 15876 30100 15886
rect 30044 15782 30100 15820
rect 30940 15204 30996 15932
rect 31052 15426 31108 17276
rect 31164 16210 31220 18396
rect 31164 16158 31166 16210
rect 31218 16158 31220 16210
rect 31164 16146 31220 16158
rect 31052 15374 31054 15426
rect 31106 15374 31108 15426
rect 31052 15362 31108 15374
rect 29820 15092 30100 15148
rect 29708 14532 29764 14542
rect 29596 14530 29764 14532
rect 29596 14478 29710 14530
rect 29762 14478 29764 14530
rect 29596 14476 29764 14478
rect 29708 14466 29764 14476
rect 29148 14418 29204 14430
rect 29148 14366 29150 14418
rect 29202 14366 29204 14418
rect 28924 13748 28980 13758
rect 28924 13654 28980 13692
rect 28364 12870 28420 12908
rect 28140 12740 28196 12750
rect 27916 12126 27918 12178
rect 27970 12126 27972 12178
rect 27692 11844 27748 11854
rect 27580 11284 27636 11294
rect 27580 10722 27636 11228
rect 27580 10670 27582 10722
rect 27634 10670 27636 10722
rect 27580 10658 27636 10670
rect 27356 10322 27412 10332
rect 27356 9940 27412 9950
rect 27356 9846 27412 9884
rect 27580 9940 27636 9950
rect 27244 9650 27300 9660
rect 27468 9492 27524 9502
rect 27132 9436 27468 9492
rect 27468 9426 27524 9436
rect 27020 9268 27076 9278
rect 27580 9268 27636 9884
rect 27020 9266 27636 9268
rect 27020 9214 27022 9266
rect 27074 9214 27582 9266
rect 27634 9214 27636 9266
rect 27020 9212 27636 9214
rect 27020 9202 27076 9212
rect 27580 9202 27636 9212
rect 27580 9044 27636 9054
rect 27580 8596 27636 8988
rect 27580 8530 27636 8540
rect 27020 8372 27076 8382
rect 27692 8372 27748 11788
rect 27804 11620 27860 11630
rect 27916 11620 27972 12126
rect 28028 12738 28196 12740
rect 28028 12686 28142 12738
rect 28194 12686 28196 12738
rect 28028 12684 28196 12686
rect 28028 12180 28084 12684
rect 28140 12674 28196 12684
rect 28476 12738 28532 12750
rect 28476 12686 28478 12738
rect 28530 12686 28532 12738
rect 28028 12114 28084 12124
rect 28252 12290 28308 12302
rect 28252 12238 28254 12290
rect 28306 12238 28308 12290
rect 28252 12180 28308 12238
rect 28252 12114 28308 12124
rect 28476 12178 28532 12686
rect 29148 12740 29204 14366
rect 29596 14308 29652 14318
rect 29596 14306 29764 14308
rect 29596 14254 29598 14306
rect 29650 14254 29764 14306
rect 29596 14252 29764 14254
rect 29596 14242 29652 14252
rect 29484 13860 29540 13870
rect 29484 13858 29652 13860
rect 29484 13806 29486 13858
rect 29538 13806 29652 13858
rect 29484 13804 29652 13806
rect 29484 13794 29540 13804
rect 29260 13748 29316 13758
rect 29260 13746 29428 13748
rect 29260 13694 29262 13746
rect 29314 13694 29428 13746
rect 29260 13692 29428 13694
rect 29260 13682 29316 13692
rect 29148 12674 29204 12684
rect 29372 12628 29428 13692
rect 29484 13634 29540 13646
rect 29484 13582 29486 13634
rect 29538 13582 29540 13634
rect 29484 13186 29540 13582
rect 29484 13134 29486 13186
rect 29538 13134 29540 13186
rect 29484 13122 29540 13134
rect 29596 13188 29652 13804
rect 29596 13122 29652 13132
rect 29708 13076 29764 14252
rect 29932 13748 29988 13758
rect 29932 13186 29988 13692
rect 29932 13134 29934 13186
rect 29986 13134 29988 13186
rect 29932 13122 29988 13134
rect 29708 13010 29764 13020
rect 29036 12292 29092 12302
rect 29036 12198 29092 12236
rect 28476 12126 28478 12178
rect 28530 12126 28532 12178
rect 28476 11844 28532 12126
rect 29372 12180 29428 12572
rect 29596 12962 29652 12974
rect 29596 12910 29598 12962
rect 29650 12910 29652 12962
rect 29484 12180 29540 12190
rect 29372 12178 29540 12180
rect 29372 12126 29486 12178
rect 29538 12126 29540 12178
rect 29372 12124 29540 12126
rect 29484 12114 29540 12124
rect 29596 12180 29652 12910
rect 29596 12114 29652 12124
rect 29820 12962 29876 12974
rect 29820 12910 29822 12962
rect 29874 12910 29876 12962
rect 28476 11778 28532 11788
rect 29484 11956 29540 11966
rect 27804 11618 27972 11620
rect 27804 11566 27806 11618
rect 27858 11566 27972 11618
rect 27804 11564 27972 11566
rect 27804 11554 27860 11564
rect 27020 8370 27748 8372
rect 27020 8318 27022 8370
rect 27074 8318 27748 8370
rect 27020 8316 27748 8318
rect 27020 8306 27076 8316
rect 27692 8258 27748 8316
rect 27692 8206 27694 8258
rect 27746 8206 27748 8258
rect 27692 8194 27748 8206
rect 27804 11396 27860 11406
rect 27804 10724 27860 11340
rect 29484 11394 29540 11900
rect 29820 11956 29876 12910
rect 29932 12180 29988 12190
rect 29932 12086 29988 12124
rect 29820 11890 29876 11900
rect 30044 11620 30100 15092
rect 30940 15092 31220 15204
rect 31388 15148 31444 19516
rect 31948 19346 32004 19740
rect 31948 19294 31950 19346
rect 32002 19294 32004 19346
rect 31948 19282 32004 19294
rect 31276 15092 31444 15148
rect 31500 18564 31556 18574
rect 31500 15428 31556 18508
rect 32060 18452 32116 21532
rect 33964 21586 34020 21756
rect 33964 21534 33966 21586
rect 34018 21534 34020 21586
rect 33964 21522 34020 21534
rect 34188 21586 34244 22092
rect 34636 21812 34692 22542
rect 35308 22596 35364 22606
rect 35084 22484 35140 22494
rect 35084 22390 35140 22428
rect 34748 22372 34804 22382
rect 34748 22278 34804 22316
rect 35308 22258 35364 22540
rect 35644 22372 35700 22990
rect 35644 22306 35700 22316
rect 35308 22206 35310 22258
rect 35362 22206 35364 22258
rect 35308 22194 35364 22206
rect 35196 22148 35252 22158
rect 35196 22054 35252 22092
rect 34188 21534 34190 21586
rect 34242 21534 34244 21586
rect 34188 21522 34244 21534
rect 34412 21756 34692 21812
rect 34412 21586 34468 21756
rect 34412 21534 34414 21586
rect 34466 21534 34468 21586
rect 34412 21522 34468 21534
rect 34524 21362 34580 21374
rect 34524 21310 34526 21362
rect 34578 21310 34580 21362
rect 34524 20188 34580 21310
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34524 20132 34804 20188
rect 34748 20130 34804 20132
rect 34748 20078 34750 20130
rect 34802 20078 34804 20130
rect 34748 20066 34804 20078
rect 33964 20018 34020 20030
rect 33964 19966 33966 20018
rect 34018 19966 34020 20018
rect 33964 19236 34020 19966
rect 35196 19628 35460 19638
rect 34076 19572 34132 19582
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34076 19348 34132 19516
rect 34076 19346 34468 19348
rect 34076 19294 34078 19346
rect 34130 19294 34468 19346
rect 34076 19292 34468 19294
rect 34076 19282 34132 19292
rect 33964 19170 34020 19180
rect 32060 18386 32116 18396
rect 33516 18562 33572 18574
rect 33516 18510 33518 18562
rect 33570 18510 33572 18562
rect 33516 18452 33572 18510
rect 33516 18386 33572 18396
rect 33852 18450 33908 18462
rect 33852 18398 33854 18450
rect 33906 18398 33908 18450
rect 32508 18340 32564 18350
rect 32508 18246 32564 18284
rect 33852 18340 33908 18398
rect 33516 17220 33572 17230
rect 33516 17106 33572 17164
rect 33516 17054 33518 17106
rect 33570 17054 33572 17106
rect 33516 17042 33572 17054
rect 32956 16996 33012 17006
rect 31724 16884 31780 16894
rect 31780 16828 31892 16884
rect 31724 16790 31780 16828
rect 30940 14308 30996 15092
rect 31276 14756 31332 15092
rect 31052 14700 31332 14756
rect 31052 14530 31108 14700
rect 31052 14478 31054 14530
rect 31106 14478 31108 14530
rect 31052 14466 31108 14478
rect 31276 14532 31332 14542
rect 31276 14438 31332 14476
rect 31500 14530 31556 15372
rect 31836 15314 31892 16828
rect 32956 16098 33012 16940
rect 33852 16882 33908 18284
rect 34076 18452 34132 18462
rect 34076 17666 34132 18396
rect 34188 18004 34244 18014
rect 34188 17778 34244 17948
rect 34188 17726 34190 17778
rect 34242 17726 34244 17778
rect 34188 17714 34244 17726
rect 34076 17614 34078 17666
rect 34130 17614 34132 17666
rect 34076 17602 34132 17614
rect 34412 17666 34468 19292
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35868 18004 35924 26350
rect 36204 19908 36260 31052
rect 36652 31042 36708 31052
rect 36876 31106 36932 31276
rect 36876 31054 36878 31106
rect 36930 31054 36932 31106
rect 36876 31042 36932 31054
rect 37100 30994 37156 31006
rect 37100 30942 37102 30994
rect 37154 30942 37156 30994
rect 36540 30884 36596 30894
rect 36540 30790 36596 30828
rect 36988 30212 37044 30222
rect 37100 30212 37156 30942
rect 37436 30996 37492 32732
rect 37548 31220 37604 38612
rect 38108 38162 38164 38612
rect 38108 38110 38110 38162
rect 38162 38110 38164 38162
rect 38108 38098 38164 38110
rect 38556 38162 38612 38612
rect 38556 38110 38558 38162
rect 38610 38110 38612 38162
rect 38556 38098 38612 38110
rect 38892 37826 38948 38612
rect 39676 38164 39732 38782
rect 39900 38836 39956 38846
rect 39900 38742 39956 38780
rect 39676 38098 39732 38108
rect 39788 38050 39844 38062
rect 39788 37998 39790 38050
rect 39842 37998 39844 38050
rect 38892 37774 38894 37826
rect 38946 37774 38948 37826
rect 38892 37268 38948 37774
rect 39452 37828 39508 37838
rect 39788 37828 39844 37998
rect 40012 37938 40068 39788
rect 40012 37886 40014 37938
rect 40066 37886 40068 37938
rect 40012 37874 40068 37886
rect 40236 37940 40292 40348
rect 40348 38724 40404 38734
rect 40348 38630 40404 38668
rect 40348 37940 40404 37950
rect 40236 37938 40404 37940
rect 40236 37886 40350 37938
rect 40402 37886 40404 37938
rect 40236 37884 40404 37886
rect 40348 37874 40404 37884
rect 39452 37826 39788 37828
rect 39452 37774 39454 37826
rect 39506 37774 39788 37826
rect 39452 37772 39788 37774
rect 39452 37762 39508 37772
rect 39788 37762 39844 37772
rect 38892 37202 38948 37212
rect 37996 37154 38052 37166
rect 40124 37156 40180 37166
rect 37996 37102 37998 37154
rect 38050 37102 38052 37154
rect 37772 36372 37828 36382
rect 37772 36370 37940 36372
rect 37772 36318 37774 36370
rect 37826 36318 37940 36370
rect 37772 36316 37940 36318
rect 37772 36306 37828 36316
rect 37772 35252 37828 35262
rect 37772 34916 37828 35196
rect 37660 34914 37828 34916
rect 37660 34862 37774 34914
rect 37826 34862 37828 34914
rect 37660 34860 37828 34862
rect 37660 32564 37716 34860
rect 37772 34850 37828 34860
rect 37772 34692 37828 34702
rect 37884 34692 37940 36316
rect 37996 36258 38052 37102
rect 40012 37154 40180 37156
rect 40012 37102 40126 37154
rect 40178 37102 40180 37154
rect 40012 37100 40180 37102
rect 38108 36932 38164 36942
rect 38108 36482 38164 36876
rect 40012 36596 40068 37100
rect 40124 37090 40180 37100
rect 38108 36430 38110 36482
rect 38162 36430 38164 36482
rect 38108 36418 38164 36430
rect 39340 36594 40068 36596
rect 39340 36542 40014 36594
rect 40066 36542 40068 36594
rect 39340 36540 40068 36542
rect 39340 36482 39396 36540
rect 40012 36530 40068 36540
rect 39340 36430 39342 36482
rect 39394 36430 39396 36482
rect 39340 36418 39396 36430
rect 38332 36372 38388 36382
rect 38332 36278 38388 36316
rect 39228 36372 39284 36382
rect 39228 36278 39284 36316
rect 37996 36206 37998 36258
rect 38050 36206 38052 36258
rect 37996 36194 38052 36206
rect 39116 36258 39172 36270
rect 39116 36206 39118 36258
rect 39170 36206 39172 36258
rect 38668 36036 38724 36046
rect 38444 34802 38500 34814
rect 38444 34750 38446 34802
rect 38498 34750 38500 34802
rect 37828 34636 37940 34692
rect 38220 34692 38276 34702
rect 37772 34626 37828 34636
rect 37772 34130 37828 34142
rect 37772 34078 37774 34130
rect 37826 34078 37828 34130
rect 37772 33684 37828 34078
rect 37828 33628 38052 33684
rect 37772 33618 37828 33628
rect 37996 33458 38052 33628
rect 37996 33406 37998 33458
rect 38050 33406 38052 33458
rect 37996 33348 38052 33406
rect 37996 33282 38052 33292
rect 38220 33346 38276 34636
rect 38444 33458 38500 34750
rect 38444 33406 38446 33458
rect 38498 33406 38500 33458
rect 38444 33394 38500 33406
rect 38220 33294 38222 33346
rect 38274 33294 38276 33346
rect 38220 33282 38276 33294
rect 38668 33346 38724 35980
rect 39116 34244 39172 36206
rect 39564 36260 39620 36270
rect 39564 36166 39620 36204
rect 40124 36260 40180 36270
rect 40460 36260 40516 40572
rect 40684 40562 40740 40572
rect 40572 40180 40628 40190
rect 40572 39060 40628 40124
rect 40572 37380 40628 39004
rect 40684 40068 40740 40078
rect 40684 38668 40740 40012
rect 40796 39060 40852 42028
rect 40908 41970 40964 41982
rect 40908 41918 40910 41970
rect 40962 41918 40964 41970
rect 40908 40628 40964 41918
rect 41020 41972 41076 41982
rect 41020 41878 41076 41916
rect 41132 41410 41188 42252
rect 41132 41358 41134 41410
rect 41186 41358 41188 41410
rect 41132 41346 41188 41358
rect 41244 41970 41300 41982
rect 41244 41918 41246 41970
rect 41298 41918 41300 41970
rect 41132 41076 41188 41086
rect 40908 40572 41076 40628
rect 40908 40402 40964 40414
rect 40908 40350 40910 40402
rect 40962 40350 40964 40402
rect 40908 40180 40964 40350
rect 40908 40114 40964 40124
rect 41020 39956 41076 40572
rect 41132 40626 41188 41020
rect 41132 40574 41134 40626
rect 41186 40574 41188 40626
rect 41132 40562 41188 40574
rect 41244 40628 41300 41918
rect 41356 41972 41412 41982
rect 41356 41878 41412 41916
rect 41468 41188 41524 43598
rect 42364 43428 42420 43438
rect 42364 43334 42420 43372
rect 41804 43316 41860 43326
rect 41692 43314 41860 43316
rect 41692 43262 41806 43314
rect 41858 43262 41860 43314
rect 41692 43260 41860 43262
rect 41692 41748 41748 43260
rect 41804 43250 41860 43260
rect 42140 43314 42196 43326
rect 42140 43262 42142 43314
rect 42194 43262 42196 43314
rect 41916 42868 41972 42878
rect 41972 42812 42084 42868
rect 41916 42774 41972 42812
rect 42028 42194 42084 42812
rect 42028 42142 42030 42194
rect 42082 42142 42084 42194
rect 42028 42130 42084 42142
rect 41804 42084 41860 42094
rect 41804 41990 41860 42028
rect 41916 41972 41972 41982
rect 41916 41878 41972 41916
rect 41692 41692 41860 41748
rect 41692 41188 41748 41198
rect 41468 41186 41748 41188
rect 41468 41134 41694 41186
rect 41746 41134 41748 41186
rect 41468 41132 41748 41134
rect 41692 41122 41748 41132
rect 41244 40562 41300 40572
rect 41692 40852 41748 40862
rect 41468 40516 41524 40526
rect 41468 40422 41524 40460
rect 41244 40404 41300 40414
rect 41244 40310 41300 40348
rect 40908 39900 41076 39956
rect 40908 39284 40964 39900
rect 41020 39732 41076 39742
rect 41020 39730 41188 39732
rect 41020 39678 41022 39730
rect 41074 39678 41188 39730
rect 41020 39676 41188 39678
rect 41020 39666 41076 39676
rect 40908 39218 40964 39228
rect 40908 39060 40964 39070
rect 40796 39004 40908 39060
rect 40908 38966 40964 39004
rect 41132 38948 41188 39676
rect 41692 39618 41748 40796
rect 41804 40404 41860 41692
rect 42140 40628 42196 43262
rect 42812 42978 42868 44156
rect 43820 43764 43876 43774
rect 42812 42926 42814 42978
rect 42866 42926 42868 42978
rect 42812 42914 42868 42926
rect 42924 43538 42980 43550
rect 42924 43486 42926 43538
rect 42978 43486 42980 43538
rect 42476 42756 42532 42766
rect 42252 42644 42308 42654
rect 42252 42550 42308 42588
rect 42364 41970 42420 41982
rect 42364 41918 42366 41970
rect 42418 41918 42420 41970
rect 42364 41748 42420 41918
rect 42364 41682 42420 41692
rect 42140 40562 42196 40572
rect 41804 40348 41972 40404
rect 41804 40178 41860 40190
rect 41804 40126 41806 40178
rect 41858 40126 41860 40178
rect 41804 40068 41860 40126
rect 41804 40002 41860 40012
rect 41916 39732 41972 40348
rect 42140 40292 42196 40302
rect 42140 40198 42196 40236
rect 42364 40290 42420 40302
rect 42364 40238 42366 40290
rect 42418 40238 42420 40290
rect 41692 39566 41694 39618
rect 41746 39566 41748 39618
rect 41692 39554 41748 39566
rect 41804 39676 41972 39732
rect 41132 38854 41188 38892
rect 41356 38946 41412 38958
rect 41356 38894 41358 38946
rect 41410 38894 41412 38946
rect 41020 38836 41076 38846
rect 41020 38742 41076 38780
rect 41356 38724 41412 38894
rect 41412 38668 41524 38724
rect 40684 38612 41076 38668
rect 41356 38658 41412 38668
rect 40908 38164 40964 38174
rect 40572 37314 40628 37324
rect 40684 37938 40740 37950
rect 40684 37886 40686 37938
rect 40738 37886 40740 37938
rect 40684 37044 40740 37886
rect 40684 36978 40740 36988
rect 40572 36706 40628 36718
rect 40572 36654 40574 36706
rect 40626 36654 40628 36706
rect 40572 36594 40628 36654
rect 40572 36542 40574 36594
rect 40626 36542 40628 36594
rect 40572 36530 40628 36542
rect 40124 36258 40516 36260
rect 40124 36206 40126 36258
rect 40178 36206 40516 36258
rect 40124 36204 40516 36206
rect 40124 36036 40180 36204
rect 40124 35970 40180 35980
rect 40908 35140 40964 38108
rect 41020 38050 41076 38612
rect 41020 37998 41022 38050
rect 41074 37998 41076 38050
rect 41020 37986 41076 37998
rect 41356 37940 41412 37950
rect 41356 37846 41412 37884
rect 41468 37716 41524 38668
rect 41804 38668 41860 39676
rect 41916 39060 41972 39070
rect 41916 38966 41972 39004
rect 42140 38836 42196 38846
rect 42364 38836 42420 40238
rect 42476 40292 42532 42700
rect 42812 41970 42868 41982
rect 42812 41918 42814 41970
rect 42866 41918 42868 41970
rect 42476 40226 42532 40236
rect 42700 40402 42756 40414
rect 42700 40350 42702 40402
rect 42754 40350 42756 40402
rect 42476 39396 42532 39406
rect 42532 39340 42644 39396
rect 42476 39330 42532 39340
rect 42140 38834 42420 38836
rect 42140 38782 42142 38834
rect 42194 38782 42420 38834
rect 42140 38780 42420 38782
rect 42476 39172 42532 39182
rect 42476 38834 42532 39116
rect 42476 38782 42478 38834
rect 42530 38782 42532 38834
rect 42028 38722 42084 38734
rect 42028 38670 42030 38722
rect 42082 38670 42084 38722
rect 41804 38612 41972 38668
rect 41692 38052 41748 38062
rect 41692 37958 41748 37996
rect 41132 37660 41524 37716
rect 41020 37268 41076 37278
rect 41020 36706 41076 37212
rect 41020 36654 41022 36706
rect 41074 36654 41076 36706
rect 41020 36260 41076 36654
rect 41132 36372 41188 37660
rect 41692 37380 41748 37390
rect 41580 37324 41692 37380
rect 41580 36482 41636 37324
rect 41692 37314 41748 37324
rect 41692 37154 41748 37166
rect 41692 37102 41694 37154
rect 41746 37102 41748 37154
rect 41692 36596 41748 37102
rect 41804 36596 41860 36606
rect 41692 36594 41860 36596
rect 41692 36542 41806 36594
rect 41858 36542 41860 36594
rect 41692 36540 41860 36542
rect 41804 36530 41860 36540
rect 41580 36430 41582 36482
rect 41634 36430 41636 36482
rect 41580 36418 41636 36430
rect 41132 36316 41524 36372
rect 41020 36258 41188 36260
rect 41020 36206 41022 36258
rect 41074 36206 41188 36258
rect 41020 36204 41188 36206
rect 41020 36194 41076 36204
rect 41132 35586 41188 36204
rect 41468 35924 41524 36316
rect 41804 36260 41860 36270
rect 41580 35924 41636 35934
rect 41468 35922 41636 35924
rect 41468 35870 41582 35922
rect 41634 35870 41636 35922
rect 41468 35868 41636 35870
rect 41580 35858 41636 35868
rect 41132 35534 41134 35586
rect 41186 35534 41188 35586
rect 41020 35140 41076 35150
rect 40908 35138 41076 35140
rect 40908 35086 41022 35138
rect 41074 35086 41076 35138
rect 40908 35084 41076 35086
rect 40124 35028 40180 35038
rect 39116 34178 39172 34188
rect 39788 34244 39844 34254
rect 38668 33294 38670 33346
rect 38722 33294 38724 33346
rect 38668 33282 38724 33294
rect 39228 33348 39284 33358
rect 39228 33254 39284 33292
rect 38892 33234 38948 33246
rect 38892 33182 38894 33234
rect 38946 33182 38948 33234
rect 38892 33012 38948 33182
rect 38892 32946 38948 32956
rect 39116 33236 39172 33246
rect 38220 32788 38276 32798
rect 38220 32694 38276 32732
rect 38892 32788 38948 32798
rect 38892 32694 38948 32732
rect 38556 32676 38612 32686
rect 38556 32582 38612 32620
rect 37660 32562 38164 32564
rect 37660 32510 37662 32562
rect 37714 32510 38164 32562
rect 37660 32508 38164 32510
rect 37660 32498 37716 32508
rect 38108 31890 38164 32508
rect 38108 31838 38110 31890
rect 38162 31838 38164 31890
rect 38108 31826 38164 31838
rect 39116 31780 39172 33180
rect 39228 32788 39284 32798
rect 39228 32694 39284 32732
rect 39788 32786 39844 34188
rect 40124 34018 40180 34972
rect 40572 35026 40628 35038
rect 40572 34974 40574 35026
rect 40626 34974 40628 35026
rect 40572 34804 40628 34974
rect 40908 34804 40964 34814
rect 40572 34802 40964 34804
rect 40572 34750 40910 34802
rect 40962 34750 40964 34802
rect 40572 34748 40964 34750
rect 40572 34132 40628 34748
rect 40908 34738 40964 34748
rect 40124 33966 40126 34018
rect 40178 33966 40180 34018
rect 40124 33954 40180 33966
rect 40236 34076 40628 34132
rect 39788 32734 39790 32786
rect 39842 32734 39844 32786
rect 39788 32722 39844 32734
rect 39900 33012 39956 33022
rect 39900 32786 39956 32956
rect 39900 32734 39902 32786
rect 39954 32734 39956 32786
rect 39900 32722 39956 32734
rect 40012 32788 40068 32798
rect 40236 32788 40292 34076
rect 40012 32786 40292 32788
rect 40012 32734 40014 32786
rect 40066 32734 40292 32786
rect 40012 32732 40292 32734
rect 40908 33012 40964 33022
rect 40012 32722 40068 32732
rect 40460 32676 40516 32686
rect 40460 32562 40516 32620
rect 40460 32510 40462 32562
rect 40514 32510 40516 32562
rect 40460 32498 40516 32510
rect 40908 32674 40964 32956
rect 40908 32622 40910 32674
rect 40962 32622 40964 32674
rect 40908 32564 40964 32622
rect 41020 32676 41076 35084
rect 41132 35028 41188 35534
rect 41804 35252 41860 36204
rect 41916 35924 41972 38612
rect 42028 37492 42084 38670
rect 42140 38668 42196 38780
rect 42476 38724 42532 38782
rect 42140 38612 42308 38668
rect 42476 38658 42532 38668
rect 42028 37436 42196 37492
rect 42140 36482 42196 37436
rect 42252 37156 42308 38612
rect 42252 37090 42308 37100
rect 42140 36430 42142 36482
rect 42194 36430 42196 36482
rect 42140 36418 42196 36430
rect 41916 35858 41972 35868
rect 42028 36370 42084 36382
rect 42028 36318 42030 36370
rect 42082 36318 42084 36370
rect 41804 35186 41860 35196
rect 41468 35028 41524 35038
rect 41132 34972 41468 35028
rect 41468 34934 41524 34972
rect 42028 34244 42084 36318
rect 42140 35700 42196 35710
rect 42140 35606 42196 35644
rect 42588 35700 42644 39340
rect 42700 37940 42756 40350
rect 42812 39844 42868 41918
rect 42924 41860 42980 43486
rect 43708 42868 43764 42878
rect 43708 42774 43764 42812
rect 43484 42756 43540 42766
rect 43484 42662 43540 42700
rect 43148 42532 43204 42542
rect 43148 42438 43204 42476
rect 42924 41794 42980 41804
rect 43820 41524 43876 43708
rect 43932 42308 43988 44380
rect 44044 42980 44100 47740
rect 44380 45220 44436 49200
rect 44604 46116 44660 46126
rect 44604 46022 44660 46060
rect 44380 45154 44436 45164
rect 44156 45108 44212 45118
rect 44156 45014 44212 45052
rect 44716 43316 44772 49756
rect 45024 49200 45136 50000
rect 45696 49200 45808 50000
rect 45052 44884 45108 49200
rect 45052 44818 45108 44828
rect 45164 49140 45220 49150
rect 45164 44772 45220 49084
rect 45164 44706 45220 44716
rect 45276 47124 45332 47134
rect 44828 44322 44884 44334
rect 44828 44270 44830 44322
rect 44882 44270 44884 44322
rect 44828 43540 44884 44270
rect 44828 43474 44884 43484
rect 44716 43250 44772 43260
rect 44940 43426 44996 43438
rect 44940 43374 44942 43426
rect 44994 43374 44996 43426
rect 44044 42914 44100 42924
rect 44828 42756 44884 42766
rect 44828 42642 44884 42700
rect 44828 42590 44830 42642
rect 44882 42590 44884 42642
rect 44828 42578 44884 42590
rect 44156 42530 44212 42542
rect 44156 42478 44158 42530
rect 44210 42478 44212 42530
rect 43932 42242 43988 42252
rect 44044 42420 44100 42430
rect 43596 41468 43876 41524
rect 43036 40628 43092 40638
rect 43092 40572 43204 40628
rect 43036 40562 43092 40572
rect 42812 39778 42868 39788
rect 43036 40292 43092 40302
rect 42812 38948 42868 38958
rect 42812 38854 42868 38892
rect 43036 38834 43092 40236
rect 43036 38782 43038 38834
rect 43090 38782 43092 38834
rect 43036 38770 43092 38782
rect 42700 37874 42756 37884
rect 43036 36708 43092 36718
rect 43148 36708 43204 40572
rect 43596 39842 43652 41468
rect 44044 41410 44100 42364
rect 44044 41358 44046 41410
rect 44098 41358 44100 41410
rect 44044 41346 44100 41358
rect 44156 41188 44212 42478
rect 44940 41748 44996 43374
rect 45164 42642 45220 42654
rect 45164 42590 45166 42642
rect 45218 42590 45220 42642
rect 44940 41682 44996 41692
rect 45052 41746 45108 41758
rect 45052 41694 45054 41746
rect 45106 41694 45108 41746
rect 44940 41188 44996 41198
rect 44156 41186 44996 41188
rect 44156 41134 44942 41186
rect 44994 41134 44996 41186
rect 44156 41132 44996 41134
rect 43596 39790 43598 39842
rect 43650 39790 43652 39842
rect 43596 39778 43652 39790
rect 44828 39396 44884 39406
rect 44716 39394 44884 39396
rect 44716 39342 44830 39394
rect 44882 39342 44884 39394
rect 44716 39340 44884 39342
rect 44268 39172 44324 39182
rect 43708 38722 43764 38734
rect 43708 38670 43710 38722
rect 43762 38670 43764 38722
rect 43372 38610 43428 38622
rect 43372 38558 43374 38610
rect 43426 38558 43428 38610
rect 43372 38052 43428 38558
rect 43596 38276 43652 38286
rect 43596 38182 43652 38220
rect 43372 37986 43428 37996
rect 43708 36932 43764 38670
rect 43820 37156 43876 37166
rect 43820 37062 43876 37100
rect 44268 37154 44324 39116
rect 44604 38948 44660 38958
rect 44604 37492 44660 38892
rect 44716 37604 44772 39340
rect 44828 39330 44884 39340
rect 44940 38724 44996 41132
rect 45052 41188 45108 41694
rect 45052 41122 45108 41132
rect 45052 40178 45108 40190
rect 45052 40126 45054 40178
rect 45106 40126 45108 40178
rect 45052 39060 45108 40126
rect 45164 39620 45220 42590
rect 45276 41412 45332 47068
rect 45388 44996 45444 45006
rect 45388 44902 45444 44940
rect 45724 44660 45780 49200
rect 47180 46452 47236 46462
rect 45724 44594 45780 44604
rect 46508 45666 46564 45678
rect 46508 45614 46510 45666
rect 46562 45614 46564 45666
rect 45836 44548 45892 44558
rect 45836 44454 45892 44492
rect 46508 43708 46564 45614
rect 46060 43652 46564 43708
rect 46844 45666 46900 45678
rect 46844 45614 46846 45666
rect 46898 45614 46900 45666
rect 46844 43652 46900 45614
rect 47180 45330 47236 46396
rect 47404 45892 47460 45902
rect 47404 45890 48020 45892
rect 47404 45838 47406 45890
rect 47458 45838 48020 45890
rect 47404 45836 48020 45838
rect 47404 45826 47460 45836
rect 47180 45278 47182 45330
rect 47234 45278 47236 45330
rect 47180 45266 47236 45278
rect 47516 45666 47572 45678
rect 47516 45614 47518 45666
rect 47570 45614 47572 45666
rect 47516 45220 47572 45614
rect 47404 45164 47572 45220
rect 47628 45666 47684 45678
rect 47628 45614 47630 45666
rect 47682 45614 47684 45666
rect 45836 43538 45892 43550
rect 45836 43486 45838 43538
rect 45890 43486 45892 43538
rect 45612 42756 45668 42766
rect 45276 41346 45332 41356
rect 45388 42754 45668 42756
rect 45388 42702 45614 42754
rect 45666 42702 45668 42754
rect 45388 42700 45668 42702
rect 45388 40404 45444 42700
rect 45612 42690 45668 42700
rect 45836 42196 45892 43486
rect 45164 39526 45220 39564
rect 45276 40348 45444 40404
rect 45500 42140 45892 42196
rect 45052 38994 45108 39004
rect 45276 38668 45332 40348
rect 44940 38658 44996 38668
rect 45164 38612 45332 38668
rect 45388 38724 45444 38734
rect 44828 38052 44884 38062
rect 44828 37958 44884 37996
rect 45164 37938 45220 38612
rect 45164 37886 45166 37938
rect 45218 37886 45220 37938
rect 45164 37874 45220 37886
rect 44716 37548 45108 37604
rect 44604 37436 44884 37492
rect 44716 37268 44772 37278
rect 44268 37102 44270 37154
rect 44322 37102 44324 37154
rect 44268 37042 44324 37102
rect 44268 36990 44270 37042
rect 44322 36990 44324 37042
rect 44268 36978 44324 36990
rect 44380 37266 44772 37268
rect 44380 37214 44718 37266
rect 44770 37214 44772 37266
rect 44380 37212 44772 37214
rect 43036 36706 43204 36708
rect 43036 36654 43038 36706
rect 43090 36654 43204 36706
rect 43036 36652 43204 36654
rect 43484 36876 43764 36932
rect 43036 36642 43092 36652
rect 42812 36370 42868 36382
rect 42812 36318 42814 36370
rect 42866 36318 42868 36370
rect 42812 36148 42868 36318
rect 43372 36260 43428 36270
rect 43372 36166 43428 36204
rect 42812 36082 42868 36092
rect 43484 36148 43540 36876
rect 44380 36708 44436 37212
rect 44716 37202 44772 37212
rect 44156 36652 44436 36708
rect 44492 37042 44548 37054
rect 44492 36990 44494 37042
rect 44546 36990 44548 37042
rect 44156 36594 44212 36652
rect 44156 36542 44158 36594
rect 44210 36542 44212 36594
rect 44156 36530 44212 36542
rect 43484 36082 43540 36092
rect 43596 36482 43652 36494
rect 43820 36484 43876 36494
rect 43596 36430 43598 36482
rect 43650 36430 43652 36482
rect 43596 36372 43652 36430
rect 42924 35924 42980 35934
rect 42924 35830 42980 35868
rect 43260 35924 43316 35934
rect 43260 35830 43316 35868
rect 43596 35922 43652 36316
rect 43596 35870 43598 35922
rect 43650 35870 43652 35922
rect 43596 35858 43652 35870
rect 43708 36428 43820 36484
rect 43708 35700 43764 36428
rect 43820 36418 43876 36428
rect 44044 36258 44100 36270
rect 44044 36206 44046 36258
rect 44098 36206 44100 36258
rect 44044 36036 44100 36206
rect 44044 35970 44100 35980
rect 44268 36258 44324 36270
rect 44268 36206 44270 36258
rect 44322 36206 44324 36258
rect 42588 35606 42644 35644
rect 43596 35644 43764 35700
rect 43932 35700 43988 35710
rect 44268 35700 44324 36206
rect 43932 35698 44100 35700
rect 43932 35646 43934 35698
rect 43986 35646 44100 35698
rect 43932 35644 44100 35646
rect 42364 35588 42420 35598
rect 42364 35026 42420 35532
rect 43596 35138 43652 35644
rect 43932 35634 43988 35644
rect 43596 35086 43598 35138
rect 43650 35086 43652 35138
rect 43596 35074 43652 35086
rect 42364 34974 42366 35026
rect 42418 34974 42420 35026
rect 42364 34962 42420 34974
rect 42700 35028 42756 35038
rect 42700 34934 42756 34972
rect 43148 34916 43204 34926
rect 43148 34822 43204 34860
rect 43932 34916 43988 34926
rect 43932 34822 43988 34860
rect 43484 34804 43540 34814
rect 43484 34802 43652 34804
rect 43484 34750 43486 34802
rect 43538 34750 43652 34802
rect 43484 34748 43652 34750
rect 43484 34738 43540 34748
rect 42028 34188 42420 34244
rect 41468 34132 41524 34142
rect 41468 34130 41636 34132
rect 41468 34078 41470 34130
rect 41522 34078 41636 34130
rect 41468 34076 41636 34078
rect 41468 34066 41524 34076
rect 41580 33458 41636 34076
rect 42140 34020 42196 34030
rect 42140 34018 42308 34020
rect 42140 33966 42142 34018
rect 42194 33966 42308 34018
rect 42140 33964 42308 33966
rect 42140 33954 42196 33964
rect 41580 33406 41582 33458
rect 41634 33406 41636 33458
rect 41580 33236 41636 33406
rect 42252 33458 42308 33964
rect 42252 33406 42254 33458
rect 42306 33406 42308 33458
rect 42252 33394 42308 33406
rect 42364 33348 42420 34188
rect 42700 33348 42756 33358
rect 43372 33348 43428 33358
rect 42364 33346 42644 33348
rect 42364 33294 42366 33346
rect 42418 33294 42644 33346
rect 42364 33292 42644 33294
rect 42364 33282 42420 33292
rect 41580 33170 41636 33180
rect 42140 33234 42196 33246
rect 42140 33182 42142 33234
rect 42194 33182 42196 33234
rect 42140 33012 42196 33182
rect 42140 32946 42196 32956
rect 41804 32788 41860 32798
rect 41804 32694 41860 32732
rect 41020 32620 41188 32676
rect 40908 32498 40964 32508
rect 41132 32562 41188 32620
rect 41132 32510 41134 32562
rect 41186 32510 41188 32562
rect 41132 32498 41188 32510
rect 41356 32564 41412 32574
rect 41356 32470 41412 32508
rect 41916 32564 41972 32574
rect 41916 32470 41972 32508
rect 42028 32562 42084 32574
rect 42028 32510 42030 32562
rect 42082 32510 42084 32562
rect 41020 32450 41076 32462
rect 41020 32398 41022 32450
rect 41074 32398 41076 32450
rect 39900 32004 39956 32014
rect 39900 31890 39956 31948
rect 41020 32004 41076 32398
rect 41020 31938 41076 31948
rect 42028 32228 42084 32510
rect 42364 32564 42420 32574
rect 42364 32470 42420 32508
rect 42588 32452 42644 33292
rect 42700 33346 43428 33348
rect 42700 33294 42702 33346
rect 42754 33294 43374 33346
rect 43426 33294 43428 33346
rect 42700 33292 43428 33294
rect 42700 33282 42756 33292
rect 43372 33282 43428 33292
rect 43484 33348 43540 33358
rect 43484 33254 43540 33292
rect 43260 33122 43316 33134
rect 43260 33070 43262 33122
rect 43314 33070 43316 33122
rect 42924 33012 42980 33022
rect 42700 32452 42756 32462
rect 42588 32450 42756 32452
rect 42588 32398 42702 32450
rect 42754 32398 42756 32450
rect 42588 32396 42756 32398
rect 42700 32386 42756 32396
rect 42812 32450 42868 32462
rect 42812 32398 42814 32450
rect 42866 32398 42868 32450
rect 42812 32228 42868 32398
rect 42924 32452 42980 32956
rect 43260 32788 43316 33070
rect 43596 32900 43652 34748
rect 43932 33572 43988 33582
rect 43932 33348 43988 33516
rect 43596 32834 43652 32844
rect 43708 33346 43988 33348
rect 43708 33294 43934 33346
rect 43986 33294 43988 33346
rect 43708 33292 43988 33294
rect 43260 32722 43316 32732
rect 43708 32786 43764 33292
rect 43932 33282 43988 33292
rect 44044 32788 44100 35644
rect 44268 35634 44324 35644
rect 44492 35810 44548 36990
rect 44492 35758 44494 35810
rect 44546 35758 44548 35810
rect 44268 34804 44324 34814
rect 44268 34710 44324 34748
rect 44268 34018 44324 34030
rect 44268 33966 44270 34018
rect 44322 33966 44324 34018
rect 44156 33796 44212 33806
rect 44156 33124 44212 33740
rect 44268 33348 44324 33966
rect 44268 33282 44324 33292
rect 44268 33124 44324 33134
rect 44156 33122 44324 33124
rect 44156 33070 44270 33122
rect 44322 33070 44324 33122
rect 44156 33068 44324 33070
rect 44268 33012 44324 33068
rect 44268 32946 44324 32956
rect 43708 32734 43710 32786
rect 43762 32734 43764 32786
rect 43708 32564 43764 32734
rect 43708 32498 43764 32508
rect 43820 32786 44100 32788
rect 43820 32734 44046 32786
rect 44098 32734 44100 32786
rect 43820 32732 44100 32734
rect 42924 32386 42980 32396
rect 42028 32172 42868 32228
rect 39900 31838 39902 31890
rect 39954 31838 39956 31890
rect 39900 31826 39956 31838
rect 42028 31890 42084 32172
rect 42028 31838 42030 31890
rect 42082 31838 42084 31890
rect 42028 31826 42084 31838
rect 43820 31780 43876 32732
rect 44044 32722 44100 32732
rect 44156 31892 44212 31902
rect 44156 31798 44212 31836
rect 38780 31778 39172 31780
rect 38780 31726 39118 31778
rect 39170 31726 39172 31778
rect 38780 31724 39172 31726
rect 37884 31220 37940 31230
rect 37548 31218 37940 31220
rect 37548 31166 37886 31218
rect 37938 31166 37940 31218
rect 37548 31164 37940 31166
rect 37884 31154 37940 31164
rect 37996 31106 38052 31118
rect 37996 31054 37998 31106
rect 38050 31054 38052 31106
rect 37548 30996 37604 31006
rect 37436 30994 37604 30996
rect 37436 30942 37550 30994
rect 37602 30942 37604 30994
rect 37436 30940 37604 30942
rect 37548 30930 37604 30940
rect 37996 30884 38052 31054
rect 37996 30818 38052 30828
rect 36988 30210 37156 30212
rect 36988 30158 36990 30210
rect 37042 30158 37156 30210
rect 36988 30156 37156 30158
rect 37212 30772 37268 30782
rect 37212 30210 37268 30716
rect 37772 30772 37828 30782
rect 37772 30678 37828 30716
rect 37212 30158 37214 30210
rect 37266 30158 37268 30210
rect 36988 29876 37044 30156
rect 37212 30146 37268 30158
rect 38780 30210 38836 31724
rect 39116 31714 39172 31724
rect 43260 31724 43820 31780
rect 42588 31668 42644 31678
rect 42924 31668 42980 31678
rect 42644 31666 42980 31668
rect 42644 31614 42926 31666
rect 42978 31614 42980 31666
rect 42644 31612 42980 31614
rect 42588 31574 42644 31612
rect 42924 31602 42980 31612
rect 43260 31666 43316 31724
rect 43820 31686 43876 31724
rect 43260 31614 43262 31666
rect 43314 31614 43316 31666
rect 43260 31602 43316 31614
rect 44492 31220 44548 35758
rect 44604 37044 44660 37054
rect 44604 35140 44660 36988
rect 44716 36148 44772 36158
rect 44716 35922 44772 36092
rect 44716 35870 44718 35922
rect 44770 35870 44772 35922
rect 44716 35858 44772 35870
rect 44828 35922 44884 37436
rect 44940 37266 44996 37278
rect 44940 37214 44942 37266
rect 44994 37214 44996 37266
rect 44940 36484 44996 37214
rect 44940 36418 44996 36428
rect 44940 36260 44996 36270
rect 44940 36166 44996 36204
rect 44828 35870 44830 35922
rect 44882 35870 44884 35922
rect 44828 35858 44884 35870
rect 44940 35700 44996 35710
rect 44940 35606 44996 35644
rect 44716 35252 44772 35262
rect 44772 35196 44884 35252
rect 44716 35186 44772 35196
rect 44604 35074 44660 35084
rect 44716 34356 44772 34366
rect 44716 34262 44772 34300
rect 44828 34132 44884 35196
rect 45052 34914 45108 37548
rect 45276 37380 45332 37390
rect 45276 37286 45332 37324
rect 45164 37154 45220 37166
rect 45164 37102 45166 37154
rect 45218 37102 45220 37154
rect 45164 35812 45220 37102
rect 45276 36372 45332 36382
rect 45276 36278 45332 36316
rect 45164 35746 45220 35756
rect 45388 35698 45444 38668
rect 45500 35924 45556 42140
rect 45724 41970 45780 41982
rect 45724 41918 45726 41970
rect 45778 41918 45780 41970
rect 45612 41076 45668 41086
rect 45612 40982 45668 41020
rect 45500 35858 45556 35868
rect 45612 36482 45668 36494
rect 45612 36430 45614 36482
rect 45666 36430 45668 36482
rect 45388 35646 45390 35698
rect 45442 35646 45444 35698
rect 45052 34862 45054 34914
rect 45106 34862 45108 34914
rect 45052 34850 45108 34862
rect 45276 35140 45332 35150
rect 45276 34802 45332 35084
rect 45388 35028 45444 35646
rect 45612 35588 45668 36430
rect 45724 36372 45780 41918
rect 45948 40628 46004 40638
rect 45948 40404 46004 40572
rect 45948 40310 46004 40348
rect 45836 38836 45892 38846
rect 45836 38742 45892 38780
rect 46060 38050 46116 43652
rect 46844 43586 46900 43596
rect 47180 43652 47236 43662
rect 46620 39506 46676 39518
rect 46620 39454 46622 39506
rect 46674 39454 46676 39506
rect 46508 38834 46564 38846
rect 46508 38782 46510 38834
rect 46562 38782 46564 38834
rect 46508 38724 46564 38782
rect 46508 38658 46564 38668
rect 46060 37998 46062 38050
rect 46114 37998 46116 38050
rect 46060 37986 46116 37998
rect 45724 36306 45780 36316
rect 45836 37266 45892 37278
rect 45836 37214 45838 37266
rect 45890 37214 45892 37266
rect 45612 35522 45668 35532
rect 45388 34962 45444 34972
rect 45276 34750 45278 34802
rect 45330 34750 45332 34802
rect 45276 34738 45332 34750
rect 45836 34804 45892 37214
rect 45836 34738 45892 34748
rect 45948 37156 46004 37166
rect 45948 34580 46004 37100
rect 46620 37044 46676 39454
rect 47180 39172 47236 43596
rect 47404 40516 47460 45164
rect 47404 40450 47460 40460
rect 47516 44994 47572 45006
rect 47516 44942 47518 44994
rect 47570 44942 47572 44994
rect 47180 39106 47236 39116
rect 47292 40404 47348 40414
rect 47292 40292 47348 40348
rect 47516 40292 47572 44942
rect 47628 43428 47684 45614
rect 47852 45666 47908 45678
rect 47852 45614 47854 45666
rect 47906 45614 47908 45666
rect 47740 44212 47796 44222
rect 47740 44118 47796 44156
rect 47852 43652 47908 45614
rect 47964 44772 48020 45836
rect 48076 45108 48132 45118
rect 48076 45106 48468 45108
rect 48076 45054 48078 45106
rect 48130 45054 48468 45106
rect 48076 45052 48468 45054
rect 48076 45042 48132 45052
rect 47964 44716 48356 44772
rect 47852 43586 47908 43596
rect 48076 44098 48132 44110
rect 48076 44046 48078 44098
rect 48130 44046 48132 44098
rect 47684 43372 47796 43428
rect 47628 43362 47684 43372
rect 47292 40236 47572 40292
rect 47628 41858 47684 41870
rect 47628 41806 47630 41858
rect 47682 41806 47684 41858
rect 46844 38834 46900 38846
rect 46844 38782 46846 38834
rect 46898 38782 46900 38834
rect 46844 37380 46900 38782
rect 47068 38836 47124 38846
rect 47068 38742 47124 38780
rect 47180 38834 47236 38846
rect 47180 38782 47182 38834
rect 47234 38782 47236 38834
rect 46844 37314 46900 37324
rect 47180 37156 47236 38782
rect 47292 38724 47348 40236
rect 47516 38948 47572 38958
rect 47516 38854 47572 38892
rect 47292 38668 47572 38724
rect 47180 37090 47236 37100
rect 47404 37938 47460 37950
rect 47404 37886 47406 37938
rect 47458 37886 47460 37938
rect 46620 36978 46676 36988
rect 47404 36372 47460 37886
rect 47404 36306 47460 36316
rect 47292 36036 47348 36046
rect 46060 35812 46116 35822
rect 46060 35718 46116 35756
rect 47180 35700 47236 35710
rect 45612 34524 46004 34580
rect 46956 35026 47012 35038
rect 46956 34974 46958 35026
rect 47010 34974 47012 35026
rect 44828 33572 44884 34076
rect 44940 34130 44996 34142
rect 44940 34078 44942 34130
rect 44994 34078 44996 34130
rect 44940 33796 44996 34078
rect 44940 33730 44996 33740
rect 45388 34130 45444 34142
rect 45388 34078 45390 34130
rect 45442 34078 45444 34130
rect 44940 33572 44996 33582
rect 44828 33570 44996 33572
rect 44828 33518 44942 33570
rect 44994 33518 44996 33570
rect 44828 33516 44996 33518
rect 44940 33506 44996 33516
rect 45388 33572 45444 34078
rect 45388 33506 45444 33516
rect 45500 33460 45556 33470
rect 44828 33348 44884 33358
rect 44828 33254 44884 33292
rect 45388 33346 45444 33358
rect 45388 33294 45390 33346
rect 45442 33294 45444 33346
rect 45388 33236 45444 33294
rect 45164 32564 45220 32574
rect 45164 32450 45220 32508
rect 45164 32398 45166 32450
rect 45218 32398 45220 32450
rect 45164 31892 45220 32398
rect 45164 31826 45220 31836
rect 44492 31154 44548 31164
rect 44716 31780 44772 31790
rect 44716 31218 44772 31724
rect 44716 31166 44718 31218
rect 44770 31166 44772 31218
rect 44716 31154 44772 31166
rect 45388 31778 45444 33180
rect 45500 32674 45556 33404
rect 45500 32622 45502 32674
rect 45554 32622 45556 32674
rect 45500 32610 45556 32622
rect 45612 32786 45668 34524
rect 45836 34356 45892 34366
rect 46956 34356 47012 34974
rect 45836 34354 46788 34356
rect 45836 34302 45838 34354
rect 45890 34302 46788 34354
rect 45836 34300 46788 34302
rect 45836 34290 45892 34300
rect 46284 34188 46564 34244
rect 45724 34130 45780 34142
rect 45724 34078 45726 34130
rect 45778 34078 45780 34130
rect 45724 33460 45780 34078
rect 45724 33394 45780 33404
rect 45948 34130 46004 34142
rect 45948 34078 45950 34130
rect 46002 34078 46004 34130
rect 45612 32734 45614 32786
rect 45666 32734 45668 32786
rect 45388 31726 45390 31778
rect 45442 31726 45444 31778
rect 45052 31108 45108 31118
rect 45052 31014 45108 31052
rect 42140 30324 42196 30334
rect 38780 30158 38782 30210
rect 38834 30158 38836 30210
rect 38780 30146 38836 30158
rect 41468 30322 42196 30324
rect 41468 30270 42142 30322
rect 42194 30270 42196 30322
rect 41468 30268 42196 30270
rect 37660 30098 37716 30110
rect 37660 30046 37662 30098
rect 37714 30046 37716 30098
rect 36988 29810 37044 29820
rect 37324 29986 37380 29998
rect 37324 29934 37326 29986
rect 37378 29934 37380 29986
rect 37324 29764 37380 29934
rect 37436 29988 37492 29998
rect 37436 29894 37492 29932
rect 37324 29698 37380 29708
rect 36764 29540 36820 29550
rect 36764 29426 36820 29484
rect 36764 29374 36766 29426
rect 36818 29374 36820 29426
rect 36764 29362 36820 29374
rect 37436 29540 37492 29550
rect 37100 29314 37156 29326
rect 37100 29262 37102 29314
rect 37154 29262 37156 29314
rect 36876 29202 36932 29214
rect 36876 29150 36878 29202
rect 36930 29150 36932 29202
rect 36876 27860 36932 29150
rect 37100 28642 37156 29262
rect 37100 28590 37102 28642
rect 37154 28590 37156 28642
rect 37100 28420 37156 28590
rect 37436 28868 37492 29484
rect 37436 28642 37492 28812
rect 37660 28756 37716 30046
rect 39452 30100 39508 30110
rect 39452 30006 39508 30044
rect 41132 30100 41188 30110
rect 37660 28690 37716 28700
rect 37884 29708 38500 29764
rect 37436 28590 37438 28642
rect 37490 28590 37492 28642
rect 37436 28578 37492 28590
rect 37100 28354 37156 28364
rect 37548 28084 37604 28094
rect 37884 28084 37940 29708
rect 38444 29652 38500 29708
rect 38556 29652 38612 29662
rect 38444 29650 38612 29652
rect 38444 29598 38558 29650
rect 38610 29598 38612 29650
rect 38444 29596 38612 29598
rect 38556 29586 38612 29596
rect 38332 29538 38388 29550
rect 38332 29486 38334 29538
rect 38386 29486 38388 29538
rect 38220 29428 38276 29438
rect 38220 29334 38276 29372
rect 38332 28980 38388 29486
rect 41132 29538 41188 30044
rect 41132 29486 41134 29538
rect 41186 29486 41188 29538
rect 41132 29474 41188 29486
rect 41356 29988 41412 29998
rect 38332 28868 38388 28924
rect 38108 28812 38388 28868
rect 38892 29426 38948 29438
rect 38892 29374 38894 29426
rect 38946 29374 38948 29426
rect 37996 28644 38052 28654
rect 37996 28550 38052 28588
rect 37548 28082 37940 28084
rect 37548 28030 37550 28082
rect 37602 28030 37940 28082
rect 37548 28028 37940 28030
rect 37548 28018 37604 28028
rect 37436 27972 37492 27982
rect 37436 27878 37492 27916
rect 37884 27970 37940 28028
rect 37996 28084 38052 28094
rect 38108 28084 38164 28812
rect 38892 28644 38948 29374
rect 40348 29314 40404 29326
rect 40348 29262 40350 29314
rect 40402 29262 40404 29314
rect 40348 29204 40404 29262
rect 41244 29204 41300 29214
rect 40348 29202 41300 29204
rect 40348 29150 41246 29202
rect 41298 29150 41300 29202
rect 40348 29148 41300 29150
rect 38668 28530 38724 28542
rect 38668 28478 38670 28530
rect 38722 28478 38724 28530
rect 37996 28082 38164 28084
rect 37996 28030 37998 28082
rect 38050 28030 38164 28082
rect 37996 28028 38164 28030
rect 38220 28084 38276 28094
rect 38668 28084 38724 28478
rect 38892 28532 38948 28588
rect 39564 28644 39620 28654
rect 39564 28642 39844 28644
rect 39564 28590 39566 28642
rect 39618 28590 39844 28642
rect 39564 28588 39844 28590
rect 39564 28578 39620 28588
rect 39004 28532 39060 28542
rect 38892 28530 39060 28532
rect 38892 28478 39006 28530
rect 39058 28478 39060 28530
rect 38892 28476 39060 28478
rect 39004 28466 39060 28476
rect 38220 28082 38724 28084
rect 38220 28030 38222 28082
rect 38274 28030 38724 28082
rect 38220 28028 38724 28030
rect 39452 28418 39508 28430
rect 39452 28366 39454 28418
rect 39506 28366 39508 28418
rect 37996 28018 38052 28028
rect 38220 28018 38276 28028
rect 37884 27918 37886 27970
rect 37938 27918 37940 27970
rect 37884 27906 37940 27918
rect 36876 27794 36932 27804
rect 38444 27860 38500 27870
rect 36876 27636 36932 27646
rect 36428 27074 36484 27086
rect 36428 27022 36430 27074
rect 36482 27022 36484 27074
rect 36428 26852 36484 27022
rect 36428 26786 36484 26796
rect 36876 26290 36932 27580
rect 36876 26238 36878 26290
rect 36930 26238 36932 26290
rect 36876 26226 36932 26238
rect 36988 26404 37044 26414
rect 36428 25618 36484 25630
rect 36428 25566 36430 25618
rect 36482 25566 36484 25618
rect 36428 25508 36484 25566
rect 36428 25442 36484 25452
rect 36988 25282 37044 26348
rect 38444 26290 38500 27804
rect 39116 27860 39172 27870
rect 39116 27858 39284 27860
rect 39116 27806 39118 27858
rect 39170 27806 39284 27858
rect 39116 27804 39284 27806
rect 39116 27794 39172 27804
rect 38668 27636 38724 27646
rect 38668 27542 38724 27580
rect 38444 26238 38446 26290
rect 38498 26238 38500 26290
rect 38444 26226 38500 26238
rect 38556 27074 38612 27086
rect 38556 27022 38558 27074
rect 38610 27022 38612 27074
rect 37324 25508 37380 25518
rect 37324 25414 37380 25452
rect 38108 25508 38164 25518
rect 38108 25414 38164 25452
rect 38444 25506 38500 25518
rect 38444 25454 38446 25506
rect 38498 25454 38500 25506
rect 36988 25230 36990 25282
rect 37042 25230 37044 25282
rect 36988 24836 37044 25230
rect 38220 25284 38276 25294
rect 38108 24948 38164 24958
rect 38108 24854 38164 24892
rect 38220 24946 38276 25228
rect 38220 24894 38222 24946
rect 38274 24894 38276 24946
rect 38220 24882 38276 24894
rect 37436 24836 37492 24846
rect 36988 24834 37492 24836
rect 36988 24782 37438 24834
rect 37490 24782 37492 24834
rect 36988 24780 37492 24782
rect 37436 24770 37492 24780
rect 37548 24834 37604 24846
rect 37548 24782 37550 24834
rect 37602 24782 37604 24834
rect 37548 24724 37604 24782
rect 37772 24836 37828 24846
rect 37772 24742 37828 24780
rect 37548 24658 37604 24668
rect 38444 24724 38500 25454
rect 38556 25396 38612 27022
rect 39116 26852 39172 26862
rect 39004 26292 39060 26302
rect 39004 26198 39060 26236
rect 39116 25618 39172 26796
rect 39228 26514 39284 27804
rect 39340 27858 39396 27870
rect 39340 27806 39342 27858
rect 39394 27806 39396 27858
rect 39340 26908 39396 27806
rect 39452 27748 39508 28366
rect 39564 27748 39620 27758
rect 39452 27746 39620 27748
rect 39452 27694 39566 27746
rect 39618 27694 39620 27746
rect 39452 27692 39620 27694
rect 39564 27076 39620 27692
rect 39788 27636 39844 28588
rect 40348 28084 40404 29148
rect 41244 29138 41300 29148
rect 41356 28980 41412 29932
rect 41468 29426 41524 30268
rect 42140 30258 42196 30268
rect 42252 30098 42308 30110
rect 42252 30046 42254 30098
rect 42306 30046 42308 30098
rect 41468 29374 41470 29426
rect 41522 29374 41524 29426
rect 41468 29362 41524 29374
rect 41692 29986 41748 29998
rect 41692 29934 41694 29986
rect 41746 29934 41748 29986
rect 41580 29204 41636 29214
rect 41580 29110 41636 29148
rect 41356 28924 41524 28980
rect 41468 28530 41524 28924
rect 41468 28478 41470 28530
rect 41522 28478 41524 28530
rect 41468 28466 41524 28478
rect 41692 28642 41748 29934
rect 42140 29988 42196 29998
rect 42252 29988 42308 30046
rect 42476 30100 42532 30110
rect 42476 30006 42532 30044
rect 44044 30100 44100 30110
rect 42196 29932 42308 29988
rect 42140 29922 42196 29932
rect 42252 29428 42308 29932
rect 44044 29652 44100 30044
rect 44156 29986 44212 29998
rect 44156 29934 44158 29986
rect 44210 29934 44212 29986
rect 44156 29764 44212 29934
rect 44156 29708 44772 29764
rect 42476 29596 43764 29652
rect 42476 29538 42532 29596
rect 42476 29486 42478 29538
rect 42530 29486 42532 29538
rect 42476 29474 42532 29486
rect 42252 29362 42308 29372
rect 42588 29426 42644 29438
rect 42588 29374 42590 29426
rect 42642 29374 42644 29426
rect 41692 28590 41694 28642
rect 41746 28590 41748 28642
rect 40348 28018 40404 28028
rect 40012 27972 40068 27982
rect 40012 27878 40068 27916
rect 40124 27972 40180 27982
rect 41356 27972 41412 27982
rect 40124 27970 40292 27972
rect 40124 27918 40126 27970
rect 40178 27918 40292 27970
rect 40124 27916 40292 27918
rect 40124 27906 40180 27916
rect 40124 27636 40180 27646
rect 39788 27634 40180 27636
rect 39788 27582 40126 27634
rect 40178 27582 40180 27634
rect 39788 27580 40180 27582
rect 40124 27570 40180 27580
rect 40236 27300 40292 27916
rect 41244 27970 41412 27972
rect 41244 27918 41358 27970
rect 41410 27918 41412 27970
rect 41244 27916 41412 27918
rect 41244 27412 41300 27916
rect 41356 27906 41412 27916
rect 41468 27860 41524 27870
rect 41468 27766 41524 27804
rect 41356 27636 41412 27646
rect 41356 27634 41636 27636
rect 41356 27582 41358 27634
rect 41410 27582 41636 27634
rect 41356 27580 41636 27582
rect 41356 27570 41412 27580
rect 41244 27356 41412 27412
rect 40124 27244 40292 27300
rect 39900 27076 39956 27086
rect 39564 27074 39956 27076
rect 39564 27022 39902 27074
rect 39954 27022 39956 27074
rect 39564 27020 39956 27022
rect 39900 27010 39956 27020
rect 40124 26908 40180 27244
rect 40908 27076 40964 27086
rect 39340 26852 39732 26908
rect 40124 26852 40292 26908
rect 39228 26462 39230 26514
rect 39282 26462 39284 26514
rect 39228 26450 39284 26462
rect 39116 25566 39118 25618
rect 39170 25566 39172 25618
rect 39116 25554 39172 25566
rect 39340 26290 39396 26302
rect 39564 26292 39620 26302
rect 39340 26238 39342 26290
rect 39394 26238 39396 26290
rect 39228 25508 39284 25518
rect 39228 25414 39284 25452
rect 38556 25330 38612 25340
rect 38780 25394 38836 25406
rect 38780 25342 38782 25394
rect 38834 25342 38836 25394
rect 38332 24498 38388 24510
rect 38332 24446 38334 24498
rect 38386 24446 38388 24498
rect 38108 23714 38164 23726
rect 38108 23662 38110 23714
rect 38162 23662 38164 23714
rect 38108 23156 38164 23662
rect 38332 23380 38388 24446
rect 38444 23604 38500 24668
rect 38668 25172 38724 25182
rect 38556 23604 38612 23614
rect 38444 23548 38556 23604
rect 38556 23538 38612 23548
rect 38332 23286 38388 23324
rect 38108 23090 38164 23100
rect 38220 23154 38276 23166
rect 38220 23102 38222 23154
rect 38274 23102 38276 23154
rect 37772 23042 37828 23054
rect 37772 22990 37774 23042
rect 37826 22990 37828 23042
rect 37772 22932 37828 22990
rect 38220 22932 38276 23102
rect 38444 23156 38500 23166
rect 38444 23154 38612 23156
rect 38444 23102 38446 23154
rect 38498 23102 38612 23154
rect 38444 23100 38612 23102
rect 38444 23090 38500 23100
rect 37772 22876 38276 22932
rect 36204 19842 36260 19852
rect 36876 22596 36932 22606
rect 36876 20916 36932 22540
rect 37996 22370 38052 22876
rect 37996 22318 37998 22370
rect 38050 22318 38052 22370
rect 37996 22306 38052 22318
rect 37772 22260 37828 22270
rect 37772 22166 37828 22204
rect 38444 22260 38500 22270
rect 38444 22166 38500 22204
rect 38556 22146 38612 23100
rect 38668 23154 38724 25116
rect 38780 24948 38836 25342
rect 38780 24722 38836 24892
rect 38892 25396 38948 25406
rect 38892 24946 38948 25340
rect 38892 24894 38894 24946
rect 38946 24894 38948 24946
rect 38892 24882 38948 24894
rect 39340 24836 39396 26238
rect 39340 24742 39396 24780
rect 39452 26290 39620 26292
rect 39452 26238 39566 26290
rect 39618 26238 39620 26290
rect 39452 26236 39620 26238
rect 39228 24724 39284 24734
rect 38780 24670 38782 24722
rect 38834 24670 38836 24722
rect 38780 24658 38836 24670
rect 39004 24722 39284 24724
rect 39004 24670 39230 24722
rect 39282 24670 39284 24722
rect 39004 24668 39284 24670
rect 38668 23102 38670 23154
rect 38722 23102 38724 23154
rect 38668 23090 38724 23102
rect 38780 23268 38836 23278
rect 38780 22370 38836 23212
rect 38892 22932 38948 22942
rect 38892 22838 38948 22876
rect 38780 22318 38782 22370
rect 38834 22318 38836 22370
rect 38780 22306 38836 22318
rect 38556 22094 38558 22146
rect 38610 22094 38612 22146
rect 38444 21588 38500 21598
rect 38220 21140 38276 21150
rect 36876 19906 36932 20860
rect 37660 20916 37716 20926
rect 37660 20822 37716 20860
rect 37772 20916 37828 20926
rect 37996 20916 38052 20926
rect 37772 20914 37996 20916
rect 37772 20862 37774 20914
rect 37826 20862 37996 20914
rect 37772 20860 37996 20862
rect 37772 20850 37828 20860
rect 37996 20850 38052 20860
rect 37100 20804 37156 20814
rect 37100 20710 37156 20748
rect 36988 20692 37044 20702
rect 36988 20598 37044 20636
rect 38108 20692 38164 20702
rect 38108 20598 38164 20636
rect 38220 20690 38276 21084
rect 38444 20802 38500 21532
rect 38444 20750 38446 20802
rect 38498 20750 38500 20802
rect 38444 20738 38500 20750
rect 38220 20638 38222 20690
rect 38274 20638 38276 20690
rect 38220 20626 38276 20638
rect 37660 20468 37716 20478
rect 37660 20130 37716 20412
rect 37660 20078 37662 20130
rect 37714 20078 37716 20130
rect 37660 20066 37716 20078
rect 37100 20020 37156 20030
rect 36876 19854 36878 19906
rect 36930 19854 36932 19906
rect 36876 19842 36932 19854
rect 36988 20018 37156 20020
rect 36988 19966 37102 20018
rect 37154 19966 37156 20018
rect 36988 19964 37156 19966
rect 36876 19348 36932 19358
rect 36876 18450 36932 19292
rect 36876 18398 36878 18450
rect 36930 18398 36932 18450
rect 36876 18386 36932 18398
rect 35868 17938 35924 17948
rect 36092 17780 36148 17790
rect 35420 17778 36148 17780
rect 35420 17726 36094 17778
rect 36146 17726 36148 17778
rect 35420 17724 36148 17726
rect 34412 17614 34414 17666
rect 34466 17614 34468 17666
rect 34412 17602 34468 17614
rect 34748 17666 34804 17678
rect 34748 17614 34750 17666
rect 34802 17614 34804 17666
rect 34300 17444 34356 17454
rect 34076 17442 34356 17444
rect 34076 17390 34302 17442
rect 34354 17390 34356 17442
rect 34076 17388 34356 17390
rect 34076 16884 34132 17388
rect 34300 17378 34356 17388
rect 33852 16830 33854 16882
rect 33906 16830 33908 16882
rect 33852 16818 33908 16830
rect 33964 16882 34132 16884
rect 33964 16830 34078 16882
rect 34130 16830 34132 16882
rect 33964 16828 34132 16830
rect 32956 16046 32958 16098
rect 33010 16046 33012 16098
rect 32956 16034 33012 16046
rect 33292 15988 33348 15998
rect 33292 15538 33348 15932
rect 33964 15652 34020 16828
rect 34076 16818 34132 16828
rect 34300 16884 34356 16894
rect 34300 16210 34356 16828
rect 34636 16884 34692 16894
rect 34636 16790 34692 16828
rect 34300 16158 34302 16210
rect 34354 16158 34356 16210
rect 34300 16146 34356 16158
rect 33740 15596 34020 15652
rect 33292 15486 33294 15538
rect 33346 15486 33348 15538
rect 33292 15474 33348 15486
rect 33404 15540 33460 15550
rect 33404 15446 33460 15484
rect 32172 15428 32228 15438
rect 32172 15334 32228 15372
rect 31836 15262 31838 15314
rect 31890 15262 31892 15314
rect 31836 15148 31892 15262
rect 32396 15316 32452 15326
rect 32396 15222 32452 15260
rect 33180 15314 33236 15326
rect 33180 15262 33182 15314
rect 33234 15262 33236 15314
rect 31836 15092 32228 15148
rect 31500 14478 31502 14530
rect 31554 14478 31556 14530
rect 31500 14466 31556 14478
rect 32172 14642 32228 15092
rect 32172 14590 32174 14642
rect 32226 14590 32228 14642
rect 31724 14418 31780 14430
rect 31724 14366 31726 14418
rect 31778 14366 31780 14418
rect 31388 14308 31444 14318
rect 30940 14306 31444 14308
rect 30940 14254 31390 14306
rect 31442 14254 31444 14306
rect 30940 14252 31444 14254
rect 31388 14242 31444 14252
rect 31052 13860 31108 13870
rect 31052 13766 31108 13804
rect 31500 13748 31556 13758
rect 31500 13654 31556 13692
rect 31612 13746 31668 13758
rect 31612 13694 31614 13746
rect 31666 13694 31668 13746
rect 31388 13188 31444 13198
rect 31052 12964 31108 12974
rect 30492 12290 30548 12302
rect 30492 12238 30494 12290
rect 30546 12238 30548 12290
rect 30156 12066 30212 12078
rect 30156 12014 30158 12066
rect 30210 12014 30212 12066
rect 30156 11732 30212 12014
rect 30492 11956 30548 12238
rect 31052 12180 31108 12908
rect 31388 12404 31444 13132
rect 31612 13188 31668 13694
rect 31612 13122 31668 13132
rect 31388 12310 31444 12348
rect 31276 12292 31332 12302
rect 31276 12198 31332 12236
rect 30492 11890 30548 11900
rect 30940 12178 31108 12180
rect 30940 12126 31054 12178
rect 31106 12126 31108 12178
rect 30940 12124 31108 12126
rect 30156 11676 30548 11732
rect 29820 11564 30100 11620
rect 30492 11618 30548 11676
rect 30492 11566 30494 11618
rect 30546 11566 30548 11618
rect 29708 11396 29764 11406
rect 29484 11342 29486 11394
rect 29538 11342 29540 11394
rect 27916 11284 27972 11294
rect 29484 11284 29540 11342
rect 27916 11282 28084 11284
rect 27916 11230 27918 11282
rect 27970 11230 28084 11282
rect 27916 11228 28084 11230
rect 27916 11218 27972 11228
rect 27804 10610 27860 10668
rect 27804 10558 27806 10610
rect 27858 10558 27860 10610
rect 26908 7522 26964 7532
rect 26180 7196 26292 7252
rect 27244 7476 27300 7486
rect 25788 6804 25844 6814
rect 25676 6802 25844 6804
rect 25676 6750 25790 6802
rect 25842 6750 25844 6802
rect 25676 6748 25844 6750
rect 25788 6738 25844 6748
rect 26124 6690 26180 7196
rect 26236 6804 26292 6814
rect 26236 6710 26292 6748
rect 26124 6638 26126 6690
rect 26178 6638 26180 6690
rect 26124 6626 26180 6638
rect 26796 6692 26852 6702
rect 26796 6598 26852 6636
rect 24108 5404 24612 5460
rect 23660 5234 23716 5246
rect 23660 5182 23662 5234
rect 23714 5182 23716 5234
rect 23324 5068 23492 5124
rect 22316 5012 22372 5022
rect 22204 4900 22260 4910
rect 22316 4900 22372 4956
rect 22204 4898 22372 4900
rect 22204 4846 22206 4898
rect 22258 4846 22372 4898
rect 22204 4844 22372 4846
rect 22428 4900 22484 4910
rect 22204 4834 22260 4844
rect 22428 4806 22484 4844
rect 23324 4898 23380 4910
rect 23324 4846 23326 4898
rect 23378 4846 23380 4898
rect 21420 4338 21588 4340
rect 21420 4286 21422 4338
rect 21474 4286 21588 4338
rect 21420 4284 21588 4286
rect 21420 4274 21476 4284
rect 22092 4228 22148 4238
rect 22092 4134 22148 4172
rect 21868 3668 21924 3678
rect 21868 3574 21924 3612
rect 20188 3332 21252 3388
rect 21532 3556 21588 3566
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 21532 800 21588 3500
rect 23324 3388 23380 4846
rect 23436 4564 23492 5068
rect 23660 4900 23716 5182
rect 24108 5122 24164 5404
rect 24108 5070 24110 5122
rect 24162 5070 24164 5122
rect 24108 5058 24164 5070
rect 23660 4834 23716 4844
rect 23436 4508 23716 4564
rect 23660 3442 23716 4508
rect 24220 4226 24276 5404
rect 24220 4174 24222 4226
rect 24274 4174 24276 4226
rect 24220 4162 24276 4174
rect 24332 5236 24388 5246
rect 23660 3390 23662 3442
rect 23714 3390 23716 3442
rect 23324 3332 23604 3388
rect 23660 3378 23716 3390
rect 23884 3554 23940 3566
rect 23884 3502 23886 3554
rect 23938 3502 23940 3554
rect 23548 2772 23604 3332
rect 23884 2772 23940 3502
rect 23548 2716 23940 2772
rect 23548 800 23604 2716
rect 24332 2436 24388 5180
rect 24556 5122 24612 5404
rect 24556 5070 24558 5122
rect 24610 5070 24612 5122
rect 24556 5058 24612 5070
rect 24780 5852 25060 5908
rect 26348 6466 26404 6478
rect 26348 6414 26350 6466
rect 26402 6414 26404 6466
rect 26348 6244 26404 6414
rect 27244 6468 27300 7420
rect 27580 7364 27636 7374
rect 27804 7364 27860 10558
rect 27916 10612 27972 10622
rect 27916 9826 27972 10556
rect 27916 9774 27918 9826
rect 27970 9774 27972 9826
rect 27916 9762 27972 9774
rect 27916 9044 27972 9054
rect 28028 9044 28084 11228
rect 29484 11218 29540 11228
rect 29596 11394 29764 11396
rect 29596 11342 29710 11394
rect 29762 11342 29764 11394
rect 29596 11340 29764 11342
rect 29596 10948 29652 11340
rect 29708 11330 29764 11340
rect 29148 10892 29652 10948
rect 29148 10834 29204 10892
rect 29148 10782 29150 10834
rect 29202 10782 29204 10834
rect 29148 10770 29204 10782
rect 28924 10724 28980 10734
rect 28924 10630 28980 10668
rect 28364 10612 28420 10622
rect 28812 10612 28868 10622
rect 28420 10610 28868 10612
rect 28420 10558 28814 10610
rect 28866 10558 28868 10610
rect 28420 10556 28868 10558
rect 28364 10518 28420 10556
rect 28252 9940 28308 9950
rect 28252 9846 28308 9884
rect 28364 9716 28420 9726
rect 28364 9622 28420 9660
rect 28252 9380 28308 9390
rect 28252 9266 28308 9324
rect 28252 9214 28254 9266
rect 28306 9214 28308 9266
rect 28252 9202 28308 9214
rect 28476 9044 28532 10556
rect 28812 10546 28868 10556
rect 27972 8988 28084 9044
rect 28252 9042 28532 9044
rect 28252 8990 28478 9042
rect 28530 8990 28532 9042
rect 28252 8988 28532 8990
rect 27916 8978 27972 8988
rect 28252 8708 28308 8988
rect 28476 8978 28532 8988
rect 28700 10164 28756 10174
rect 28700 9154 28756 10108
rect 29596 9828 29652 9838
rect 29596 9734 29652 9772
rect 29484 9268 29540 9278
rect 29820 9268 29876 11564
rect 30492 11554 30548 11566
rect 30044 11396 30100 11406
rect 30044 11302 30100 11340
rect 30716 11396 30772 11406
rect 30940 11396 30996 12124
rect 31052 12114 31108 12124
rect 31724 11956 31780 14366
rect 31836 13972 31892 13982
rect 31836 13746 31892 13916
rect 31836 13694 31838 13746
rect 31890 13694 31892 13746
rect 31836 13682 31892 13694
rect 32060 13188 32116 13198
rect 32060 13074 32116 13132
rect 32060 13022 32062 13074
rect 32114 13022 32116 13074
rect 32060 13010 32116 13022
rect 31948 12852 32004 12862
rect 31948 12758 32004 12796
rect 31724 11890 31780 11900
rect 31836 12292 31892 12302
rect 30716 11302 30772 11340
rect 30828 11394 30996 11396
rect 30828 11342 30942 11394
rect 30994 11342 30996 11394
rect 30828 11340 30996 11342
rect 30716 10836 30772 10846
rect 30828 10836 30884 11340
rect 30940 11330 30996 11340
rect 31052 11396 31108 11406
rect 31052 11302 31108 11340
rect 31724 11396 31780 11406
rect 31724 11302 31780 11340
rect 30716 10834 30884 10836
rect 30716 10782 30718 10834
rect 30770 10782 30884 10834
rect 30716 10780 30884 10782
rect 31164 11170 31220 11182
rect 31164 11118 31166 11170
rect 31218 11118 31220 11170
rect 30716 10770 30772 10780
rect 31164 10724 31220 11118
rect 31836 10836 31892 12236
rect 32060 10836 32116 10846
rect 31164 10658 31220 10668
rect 31612 10834 32116 10836
rect 31612 10782 32062 10834
rect 32114 10782 32116 10834
rect 31612 10780 32116 10782
rect 29932 10612 29988 10622
rect 29932 9938 29988 10556
rect 30716 10610 30772 10622
rect 30716 10558 30718 10610
rect 30770 10558 30772 10610
rect 30716 10164 30772 10558
rect 30716 10098 30772 10108
rect 29932 9886 29934 9938
rect 29986 9886 29988 9938
rect 29932 9874 29988 9886
rect 30940 9828 30996 9838
rect 30940 9734 30996 9772
rect 30268 9716 30324 9726
rect 29484 9266 29876 9268
rect 29484 9214 29486 9266
rect 29538 9214 29876 9266
rect 29484 9212 29876 9214
rect 29484 9202 29540 9212
rect 28700 9102 28702 9154
rect 28754 9102 28756 9154
rect 27916 8652 28308 8708
rect 27916 8370 27972 8652
rect 27916 8318 27918 8370
rect 27970 8318 27972 8370
rect 27916 8306 27972 8318
rect 28028 8484 28084 8494
rect 28028 7474 28084 8428
rect 28476 7588 28532 7598
rect 28476 7494 28532 7532
rect 28700 7476 28756 9102
rect 29820 9042 29876 9212
rect 30156 9714 30324 9716
rect 30156 9662 30270 9714
rect 30322 9662 30324 9714
rect 30156 9660 30324 9662
rect 30156 9154 30212 9660
rect 30268 9650 30324 9660
rect 31052 9716 31108 9726
rect 31052 9714 31556 9716
rect 31052 9662 31054 9714
rect 31106 9662 31556 9714
rect 31052 9660 31556 9662
rect 31052 9650 31108 9660
rect 31500 9380 31556 9660
rect 31612 9602 31668 10780
rect 32060 10770 32116 10780
rect 31612 9550 31614 9602
rect 31666 9550 31668 9602
rect 31612 9538 31668 9550
rect 31836 9826 31892 9838
rect 31836 9774 31838 9826
rect 31890 9774 31892 9826
rect 31836 9380 31892 9774
rect 31500 9324 31892 9380
rect 30156 9102 30158 9154
rect 30210 9102 30212 9154
rect 30156 9090 30212 9102
rect 29820 8990 29822 9042
rect 29874 8990 29876 9042
rect 29148 8260 29204 8270
rect 28028 7422 28030 7474
rect 28082 7422 28084 7474
rect 27580 7362 27972 7364
rect 27580 7310 27582 7362
rect 27634 7310 27972 7362
rect 27580 7308 27972 7310
rect 27580 7298 27636 7308
rect 27356 6692 27412 6702
rect 27916 6692 27972 7308
rect 28028 7028 28084 7422
rect 28588 7474 28756 7476
rect 28588 7422 28702 7474
rect 28754 7422 28756 7474
rect 28588 7420 28756 7422
rect 28028 6972 28420 7028
rect 28028 6692 28084 6702
rect 27916 6690 28084 6692
rect 27916 6638 28030 6690
rect 28082 6638 28084 6690
rect 27916 6636 28084 6638
rect 27356 6598 27412 6636
rect 28028 6626 28084 6636
rect 27804 6468 27860 6478
rect 27244 6412 27412 6468
rect 24780 4900 24836 5852
rect 25228 5796 25284 5806
rect 24780 4834 24836 4844
rect 24892 5794 25284 5796
rect 24892 5742 25230 5794
rect 25282 5742 25284 5794
rect 24892 5740 25284 5742
rect 24668 3554 24724 3566
rect 24668 3502 24670 3554
rect 24722 3502 24724 3554
rect 24668 3444 24724 3502
rect 24668 3378 24724 3388
rect 24892 3442 24948 5740
rect 25228 5730 25284 5740
rect 25900 5794 25956 5806
rect 25900 5742 25902 5794
rect 25954 5742 25956 5794
rect 25340 5684 25396 5694
rect 25340 5590 25396 5628
rect 25452 5236 25508 5246
rect 25452 5142 25508 5180
rect 25452 4226 25508 4238
rect 25452 4174 25454 4226
rect 25506 4174 25508 4226
rect 25452 3556 25508 4174
rect 25452 3490 25508 3500
rect 25564 3666 25620 3678
rect 25564 3614 25566 3666
rect 25618 3614 25620 3666
rect 24892 3390 24894 3442
rect 24946 3390 24948 3442
rect 24892 3378 24948 3390
rect 24220 2380 24388 2436
rect 24220 800 24276 2380
rect 25564 800 25620 3614
rect 25900 3444 25956 5742
rect 26348 5012 26404 6188
rect 26572 6020 26628 6030
rect 26572 5906 26628 5964
rect 26572 5854 26574 5906
rect 26626 5854 26628 5906
rect 26572 5842 26628 5854
rect 26796 6018 26852 6030
rect 26796 5966 26798 6018
rect 26850 5966 26852 6018
rect 26796 5124 26852 5966
rect 27132 6020 27188 6030
rect 27132 5926 27188 5964
rect 26796 5058 26852 5068
rect 27244 5684 27300 5694
rect 27244 5122 27300 5628
rect 27244 5070 27246 5122
rect 27298 5070 27300 5122
rect 27244 5058 27300 5070
rect 26348 4946 26404 4956
rect 26908 5012 26964 5022
rect 25900 3332 26292 3388
rect 26236 800 26292 3332
rect 26908 800 26964 4956
rect 27356 3554 27412 6412
rect 27804 6374 27860 6412
rect 27916 6466 27972 6478
rect 27916 6414 27918 6466
rect 27970 6414 27972 6466
rect 27468 5908 27524 5918
rect 27804 5908 27860 5918
rect 27468 5906 27860 5908
rect 27468 5854 27470 5906
rect 27522 5854 27806 5906
rect 27858 5854 27860 5906
rect 27468 5852 27860 5854
rect 27468 5842 27524 5852
rect 27692 5124 27748 5134
rect 27692 5030 27748 5068
rect 27580 4898 27636 4910
rect 27580 4846 27582 4898
rect 27634 4846 27636 4898
rect 27580 4450 27636 4846
rect 27804 4900 27860 5852
rect 27916 5122 27972 6414
rect 28140 6468 28196 6478
rect 28140 6130 28196 6412
rect 28140 6078 28142 6130
rect 28194 6078 28196 6130
rect 28140 6066 28196 6078
rect 27916 5070 27918 5122
rect 27970 5070 27972 5122
rect 27916 5058 27972 5070
rect 28252 4900 28308 4910
rect 27804 4898 28308 4900
rect 27804 4846 28254 4898
rect 28306 4846 28308 4898
rect 27804 4844 28308 4846
rect 28252 4834 28308 4844
rect 28364 4676 28420 6972
rect 28476 6466 28532 6478
rect 28476 6414 28478 6466
rect 28530 6414 28532 6466
rect 28476 5122 28532 6414
rect 28476 5070 28478 5122
rect 28530 5070 28532 5122
rect 28476 5012 28532 5070
rect 28476 4946 28532 4956
rect 28588 4900 28644 7420
rect 28700 7410 28756 7420
rect 29036 8258 29204 8260
rect 29036 8206 29150 8258
rect 29202 8206 29204 8258
rect 29036 8204 29204 8206
rect 29036 6132 29092 8204
rect 29148 8194 29204 8204
rect 29820 7700 29876 8990
rect 29932 8930 29988 8942
rect 29932 8878 29934 8930
rect 29986 8878 29988 8930
rect 29932 8370 29988 8878
rect 29932 8318 29934 8370
rect 29986 8318 29988 8370
rect 29932 8306 29988 8318
rect 31836 8372 31892 9324
rect 32172 8484 32228 14590
rect 33180 14530 33236 15262
rect 33180 14478 33182 14530
rect 33234 14478 33236 14530
rect 33180 14466 33236 14478
rect 32844 14418 32900 14430
rect 32844 14366 32846 14418
rect 32898 14366 32900 14418
rect 32844 14084 32900 14366
rect 32956 14420 33012 14430
rect 32956 14326 33012 14364
rect 32844 14018 32900 14028
rect 32396 13972 32452 13982
rect 32396 13878 32452 13916
rect 32284 13076 32340 13086
rect 32284 12962 32340 13020
rect 32732 13076 32788 13086
rect 33516 13076 33572 13086
rect 32788 13020 32900 13076
rect 32732 13010 32788 13020
rect 32284 12910 32286 12962
rect 32338 12910 32340 12962
rect 32284 12898 32340 12910
rect 32508 12852 32564 12862
rect 32508 12850 32676 12852
rect 32508 12798 32510 12850
rect 32562 12798 32676 12850
rect 32508 12796 32676 12798
rect 32508 12786 32564 12796
rect 32284 12290 32340 12302
rect 32284 12238 32286 12290
rect 32338 12238 32340 12290
rect 32284 11956 32340 12238
rect 32508 12180 32564 12190
rect 32508 12086 32564 12124
rect 32284 11890 32340 11900
rect 32620 11284 32676 12796
rect 32732 12404 32788 12414
rect 32732 11394 32788 12348
rect 32732 11342 32734 11394
rect 32786 11342 32788 11394
rect 32732 11330 32788 11342
rect 32620 11218 32676 11228
rect 32396 10724 32452 10734
rect 32284 9714 32340 9726
rect 32284 9662 32286 9714
rect 32338 9662 32340 9714
rect 32284 9604 32340 9662
rect 32396 9714 32452 10668
rect 32844 10388 32900 13020
rect 33572 13020 33684 13076
rect 33516 13010 33572 13020
rect 33180 12852 33236 12862
rect 33236 12796 33460 12852
rect 33180 12786 33236 12796
rect 33180 11284 33236 11294
rect 33404 11284 33460 12796
rect 33516 12404 33572 12414
rect 33516 11506 33572 12348
rect 33516 11454 33518 11506
rect 33570 11454 33572 11506
rect 33516 11442 33572 11454
rect 33628 11394 33684 13020
rect 33740 12180 33796 15596
rect 34188 15540 34244 15550
rect 33964 15538 34244 15540
rect 33964 15486 34190 15538
rect 34242 15486 34244 15538
rect 33964 15484 34244 15486
rect 33852 15316 33908 15326
rect 33964 15316 34020 15484
rect 34188 15474 34244 15484
rect 33852 15314 34020 15316
rect 33852 15262 33854 15314
rect 33906 15262 34020 15314
rect 33852 15260 34020 15262
rect 34076 15314 34132 15326
rect 34076 15262 34078 15314
rect 34130 15262 34132 15314
rect 33852 15250 33908 15260
rect 34076 14308 34132 15262
rect 34412 15314 34468 15326
rect 34412 15262 34414 15314
rect 34466 15262 34468 15314
rect 34412 14420 34468 15262
rect 34636 15314 34692 15326
rect 34636 15262 34638 15314
rect 34690 15262 34692 15314
rect 34636 14644 34692 15262
rect 34636 14578 34692 14588
rect 34748 14532 34804 17614
rect 35420 16994 35476 17724
rect 36092 17714 36148 17724
rect 36204 17780 36260 17790
rect 35420 16942 35422 16994
rect 35474 16942 35476 16994
rect 35420 16930 35476 16942
rect 35756 17556 35812 17566
rect 36204 17556 36260 17724
rect 35756 17554 36260 17556
rect 35756 17502 35758 17554
rect 35810 17502 36206 17554
rect 36258 17502 36260 17554
rect 35756 17500 36260 17502
rect 35756 16660 35812 17500
rect 36204 17490 36260 17500
rect 36428 17554 36484 17566
rect 36428 17502 36430 17554
rect 36482 17502 36484 17554
rect 35756 16594 35812 16604
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35980 16324 36036 16334
rect 35980 16098 36036 16268
rect 36428 16210 36484 17502
rect 36428 16158 36430 16210
rect 36482 16158 36484 16210
rect 36428 16146 36484 16158
rect 35980 16046 35982 16098
rect 36034 16046 36036 16098
rect 35980 16034 36036 16046
rect 36316 16098 36372 16110
rect 36316 16046 36318 16098
rect 36370 16046 36372 16098
rect 36204 15876 36260 15886
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35644 14644 35700 14654
rect 35644 14550 35700 14588
rect 34748 14466 34804 14476
rect 35196 14530 35252 14542
rect 35420 14532 35476 14542
rect 35196 14478 35198 14530
rect 35250 14478 35252 14530
rect 34412 14326 34468 14364
rect 34860 14418 34916 14430
rect 34860 14366 34862 14418
rect 34914 14366 34916 14418
rect 34076 14242 34132 14252
rect 34300 14196 34356 14206
rect 33852 13748 33908 13758
rect 33852 13746 34020 13748
rect 33852 13694 33854 13746
rect 33906 13694 34020 13746
rect 33852 13692 34020 13694
rect 33852 13682 33908 13692
rect 33964 12292 34020 13692
rect 33740 12124 33908 12180
rect 33628 11342 33630 11394
rect 33682 11342 33684 11394
rect 33628 11330 33684 11342
rect 33740 11956 33796 11966
rect 33516 11284 33572 11294
rect 33180 11190 33236 11228
rect 33292 11282 33572 11284
rect 33292 11230 33518 11282
rect 33570 11230 33572 11282
rect 33292 11228 33572 11230
rect 32732 10332 32900 10388
rect 33068 10724 33124 10734
rect 32396 9662 32398 9714
rect 32450 9662 32452 9714
rect 32396 9650 32452 9662
rect 32620 9716 32676 9726
rect 32620 9622 32676 9660
rect 32284 9538 32340 9548
rect 32172 8428 32564 8484
rect 32060 8372 32116 8382
rect 31836 8370 32116 8372
rect 31836 8318 32062 8370
rect 32114 8318 32116 8370
rect 31836 8316 32116 8318
rect 32060 8306 32116 8316
rect 29820 7634 29876 7644
rect 29148 7588 29204 7598
rect 29148 6690 29204 7532
rect 32060 6804 32116 6814
rect 32172 6804 32228 8428
rect 32508 8370 32564 8428
rect 32508 8318 32510 8370
rect 32562 8318 32564 8370
rect 32508 8306 32564 8318
rect 32060 6802 32228 6804
rect 32060 6750 32062 6802
rect 32114 6750 32228 6802
rect 32060 6748 32228 6750
rect 32060 6738 32116 6748
rect 29148 6638 29150 6690
rect 29202 6638 29204 6690
rect 29148 6626 29204 6638
rect 29260 6692 29316 6702
rect 29596 6692 29652 6702
rect 29260 6690 29540 6692
rect 29260 6638 29262 6690
rect 29314 6638 29540 6690
rect 29260 6636 29540 6638
rect 29260 6626 29316 6636
rect 29372 6468 29428 6478
rect 29372 6374 29428 6412
rect 29260 6132 29316 6142
rect 29036 6076 29260 6132
rect 28588 4834 28644 4844
rect 28700 5794 28756 5806
rect 28700 5742 28702 5794
rect 28754 5742 28756 5794
rect 27580 4398 27582 4450
rect 27634 4398 27636 4450
rect 27580 4386 27636 4398
rect 28140 4620 28420 4676
rect 27356 3502 27358 3554
rect 27410 3502 27412 3554
rect 27356 3490 27412 3502
rect 27580 3668 27636 3678
rect 27580 800 27636 3612
rect 28140 3556 28196 4620
rect 28700 4564 28756 5742
rect 28812 5684 28868 5694
rect 28812 5682 29092 5684
rect 28812 5630 28814 5682
rect 28866 5630 29092 5682
rect 28812 5628 29092 5630
rect 28812 5618 28868 5628
rect 29036 5122 29092 5628
rect 29036 5070 29038 5122
rect 29090 5070 29092 5122
rect 29036 5058 29092 5070
rect 29148 4900 29204 6076
rect 29260 6038 29316 6076
rect 29372 5684 29428 5694
rect 29372 5124 29428 5628
rect 29484 5460 29540 6636
rect 29596 6578 29652 6636
rect 29596 6526 29598 6578
rect 29650 6526 29652 6578
rect 29596 6514 29652 6526
rect 30156 6692 30212 6702
rect 30156 6578 30212 6636
rect 30716 6692 30772 6702
rect 30716 6598 30772 6636
rect 31388 6692 31444 6702
rect 31388 6598 31444 6636
rect 30156 6526 30158 6578
rect 30210 6526 30212 6578
rect 30156 6514 30212 6526
rect 30492 6466 30548 6478
rect 30492 6414 30494 6466
rect 30546 6414 30548 6466
rect 29932 6020 29988 6030
rect 29932 5926 29988 5964
rect 30492 6020 30548 6414
rect 31164 6468 31220 6478
rect 31164 6374 31220 6412
rect 31276 6466 31332 6478
rect 31276 6414 31278 6466
rect 31330 6414 31332 6466
rect 30492 5954 30548 5964
rect 30604 6300 30884 6356
rect 30604 5460 30660 6300
rect 29484 5404 29652 5460
rect 29372 5058 29428 5068
rect 29596 5122 29652 5404
rect 30268 5404 30660 5460
rect 30716 6132 30772 6142
rect 30268 5346 30324 5404
rect 30268 5294 30270 5346
rect 30322 5294 30324 5346
rect 30268 5282 30324 5294
rect 29596 5070 29598 5122
rect 29650 5070 29652 5122
rect 29596 5058 29652 5070
rect 30716 5122 30772 6076
rect 30828 5906 30884 6300
rect 30828 5854 30830 5906
rect 30882 5854 30884 5906
rect 30828 5842 30884 5854
rect 31164 6130 31220 6142
rect 31164 6078 31166 6130
rect 31218 6078 31220 6130
rect 31164 5236 31220 6078
rect 31276 6132 31332 6414
rect 32172 6132 32228 6748
rect 31276 6076 31444 6132
rect 31276 5906 31332 5918
rect 31276 5854 31278 5906
rect 31330 5854 31332 5906
rect 31276 5684 31332 5854
rect 31388 5906 31444 6076
rect 32172 6066 32228 6076
rect 32508 7364 32564 7374
rect 32508 6020 32564 7308
rect 32732 6692 32788 10332
rect 33068 9826 33124 10668
rect 33068 9774 33070 9826
rect 33122 9774 33124 9826
rect 33068 9762 33124 9774
rect 33292 9828 33348 11228
rect 33516 11218 33572 11228
rect 33740 11060 33796 11900
rect 32956 9714 33012 9726
rect 32956 9662 32958 9714
rect 33010 9662 33012 9714
rect 32844 9380 32900 9390
rect 32844 8370 32900 9324
rect 32956 9268 33012 9662
rect 33180 9714 33236 9726
rect 33180 9662 33182 9714
rect 33234 9662 33236 9714
rect 33180 9604 33236 9662
rect 33180 9538 33236 9548
rect 33180 9268 33236 9278
rect 32956 9212 33180 9268
rect 33180 9154 33236 9212
rect 33180 9102 33182 9154
rect 33234 9102 33236 9154
rect 33180 9090 33236 9102
rect 33068 8932 33124 8942
rect 33292 8932 33348 9772
rect 33068 8930 33348 8932
rect 33068 8878 33070 8930
rect 33122 8878 33348 8930
rect 33068 8876 33348 8878
rect 33516 11004 33796 11060
rect 33068 8866 33124 8876
rect 32844 8318 32846 8370
rect 32898 8318 32900 8370
rect 32844 8306 32900 8318
rect 33404 7700 33460 7710
rect 33516 7700 33572 11004
rect 33852 10164 33908 12124
rect 33964 12178 34020 12236
rect 33964 12126 33966 12178
rect 34018 12126 34020 12178
rect 33964 12114 34020 12126
rect 34076 13746 34132 13758
rect 34076 13694 34078 13746
rect 34130 13694 34132 13746
rect 34076 11956 34132 13694
rect 34300 13746 34356 14140
rect 34636 13972 34692 13982
rect 34860 13972 34916 14366
rect 34972 14420 35028 14430
rect 35196 14420 35252 14478
rect 34972 14418 35140 14420
rect 34972 14366 34974 14418
rect 35026 14366 35140 14418
rect 34972 14364 35140 14366
rect 34972 14354 35028 14364
rect 34636 13970 34916 13972
rect 34636 13918 34638 13970
rect 34690 13918 34916 13970
rect 34636 13916 34916 13918
rect 34636 13906 34692 13916
rect 35084 13858 35140 14364
rect 35196 14354 35252 14364
rect 35308 14530 35476 14532
rect 35308 14478 35422 14530
rect 35474 14478 35476 14530
rect 35308 14476 35476 14478
rect 35308 13970 35364 14476
rect 35420 14466 35476 14476
rect 35532 14532 35588 14542
rect 35308 13918 35310 13970
rect 35362 13918 35364 13970
rect 35308 13906 35364 13918
rect 35084 13806 35086 13858
rect 35138 13806 35140 13858
rect 34300 13694 34302 13746
rect 34354 13694 34356 13746
rect 34300 13682 34356 13694
rect 34412 13748 34468 13758
rect 34972 13748 35028 13758
rect 34412 13746 35028 13748
rect 34412 13694 34414 13746
rect 34466 13694 34974 13746
rect 35026 13694 35028 13746
rect 34412 13692 35028 13694
rect 34412 13188 34468 13692
rect 34972 13682 35028 13692
rect 34300 13132 34468 13188
rect 34300 12402 34356 13132
rect 34300 12350 34302 12402
rect 34354 12350 34356 12402
rect 34300 12338 34356 12350
rect 34076 11890 34132 11900
rect 34188 12292 34244 12302
rect 34188 11620 34244 12236
rect 34860 12292 34916 12302
rect 34860 12198 34916 12236
rect 34412 12180 34468 12190
rect 34468 12124 34692 12180
rect 34412 12086 34468 12124
rect 34412 11956 34468 11966
rect 34300 11620 34356 11630
rect 34188 11618 34356 11620
rect 34188 11566 34302 11618
rect 34354 11566 34356 11618
rect 34188 11564 34356 11566
rect 34300 11554 34356 11564
rect 34412 11506 34468 11900
rect 34412 11454 34414 11506
rect 34466 11454 34468 11506
rect 34412 10164 34468 11454
rect 34524 10612 34580 10622
rect 34524 10518 34580 10556
rect 33852 10098 33908 10108
rect 34300 10108 34468 10164
rect 33628 9940 33684 9950
rect 33628 9846 33684 9884
rect 34188 9828 34244 9838
rect 34188 9734 34244 9772
rect 33964 9716 34020 9726
rect 33964 9622 34020 9660
rect 33628 8930 33684 8942
rect 33628 8878 33630 8930
rect 33682 8878 33684 8930
rect 33628 8820 33684 8878
rect 33628 8754 33684 8764
rect 33404 7698 33572 7700
rect 33404 7646 33406 7698
rect 33458 7646 33572 7698
rect 33404 7644 33572 7646
rect 33404 7634 33460 7644
rect 34188 7586 34244 7598
rect 34188 7534 34190 7586
rect 34242 7534 34244 7586
rect 33852 7474 33908 7486
rect 33852 7422 33854 7474
rect 33906 7422 33908 7474
rect 32732 6598 32788 6636
rect 33516 7362 33572 7374
rect 33516 7310 33518 7362
rect 33570 7310 33572 7362
rect 33292 6466 33348 6478
rect 33292 6414 33294 6466
rect 33346 6414 33348 6466
rect 33292 6356 33348 6414
rect 33516 6356 33572 7310
rect 33852 7364 33908 7422
rect 33852 7298 33908 7308
rect 33852 6916 33908 6926
rect 33852 6578 33908 6860
rect 34188 6916 34244 7534
rect 34188 6850 34244 6860
rect 34300 6692 34356 10108
rect 34412 9940 34468 9950
rect 34412 9846 34468 9884
rect 34524 9826 34580 9838
rect 34524 9774 34526 9826
rect 34578 9774 34580 9826
rect 34524 9604 34580 9774
rect 34524 8820 34580 9548
rect 34636 9380 34692 12124
rect 35084 11956 35140 13806
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35420 12180 35476 12190
rect 35532 12180 35588 14476
rect 35868 14420 35924 14430
rect 35868 13636 35924 14364
rect 36092 14418 36148 14430
rect 36092 14366 36094 14418
rect 36146 14366 36148 14418
rect 36092 14196 36148 14366
rect 36092 14130 36148 14140
rect 36092 13972 36148 13982
rect 36204 13972 36260 15820
rect 36092 13970 36260 13972
rect 36092 13918 36094 13970
rect 36146 13918 36260 13970
rect 36092 13916 36260 13918
rect 36316 15428 36372 16046
rect 36988 15876 37044 19964
rect 37100 19954 37156 19964
rect 37436 20018 37492 20030
rect 37436 19966 37438 20018
rect 37490 19966 37492 20018
rect 37324 19908 37380 19918
rect 37324 19814 37380 19852
rect 37100 19012 37156 19022
rect 37436 19012 37492 19966
rect 37100 19010 37492 19012
rect 37100 18958 37102 19010
rect 37154 18958 37492 19010
rect 37100 18956 37492 18958
rect 38444 19012 38500 19022
rect 37100 18116 37156 18956
rect 37660 18564 37716 18574
rect 37548 18340 37604 18350
rect 37100 18050 37156 18060
rect 37436 18338 37604 18340
rect 37436 18286 37550 18338
rect 37602 18286 37604 18338
rect 37436 18284 37604 18286
rect 37212 17442 37268 17454
rect 37212 17390 37214 17442
rect 37266 17390 37268 17442
rect 37212 16996 37268 17390
rect 37212 16930 37268 16940
rect 36988 15810 37044 15820
rect 37100 16212 37156 16222
rect 37100 15540 37156 16156
rect 37100 15538 37380 15540
rect 37100 15486 37102 15538
rect 37154 15486 37380 15538
rect 37100 15484 37380 15486
rect 37100 15474 37156 15484
rect 36092 13906 36148 13916
rect 35868 13570 35924 13580
rect 35980 13746 36036 13758
rect 36204 13748 36260 13758
rect 35980 13694 35982 13746
rect 36034 13694 36036 13746
rect 35756 13076 35812 13086
rect 35420 12178 35700 12180
rect 35420 12126 35422 12178
rect 35474 12126 35700 12178
rect 35420 12124 35700 12126
rect 35420 12114 35476 12124
rect 35084 11900 35588 11956
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34972 11620 35028 11630
rect 34748 10724 34804 10734
rect 34748 10630 34804 10668
rect 34972 9716 35028 11564
rect 35084 10610 35140 10622
rect 35084 10558 35086 10610
rect 35138 10558 35140 10610
rect 35084 9940 35140 10558
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35420 10052 35476 10062
rect 35084 9884 35364 9940
rect 35084 9716 35140 9726
rect 34972 9714 35140 9716
rect 34972 9662 35086 9714
rect 35138 9662 35140 9714
rect 34972 9660 35140 9662
rect 35084 9650 35140 9660
rect 34748 9604 34804 9614
rect 34748 9602 35028 9604
rect 34748 9550 34750 9602
rect 34802 9550 35028 9602
rect 34748 9548 35028 9550
rect 34748 9538 34804 9548
rect 34692 9324 34916 9380
rect 34636 9286 34692 9324
rect 34860 9266 34916 9324
rect 34860 9214 34862 9266
rect 34914 9214 34916 9266
rect 34860 9202 34916 9214
rect 34524 8754 34580 8764
rect 34972 8370 35028 9548
rect 35196 9268 35252 9884
rect 35308 9826 35364 9884
rect 35308 9774 35310 9826
rect 35362 9774 35364 9826
rect 35308 9762 35364 9774
rect 35420 9716 35476 9996
rect 35532 9938 35588 11900
rect 35644 11620 35700 12124
rect 35644 11554 35700 11564
rect 35644 11394 35700 11406
rect 35644 11342 35646 11394
rect 35698 11342 35700 11394
rect 35644 10386 35700 11342
rect 35756 11170 35812 13020
rect 35980 12404 36036 13694
rect 35980 12338 36036 12348
rect 36092 13746 36260 13748
rect 36092 13694 36206 13746
rect 36258 13694 36260 13746
rect 36092 13692 36260 13694
rect 36092 12402 36148 13692
rect 36204 13682 36260 13692
rect 36316 13076 36372 15372
rect 37324 15316 37380 15484
rect 37436 15538 37492 18284
rect 37548 18274 37604 18284
rect 37660 17668 37716 18508
rect 37548 17666 37716 17668
rect 37548 17614 37662 17666
rect 37714 17614 37716 17666
rect 37548 17612 37716 17614
rect 37548 16770 37604 17612
rect 37660 17602 37716 17612
rect 38220 17668 38276 17678
rect 38444 17668 38500 18956
rect 38220 17666 38500 17668
rect 38220 17614 38222 17666
rect 38274 17614 38500 17666
rect 38220 17612 38500 17614
rect 38556 18452 38612 22094
rect 38892 21812 38948 21822
rect 39004 21812 39060 24668
rect 39228 24658 39284 24668
rect 39228 23380 39284 23390
rect 39228 23266 39284 23324
rect 39228 23214 39230 23266
rect 39282 23214 39284 23266
rect 39228 23202 39284 23214
rect 39340 23380 39396 23390
rect 39452 23380 39508 26236
rect 39564 26226 39620 26236
rect 39676 23380 39732 26852
rect 39788 26290 39844 26302
rect 39788 26238 39790 26290
rect 39842 26238 39844 26290
rect 39788 24948 39844 26238
rect 39900 26290 39956 26302
rect 39900 26238 39902 26290
rect 39954 26238 39956 26290
rect 39900 25284 39956 26238
rect 40236 26180 40292 26852
rect 40572 26850 40628 26862
rect 40572 26798 40574 26850
rect 40626 26798 40628 26850
rect 40572 26292 40628 26798
rect 40572 26226 40628 26236
rect 40236 26114 40292 26124
rect 39900 25218 39956 25228
rect 39788 24882 39844 24892
rect 40908 24722 40964 27020
rect 41132 26964 41188 26974
rect 41132 25508 41188 26908
rect 40908 24670 40910 24722
rect 40962 24670 40964 24722
rect 40908 24658 40964 24670
rect 41020 24948 41076 24958
rect 41020 24610 41076 24892
rect 41020 24558 41022 24610
rect 41074 24558 41076 24610
rect 41020 24546 41076 24558
rect 41132 24946 41188 25452
rect 41132 24894 41134 24946
rect 41186 24894 41188 24946
rect 41132 24050 41188 24894
rect 41132 23998 41134 24050
rect 41186 23998 41188 24050
rect 41132 23986 41188 23998
rect 41244 26290 41300 26302
rect 41244 26238 41246 26290
rect 41298 26238 41300 26290
rect 39340 23378 39508 23380
rect 39340 23326 39342 23378
rect 39394 23326 39508 23378
rect 39340 23324 39508 23326
rect 39564 23324 39732 23380
rect 39340 23268 39396 23324
rect 39340 23202 39396 23212
rect 38892 21810 39060 21812
rect 38892 21758 38894 21810
rect 38946 21758 39060 21810
rect 38892 21756 39060 21758
rect 39340 22930 39396 22942
rect 39340 22878 39342 22930
rect 39394 22878 39396 22930
rect 38892 21746 38948 21756
rect 38780 21588 38836 21598
rect 38780 21586 38948 21588
rect 38780 21534 38782 21586
rect 38834 21534 38948 21586
rect 38780 21532 38948 21534
rect 38780 21522 38836 21532
rect 38780 21140 38836 21150
rect 38780 20914 38836 21084
rect 38780 20862 38782 20914
rect 38834 20862 38836 20914
rect 38780 20850 38836 20862
rect 38668 20804 38724 20814
rect 38892 20804 38948 21532
rect 39004 21586 39060 21598
rect 39004 21534 39006 21586
rect 39058 21534 39060 21586
rect 39004 21140 39060 21534
rect 39228 21588 39284 21598
rect 39340 21588 39396 22878
rect 39452 21588 39508 21598
rect 39340 21586 39508 21588
rect 39340 21534 39454 21586
rect 39506 21534 39508 21586
rect 39340 21532 39508 21534
rect 39228 21474 39284 21532
rect 39452 21522 39508 21532
rect 39228 21422 39230 21474
rect 39282 21422 39284 21474
rect 39228 21364 39284 21422
rect 39564 21364 39620 23324
rect 41244 23268 41300 26238
rect 41356 26292 41412 27356
rect 41468 26964 41524 27002
rect 41468 26898 41524 26908
rect 41356 26226 41412 26236
rect 41580 26290 41636 27580
rect 41692 26908 41748 28590
rect 42028 29204 42084 29214
rect 41692 26852 41860 26908
rect 41580 26238 41582 26290
rect 41634 26238 41636 26290
rect 41580 26226 41636 26238
rect 41580 25508 41636 25518
rect 41580 25414 41636 25452
rect 41804 25506 41860 26852
rect 41804 25454 41806 25506
rect 41858 25454 41860 25506
rect 41356 24948 41412 24958
rect 41356 24854 41412 24892
rect 41804 24948 41860 25454
rect 41804 24882 41860 24892
rect 41916 25394 41972 25406
rect 41916 25342 41918 25394
rect 41970 25342 41972 25394
rect 41580 24724 41636 24734
rect 41580 24722 41748 24724
rect 41580 24670 41582 24722
rect 41634 24670 41748 24722
rect 41580 24668 41748 24670
rect 41580 24658 41636 24668
rect 41580 23940 41636 23950
rect 41580 23846 41636 23884
rect 41132 23212 41300 23268
rect 39228 21308 39620 21364
rect 39676 23156 39732 23166
rect 39676 22370 39732 23100
rect 39676 22318 39678 22370
rect 39730 22318 39732 22370
rect 39676 22148 39732 22318
rect 40460 22260 40516 22270
rect 40460 22258 40964 22260
rect 40460 22206 40462 22258
rect 40514 22206 40964 22258
rect 40460 22204 40964 22206
rect 40460 22194 40516 22204
rect 39004 21074 39060 21084
rect 39564 21028 39620 21038
rect 39116 20916 39172 20926
rect 38892 20748 39060 20804
rect 38668 20132 38724 20748
rect 38892 20578 38948 20590
rect 38892 20526 38894 20578
rect 38946 20526 38948 20578
rect 38892 20356 38948 20526
rect 38892 20290 38948 20300
rect 39004 20468 39060 20748
rect 39116 20802 39172 20860
rect 39116 20750 39118 20802
rect 39170 20750 39172 20802
rect 39116 20738 39172 20750
rect 39564 20802 39620 20972
rect 39564 20750 39566 20802
rect 39618 20750 39620 20802
rect 39564 20738 39620 20750
rect 39004 20244 39060 20412
rect 39340 20690 39396 20702
rect 39340 20638 39342 20690
rect 39394 20638 39396 20690
rect 39228 20356 39284 20366
rect 39116 20244 39172 20254
rect 39004 20242 39172 20244
rect 39004 20190 39118 20242
rect 39170 20190 39172 20242
rect 39004 20188 39172 20190
rect 39116 20178 39172 20188
rect 39228 20242 39284 20300
rect 39228 20190 39230 20242
rect 39282 20190 39284 20242
rect 38668 20076 39060 20132
rect 39004 20018 39060 20076
rect 39004 19966 39006 20018
rect 39058 19966 39060 20018
rect 39004 19954 39060 19966
rect 38780 19236 38836 19246
rect 38780 19142 38836 19180
rect 37884 17444 37940 17454
rect 37884 17442 38052 17444
rect 37884 17390 37886 17442
rect 37938 17390 38052 17442
rect 37884 17388 38052 17390
rect 37884 17378 37940 17388
rect 37548 16718 37550 16770
rect 37602 16718 37604 16770
rect 37548 16706 37604 16718
rect 37996 16884 38052 17388
rect 38220 16996 38276 17612
rect 38556 17220 38612 18396
rect 39228 18228 39284 20190
rect 39228 18162 39284 18172
rect 39228 18004 39284 18014
rect 38556 17164 38836 17220
rect 38220 16930 38276 16940
rect 38780 16994 38836 17164
rect 39228 17106 39284 17948
rect 39340 17556 39396 20638
rect 39676 19348 39732 22092
rect 40348 21812 40404 21822
rect 40348 21474 40404 21756
rect 40348 21422 40350 21474
rect 40402 21422 40404 21474
rect 40012 20972 40292 21028
rect 40012 20802 40068 20972
rect 40012 20750 40014 20802
rect 40066 20750 40068 20802
rect 40012 20738 40068 20750
rect 40124 20802 40180 20814
rect 40124 20750 40126 20802
rect 40178 20750 40180 20802
rect 39788 20692 39844 20702
rect 39788 20598 39844 20636
rect 40012 20468 40068 20478
rect 40124 20468 40180 20750
rect 40068 20412 40180 20468
rect 40012 20402 40068 20412
rect 39900 19348 39956 19358
rect 39732 19346 40180 19348
rect 39732 19294 39902 19346
rect 39954 19294 40180 19346
rect 39732 19292 40180 19294
rect 39676 19254 39732 19292
rect 39900 19282 39956 19292
rect 40012 19012 40068 19022
rect 39676 18338 39732 18350
rect 39676 18286 39678 18338
rect 39730 18286 39732 18338
rect 39676 17780 39732 18286
rect 39676 17714 39732 17724
rect 39340 17490 39396 17500
rect 39228 17054 39230 17106
rect 39282 17054 39284 17106
rect 39228 17042 39284 17054
rect 38780 16942 38782 16994
rect 38834 16942 38836 16994
rect 38780 16930 38836 16942
rect 39788 16994 39844 17006
rect 39788 16942 39790 16994
rect 39842 16942 39844 16994
rect 37996 16210 38052 16828
rect 39004 16884 39060 16894
rect 38108 16324 38164 16334
rect 38108 16230 38164 16268
rect 38556 16212 38612 16222
rect 37996 16158 37998 16210
rect 38050 16158 38052 16210
rect 37996 15652 38052 16158
rect 38220 16210 38612 16212
rect 38220 16158 38558 16210
rect 38610 16158 38612 16210
rect 38220 16156 38612 16158
rect 37996 15596 38164 15652
rect 37436 15486 37438 15538
rect 37490 15486 37492 15538
rect 37436 15474 37492 15486
rect 37436 15316 37492 15326
rect 37324 15314 37492 15316
rect 37324 15262 37438 15314
rect 37490 15262 37492 15314
rect 37324 15260 37492 15262
rect 37436 15250 37492 15260
rect 37996 15314 38052 15326
rect 37996 15262 37998 15314
rect 38050 15262 38052 15314
rect 37772 15204 37828 15214
rect 37100 15092 37156 15102
rect 36428 13972 36484 13982
rect 36428 13878 36484 13916
rect 37100 13972 37156 15036
rect 37772 15090 37828 15148
rect 37772 15038 37774 15090
rect 37826 15038 37828 15090
rect 37772 15026 37828 15038
rect 37100 13878 37156 13916
rect 37548 14196 37604 14206
rect 37548 13970 37604 14140
rect 37548 13918 37550 13970
rect 37602 13918 37604 13970
rect 37548 13906 37604 13918
rect 37884 13858 37940 13870
rect 37884 13806 37886 13858
rect 37938 13806 37940 13858
rect 37772 13748 37828 13758
rect 37884 13748 37940 13806
rect 37996 13860 38052 15262
rect 38108 14530 38164 15596
rect 38220 15426 38276 16156
rect 38556 16146 38612 16156
rect 38220 15374 38222 15426
rect 38274 15374 38276 15426
rect 38220 14644 38276 15374
rect 38444 15986 38500 15998
rect 38444 15934 38446 15986
rect 38498 15934 38500 15986
rect 38220 14578 38276 14588
rect 38332 15316 38388 15326
rect 38108 14478 38110 14530
rect 38162 14478 38164 14530
rect 38108 14466 38164 14478
rect 38220 14420 38276 14430
rect 38332 14420 38388 15260
rect 38444 14530 38500 15934
rect 38556 15428 38612 15438
rect 38556 15334 38612 15372
rect 38892 15428 38948 15438
rect 39004 15428 39060 16828
rect 39340 16884 39396 16894
rect 39788 16884 39844 16942
rect 39340 16882 39788 16884
rect 39340 16830 39342 16882
rect 39394 16830 39788 16882
rect 39340 16828 39788 16830
rect 39116 16772 39172 16782
rect 39116 16678 39172 16716
rect 38892 15426 39060 15428
rect 38892 15374 38894 15426
rect 38946 15374 39060 15426
rect 38892 15372 39060 15374
rect 38892 15362 38948 15372
rect 39116 15316 39172 15326
rect 39340 15316 39396 16828
rect 39788 16790 39844 16828
rect 39172 15260 39396 15316
rect 38668 15204 38724 15242
rect 39116 15222 39172 15260
rect 38668 15138 38724 15148
rect 38444 14478 38446 14530
rect 38498 14478 38500 14530
rect 38444 14466 38500 14478
rect 39900 14644 39956 14654
rect 38220 14418 38388 14420
rect 38220 14366 38222 14418
rect 38274 14366 38388 14418
rect 38220 14364 38388 14366
rect 38668 14420 38724 14430
rect 38220 14354 38276 14364
rect 37996 13794 38052 13804
rect 38668 13858 38724 14364
rect 38668 13806 38670 13858
rect 38722 13806 38724 13858
rect 38668 13794 38724 13806
rect 38892 13860 38948 13870
rect 37772 13746 37940 13748
rect 37772 13694 37774 13746
rect 37826 13694 37940 13746
rect 37772 13692 37940 13694
rect 38220 13746 38276 13758
rect 38220 13694 38222 13746
rect 38274 13694 38276 13746
rect 37772 13682 37828 13692
rect 38108 13636 38164 13646
rect 38220 13636 38276 13694
rect 38332 13636 38388 13646
rect 38220 13634 38388 13636
rect 38220 13582 38334 13634
rect 38386 13582 38388 13634
rect 38220 13580 38388 13582
rect 36316 13010 36372 13020
rect 37436 13522 37492 13534
rect 37436 13470 37438 13522
rect 37490 13470 37492 13522
rect 37100 12404 37156 12414
rect 36092 12350 36094 12402
rect 36146 12350 36148 12402
rect 36092 12338 36148 12350
rect 36988 12348 37100 12404
rect 37156 12348 37380 12404
rect 35868 12292 35924 12302
rect 35868 11394 35924 12236
rect 36988 12290 37044 12348
rect 37100 12338 37156 12348
rect 36988 12238 36990 12290
rect 37042 12238 37044 12290
rect 36988 12226 37044 12238
rect 36204 12180 36260 12190
rect 36316 12180 36372 12190
rect 36204 12178 36316 12180
rect 36204 12126 36206 12178
rect 36258 12126 36316 12178
rect 36204 12124 36316 12126
rect 36204 12114 36260 12124
rect 35868 11342 35870 11394
rect 35922 11342 35924 11394
rect 35868 11330 35924 11342
rect 35756 11118 35758 11170
rect 35810 11118 35812 11170
rect 35756 11106 35812 11118
rect 35644 10334 35646 10386
rect 35698 10334 35700 10386
rect 35644 10322 35700 10334
rect 35756 10610 35812 10622
rect 35756 10558 35758 10610
rect 35810 10558 35812 10610
rect 35532 9886 35534 9938
rect 35586 9886 35588 9938
rect 35532 9874 35588 9886
rect 35756 9828 35812 10558
rect 35756 9734 35812 9772
rect 35532 9716 35588 9726
rect 35420 9714 35588 9716
rect 35420 9662 35534 9714
rect 35586 9662 35588 9714
rect 35420 9660 35588 9662
rect 35532 9650 35588 9660
rect 35196 9174 35252 9212
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 34972 8318 34974 8370
rect 35026 8318 35028 8370
rect 34972 8306 35028 8318
rect 35756 8258 35812 8270
rect 35756 8206 35758 8258
rect 35810 8206 35812 8258
rect 35756 8036 35812 8206
rect 36204 8036 36260 8046
rect 35756 8034 36260 8036
rect 35756 7982 36206 8034
rect 36258 7982 36260 8034
rect 35756 7980 36260 7982
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 36092 7028 36148 7038
rect 35196 6804 35252 6814
rect 34300 6690 34916 6692
rect 34300 6638 34302 6690
rect 34354 6638 34916 6690
rect 34300 6636 34916 6638
rect 34300 6626 34356 6636
rect 33852 6526 33854 6578
rect 33906 6526 33908 6578
rect 33852 6514 33908 6526
rect 34076 6468 34132 6478
rect 34076 6374 34132 6412
rect 34188 6466 34244 6478
rect 34188 6414 34190 6466
rect 34242 6414 34244 6466
rect 33292 6300 33684 6356
rect 33292 6132 33348 6142
rect 33292 6038 33348 6076
rect 32508 5954 32564 5964
rect 33516 5908 33572 5918
rect 31388 5854 31390 5906
rect 31442 5854 31444 5906
rect 31388 5842 31444 5854
rect 33404 5906 33572 5908
rect 33404 5854 33518 5906
rect 33570 5854 33572 5906
rect 33404 5852 33572 5854
rect 31276 5618 31332 5628
rect 31948 5794 32004 5806
rect 31948 5742 31950 5794
rect 32002 5742 32004 5794
rect 31388 5236 31444 5246
rect 31164 5234 31444 5236
rect 31164 5182 31390 5234
rect 31442 5182 31444 5234
rect 31164 5180 31444 5182
rect 31388 5170 31444 5180
rect 30716 5070 30718 5122
rect 30770 5070 30772 5122
rect 30716 5058 30772 5070
rect 30156 5012 30212 5022
rect 30156 4918 30212 4956
rect 28700 4498 28756 4508
rect 28812 4844 29204 4900
rect 29372 4898 29428 4910
rect 29372 4846 29374 4898
rect 29426 4846 29428 4898
rect 28364 4340 28420 4350
rect 28812 4340 28868 4844
rect 29372 4452 29428 4846
rect 31612 4900 31668 4910
rect 31276 4564 31332 4574
rect 29484 4452 29540 4462
rect 29372 4450 29540 4452
rect 29372 4398 29486 4450
rect 29538 4398 29540 4450
rect 29372 4396 29540 4398
rect 29484 4386 29540 4396
rect 28364 4338 28868 4340
rect 28364 4286 28366 4338
rect 28418 4286 28814 4338
rect 28866 4286 28868 4338
rect 28364 4284 28868 4286
rect 28364 4274 28420 4284
rect 28812 4274 28868 4284
rect 30940 4340 30996 4350
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 28140 3490 28196 3500
rect 28588 3556 28644 3566
rect 28588 3462 28644 3500
rect 28924 3556 28980 3566
rect 28924 800 28980 3500
rect 29596 3444 29652 3454
rect 29596 800 29652 3388
rect 30940 800 30996 4284
rect 31276 3442 31332 4508
rect 31612 4228 31668 4844
rect 31948 4228 32004 5742
rect 32396 5794 32452 5806
rect 32396 5742 32398 5794
rect 32450 5742 32452 5794
rect 32172 5012 32228 5022
rect 32172 4562 32228 4956
rect 32172 4510 32174 4562
rect 32226 4510 32228 4562
rect 32172 4498 32228 4510
rect 32396 4340 32452 5742
rect 32396 4246 32452 4284
rect 32956 5236 33012 5246
rect 31612 4134 31668 4172
rect 31724 4172 32004 4228
rect 32172 4228 32228 4238
rect 31612 3556 31668 3566
rect 31724 3556 31780 4172
rect 31668 3500 31780 3556
rect 32172 3554 32228 4172
rect 32172 3502 32174 3554
rect 32226 3502 32228 3554
rect 31612 3462 31668 3500
rect 32172 3490 32228 3502
rect 31276 3390 31278 3442
rect 31330 3390 31332 3442
rect 31276 3378 31332 3390
rect 32956 800 33012 5180
rect 33404 4562 33460 5852
rect 33516 5842 33572 5852
rect 33516 5236 33572 5246
rect 33628 5236 33684 6300
rect 33740 6132 33796 6142
rect 33796 6076 33908 6132
rect 33740 6066 33796 6076
rect 33740 5796 33796 5806
rect 33740 5702 33796 5740
rect 33852 5572 33908 6076
rect 34188 6018 34244 6414
rect 34748 6466 34804 6478
rect 34748 6414 34750 6466
rect 34802 6414 34804 6466
rect 34748 6132 34804 6414
rect 34748 6066 34804 6076
rect 34188 5966 34190 6018
rect 34242 5966 34244 6018
rect 34188 5954 34244 5966
rect 33964 5906 34020 5918
rect 33964 5854 33966 5906
rect 34018 5854 34020 5906
rect 33964 5684 34020 5854
rect 34636 5908 34692 5918
rect 34636 5814 34692 5852
rect 34300 5796 34356 5806
rect 34748 5796 34804 5806
rect 34356 5740 34580 5796
rect 34300 5730 34356 5740
rect 33964 5618 34020 5628
rect 33516 5234 33684 5236
rect 33516 5182 33518 5234
rect 33570 5182 33684 5234
rect 33516 5180 33684 5182
rect 33740 5516 33908 5572
rect 33516 5124 33572 5180
rect 33516 5058 33572 5068
rect 33404 4510 33406 4562
rect 33458 4510 33460 4562
rect 33404 4498 33460 4510
rect 33740 4338 33796 5516
rect 33852 5124 33908 5134
rect 33852 5030 33908 5068
rect 34524 4450 34580 5740
rect 34748 5702 34804 5740
rect 34860 5460 34916 6636
rect 34972 6468 35028 6478
rect 34972 6018 35028 6412
rect 34972 5966 34974 6018
rect 35026 5966 35028 6018
rect 34972 5954 35028 5966
rect 35196 6018 35252 6748
rect 35980 6804 36036 6814
rect 35980 6710 36036 6748
rect 36092 6690 36148 6972
rect 36092 6638 36094 6690
rect 36146 6638 36148 6690
rect 36092 6626 36148 6638
rect 35532 6578 35588 6590
rect 35532 6526 35534 6578
rect 35586 6526 35588 6578
rect 35420 6468 35476 6478
rect 35420 6374 35476 6412
rect 35196 5966 35198 6018
rect 35250 5966 35252 6018
rect 35196 5954 35252 5966
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 34860 5404 35028 5460
rect 35196 5450 35460 5460
rect 34860 5236 34916 5246
rect 34860 5142 34916 5180
rect 34972 5012 35028 5404
rect 34972 4946 35028 4956
rect 35532 4564 35588 6526
rect 35868 6468 35924 6478
rect 35868 6374 35924 6412
rect 35644 6132 35700 6142
rect 35644 5906 35700 6076
rect 36204 6132 36260 7980
rect 36316 7028 36372 12124
rect 36428 12178 36484 12190
rect 36428 12126 36430 12178
rect 36482 12126 36484 12178
rect 36428 11172 36484 12126
rect 36764 12178 36820 12190
rect 36764 12126 36766 12178
rect 36818 12126 36820 12178
rect 36764 11956 36820 12126
rect 37212 12180 37268 12190
rect 37212 12086 37268 12124
rect 36764 11890 36820 11900
rect 37100 12066 37156 12078
rect 37100 12014 37102 12066
rect 37154 12014 37156 12066
rect 36428 11106 36484 11116
rect 36540 11620 36596 11630
rect 36540 10722 36596 11564
rect 37100 11396 37156 12014
rect 37212 11396 37268 11406
rect 37100 11394 37268 11396
rect 37100 11342 37214 11394
rect 37266 11342 37268 11394
rect 37100 11340 37268 11342
rect 37212 11330 37268 11340
rect 36876 11284 36932 11294
rect 36876 11190 36932 11228
rect 37100 11172 37156 11182
rect 36988 11116 37100 11172
rect 36876 10836 36932 10846
rect 36988 10836 37044 11116
rect 37100 11078 37156 11116
rect 37324 10836 37380 12348
rect 37436 12180 37492 13470
rect 37996 12404 38052 12414
rect 37996 12310 38052 12348
rect 38108 12402 38164 13580
rect 38108 12350 38110 12402
rect 38162 12350 38164 12402
rect 38108 12338 38164 12350
rect 37772 12180 37828 12190
rect 37436 12178 37716 12180
rect 37436 12126 37438 12178
rect 37490 12126 37716 12178
rect 37436 12124 37716 12126
rect 37436 12114 37492 12124
rect 37660 11956 37716 12124
rect 37772 12086 37828 12124
rect 38220 12180 38276 12190
rect 38332 12180 38388 13580
rect 38220 12178 38388 12180
rect 38220 12126 38222 12178
rect 38274 12126 38388 12178
rect 38220 12124 38388 12126
rect 38444 12292 38500 12302
rect 38444 12178 38500 12236
rect 38444 12126 38446 12178
rect 38498 12126 38500 12178
rect 37996 11956 38052 11966
rect 37660 11900 37996 11956
rect 37996 11618 38052 11900
rect 37996 11566 37998 11618
rect 38050 11566 38052 11618
rect 37996 11554 38052 11566
rect 38108 11282 38164 11294
rect 38108 11230 38110 11282
rect 38162 11230 38164 11282
rect 38108 10836 38164 11230
rect 36876 10834 37044 10836
rect 36876 10782 36878 10834
rect 36930 10782 37044 10834
rect 36876 10780 37044 10782
rect 37100 10780 37380 10836
rect 37772 10780 38164 10836
rect 36876 10770 36932 10780
rect 36540 10670 36542 10722
rect 36594 10670 36596 10722
rect 36540 10658 36596 10670
rect 36764 10610 36820 10622
rect 36764 10558 36766 10610
rect 36818 10558 36820 10610
rect 36652 10052 36708 10062
rect 36652 8820 36708 9996
rect 36764 9604 36820 10558
rect 36988 10610 37044 10622
rect 36988 10558 36990 10610
rect 37042 10558 37044 10610
rect 36988 10052 37044 10558
rect 36988 9986 37044 9996
rect 36988 9604 37044 9614
rect 36764 9602 37044 9604
rect 36764 9550 36990 9602
rect 37042 9550 37044 9602
rect 36764 9548 37044 9550
rect 36876 8932 36932 9548
rect 36988 9538 37044 9548
rect 36988 9268 37044 9278
rect 37100 9268 37156 10780
rect 37212 10612 37268 10622
rect 37772 10612 37828 10780
rect 38220 10724 38276 12124
rect 38444 12114 38500 12126
rect 38780 12180 38836 12190
rect 38780 12086 38836 12124
rect 38444 10836 38500 10846
rect 38444 10742 38500 10780
rect 38892 10836 38948 13804
rect 39788 13860 39844 13870
rect 39788 13766 39844 13804
rect 39900 13858 39956 14588
rect 40012 14420 40068 18956
rect 40124 18674 40180 19292
rect 40124 18622 40126 18674
rect 40178 18622 40180 18674
rect 40124 18610 40180 18622
rect 40236 18004 40292 20972
rect 40236 17938 40292 17948
rect 40348 17892 40404 21422
rect 40796 21476 40852 21486
rect 40684 20804 40740 20814
rect 40684 20690 40740 20748
rect 40796 20802 40852 21420
rect 40908 21474 40964 22204
rect 41020 21812 41076 21822
rect 41020 21718 41076 21756
rect 40908 21422 40910 21474
rect 40962 21422 40964 21474
rect 40908 21410 40964 21422
rect 41132 21028 41188 23212
rect 41244 23044 41300 23054
rect 41244 21698 41300 22988
rect 41244 21646 41246 21698
rect 41298 21646 41300 21698
rect 41244 21634 41300 21646
rect 41692 22932 41748 24668
rect 41916 23604 41972 25342
rect 42028 25172 42084 29148
rect 42140 28756 42196 28766
rect 42140 26066 42196 28700
rect 42588 28644 42644 29374
rect 42700 29428 42756 29438
rect 42700 29334 42756 29372
rect 42588 28578 42644 28588
rect 42700 28868 42756 28878
rect 42588 27860 42644 27870
rect 42252 27188 42308 27198
rect 42252 27074 42308 27132
rect 42588 27186 42644 27804
rect 42588 27134 42590 27186
rect 42642 27134 42644 27186
rect 42588 27122 42644 27134
rect 42252 27022 42254 27074
rect 42306 27022 42308 27074
rect 42252 26290 42308 27022
rect 42364 26964 42420 27002
rect 42364 26898 42420 26908
rect 42700 26908 42756 28812
rect 42812 27300 42868 27310
rect 42812 27074 42868 27244
rect 43036 27298 43092 29596
rect 43036 27246 43038 27298
rect 43090 27246 43092 27298
rect 43036 27234 43092 27246
rect 43148 29428 43204 29438
rect 42812 27022 42814 27074
rect 42866 27022 42868 27074
rect 42812 27010 42868 27022
rect 42700 26852 42868 26908
rect 42252 26238 42254 26290
rect 42306 26238 42308 26290
rect 42252 26226 42308 26238
rect 42588 26292 42644 26302
rect 42140 26014 42142 26066
rect 42194 26014 42196 26066
rect 42140 26002 42196 26014
rect 42476 26180 42532 26190
rect 42476 25508 42532 26124
rect 42588 25620 42644 26236
rect 42588 25554 42644 25564
rect 42812 26292 42868 26852
rect 42924 26292 42980 26302
rect 42812 26290 42980 26292
rect 42812 26238 42926 26290
rect 42978 26238 42980 26290
rect 42812 26236 42980 26238
rect 42028 25116 42196 25172
rect 42028 24948 42084 24958
rect 42028 24854 42084 24892
rect 42028 24612 42084 24622
rect 42028 24050 42084 24556
rect 42028 23998 42030 24050
rect 42082 23998 42084 24050
rect 42028 23986 42084 23998
rect 42140 23716 42196 25116
rect 42252 24948 42308 24958
rect 42252 24946 42420 24948
rect 42252 24894 42254 24946
rect 42306 24894 42420 24946
rect 42252 24892 42420 24894
rect 42252 24882 42308 24892
rect 42252 23716 42308 23726
rect 42140 23660 42252 23716
rect 42252 23650 42308 23660
rect 41916 23548 42084 23604
rect 40796 20750 40798 20802
rect 40850 20750 40852 20802
rect 40796 20738 40852 20750
rect 40908 20972 41188 21028
rect 40684 20638 40686 20690
rect 40738 20638 40740 20690
rect 40684 20626 40740 20638
rect 40460 20580 40516 20590
rect 40908 20580 40964 20972
rect 40460 20486 40516 20524
rect 40796 20524 40964 20580
rect 41692 20802 41748 22876
rect 42028 21810 42084 23548
rect 42252 23492 42308 23502
rect 42028 21758 42030 21810
rect 42082 21758 42084 21810
rect 41804 21586 41860 21598
rect 41804 21534 41806 21586
rect 41858 21534 41860 21586
rect 41804 21140 41860 21534
rect 41916 21476 41972 21486
rect 41916 21382 41972 21420
rect 41804 21074 41860 21084
rect 41804 20916 41860 20926
rect 41804 20914 41972 20916
rect 41804 20862 41806 20914
rect 41858 20862 41972 20914
rect 41804 20860 41972 20862
rect 41804 20850 41860 20860
rect 41692 20750 41694 20802
rect 41746 20750 41748 20802
rect 41692 20580 41748 20750
rect 40348 17826 40404 17836
rect 40124 17780 40180 17790
rect 40124 17106 40180 17724
rect 40124 17054 40126 17106
rect 40178 17054 40180 17106
rect 40124 17042 40180 17054
rect 40236 17778 40292 17790
rect 40236 17726 40238 17778
rect 40290 17726 40292 17778
rect 40236 15148 40292 17726
rect 40796 16660 40852 20524
rect 41692 20514 41748 20524
rect 41804 20690 41860 20702
rect 41804 20638 41806 20690
rect 41858 20638 41860 20690
rect 41804 20130 41860 20638
rect 41804 20078 41806 20130
rect 41858 20078 41860 20130
rect 41804 20066 41860 20078
rect 41804 19124 41860 19134
rect 41132 18564 41188 18574
rect 41020 18562 41188 18564
rect 41020 18510 41134 18562
rect 41186 18510 41188 18562
rect 41020 18508 41188 18510
rect 41020 18452 41076 18508
rect 41132 18498 41188 18508
rect 41020 18386 41076 18396
rect 41468 18452 41524 18462
rect 41804 18452 41860 19068
rect 41916 19010 41972 20860
rect 42028 20020 42084 21758
rect 42140 23436 42252 23492
rect 42140 20804 42196 23436
rect 42252 23426 42308 23436
rect 42252 23044 42308 23054
rect 42252 22950 42308 22988
rect 42364 21586 42420 24892
rect 42476 24722 42532 25452
rect 42476 24670 42478 24722
rect 42530 24670 42532 24722
rect 42476 24658 42532 24670
rect 42700 24612 42756 24622
rect 42812 24612 42868 26236
rect 42924 26226 42980 26236
rect 43148 26290 43204 29372
rect 43708 29428 43764 29596
rect 44044 29650 44660 29652
rect 44044 29598 44046 29650
rect 44098 29598 44660 29650
rect 44044 29596 44660 29598
rect 44044 29586 44100 29596
rect 44380 29428 44436 29438
rect 43708 29426 43876 29428
rect 43708 29374 43710 29426
rect 43762 29374 43876 29426
rect 43708 29372 43876 29374
rect 43708 29362 43764 29372
rect 43484 29314 43540 29326
rect 43484 29262 43486 29314
rect 43538 29262 43540 29314
rect 43148 26238 43150 26290
rect 43202 26238 43204 26290
rect 43148 26226 43204 26238
rect 43260 28644 43316 28654
rect 43484 28644 43540 29262
rect 43316 28588 43540 28644
rect 43820 28866 43876 29372
rect 43820 28814 43822 28866
rect 43874 28814 43876 28866
rect 43260 25506 43316 28588
rect 43484 28084 43540 28094
rect 43484 27990 43540 28028
rect 43820 27858 43876 28814
rect 44156 29426 44436 29428
rect 44156 29374 44382 29426
rect 44434 29374 44436 29426
rect 44156 29372 44436 29374
rect 44156 28866 44212 29372
rect 44380 29362 44436 29372
rect 44604 29426 44660 29596
rect 44604 29374 44606 29426
rect 44658 29374 44660 29426
rect 44604 29362 44660 29374
rect 44156 28814 44158 28866
rect 44210 28814 44212 28866
rect 44156 28802 44212 28814
rect 44716 29204 44772 29708
rect 45388 29428 45444 31726
rect 45500 32452 45556 32462
rect 45500 31106 45556 32396
rect 45500 31054 45502 31106
rect 45554 31054 45556 31106
rect 45500 31042 45556 31054
rect 45612 30996 45668 32734
rect 45948 32788 46004 34078
rect 46284 34130 46340 34188
rect 46284 34078 46286 34130
rect 46338 34078 46340 34130
rect 46284 34066 46340 34078
rect 46396 34018 46452 34030
rect 46396 33966 46398 34018
rect 46450 33966 46452 34018
rect 46396 33572 46452 33966
rect 46060 33516 46452 33572
rect 46060 33458 46116 33516
rect 46060 33406 46062 33458
rect 46114 33406 46116 33458
rect 46060 33394 46116 33406
rect 45948 32694 46004 32732
rect 46172 32900 46228 32910
rect 46172 32786 46228 32844
rect 46508 32788 46564 34188
rect 46620 34132 46676 34142
rect 46620 34038 46676 34076
rect 46732 34130 46788 34300
rect 46956 34290 47012 34300
rect 46732 34078 46734 34130
rect 46786 34078 46788 34130
rect 46732 34066 46788 34078
rect 47068 33124 47124 33134
rect 46172 32734 46174 32786
rect 46226 32734 46228 32786
rect 46172 32722 46228 32734
rect 46396 32732 46564 32788
rect 46844 33012 46900 33022
rect 46844 32786 46900 32956
rect 46844 32734 46846 32786
rect 46898 32734 46900 32786
rect 46060 32452 46116 32462
rect 46396 32452 46452 32732
rect 46844 32722 46900 32734
rect 46060 32450 46228 32452
rect 46060 32398 46062 32450
rect 46114 32398 46228 32450
rect 46060 32396 46228 32398
rect 46060 32386 46116 32396
rect 46060 31668 46116 31678
rect 45724 31666 46116 31668
rect 45724 31614 46062 31666
rect 46114 31614 46116 31666
rect 45724 31612 46116 31614
rect 45724 31218 45780 31612
rect 46060 31602 46116 31612
rect 45724 31166 45726 31218
rect 45778 31166 45780 31218
rect 45724 31154 45780 31166
rect 46060 31108 46116 31118
rect 46172 31108 46228 32396
rect 46396 32386 46452 32396
rect 46508 32564 46564 32574
rect 47068 32564 47124 33068
rect 46060 31106 46228 31108
rect 46060 31054 46062 31106
rect 46114 31054 46228 31106
rect 46060 31052 46228 31054
rect 46060 31042 46116 31052
rect 45724 30996 45780 31006
rect 45612 30994 45780 30996
rect 45612 30942 45726 30994
rect 45778 30942 45780 30994
rect 45612 30940 45780 30942
rect 45724 30930 45780 30940
rect 45388 29426 45556 29428
rect 45388 29374 45390 29426
rect 45442 29374 45556 29426
rect 45388 29372 45556 29374
rect 45388 29362 45444 29372
rect 44940 29316 44996 29326
rect 44940 29222 44996 29260
rect 44828 29204 44884 29214
rect 44716 29202 44884 29204
rect 44716 29150 44830 29202
rect 44882 29150 44884 29202
rect 44716 29148 44884 29150
rect 44044 28644 44100 28654
rect 44044 28530 44100 28588
rect 44044 28478 44046 28530
rect 44098 28478 44100 28530
rect 44044 28466 44100 28478
rect 43820 27806 43822 27858
rect 43874 27806 43876 27858
rect 43820 27794 43876 27806
rect 44268 28084 44324 28094
rect 44716 28084 44772 29148
rect 44828 29138 44884 29148
rect 44828 28644 44884 28654
rect 45276 28644 45332 28654
rect 44828 28550 44884 28588
rect 44940 28588 45276 28644
rect 44324 28028 44772 28084
rect 44268 27858 44324 28028
rect 44828 27972 44884 27982
rect 44940 27972 44996 28588
rect 45276 28550 45332 28588
rect 44828 27970 44996 27972
rect 44828 27918 44830 27970
rect 44882 27918 44996 27970
rect 44828 27916 44996 27918
rect 44828 27906 44884 27916
rect 44268 27806 44270 27858
rect 44322 27806 44324 27858
rect 44268 27794 44324 27806
rect 45388 27860 45444 27870
rect 45500 27860 45556 29372
rect 46060 29316 46116 29326
rect 46060 29222 46116 29260
rect 45388 27858 45556 27860
rect 45388 27806 45390 27858
rect 45442 27806 45556 27858
rect 45388 27804 45556 27806
rect 45724 28980 45780 28990
rect 45724 28754 45780 28924
rect 45724 28702 45726 28754
rect 45778 28702 45780 28754
rect 44380 27748 44436 27758
rect 44380 27654 44436 27692
rect 44044 27634 44100 27646
rect 44044 27582 44046 27634
rect 44098 27582 44100 27634
rect 43596 27300 43652 27310
rect 43596 27186 43652 27244
rect 43596 27134 43598 27186
rect 43650 27134 43652 27186
rect 43596 27122 43652 27134
rect 44044 27186 44100 27582
rect 44716 27636 44772 27646
rect 44716 27634 45220 27636
rect 44716 27582 44718 27634
rect 44770 27582 45220 27634
rect 44716 27580 45220 27582
rect 44716 27570 44772 27580
rect 44268 27300 44324 27310
rect 44044 27134 44046 27186
rect 44098 27134 44100 27186
rect 44044 27122 44100 27134
rect 44156 27244 44268 27300
rect 43260 25454 43262 25506
rect 43314 25454 43316 25506
rect 43260 25442 43316 25454
rect 43372 27076 43428 27086
rect 43372 24948 43428 27020
rect 43932 27076 43988 27086
rect 43932 26982 43988 27020
rect 44156 26962 44212 27244
rect 44268 27234 44324 27244
rect 45164 27298 45220 27580
rect 45164 27246 45166 27298
rect 45218 27246 45220 27298
rect 44828 27188 44884 27198
rect 44828 27094 44884 27132
rect 44156 26910 44158 26962
rect 44210 26910 44212 26962
rect 43932 26180 43988 26190
rect 43932 26086 43988 26124
rect 43260 24892 43428 24948
rect 43596 25506 43652 25518
rect 43596 25454 43598 25506
rect 43650 25454 43652 25506
rect 43596 24948 43652 25454
rect 44044 25508 44100 25518
rect 43708 24948 43764 24958
rect 43596 24946 43764 24948
rect 43596 24894 43710 24946
rect 43762 24894 43764 24946
rect 43596 24892 43764 24894
rect 42756 24556 42868 24612
rect 42924 24834 42980 24846
rect 42924 24782 42926 24834
rect 42978 24782 42980 24834
rect 42700 24546 42756 24556
rect 42924 24164 42980 24782
rect 42476 24162 42980 24164
rect 42476 24110 42926 24162
rect 42978 24110 42980 24162
rect 42476 24108 42980 24110
rect 42476 23938 42532 24108
rect 42924 24098 42980 24108
rect 42476 23886 42478 23938
rect 42530 23886 42532 23938
rect 42476 23874 42532 23886
rect 43036 23826 43092 23838
rect 43036 23774 43038 23826
rect 43090 23774 43092 23826
rect 42476 23716 42532 23726
rect 42476 23154 42532 23660
rect 43036 23548 43092 23774
rect 42476 23102 42478 23154
rect 42530 23102 42532 23154
rect 42476 23090 42532 23102
rect 42588 23492 42644 23502
rect 42588 22482 42644 23436
rect 42588 22430 42590 22482
rect 42642 22430 42644 22482
rect 42588 22418 42644 22430
rect 42812 23492 43092 23548
rect 42812 22372 42868 23492
rect 42924 23156 42980 23166
rect 42924 23062 42980 23100
rect 43148 23156 43204 23166
rect 42812 22316 43092 22372
rect 43036 22260 43092 22316
rect 43148 22370 43204 23100
rect 43148 22318 43150 22370
rect 43202 22318 43204 22370
rect 43148 22306 43204 22318
rect 43036 22166 43092 22204
rect 42364 21534 42366 21586
rect 42418 21534 42420 21586
rect 42140 20748 42308 20804
rect 42028 19954 42084 19964
rect 42140 20580 42196 20590
rect 41916 18958 41918 19010
rect 41970 18958 41972 19010
rect 41916 18676 41972 18958
rect 42028 19236 42084 19246
rect 42140 19236 42196 20524
rect 42028 19234 42196 19236
rect 42028 19182 42030 19234
rect 42082 19182 42196 19234
rect 42028 19180 42196 19182
rect 42028 19012 42084 19180
rect 42028 18946 42084 18956
rect 41916 18610 41972 18620
rect 41468 18450 41860 18452
rect 41468 18398 41470 18450
rect 41522 18398 41806 18450
rect 41858 18398 41860 18450
rect 41468 18396 41860 18398
rect 41468 18386 41524 18396
rect 41804 18386 41860 18396
rect 41916 18338 41972 18350
rect 41916 18286 41918 18338
rect 41970 18286 41972 18338
rect 41020 18004 41076 18014
rect 41020 16996 41076 17948
rect 41020 16930 41076 16940
rect 41916 16996 41972 18286
rect 42252 18004 42308 20748
rect 42364 20802 42420 21534
rect 42364 20750 42366 20802
rect 42418 20750 42420 20802
rect 42364 20738 42420 20750
rect 42812 22146 42868 22158
rect 42812 22094 42814 22146
rect 42866 22094 42868 22146
rect 42812 20804 42868 22094
rect 42812 20710 42868 20748
rect 43260 20580 43316 24892
rect 43372 24724 43428 24734
rect 43372 24722 43540 24724
rect 43372 24670 43374 24722
rect 43426 24670 43540 24722
rect 43372 24668 43540 24670
rect 43372 24658 43428 24668
rect 43484 23492 43540 24668
rect 43596 23940 43652 24892
rect 43708 24882 43764 24892
rect 43596 23874 43652 23884
rect 43820 24722 43876 24734
rect 43820 24670 43822 24722
rect 43874 24670 43876 24722
rect 43820 23940 43876 24670
rect 43540 23436 43764 23492
rect 43484 23398 43540 23436
rect 43708 23266 43764 23436
rect 43708 23214 43710 23266
rect 43762 23214 43764 23266
rect 43708 23202 43764 23214
rect 43596 23156 43652 23166
rect 43596 23062 43652 23100
rect 43596 22148 43652 22158
rect 43596 22054 43652 22092
rect 43820 21586 43876 23884
rect 43820 21534 43822 21586
rect 43874 21534 43876 21586
rect 43820 21522 43876 21534
rect 44044 21474 44100 25452
rect 44156 25506 44212 26910
rect 44268 27076 44324 27086
rect 44268 26402 44324 27020
rect 44940 27076 44996 27086
rect 44940 26962 44996 27020
rect 44940 26910 44942 26962
rect 44994 26910 44996 26962
rect 44940 26898 44996 26910
rect 45164 26908 45220 27246
rect 45388 26908 45444 27804
rect 44268 26350 44270 26402
rect 44322 26350 44324 26402
rect 44268 26338 44324 26350
rect 45052 26852 45220 26908
rect 45276 26852 45444 26908
rect 44156 25454 44158 25506
rect 44210 25454 44212 25506
rect 44156 25442 44212 25454
rect 45052 25508 45108 26852
rect 45164 26292 45220 26302
rect 45276 26292 45332 26852
rect 45164 26290 45332 26292
rect 45164 26238 45166 26290
rect 45218 26238 45332 26290
rect 45164 26236 45332 26238
rect 45164 26226 45220 26236
rect 45724 25732 45780 28702
rect 46172 28642 46228 28654
rect 46172 28590 46174 28642
rect 46226 28590 46228 28642
rect 46060 27748 46116 27758
rect 46060 27654 46116 27692
rect 46060 27076 46116 27086
rect 46172 27076 46228 28590
rect 46116 27020 46228 27076
rect 46060 26982 46116 27020
rect 46508 26908 46564 32508
rect 46620 32562 47124 32564
rect 46620 32510 47070 32562
rect 47122 32510 47124 32562
rect 46620 32508 47124 32510
rect 46620 31218 46676 32508
rect 47068 32498 47124 32508
rect 46620 31166 46622 31218
rect 46674 31166 46676 31218
rect 46620 31154 46676 31166
rect 47068 31220 47124 31230
rect 47180 31220 47236 35644
rect 47292 34242 47348 35980
rect 47292 34190 47294 34242
rect 47346 34190 47348 34242
rect 47292 34178 47348 34190
rect 47516 34130 47572 38668
rect 47628 38388 47684 41806
rect 47740 41298 47796 43372
rect 47740 41246 47742 41298
rect 47794 41246 47796 41298
rect 47740 41234 47796 41246
rect 47852 43426 47908 43438
rect 47852 43374 47854 43426
rect 47906 43374 47908 43426
rect 47852 40404 47908 43374
rect 47852 40338 47908 40348
rect 47964 42866 48020 42878
rect 47964 42814 47966 42866
rect 48018 42814 48020 42866
rect 47628 38322 47684 38332
rect 47740 40290 47796 40302
rect 47740 40238 47742 40290
rect 47794 40238 47796 40290
rect 47740 37716 47796 40238
rect 47964 39732 48020 42814
rect 47964 39666 48020 39676
rect 48076 39618 48132 44046
rect 48188 41412 48244 41422
rect 48188 41318 48244 41356
rect 48076 39566 48078 39618
rect 48130 39566 48132 39618
rect 48076 39554 48132 39566
rect 48188 38948 48244 38958
rect 48076 38946 48244 38948
rect 48076 38894 48190 38946
rect 48242 38894 48244 38946
rect 48076 38892 48244 38894
rect 47740 37650 47796 37660
rect 47852 38834 47908 38846
rect 47852 38782 47854 38834
rect 47906 38782 47908 38834
rect 47740 37154 47796 37166
rect 47740 37102 47742 37154
rect 47794 37102 47796 37154
rect 47740 35700 47796 37102
rect 47740 35634 47796 35644
rect 47516 34078 47518 34130
rect 47570 34078 47572 34130
rect 47516 34066 47572 34078
rect 47628 35140 47684 35150
rect 47628 32674 47684 35084
rect 47852 34354 47908 38782
rect 47964 36594 48020 36606
rect 47964 36542 47966 36594
rect 48018 36542 48020 36594
rect 47964 35028 48020 36542
rect 47964 34962 48020 34972
rect 48076 34914 48132 38892
rect 48188 38882 48244 38892
rect 48188 36036 48244 36046
rect 48188 35586 48244 35980
rect 48300 35812 48356 44716
rect 48300 35746 48356 35756
rect 48412 37828 48468 45052
rect 48188 35534 48190 35586
rect 48242 35534 48244 35586
rect 48188 35522 48244 35534
rect 48076 34862 48078 34914
rect 48130 34862 48132 34914
rect 48076 34850 48132 34862
rect 48412 34692 48468 37772
rect 47852 34302 47854 34354
rect 47906 34302 47908 34354
rect 47852 34290 47908 34302
rect 48076 34636 48468 34692
rect 47628 32622 47630 32674
rect 47682 32622 47684 32674
rect 47628 32610 47684 32622
rect 47964 32676 48020 32686
rect 48076 32676 48132 34636
rect 48188 33460 48244 33470
rect 48188 33366 48244 33404
rect 47964 32674 48132 32676
rect 47964 32622 47966 32674
rect 48018 32622 48132 32674
rect 47964 32620 48132 32622
rect 48188 32900 48244 32910
rect 47068 31218 47236 31220
rect 47068 31166 47070 31218
rect 47122 31166 47236 31218
rect 47068 31164 47236 31166
rect 47516 31220 47572 31230
rect 47964 31220 48020 32620
rect 48188 31890 48244 32844
rect 48188 31838 48190 31890
rect 48242 31838 48244 31890
rect 48188 31826 48244 31838
rect 48188 31220 48244 31230
rect 47964 31218 48244 31220
rect 47964 31166 48190 31218
rect 48242 31166 48244 31218
rect 47964 31164 48244 31166
rect 47068 31154 47124 31164
rect 47516 31126 47572 31164
rect 48188 31154 48244 31164
rect 47740 31108 47796 31118
rect 46508 26852 46788 26908
rect 45836 26180 45892 26190
rect 45836 26178 46452 26180
rect 45836 26126 45838 26178
rect 45890 26126 46452 26178
rect 45836 26124 46452 26126
rect 45836 26114 45892 26124
rect 45724 25676 45892 25732
rect 45612 25620 45668 25630
rect 45612 25526 45668 25564
rect 45052 25442 45108 25452
rect 45276 25506 45332 25518
rect 45276 25454 45278 25506
rect 45330 25454 45332 25506
rect 44156 25284 44212 25294
rect 45052 25284 45108 25294
rect 44156 25282 45108 25284
rect 44156 25230 44158 25282
rect 44210 25230 45054 25282
rect 45106 25230 45108 25282
rect 44156 25228 45108 25230
rect 44156 25218 44212 25228
rect 44828 24164 44884 24174
rect 44604 23492 44660 23502
rect 44660 23436 44772 23492
rect 44604 23426 44660 23436
rect 44492 23044 44548 23054
rect 44044 21422 44046 21474
rect 44098 21422 44100 21474
rect 44044 21410 44100 21422
rect 44156 22148 44212 22158
rect 44492 22148 44548 22988
rect 44716 22484 44772 23436
rect 44828 23266 44884 24108
rect 44940 23828 44996 23838
rect 44940 23378 44996 23772
rect 44940 23326 44942 23378
rect 44994 23326 44996 23378
rect 44940 23314 44996 23326
rect 44828 23214 44830 23266
rect 44882 23214 44884 23266
rect 44828 23202 44884 23214
rect 45052 22820 45108 25228
rect 45276 23940 45332 25454
rect 45724 25508 45780 25546
rect 45724 25442 45780 25452
rect 45836 25394 45892 25676
rect 45836 25342 45838 25394
rect 45890 25342 45892 25394
rect 45724 25284 45780 25294
rect 45612 24836 45668 24846
rect 45612 24742 45668 24780
rect 45724 24724 45780 25228
rect 45836 24948 45892 25342
rect 45836 24882 45892 24892
rect 46396 24946 46452 26124
rect 46396 24894 46398 24946
rect 46450 24894 46452 24946
rect 46396 24882 46452 24894
rect 45836 24724 45892 24734
rect 45724 24722 45892 24724
rect 45724 24670 45838 24722
rect 45890 24670 45892 24722
rect 45724 24668 45892 24670
rect 45836 24658 45892 24668
rect 45948 24724 46004 24734
rect 46172 24724 46228 24734
rect 45948 24722 46228 24724
rect 45948 24670 45950 24722
rect 46002 24670 46174 24722
rect 46226 24670 46228 24722
rect 45948 24668 46228 24670
rect 45948 24658 46004 24668
rect 46172 24658 46228 24668
rect 46508 24722 46564 24734
rect 46508 24670 46510 24722
rect 46562 24670 46564 24722
rect 45276 23716 45332 23884
rect 46508 23940 46564 24670
rect 46732 24612 46788 26852
rect 46956 25396 47012 25406
rect 46956 25302 47012 25340
rect 47516 25396 47572 25406
rect 47180 25284 47236 25294
rect 47068 25282 47236 25284
rect 47068 25230 47182 25282
rect 47234 25230 47236 25282
rect 47068 25228 47236 25230
rect 46844 24724 46900 24734
rect 46844 24630 46900 24668
rect 46732 24546 46788 24556
rect 47068 24164 47124 25228
rect 47180 25218 47236 25228
rect 47180 24948 47236 24958
rect 47180 24854 47236 24892
rect 47292 24724 47348 24734
rect 47292 24630 47348 24668
rect 47404 24722 47460 24734
rect 47404 24670 47406 24722
rect 47458 24670 47460 24722
rect 47068 24098 47124 24108
rect 46732 23940 46788 23950
rect 47180 23940 47236 23950
rect 46508 23938 46676 23940
rect 46508 23886 46510 23938
rect 46562 23886 46676 23938
rect 46508 23884 46676 23886
rect 46508 23874 46564 23884
rect 46172 23828 46228 23838
rect 46172 23734 46228 23772
rect 45276 23650 45332 23660
rect 45836 23714 45892 23726
rect 45836 23662 45838 23714
rect 45890 23662 45892 23714
rect 45500 23604 45556 23614
rect 45276 23154 45332 23166
rect 45276 23102 45278 23154
rect 45330 23102 45332 23154
rect 45276 23044 45332 23102
rect 45276 22978 45332 22988
rect 44940 22764 45108 22820
rect 44828 22484 44884 22494
rect 44716 22482 44884 22484
rect 44716 22430 44830 22482
rect 44882 22430 44884 22482
rect 44716 22428 44884 22430
rect 44828 22418 44884 22428
rect 44212 22092 44548 22148
rect 43932 21362 43988 21374
rect 43932 21310 43934 21362
rect 43986 21310 43988 21362
rect 43596 21140 43652 21150
rect 43596 20914 43652 21084
rect 43596 20862 43598 20914
rect 43650 20862 43652 20914
rect 43596 20850 43652 20862
rect 43708 20802 43764 20814
rect 43708 20750 43710 20802
rect 43762 20750 43764 20802
rect 43260 20514 43316 20524
rect 43484 20690 43540 20702
rect 43484 20638 43486 20690
rect 43538 20638 43540 20690
rect 43260 20020 43316 20030
rect 43148 20018 43316 20020
rect 43148 19966 43262 20018
rect 43314 19966 43316 20018
rect 43148 19964 43316 19966
rect 42924 19346 42980 19358
rect 42924 19294 42926 19346
rect 42978 19294 42980 19346
rect 42700 19124 42756 19134
rect 42700 19030 42756 19068
rect 42924 18564 42980 19294
rect 42700 18452 42756 18462
rect 42588 18338 42644 18350
rect 42588 18286 42590 18338
rect 42642 18286 42644 18338
rect 42588 18116 42644 18286
rect 42588 18050 42644 18060
rect 42140 17948 42308 18004
rect 42140 17220 42196 17948
rect 42700 17890 42756 18396
rect 42924 18450 42980 18508
rect 42924 18398 42926 18450
rect 42978 18398 42980 18450
rect 42924 18386 42980 18398
rect 43036 19234 43092 19246
rect 43036 19182 43038 19234
rect 43090 19182 43092 19234
rect 42700 17838 42702 17890
rect 42754 17838 42756 17890
rect 42700 17826 42756 17838
rect 42252 17780 42308 17790
rect 42252 17686 42308 17724
rect 43036 17780 43092 19182
rect 43148 18226 43204 19964
rect 43260 19954 43316 19964
rect 43484 19460 43540 20638
rect 43484 19394 43540 19404
rect 43596 19906 43652 19918
rect 43596 19854 43598 19906
rect 43650 19854 43652 19906
rect 43148 18174 43150 18226
rect 43202 18174 43204 18226
rect 43148 18162 43204 18174
rect 43484 18450 43540 18462
rect 43484 18398 43486 18450
rect 43538 18398 43540 18450
rect 43036 17666 43092 17724
rect 43036 17614 43038 17666
rect 43090 17614 43092 17666
rect 43036 17602 43092 17614
rect 43148 18004 43204 18014
rect 43148 17666 43204 17948
rect 43484 17780 43540 18398
rect 43484 17714 43540 17724
rect 43148 17614 43150 17666
rect 43202 17614 43204 17666
rect 43148 17602 43204 17614
rect 43596 17556 43652 19854
rect 43708 19348 43764 20750
rect 43932 20802 43988 21310
rect 43932 20750 43934 20802
rect 43986 20750 43988 20802
rect 43820 20020 43876 20030
rect 43932 20020 43988 20750
rect 43820 20018 43988 20020
rect 43820 19966 43822 20018
rect 43874 19966 43988 20018
rect 43820 19964 43988 19966
rect 44156 20804 44212 22092
rect 44940 21588 44996 22764
rect 45164 22258 45220 22270
rect 45164 22206 45166 22258
rect 45218 22206 45220 22258
rect 45052 21588 45108 21598
rect 44940 21586 45108 21588
rect 44940 21534 45054 21586
rect 45106 21534 45108 21586
rect 44940 21532 45108 21534
rect 43820 19954 43876 19964
rect 43708 18452 43764 19292
rect 43932 19684 43988 19694
rect 43932 19346 43988 19628
rect 43932 19294 43934 19346
rect 43986 19294 43988 19346
rect 43932 19282 43988 19294
rect 44156 19348 44212 20748
rect 44828 20690 44884 20702
rect 44828 20638 44830 20690
rect 44882 20638 44884 20690
rect 44268 20130 44324 20142
rect 44268 20078 44270 20130
rect 44322 20078 44324 20130
rect 44268 20020 44324 20078
rect 44268 19954 44324 19964
rect 44828 19908 44884 20638
rect 44940 20578 44996 20590
rect 44940 20526 44942 20578
rect 44994 20526 44996 20578
rect 44940 20020 44996 20526
rect 44940 19954 44996 19964
rect 44828 19842 44884 19852
rect 44716 19460 44772 19470
rect 44268 19348 44324 19358
rect 44156 19346 44324 19348
rect 44156 19294 44270 19346
rect 44322 19294 44324 19346
rect 44156 19292 44324 19294
rect 44268 18788 44324 19292
rect 44268 18722 44324 18732
rect 44268 18564 44324 18574
rect 44604 18564 44660 18574
rect 44268 18562 44436 18564
rect 44268 18510 44270 18562
rect 44322 18510 44436 18562
rect 44268 18508 44436 18510
rect 44268 18498 44324 18508
rect 44044 18452 44100 18462
rect 43708 18450 44100 18452
rect 43708 18398 44046 18450
rect 44098 18398 44100 18450
rect 43708 18396 44100 18398
rect 44044 18386 44100 18396
rect 43484 17500 43652 17556
rect 43932 17948 44212 18004
rect 42364 17444 42420 17454
rect 43036 17444 43092 17454
rect 42364 17442 42868 17444
rect 42364 17390 42366 17442
rect 42418 17390 42868 17442
rect 42364 17388 42868 17390
rect 42364 17378 42420 17388
rect 42140 17164 42532 17220
rect 41916 16930 41972 16940
rect 40908 16884 40964 16894
rect 40908 16790 40964 16828
rect 42140 16882 42196 16894
rect 42364 16884 42420 16894
rect 42140 16830 42142 16882
rect 42194 16830 42196 16882
rect 41020 16772 41076 16782
rect 40796 16604 40964 16660
rect 40908 16210 40964 16604
rect 40908 16158 40910 16210
rect 40962 16158 40964 16210
rect 40908 16146 40964 16158
rect 40796 16098 40852 16110
rect 40796 16046 40798 16098
rect 40850 16046 40852 16098
rect 40460 15988 40516 15998
rect 40460 15894 40516 15932
rect 40796 15538 40852 16046
rect 40796 15486 40798 15538
rect 40850 15486 40852 15538
rect 40796 15474 40852 15486
rect 41020 15314 41076 16716
rect 41356 16772 41412 16782
rect 41356 15426 41412 16716
rect 41468 16770 41524 16782
rect 41468 16718 41470 16770
rect 41522 16718 41524 16770
rect 41468 16098 41524 16718
rect 42140 16772 42196 16830
rect 42140 16706 42196 16716
rect 42252 16882 42420 16884
rect 42252 16830 42366 16882
rect 42418 16830 42420 16882
rect 42252 16828 42420 16830
rect 42252 16324 42308 16828
rect 42364 16818 42420 16828
rect 42028 16268 42308 16324
rect 41468 16046 41470 16098
rect 41522 16046 41524 16098
rect 41468 16034 41524 16046
rect 41916 16212 41972 16222
rect 41916 16098 41972 16156
rect 41916 16046 41918 16098
rect 41970 16046 41972 16098
rect 41916 16034 41972 16046
rect 42028 15538 42084 16268
rect 42364 16212 42420 16222
rect 42364 16118 42420 16156
rect 42028 15486 42030 15538
rect 42082 15486 42084 15538
rect 42028 15474 42084 15486
rect 42140 16100 42196 16110
rect 42140 15540 42196 16044
rect 42476 16098 42532 17164
rect 42812 17108 42868 17388
rect 42812 16882 42868 17052
rect 43036 17106 43092 17388
rect 43260 17442 43316 17454
rect 43260 17390 43262 17442
rect 43314 17390 43316 17442
rect 43260 17220 43316 17390
rect 43372 17444 43428 17454
rect 43372 17350 43428 17388
rect 43260 17154 43316 17164
rect 43484 17108 43540 17500
rect 43036 17054 43038 17106
rect 43090 17054 43092 17106
rect 43036 17042 43092 17054
rect 43372 17052 43540 17108
rect 42812 16830 42814 16882
rect 42866 16830 42868 16882
rect 42812 16818 42868 16830
rect 43260 16882 43316 16894
rect 43260 16830 43262 16882
rect 43314 16830 43316 16882
rect 43036 16772 43092 16782
rect 43036 16678 43092 16716
rect 43260 16324 43316 16830
rect 43260 16258 43316 16268
rect 43372 16212 43428 17052
rect 43820 16996 43876 17006
rect 43708 16940 43820 16996
rect 43484 16884 43540 16894
rect 43484 16882 43652 16884
rect 43484 16830 43486 16882
rect 43538 16830 43652 16882
rect 43484 16828 43652 16830
rect 43484 16818 43540 16828
rect 43372 16146 43428 16156
rect 43484 16660 43540 16670
rect 43484 16210 43540 16604
rect 43484 16158 43486 16210
rect 43538 16158 43540 16210
rect 43484 16146 43540 16158
rect 42476 16046 42478 16098
rect 42530 16046 42532 16098
rect 42252 15988 42308 15998
rect 42476 15988 42532 16046
rect 42812 16100 42868 16110
rect 42812 16006 42868 16044
rect 42252 15986 42420 15988
rect 42252 15934 42254 15986
rect 42306 15934 42420 15986
rect 42252 15932 42420 15934
rect 42252 15922 42308 15932
rect 42364 15652 42420 15932
rect 42476 15922 42532 15932
rect 43036 15988 43092 15998
rect 42364 15596 42644 15652
rect 42252 15540 42308 15550
rect 42140 15538 42308 15540
rect 42140 15486 42254 15538
rect 42306 15486 42308 15538
rect 42140 15484 42308 15486
rect 41356 15374 41358 15426
rect 41410 15374 41412 15426
rect 41356 15362 41412 15374
rect 41692 15426 41748 15438
rect 41692 15374 41694 15426
rect 41746 15374 41748 15426
rect 41020 15262 41022 15314
rect 41074 15262 41076 15314
rect 41020 15250 41076 15262
rect 41692 15316 41748 15374
rect 41692 15250 41748 15260
rect 41804 15316 41860 15326
rect 42140 15316 42196 15484
rect 42252 15474 42308 15484
rect 41804 15314 42196 15316
rect 41804 15262 41806 15314
rect 41858 15262 42196 15314
rect 41804 15260 42196 15262
rect 42364 15316 42420 15326
rect 41804 15250 41860 15260
rect 42364 15222 42420 15260
rect 42588 15316 42644 15596
rect 43036 15538 43092 15932
rect 43036 15486 43038 15538
rect 43090 15486 43092 15538
rect 43036 15474 43092 15486
rect 43372 15874 43428 15886
rect 43372 15822 43374 15874
rect 43426 15822 43428 15874
rect 43372 15428 43428 15822
rect 42812 15316 42868 15326
rect 42588 15314 42868 15316
rect 42588 15262 42814 15314
rect 42866 15262 42868 15314
rect 42588 15260 42868 15262
rect 40236 15092 40852 15148
rect 40684 14420 40740 14430
rect 40012 14354 40068 14364
rect 40348 14364 40684 14420
rect 40348 13970 40404 14364
rect 40684 14354 40740 14364
rect 40348 13918 40350 13970
rect 40402 13918 40404 13970
rect 39900 13806 39902 13858
rect 39954 13806 39956 13858
rect 39676 13746 39732 13758
rect 39676 13694 39678 13746
rect 39730 13694 39732 13746
rect 39676 13524 39732 13694
rect 39900 13748 39956 13806
rect 39900 13682 39956 13692
rect 40124 13860 40180 13870
rect 40124 13524 40180 13804
rect 39676 13468 40180 13524
rect 40124 12962 40180 13468
rect 40124 12910 40126 12962
rect 40178 12910 40180 12962
rect 40124 12898 40180 12910
rect 40236 13300 40292 13310
rect 40236 12964 40292 13244
rect 40236 12870 40292 12908
rect 40236 12516 40292 12526
rect 38892 10770 38948 10780
rect 39116 12290 39172 12302
rect 39116 12238 39118 12290
rect 39170 12238 39172 12290
rect 39116 12180 39172 12238
rect 40236 12180 40292 12460
rect 40348 12292 40404 13918
rect 40572 13748 40628 13758
rect 40572 12962 40628 13692
rect 40572 12910 40574 12962
rect 40626 12910 40628 12962
rect 40572 12898 40628 12910
rect 40460 12738 40516 12750
rect 40460 12686 40462 12738
rect 40514 12686 40516 12738
rect 40460 12404 40516 12686
rect 40796 12516 40852 15092
rect 41468 14644 41524 14654
rect 40908 14532 40964 14542
rect 40908 13746 40964 14476
rect 41244 14420 41300 14430
rect 41244 14326 41300 14364
rect 41356 14308 41412 14318
rect 41356 14214 41412 14252
rect 41468 13972 41524 14588
rect 41580 14530 41636 14542
rect 41580 14478 41582 14530
rect 41634 14478 41636 14530
rect 41580 14420 41636 14478
rect 41580 14354 41636 14364
rect 42588 14420 42644 15260
rect 42812 15250 42868 15260
rect 43148 15316 43204 15326
rect 43148 15222 43204 15260
rect 43260 15314 43316 15326
rect 43260 15262 43262 15314
rect 43314 15262 43316 15314
rect 42588 14354 42644 14364
rect 42028 14308 42084 14318
rect 42476 14308 42532 14318
rect 42028 14306 42308 14308
rect 42028 14254 42030 14306
rect 42082 14254 42308 14306
rect 42028 14252 42308 14254
rect 42028 14242 42084 14252
rect 41356 13916 41524 13972
rect 41132 13860 41188 13870
rect 41132 13766 41188 13804
rect 40908 13694 40910 13746
rect 40962 13694 40964 13746
rect 40908 13682 40964 13694
rect 41244 13746 41300 13758
rect 41244 13694 41246 13746
rect 41298 13694 41300 13746
rect 41244 13300 41300 13694
rect 41244 13234 41300 13244
rect 41132 13076 41188 13086
rect 41356 13076 41412 13916
rect 41468 13748 41524 13758
rect 41468 13654 41524 13692
rect 41916 13748 41972 13758
rect 41916 13654 41972 13692
rect 41132 13074 41412 13076
rect 41132 13022 41134 13074
rect 41186 13022 41412 13074
rect 41132 13020 41412 13022
rect 41132 13010 41188 13020
rect 41356 12962 41412 13020
rect 42140 13522 42196 13534
rect 42140 13470 42142 13522
rect 42194 13470 42196 13522
rect 42140 13074 42196 13470
rect 42140 13022 42142 13074
rect 42194 13022 42196 13074
rect 42140 13010 42196 13022
rect 42252 13522 42308 14252
rect 42476 13746 42532 14252
rect 43260 13860 43316 15262
rect 43372 15314 43428 15372
rect 43372 15262 43374 15314
rect 43426 15262 43428 15314
rect 43372 15250 43428 15262
rect 43596 15148 43652 16828
rect 42476 13694 42478 13746
rect 42530 13694 42532 13746
rect 42476 13682 42532 13694
rect 42700 13748 42756 13758
rect 42700 13654 42756 13692
rect 42252 13470 42254 13522
rect 42306 13470 42308 13522
rect 41356 12910 41358 12962
rect 41410 12910 41412 12962
rect 41356 12898 41412 12910
rect 41356 12516 41412 12526
rect 40796 12460 41300 12516
rect 40460 12348 41188 12404
rect 40348 12236 40964 12292
rect 40236 12124 40404 12180
rect 38108 10668 38276 10724
rect 37212 10610 37828 10612
rect 37212 10558 37214 10610
rect 37266 10558 37774 10610
rect 37826 10558 37828 10610
rect 37212 10556 37828 10558
rect 37212 10546 37268 10556
rect 37324 10276 37380 10286
rect 37324 9828 37380 10220
rect 37772 10052 37828 10556
rect 37884 10610 37940 10622
rect 37884 10558 37886 10610
rect 37938 10558 37940 10610
rect 37884 10276 37940 10558
rect 37884 10210 37940 10220
rect 37996 10610 38052 10622
rect 37996 10558 37998 10610
rect 38050 10558 38052 10610
rect 37996 10052 38052 10558
rect 37772 9986 37828 9996
rect 37884 9996 38052 10052
rect 37324 9714 37380 9772
rect 37324 9662 37326 9714
rect 37378 9662 37380 9714
rect 37324 9650 37380 9662
rect 37884 9716 37940 9996
rect 36988 9266 37716 9268
rect 36988 9214 36990 9266
rect 37042 9214 37716 9266
rect 36988 9212 37716 9214
rect 36988 9202 37044 9212
rect 37660 9042 37716 9212
rect 37660 8990 37662 9042
rect 37714 8990 37716 9042
rect 37660 8978 37716 8990
rect 36876 8838 36932 8876
rect 37884 8930 37940 9660
rect 37996 9828 38052 9838
rect 37996 9714 38052 9772
rect 37996 9662 37998 9714
rect 38050 9662 38052 9714
rect 37996 9650 38052 9662
rect 37884 8878 37886 8930
rect 37938 8878 37940 8930
rect 37884 8866 37940 8878
rect 36652 8754 36708 8764
rect 37436 8820 37492 8830
rect 37436 7698 37492 8764
rect 37436 7646 37438 7698
rect 37490 7646 37492 7698
rect 37436 7634 37492 7646
rect 37548 7476 37604 7486
rect 38108 7476 38164 10668
rect 38780 10610 38836 10622
rect 38780 10558 38782 10610
rect 38834 10558 38836 10610
rect 38220 10164 38276 10174
rect 38220 9826 38276 10108
rect 38780 10164 38836 10558
rect 39116 10610 39172 12124
rect 40348 12066 40404 12124
rect 40908 12178 40964 12236
rect 40908 12126 40910 12178
rect 40962 12126 40964 12178
rect 40908 12114 40964 12126
rect 41132 12178 41188 12348
rect 41132 12126 41134 12178
rect 41186 12126 41188 12178
rect 41132 12114 41188 12126
rect 40348 12014 40350 12066
rect 40402 12014 40404 12066
rect 40348 12002 40404 12014
rect 40908 11396 40964 11406
rect 41244 11396 41300 12460
rect 41356 12178 41412 12460
rect 42252 12516 42308 13470
rect 42252 12450 42308 12460
rect 43260 12404 43316 13804
rect 43484 15092 43652 15148
rect 43708 15148 43764 16940
rect 43820 16902 43876 16940
rect 43820 16772 43876 16782
rect 43820 15986 43876 16716
rect 43820 15934 43822 15986
rect 43874 15934 43876 15986
rect 43820 15922 43876 15934
rect 43932 15988 43988 17948
rect 44044 17780 44100 17790
rect 44044 17332 44100 17724
rect 44156 17778 44212 17948
rect 44156 17726 44158 17778
rect 44210 17726 44212 17778
rect 44156 17714 44212 17726
rect 44268 17668 44324 17678
rect 44268 17574 44324 17612
rect 44156 17556 44212 17566
rect 44156 17444 44212 17500
rect 44156 17388 44324 17444
rect 44044 17276 44212 17332
rect 44044 17108 44100 17118
rect 44044 17014 44100 17052
rect 44156 16660 44212 17276
rect 44268 17106 44324 17388
rect 44268 17054 44270 17106
rect 44322 17054 44324 17106
rect 44268 17042 44324 17054
rect 44380 16770 44436 18508
rect 44604 18470 44660 18508
rect 44716 18450 44772 19404
rect 44940 19348 44996 19386
rect 44940 19282 44996 19292
rect 45052 19234 45108 21532
rect 45164 21474 45220 22206
rect 45164 21422 45166 21474
rect 45218 21422 45220 21474
rect 45164 20244 45220 21422
rect 45276 20804 45332 20814
rect 45276 20710 45332 20748
rect 45500 20580 45556 23548
rect 45836 23044 45892 23662
rect 46284 23714 46340 23726
rect 46284 23662 46286 23714
rect 46338 23662 46340 23714
rect 46284 23380 46340 23662
rect 46060 23324 46340 23380
rect 46060 23266 46116 23324
rect 46060 23214 46062 23266
rect 46114 23214 46116 23266
rect 46060 23202 46116 23214
rect 45836 22370 45892 22988
rect 45836 22318 45838 22370
rect 45890 22318 45892 22370
rect 45836 22306 45892 22318
rect 46060 21586 46116 21598
rect 46060 21534 46062 21586
rect 46114 21534 46116 21586
rect 46060 20916 46116 21534
rect 45164 20178 45220 20188
rect 45388 20524 45556 20580
rect 45948 20860 46060 20916
rect 46620 20916 46676 23884
rect 46732 23938 47236 23940
rect 46732 23886 46734 23938
rect 46786 23886 47182 23938
rect 47234 23886 47236 23938
rect 46732 23884 47236 23886
rect 46732 23874 46788 23884
rect 47180 23874 47236 23884
rect 47068 23716 47124 23726
rect 47068 23622 47124 23660
rect 47292 23716 47348 23726
rect 47404 23716 47460 24670
rect 47292 23714 47460 23716
rect 47292 23662 47294 23714
rect 47346 23662 47460 23714
rect 47292 23660 47460 23662
rect 47516 23716 47572 25340
rect 46620 20860 47012 20916
rect 45052 19182 45054 19234
rect 45106 19182 45108 19234
rect 45052 19170 45108 19182
rect 45164 19796 45220 19806
rect 45164 19122 45220 19740
rect 45164 19070 45166 19122
rect 45218 19070 45220 19122
rect 45164 19058 45220 19070
rect 44716 18398 44718 18450
rect 44770 18398 44772 18450
rect 44716 18386 44772 18398
rect 44828 18452 44884 18490
rect 44828 18386 44884 18396
rect 45164 18450 45220 18462
rect 45164 18398 45166 18450
rect 45218 18398 45220 18450
rect 44828 18228 44884 18238
rect 44828 17666 44884 18172
rect 45052 17780 45108 17790
rect 45164 17780 45220 18398
rect 45108 17724 45220 17780
rect 45052 17714 45108 17724
rect 44828 17614 44830 17666
rect 44882 17614 44884 17666
rect 44828 17602 44884 17614
rect 44940 17442 44996 17454
rect 44940 17390 44942 17442
rect 44994 17390 44996 17442
rect 44940 17108 44996 17390
rect 44492 17106 44996 17108
rect 44492 17054 44942 17106
rect 44994 17054 44996 17106
rect 44492 17052 44996 17054
rect 44492 16882 44548 17052
rect 44940 17042 44996 17052
rect 45052 17444 45108 17454
rect 44492 16830 44494 16882
rect 44546 16830 44548 16882
rect 44492 16818 44548 16830
rect 44828 16884 44884 16894
rect 45052 16884 45108 17388
rect 44828 16882 45332 16884
rect 44828 16830 44830 16882
rect 44882 16830 45332 16882
rect 44828 16828 45332 16830
rect 44828 16818 44884 16828
rect 44380 16718 44382 16770
rect 44434 16718 44436 16770
rect 44380 16706 44436 16718
rect 44156 16604 44324 16660
rect 43932 15922 43988 15932
rect 44156 15874 44212 15886
rect 44156 15822 44158 15874
rect 44210 15822 44212 15874
rect 43932 15428 43988 15466
rect 43932 15362 43988 15372
rect 44156 15316 44212 15822
rect 44268 15538 44324 16604
rect 45052 16548 45108 16558
rect 45052 16098 45108 16492
rect 45052 16046 45054 16098
rect 45106 16046 45108 16098
rect 45052 16034 45108 16046
rect 44268 15486 44270 15538
rect 44322 15486 44324 15538
rect 44268 15474 44324 15486
rect 45164 15540 45220 15550
rect 45276 15540 45332 16828
rect 45164 15538 45332 15540
rect 45164 15486 45166 15538
rect 45218 15486 45332 15538
rect 45164 15484 45332 15486
rect 44156 15250 44212 15260
rect 44380 15314 44436 15326
rect 44380 15262 44382 15314
rect 44434 15262 44436 15314
rect 44380 15204 44436 15262
rect 43708 15092 43876 15148
rect 43372 12404 43428 12414
rect 43260 12402 43428 12404
rect 43260 12350 43374 12402
rect 43426 12350 43428 12402
rect 43260 12348 43428 12350
rect 43372 12338 43428 12348
rect 41356 12126 41358 12178
rect 41410 12126 41412 12178
rect 41356 12114 41412 12126
rect 41468 11956 41524 11966
rect 41468 11954 41972 11956
rect 41468 11902 41470 11954
rect 41522 11902 41972 11954
rect 41468 11900 41972 11902
rect 41468 11890 41524 11900
rect 41916 11508 41972 11900
rect 42028 11508 42084 11518
rect 41916 11506 42084 11508
rect 41916 11454 42030 11506
rect 42082 11454 42084 11506
rect 41916 11452 42084 11454
rect 42028 11442 42084 11452
rect 40908 11394 41300 11396
rect 40908 11342 40910 11394
rect 40962 11342 41246 11394
rect 41298 11342 41300 11394
rect 40908 11340 41300 11342
rect 40908 11330 40964 11340
rect 39116 10558 39118 10610
rect 39170 10558 39172 10610
rect 39116 10546 39172 10558
rect 39228 10836 39284 10846
rect 39228 10610 39284 10780
rect 39564 10834 39620 10846
rect 39564 10782 39566 10834
rect 39618 10782 39620 10834
rect 39228 10558 39230 10610
rect 39282 10558 39284 10610
rect 39228 10546 39284 10558
rect 39340 10610 39396 10622
rect 39340 10558 39342 10610
rect 39394 10558 39396 10610
rect 38780 10098 38836 10108
rect 39228 10052 39284 10062
rect 39228 9938 39284 9996
rect 39228 9886 39230 9938
rect 39282 9886 39284 9938
rect 39228 9874 39284 9886
rect 39340 9940 39396 10558
rect 39340 9874 39396 9884
rect 39564 9940 39620 10782
rect 39564 9874 39620 9884
rect 38220 9774 38222 9826
rect 38274 9774 38276 9826
rect 38220 9762 38276 9774
rect 38556 9604 38612 9614
rect 38556 9510 38612 9548
rect 41244 9268 41300 11340
rect 43484 11172 43540 15092
rect 43708 14756 43764 14766
rect 43148 11116 43540 11172
rect 43596 13076 43652 13086
rect 41356 9940 41412 9950
rect 41356 9846 41412 9884
rect 42028 9826 42084 9838
rect 42028 9774 42030 9826
rect 42082 9774 42084 9826
rect 42028 9604 42084 9774
rect 43148 9826 43204 11116
rect 43596 10722 43652 13020
rect 43708 12292 43764 14700
rect 43708 12198 43764 12236
rect 43820 11060 43876 15092
rect 44156 15092 44436 15148
rect 45052 15204 45108 15214
rect 44156 13076 44212 15092
rect 44268 14644 44324 14654
rect 44268 14550 44324 14588
rect 45052 14530 45108 15148
rect 45164 14756 45220 15484
rect 45276 15316 45332 15326
rect 45276 15222 45332 15260
rect 45164 14690 45220 14700
rect 45052 14478 45054 14530
rect 45106 14478 45108 14530
rect 45052 14466 45108 14478
rect 44828 14420 44884 14430
rect 44828 14326 44884 14364
rect 45388 14084 45444 20524
rect 45948 20018 46004 20860
rect 46060 20850 46116 20860
rect 46060 20692 46116 20702
rect 46060 20690 46900 20692
rect 46060 20638 46062 20690
rect 46114 20638 46900 20690
rect 46060 20636 46900 20638
rect 46060 20626 46116 20636
rect 46844 20242 46900 20636
rect 46844 20190 46846 20242
rect 46898 20190 46900 20242
rect 46844 20178 46900 20190
rect 45948 19966 45950 20018
rect 46002 19966 46004 20018
rect 45948 19796 46004 19966
rect 45948 19730 46004 19740
rect 46396 20132 46452 20142
rect 46396 19906 46452 20076
rect 46620 20020 46676 20030
rect 46844 20020 46900 20030
rect 46620 19926 46676 19964
rect 46732 19964 46844 20020
rect 46396 19854 46398 19906
rect 46450 19854 46452 19906
rect 46172 19234 46228 19246
rect 46172 19182 46174 19234
rect 46226 19182 46228 19234
rect 46060 19012 46116 19022
rect 45724 19010 46116 19012
rect 45724 18958 46062 19010
rect 46114 18958 46116 19010
rect 45724 18956 46116 18958
rect 45612 18450 45668 18462
rect 45612 18398 45614 18450
rect 45666 18398 45668 18450
rect 45612 18228 45668 18398
rect 45612 18162 45668 18172
rect 45612 17780 45668 17790
rect 45500 17778 45668 17780
rect 45500 17726 45614 17778
rect 45666 17726 45668 17778
rect 45500 17724 45668 17726
rect 45500 16100 45556 17724
rect 45612 17714 45668 17724
rect 45724 17666 45780 18956
rect 46060 18946 46116 18956
rect 45836 18562 45892 18574
rect 45836 18510 45838 18562
rect 45890 18510 45892 18562
rect 45836 18452 45892 18510
rect 45836 18386 45892 18396
rect 45724 17614 45726 17666
rect 45778 17614 45780 17666
rect 45612 16882 45668 16894
rect 45612 16830 45614 16882
rect 45666 16830 45668 16882
rect 45612 16660 45668 16830
rect 45612 16594 45668 16604
rect 45500 16034 45556 16044
rect 45724 15538 45780 17614
rect 46060 18226 46116 18238
rect 46060 18174 46062 18226
rect 46114 18174 46116 18226
rect 45836 17556 45892 17566
rect 45892 17500 46004 17556
rect 45836 17490 45892 17500
rect 45836 17108 45892 17118
rect 45836 16210 45892 17052
rect 45836 16158 45838 16210
rect 45890 16158 45892 16210
rect 45836 16146 45892 16158
rect 45724 15486 45726 15538
rect 45778 15486 45780 15538
rect 45724 15474 45780 15486
rect 45612 15314 45668 15326
rect 45612 15262 45614 15314
rect 45666 15262 45668 15314
rect 45612 15204 45668 15262
rect 45612 15138 45668 15148
rect 45948 14868 46004 17500
rect 46060 17554 46116 18174
rect 46060 17502 46062 17554
rect 46114 17502 46116 17554
rect 46060 17490 46116 17502
rect 46172 16996 46228 19182
rect 46396 19012 46452 19854
rect 46732 19346 46788 19964
rect 46844 19954 46900 19964
rect 46956 20018 47012 20860
rect 47292 20244 47348 23660
rect 47516 23650 47572 23660
rect 47628 24834 47684 24846
rect 47628 24782 47630 24834
rect 47682 24782 47684 24834
rect 47628 24612 47684 24782
rect 47628 23604 47684 24556
rect 47628 23538 47684 23548
rect 47740 23940 47796 31052
rect 48188 29314 48244 29326
rect 48188 29262 48190 29314
rect 48242 29262 48244 29314
rect 48188 28644 48244 29262
rect 48188 28578 48244 28588
rect 48188 27746 48244 27758
rect 48188 27694 48190 27746
rect 48242 27694 48244 27746
rect 48188 27300 48244 27694
rect 48188 27234 48244 27244
rect 47852 27186 47908 27198
rect 47852 27134 47854 27186
rect 47906 27134 47908 27186
rect 47852 26292 47908 27134
rect 48076 27076 48132 27086
rect 48076 26514 48132 27020
rect 48076 26462 48078 26514
rect 48130 26462 48132 26514
rect 48076 26450 48132 26462
rect 47852 26226 47908 26236
rect 48188 25394 48244 25406
rect 48188 25342 48190 25394
rect 48242 25342 48244 25394
rect 47852 25284 47908 25294
rect 47852 25190 47908 25228
rect 48188 24948 48244 25342
rect 48188 24882 48244 24892
rect 48188 24612 48244 24622
rect 48188 24518 48244 24556
rect 48076 23940 48132 23950
rect 47740 23938 48132 23940
rect 47740 23886 47742 23938
rect 47794 23886 48078 23938
rect 48130 23886 48132 23938
rect 47740 23884 48132 23886
rect 46956 19966 46958 20018
rect 47010 19966 47012 20018
rect 46732 19294 46734 19346
rect 46786 19294 46788 19346
rect 46732 19282 46788 19294
rect 46620 19012 46676 19022
rect 46396 19010 46676 19012
rect 46396 18958 46622 19010
rect 46674 18958 46676 19010
rect 46396 18956 46676 18958
rect 46284 18338 46340 18350
rect 46284 18286 46286 18338
rect 46338 18286 46340 18338
rect 46284 18116 46340 18286
rect 46508 18228 46564 18238
rect 46620 18228 46676 18956
rect 46844 19012 46900 19022
rect 46844 18918 46900 18956
rect 46508 18226 46676 18228
rect 46508 18174 46510 18226
rect 46562 18174 46676 18226
rect 46508 18172 46676 18174
rect 46732 18450 46788 18462
rect 46732 18398 46734 18450
rect 46786 18398 46788 18450
rect 46508 18162 46564 18172
rect 46732 18116 46788 18398
rect 46340 18060 46452 18116
rect 46284 18050 46340 18060
rect 46396 17332 46452 18060
rect 46732 18050 46788 18060
rect 46844 18228 46900 18238
rect 46620 17668 46676 17678
rect 46620 17574 46676 17612
rect 46172 16930 46228 16940
rect 46284 17276 46452 17332
rect 46732 17442 46788 17454
rect 46732 17390 46734 17442
rect 46786 17390 46788 17442
rect 45948 14802 46004 14812
rect 46284 14644 46340 17276
rect 46732 17108 46788 17390
rect 46732 17042 46788 17052
rect 46844 16660 46900 18172
rect 46956 17668 47012 19966
rect 46956 17574 47012 17612
rect 47068 20188 47348 20244
rect 47068 19012 47124 20188
rect 47180 20020 47236 20030
rect 47180 19926 47236 19964
rect 47740 19460 47796 23884
rect 48076 23874 48132 23884
rect 48188 23044 48244 23054
rect 48188 22950 48244 22988
rect 47964 22932 48020 22942
rect 47964 22594 48020 22876
rect 47964 22542 47966 22594
rect 48018 22542 48020 22594
rect 47964 22530 48020 22542
rect 47964 21362 48020 21374
rect 47964 21310 47966 21362
rect 48018 21310 48020 21362
rect 47964 20244 48020 21310
rect 48188 20916 48244 20926
rect 48188 20822 48244 20860
rect 47964 20178 48020 20188
rect 48076 20804 48132 20814
rect 47852 20130 47908 20142
rect 47852 20078 47854 20130
rect 47906 20078 47908 20130
rect 47852 19908 47908 20078
rect 47852 19842 47908 19852
rect 48076 20018 48132 20748
rect 48076 19966 48078 20018
rect 48130 19966 48132 20018
rect 48076 19684 48132 19966
rect 48076 19618 48132 19628
rect 47404 19404 47796 19460
rect 47292 19236 47348 19246
rect 47404 19236 47460 19404
rect 47292 19234 47460 19236
rect 47292 19182 47294 19234
rect 47346 19182 47460 19234
rect 47292 19180 47460 19182
rect 47292 19170 47348 19180
rect 47068 18562 47124 18956
rect 47068 18510 47070 18562
rect 47122 18510 47124 18562
rect 46396 16604 46900 16660
rect 46396 15538 46452 16604
rect 46396 15486 46398 15538
rect 46450 15486 46452 15538
rect 46396 15474 46452 15486
rect 46620 16436 46676 16446
rect 45388 14018 45444 14028
rect 45500 14588 46340 14644
rect 44380 13972 44436 13982
rect 44380 13878 44436 13916
rect 45500 13970 45556 14588
rect 46284 14530 46340 14588
rect 46284 14478 46286 14530
rect 46338 14478 46340 14530
rect 46284 14466 46340 14478
rect 45724 14420 45780 14430
rect 45724 14326 45780 14364
rect 45500 13918 45502 13970
rect 45554 13918 45556 13970
rect 45500 13906 45556 13918
rect 45836 14306 45892 14318
rect 45836 14254 45838 14306
rect 45890 14254 45892 14306
rect 44604 13860 44660 13870
rect 44492 13804 44604 13860
rect 44268 13076 44324 13086
rect 44156 13074 44324 13076
rect 44156 13022 44270 13074
rect 44322 13022 44324 13074
rect 44156 13020 44324 13022
rect 44268 13010 44324 13020
rect 44492 12516 44548 13804
rect 44604 13794 44660 13804
rect 44716 13636 44772 13646
rect 44268 12460 44548 12516
rect 44604 13634 44772 13636
rect 44604 13582 44718 13634
rect 44770 13582 44772 13634
rect 44604 13580 44772 13582
rect 44604 12964 44660 13580
rect 44716 13570 44772 13580
rect 45276 13636 45332 13646
rect 45052 12964 45108 12974
rect 44604 12962 45108 12964
rect 44604 12910 45054 12962
rect 45106 12910 45108 12962
rect 44604 12908 45108 12910
rect 44156 12292 44212 12302
rect 44156 11506 44212 12236
rect 44268 12290 44324 12460
rect 44268 12238 44270 12290
rect 44322 12238 44324 12290
rect 44268 12226 44324 12238
rect 44380 12292 44436 12302
rect 44380 12198 44436 12236
rect 44156 11454 44158 11506
rect 44210 11454 44212 11506
rect 44156 11442 44212 11454
rect 43596 10670 43598 10722
rect 43650 10670 43652 10722
rect 43596 10658 43652 10670
rect 43708 11004 43876 11060
rect 43596 9940 43652 9950
rect 43708 9940 43764 11004
rect 43932 10948 43988 10958
rect 43820 10892 43932 10948
rect 43820 10722 43876 10892
rect 43932 10882 43988 10892
rect 44604 10836 44660 12908
rect 45052 12898 45108 12908
rect 44940 12404 44996 12414
rect 44940 12310 44996 12348
rect 45052 12292 45108 12302
rect 45052 12198 45108 12236
rect 45276 12290 45332 13580
rect 45836 13076 45892 14254
rect 45948 14308 46004 14318
rect 45948 14306 46452 14308
rect 45948 14254 45950 14306
rect 46002 14254 46452 14306
rect 45948 14252 46452 14254
rect 45948 14242 46004 14252
rect 45948 14084 46004 14094
rect 46004 14028 46116 14084
rect 45948 14018 46004 14028
rect 46060 13860 46116 14028
rect 46172 13860 46228 13870
rect 46060 13858 46228 13860
rect 46060 13806 46174 13858
rect 46226 13806 46228 13858
rect 46060 13804 46228 13806
rect 46172 13794 46228 13804
rect 45836 13010 45892 13020
rect 46060 13076 46116 13086
rect 45836 12850 45892 12862
rect 45836 12798 45838 12850
rect 45890 12798 45892 12850
rect 45836 12404 45892 12798
rect 45836 12338 45892 12348
rect 45276 12238 45278 12290
rect 45330 12238 45332 12290
rect 45276 12226 45332 12238
rect 44716 12178 44772 12190
rect 44716 12126 44718 12178
rect 44770 12126 44772 12178
rect 44716 10948 44772 12126
rect 46060 12178 46116 13020
rect 46284 12292 46340 14252
rect 46396 13970 46452 14252
rect 46396 13918 46398 13970
rect 46450 13918 46452 13970
rect 46396 13906 46452 13918
rect 46620 13970 46676 16380
rect 47068 15540 47124 18510
rect 47292 18450 47348 18462
rect 47292 18398 47294 18450
rect 47346 18398 47348 18450
rect 47180 18338 47236 18350
rect 47180 18286 47182 18338
rect 47234 18286 47236 18338
rect 47180 17666 47236 18286
rect 47292 18340 47348 18398
rect 47292 18274 47348 18284
rect 47404 18116 47460 19180
rect 47404 18050 47460 18060
rect 47516 19010 47572 19022
rect 47516 18958 47518 19010
rect 47570 18958 47572 19010
rect 47516 18452 47572 18958
rect 47180 17614 47182 17666
rect 47234 17614 47236 17666
rect 47180 17602 47236 17614
rect 47516 17220 47572 18396
rect 47852 19010 47908 19022
rect 47852 18958 47854 19010
rect 47906 18958 47908 19010
rect 47628 18340 47684 18350
rect 47628 18246 47684 18284
rect 47628 17668 47684 17678
rect 47852 17668 47908 18958
rect 47628 17554 47684 17612
rect 47628 17502 47630 17554
rect 47682 17502 47684 17554
rect 47628 17490 47684 17502
rect 47740 17666 47908 17668
rect 47740 17614 47854 17666
rect 47906 17614 47908 17666
rect 47740 17612 47908 17614
rect 47628 17220 47684 17230
rect 47516 17164 47628 17220
rect 47628 17154 47684 17164
rect 47516 15540 47572 15550
rect 47068 15538 47572 15540
rect 47068 15486 47518 15538
rect 47570 15486 47572 15538
rect 47068 15484 47572 15486
rect 47516 15474 47572 15484
rect 46956 15316 47012 15326
rect 46956 15222 47012 15260
rect 47068 15202 47124 15214
rect 47068 15150 47070 15202
rect 47122 15150 47124 15202
rect 47068 15148 47124 15150
rect 47740 15148 47796 17612
rect 47852 17602 47908 17612
rect 48076 18450 48132 18462
rect 48076 18398 48078 18450
rect 48130 18398 48132 18450
rect 47852 17220 47908 17230
rect 47852 15538 47908 17164
rect 47964 16658 48020 16670
rect 47964 16606 47966 16658
rect 48018 16606 48020 16658
rect 47964 16212 48020 16606
rect 47964 16146 48020 16156
rect 48076 16660 48132 18398
rect 48076 16210 48132 16604
rect 48076 16158 48078 16210
rect 48130 16158 48132 16210
rect 48076 16146 48132 16158
rect 48188 17556 48244 17566
rect 47852 15486 47854 15538
rect 47906 15486 47908 15538
rect 47852 15474 47908 15486
rect 47964 15988 48020 15998
rect 47964 15148 48020 15932
rect 48188 15148 48244 17500
rect 47068 15092 47460 15148
rect 47068 14420 47124 14430
rect 47068 14326 47124 14364
rect 46620 13918 46622 13970
rect 46674 13918 46676 13970
rect 46508 13636 46564 13646
rect 46508 13542 46564 13580
rect 46620 13076 46676 13918
rect 46844 14306 46900 14318
rect 46844 14254 46846 14306
rect 46898 14254 46900 14306
rect 46844 13748 46900 14254
rect 47404 14306 47460 15092
rect 47404 14254 47406 14306
rect 47458 14254 47460 14306
rect 46844 13682 46900 13692
rect 46956 14084 47012 14094
rect 46956 13746 47012 14028
rect 46956 13694 46958 13746
rect 47010 13694 47012 13746
rect 46956 13682 47012 13694
rect 46620 13010 46676 13020
rect 46060 12126 46062 12178
rect 46114 12126 46116 12178
rect 46060 12114 46116 12126
rect 46172 12236 46340 12292
rect 46060 11394 46116 11406
rect 46060 11342 46062 11394
rect 46114 11342 46116 11394
rect 44772 10892 45108 10948
rect 44716 10882 44772 10892
rect 43820 10670 43822 10722
rect 43874 10670 43876 10722
rect 43820 10658 43876 10670
rect 44156 10780 44660 10836
rect 44044 10500 44100 10510
rect 44044 10406 44100 10444
rect 43596 9938 43988 9940
rect 43596 9886 43598 9938
rect 43650 9886 43988 9938
rect 43596 9884 43988 9886
rect 43596 9874 43652 9884
rect 43148 9774 43150 9826
rect 43202 9774 43204 9826
rect 42588 9604 42644 9614
rect 42028 9548 42588 9604
rect 41356 9268 41412 9278
rect 42028 9268 42084 9548
rect 42588 9510 42644 9548
rect 41244 9266 42084 9268
rect 41244 9214 41358 9266
rect 41410 9214 42084 9266
rect 41244 9212 42084 9214
rect 38220 8932 38276 8942
rect 38220 8370 38276 8876
rect 38332 8932 38388 8942
rect 38332 8930 38500 8932
rect 38332 8878 38334 8930
rect 38386 8878 38500 8930
rect 38332 8876 38500 8878
rect 38332 8866 38388 8876
rect 38220 8318 38222 8370
rect 38274 8318 38276 8370
rect 38220 8306 38276 8318
rect 38332 7700 38388 7710
rect 38220 7476 38276 7486
rect 37548 7474 37716 7476
rect 37548 7422 37550 7474
rect 37602 7422 37716 7474
rect 37548 7420 37716 7422
rect 38108 7420 38220 7476
rect 37548 7410 37604 7420
rect 36316 6962 36372 6972
rect 37548 7028 37604 7038
rect 36540 6916 36596 6926
rect 36540 6690 36596 6860
rect 36540 6638 36542 6690
rect 36594 6638 36596 6690
rect 36540 6626 36596 6638
rect 37548 6578 37604 6972
rect 37548 6526 37550 6578
rect 37602 6526 37604 6578
rect 37548 6514 37604 6526
rect 37660 6468 37716 7420
rect 38220 7410 38276 7420
rect 38332 7364 38388 7644
rect 38444 7588 38500 8876
rect 41132 8260 41188 8270
rect 41244 8260 41300 9212
rect 41356 9202 41412 9212
rect 41580 8370 41636 9212
rect 41692 9042 41748 9212
rect 41692 8990 41694 9042
rect 41746 8990 41748 9042
rect 41692 8978 41748 8990
rect 42476 8930 42532 8942
rect 42476 8878 42478 8930
rect 42530 8878 42532 8930
rect 41580 8318 41582 8370
rect 41634 8318 41636 8370
rect 41580 8306 41636 8318
rect 42028 8596 42084 8606
rect 42028 8370 42084 8540
rect 42028 8318 42030 8370
rect 42082 8318 42084 8370
rect 42028 8306 42084 8318
rect 42476 8372 42532 8878
rect 43148 8932 43204 9774
rect 43148 8866 43204 8876
rect 43932 9828 43988 9884
rect 42588 8372 42644 8382
rect 42476 8370 42644 8372
rect 42476 8318 42590 8370
rect 42642 8318 42644 8370
rect 42476 8316 42644 8318
rect 42588 8306 42644 8316
rect 41020 8258 41300 8260
rect 41020 8206 41134 8258
rect 41186 8206 41300 8258
rect 41020 8204 41300 8206
rect 42140 8260 42196 8270
rect 42364 8260 42420 8270
rect 42140 8258 42420 8260
rect 42140 8206 42142 8258
rect 42194 8206 42366 8258
rect 42418 8206 42420 8258
rect 42140 8204 42420 8206
rect 39004 8148 39060 8158
rect 38892 7700 38948 7710
rect 38892 7606 38948 7644
rect 38668 7588 38724 7598
rect 38444 7586 38724 7588
rect 38444 7534 38670 7586
rect 38722 7534 38724 7586
rect 38444 7532 38724 7534
rect 38668 7522 38724 7532
rect 38444 7364 38500 7374
rect 38332 7362 38500 7364
rect 38332 7310 38446 7362
rect 38498 7310 38500 7362
rect 38332 7308 38500 7310
rect 38444 7298 38500 7308
rect 39004 7362 39060 8092
rect 40348 8148 40404 8158
rect 40348 8054 40404 8092
rect 39004 7310 39006 7362
rect 39058 7310 39060 7362
rect 39004 7298 39060 7310
rect 37884 6468 37940 6478
rect 37660 6466 37940 6468
rect 37660 6414 37886 6466
rect 37938 6414 37940 6466
rect 37660 6412 37940 6414
rect 36204 6066 36260 6076
rect 35644 5854 35646 5906
rect 35698 5854 35700 5906
rect 35644 5842 35700 5854
rect 36316 5796 36372 5806
rect 37884 5796 37940 6412
rect 38892 6132 38948 6142
rect 38892 6038 38948 6076
rect 40348 6132 40404 6142
rect 40348 6038 40404 6076
rect 41020 6132 41076 8204
rect 41132 8194 41188 8204
rect 42140 8194 42196 8204
rect 42364 8194 42420 8204
rect 42812 8260 42868 8270
rect 43260 8260 43316 8270
rect 42812 8166 42868 8204
rect 43148 8258 43316 8260
rect 43148 8206 43262 8258
rect 43314 8206 43316 8258
rect 43148 8204 43316 8206
rect 43036 8148 43092 8158
rect 43036 8054 43092 8092
rect 42140 8036 42196 8046
rect 41580 6692 41636 6702
rect 41804 6692 41860 6702
rect 41580 6690 41860 6692
rect 41580 6638 41582 6690
rect 41634 6638 41806 6690
rect 41858 6638 41860 6690
rect 41580 6636 41860 6638
rect 41580 6626 41636 6636
rect 41804 6626 41860 6636
rect 42140 6690 42196 7980
rect 42924 7924 42980 7934
rect 42924 7698 42980 7868
rect 42924 7646 42926 7698
rect 42978 7646 42980 7698
rect 42924 7634 42980 7646
rect 43148 7586 43204 8204
rect 43260 8194 43316 8204
rect 43932 8258 43988 9772
rect 44156 9604 44212 10780
rect 44268 10612 44324 10622
rect 44268 10610 44436 10612
rect 44268 10558 44270 10610
rect 44322 10558 44436 10610
rect 44268 10556 44436 10558
rect 44268 10546 44324 10556
rect 44380 10052 44436 10556
rect 44492 10610 44548 10780
rect 44492 10558 44494 10610
rect 44546 10558 44548 10610
rect 44492 10546 44548 10558
rect 44940 10724 44996 10734
rect 44828 10052 44884 10062
rect 44380 10050 44884 10052
rect 44380 9998 44830 10050
rect 44882 9998 44884 10050
rect 44380 9996 44884 9998
rect 44828 9986 44884 9996
rect 44940 9938 44996 10668
rect 44940 9886 44942 9938
rect 44994 9886 44996 9938
rect 44940 9874 44996 9886
rect 44156 9510 44212 9548
rect 44604 8932 44660 8942
rect 44604 8838 44660 8876
rect 43932 8206 43934 8258
rect 43986 8206 43988 8258
rect 43932 8194 43988 8206
rect 45052 8260 45108 10892
rect 45276 10610 45332 10622
rect 45276 10558 45278 10610
rect 45330 10558 45332 10610
rect 45164 10500 45220 10510
rect 45276 10500 45332 10558
rect 45220 10444 45332 10500
rect 46060 10500 46116 11342
rect 45164 10434 45220 10444
rect 46060 10434 46116 10444
rect 45612 9828 45668 9838
rect 45612 9734 45668 9772
rect 43820 8148 43876 8158
rect 45052 8148 45108 8204
rect 45388 8260 45444 8270
rect 45836 8260 45892 8270
rect 45388 8258 45836 8260
rect 45388 8206 45390 8258
rect 45442 8206 45836 8258
rect 45388 8204 45836 8206
rect 45164 8148 45220 8158
rect 45052 8146 45220 8148
rect 45052 8094 45166 8146
rect 45218 8094 45220 8146
rect 45052 8092 45220 8094
rect 43820 8054 43876 8092
rect 45164 8082 45220 8092
rect 43708 8036 43764 8046
rect 43708 7942 43764 7980
rect 43148 7534 43150 7586
rect 43202 7534 43204 7586
rect 42700 7476 42756 7486
rect 42700 7382 42756 7420
rect 42812 7362 42868 7374
rect 42812 7310 42814 7362
rect 42866 7310 42868 7362
rect 42140 6638 42142 6690
rect 42194 6638 42196 6690
rect 42140 6626 42196 6638
rect 42476 6692 42532 6702
rect 42812 6692 42868 7310
rect 43148 6916 43204 7534
rect 43596 7586 43652 7598
rect 43596 7534 43598 7586
rect 43650 7534 43652 7586
rect 43596 7476 43652 7534
rect 43596 7410 43652 7420
rect 43932 7474 43988 7486
rect 43932 7422 43934 7474
rect 43986 7422 43988 7474
rect 43148 6850 43204 6860
rect 43932 6692 43988 7422
rect 42476 6690 42868 6692
rect 42476 6638 42478 6690
rect 42530 6638 42868 6690
rect 42476 6636 42868 6638
rect 43820 6636 43932 6692
rect 42476 6626 42532 6636
rect 41020 5906 41076 6076
rect 41020 5854 41022 5906
rect 41074 5854 41076 5906
rect 41020 5842 41076 5854
rect 41468 6578 41524 6590
rect 41468 6526 41470 6578
rect 41522 6526 41524 6578
rect 38444 5796 38500 5806
rect 37884 5794 38500 5796
rect 37884 5742 38446 5794
rect 38498 5742 38500 5794
rect 37884 5740 38500 5742
rect 36316 5702 36372 5740
rect 35532 4498 35588 4508
rect 36652 5012 36708 5022
rect 34524 4398 34526 4450
rect 34578 4398 34580 4450
rect 34524 4386 34580 4398
rect 33740 4286 33742 4338
rect 33794 4286 33796 4338
rect 33740 4274 33796 4286
rect 35644 4340 35700 4350
rect 33292 4228 33348 4238
rect 33292 4134 33348 4172
rect 35084 4228 35140 4238
rect 34300 3668 34356 3678
rect 33628 3556 33684 3566
rect 33628 800 33684 3500
rect 33740 3444 33796 3482
rect 33740 3378 33796 3388
rect 34300 800 34356 3612
rect 35084 3442 35140 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35420 3556 35476 3566
rect 35420 3462 35476 3500
rect 35084 3390 35086 3442
rect 35138 3390 35140 3442
rect 35084 3378 35140 3390
rect 35644 800 35700 4284
rect 36652 4228 36708 4956
rect 37212 4900 37268 4910
rect 37212 4898 37380 4900
rect 37212 4846 37214 4898
rect 37266 4846 37380 4898
rect 37212 4844 37380 4846
rect 37212 4834 37268 4844
rect 37212 4564 37268 4574
rect 37212 4470 37268 4508
rect 37324 4340 37380 4844
rect 37436 4340 37492 4350
rect 37324 4284 37436 4340
rect 37436 4246 37492 4284
rect 36428 4226 36708 4228
rect 36428 4174 36654 4226
rect 36706 4174 36708 4226
rect 36428 4172 36708 4174
rect 36428 3554 36484 4172
rect 36652 4162 36708 4172
rect 37996 4226 38052 4238
rect 37996 4174 37998 4226
rect 38050 4174 38052 4226
rect 36988 3668 37044 3678
rect 36988 3574 37044 3612
rect 37884 3668 37940 3678
rect 36428 3502 36430 3554
rect 36482 3502 36484 3554
rect 36428 3490 36484 3502
rect 37884 3388 37940 3612
rect 37996 3556 38052 4174
rect 37996 3490 38052 3500
rect 38444 3556 38500 5740
rect 41468 5012 41524 6526
rect 42028 6468 42084 6478
rect 41692 6466 42084 6468
rect 41692 6414 42030 6466
rect 42082 6414 42084 6466
rect 41692 6412 42084 6414
rect 41692 6018 41748 6412
rect 42028 6402 42084 6412
rect 41692 5966 41694 6018
rect 41746 5966 41748 6018
rect 41692 5954 41748 5966
rect 43820 5794 43876 6636
rect 43932 6626 43988 6636
rect 45388 6580 45444 8204
rect 45836 8166 45892 8204
rect 46172 8146 46228 12236
rect 47404 10500 47460 14254
rect 47404 10406 47460 10444
rect 47516 15092 47796 15148
rect 47852 15092 48020 15148
rect 48076 15092 48244 15148
rect 47516 13634 47572 15092
rect 47852 14418 47908 15092
rect 47852 14366 47854 14418
rect 47906 14366 47908 14418
rect 47852 14354 47908 14366
rect 48076 14530 48132 15092
rect 48076 14478 48078 14530
rect 48130 14478 48132 14530
rect 48076 13972 48132 14478
rect 48076 13906 48132 13916
rect 47852 13860 47908 13870
rect 47852 13766 47908 13804
rect 47516 13582 47518 13634
rect 47570 13582 47572 13634
rect 46620 8260 46676 8270
rect 46620 8166 46676 8204
rect 47068 8260 47124 8270
rect 47516 8260 47572 13582
rect 48188 13748 48244 13758
rect 47964 13076 48020 13086
rect 47964 12982 48020 13020
rect 47964 12852 48020 12862
rect 47964 12066 48020 12796
rect 48188 12180 48244 13692
rect 48188 12114 48244 12124
rect 47964 12014 47966 12066
rect 48018 12014 48020 12066
rect 47964 12002 48020 12014
rect 47964 11508 48020 11518
rect 47964 11414 48020 11452
rect 47628 10836 47684 10846
rect 47628 9266 47684 10780
rect 48188 10836 48244 10846
rect 47852 10724 47908 10734
rect 47852 10630 47908 10668
rect 48188 10722 48244 10780
rect 48188 10670 48190 10722
rect 48242 10670 48244 10722
rect 48188 10658 48244 10670
rect 47964 9938 48020 9950
rect 47964 9886 47966 9938
rect 48018 9886 48020 9938
rect 47964 9492 48020 9886
rect 47964 9426 48020 9436
rect 47628 9214 47630 9266
rect 47682 9214 47684 9266
rect 47628 9202 47684 9214
rect 47852 9154 47908 9166
rect 47852 9102 47854 9154
rect 47906 9102 47908 9154
rect 47852 8596 47908 9102
rect 48188 9042 48244 9054
rect 48188 8990 48190 9042
rect 48242 8990 48244 9042
rect 48188 8820 48244 8990
rect 48244 8764 48356 8820
rect 48188 8754 48244 8764
rect 47852 8530 47908 8540
rect 48300 8370 48356 8764
rect 48300 8318 48302 8370
rect 48354 8318 48356 8370
rect 48300 8306 48356 8318
rect 47124 8204 47572 8260
rect 47068 8166 47124 8204
rect 46172 8094 46174 8146
rect 46226 8094 46228 8146
rect 46172 8036 46228 8094
rect 46172 7970 46228 7980
rect 45612 6692 45668 6702
rect 45612 6598 45668 6636
rect 45388 6514 45444 6524
rect 47292 6578 47348 6590
rect 47292 6526 47294 6578
rect 47346 6526 47348 6578
rect 47292 6132 47348 6526
rect 47292 6066 47348 6076
rect 43820 5742 43822 5794
rect 43874 5742 43876 5794
rect 43820 5730 43876 5742
rect 41468 4946 41524 4956
rect 42700 5012 42756 5022
rect 41244 4450 41300 4462
rect 41244 4398 41246 4450
rect 41298 4398 41300 4450
rect 40796 3668 40852 3678
rect 40796 3574 40852 3612
rect 38444 3490 38500 3500
rect 39788 3556 39844 3566
rect 39788 3462 39844 3500
rect 41244 3388 41300 4398
rect 42476 4226 42532 4238
rect 42476 4174 42478 4226
rect 42530 4174 42532 4226
rect 37660 3332 37940 3388
rect 41020 3332 41300 3388
rect 41692 3444 41748 3454
rect 37660 800 37716 3332
rect 41020 800 41076 3332
rect 41692 800 41748 3388
rect 42476 3444 42532 4174
rect 42476 3378 42532 3388
rect 42700 3442 42756 4956
rect 42700 3390 42702 3442
rect 42754 3390 42756 3442
rect 42700 3378 42756 3390
rect 42924 3554 42980 3566
rect 42924 3502 42926 3554
rect 42978 3502 42980 3554
rect 42924 3444 42980 3502
rect 42924 3378 42980 3388
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 32928 0 33040 800
rect 33600 0 33712 800
rect 34272 0 34384 800
rect 35616 0 35728 800
rect 37632 0 37744 800
rect 40992 0 41104 800
rect 41664 0 41776 800
<< via2 >>
rect 44716 49756 44772 49812
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4172 45052 4228 45108
rect 1932 42364 1988 42420
rect 1708 40908 1764 40964
rect 2044 41692 2100 41748
rect 1932 40348 1988 40404
rect 1932 39676 1988 39732
rect 2492 39452 2548 39508
rect 2380 39004 2436 39060
rect 3164 39004 3220 39060
rect 4060 39340 4116 39396
rect 3724 39004 3780 39060
rect 2604 38892 2660 38948
rect 3612 38946 3668 38948
rect 3612 38894 3614 38946
rect 3614 38894 3666 38946
rect 3666 38894 3668 38946
rect 3612 38892 3668 38894
rect 2716 38834 2772 38836
rect 2716 38782 2718 38834
rect 2718 38782 2770 38834
rect 2770 38782 2772 38834
rect 2716 38780 2772 38782
rect 3948 38668 4004 38724
rect 1932 37042 1988 37044
rect 1932 36990 1934 37042
rect 1934 36990 1986 37042
rect 1986 36990 1988 37042
rect 1932 36988 1988 36990
rect 1932 36594 1988 36596
rect 1932 36542 1934 36594
rect 1934 36542 1986 36594
rect 1986 36542 1988 36594
rect 1932 36540 1988 36542
rect 1820 35532 1876 35588
rect 1708 34300 1764 34356
rect 2044 34412 2100 34468
rect 1932 33628 1988 33684
rect 1820 33346 1876 33348
rect 1820 33294 1822 33346
rect 1822 33294 1874 33346
rect 1874 33294 1876 33346
rect 1820 33292 1876 33294
rect 1820 27858 1876 27860
rect 1820 27806 1822 27858
rect 1822 27806 1874 27858
rect 1874 27806 1876 27858
rect 1820 27804 1876 27806
rect 2492 35698 2548 35700
rect 2492 35646 2494 35698
rect 2494 35646 2546 35698
rect 2546 35646 2548 35698
rect 2492 35644 2548 35646
rect 2492 34354 2548 34356
rect 2492 34302 2494 34354
rect 2494 34302 2546 34354
rect 2546 34302 2548 34354
rect 2492 34300 2548 34302
rect 2940 32786 2996 32788
rect 2940 32734 2942 32786
rect 2942 32734 2994 32786
rect 2994 32734 2996 32786
rect 2940 32732 2996 32734
rect 3164 36988 3220 37044
rect 3948 35308 4004 35364
rect 3948 33292 4004 33348
rect 3948 32396 4004 32452
rect 3612 32284 3668 32340
rect 2828 30716 2884 30772
rect 2828 29260 2884 29316
rect 3612 31890 3668 31892
rect 3612 31838 3614 31890
rect 3614 31838 3666 31890
rect 3666 31838 3668 31890
rect 3612 31836 3668 31838
rect 3388 30380 3444 30436
rect 3948 29932 4004 29988
rect 3276 29314 3332 29316
rect 3276 29262 3278 29314
rect 3278 29262 3330 29314
rect 3330 29262 3332 29314
rect 3276 29260 3332 29262
rect 2940 28754 2996 28756
rect 2940 28702 2942 28754
rect 2942 28702 2994 28754
rect 2994 28702 2996 28754
rect 2940 28700 2996 28702
rect 3052 28812 3108 28868
rect 3724 28812 3780 28868
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4844 43538 4900 43540
rect 4844 43486 4846 43538
rect 4846 43486 4898 43538
rect 4898 43486 4900 43538
rect 4844 43484 4900 43486
rect 8764 43484 8820 43540
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 8204 42028 8260 42084
rect 6188 41916 6244 41972
rect 4956 41746 5012 41748
rect 4956 41694 4958 41746
rect 4958 41694 5010 41746
rect 5010 41694 5012 41746
rect 4956 41692 5012 41694
rect 5292 41746 5348 41748
rect 5292 41694 5294 41746
rect 5294 41694 5346 41746
rect 5346 41694 5348 41746
rect 5292 41692 5348 41694
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4284 40684 4340 40740
rect 4284 40460 4340 40516
rect 5068 40962 5124 40964
rect 5068 40910 5070 40962
rect 5070 40910 5122 40962
rect 5122 40910 5124 40962
rect 5068 40908 5124 40910
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4396 39842 4452 39844
rect 4396 39790 4398 39842
rect 4398 39790 4450 39842
rect 4450 39790 4452 39842
rect 4396 39788 4452 39790
rect 4284 38946 4340 38948
rect 4284 38894 4286 38946
rect 4286 38894 4338 38946
rect 4338 38894 4340 38946
rect 4284 38892 4340 38894
rect 4620 38946 4676 38948
rect 4620 38894 4622 38946
rect 4622 38894 4674 38946
rect 4674 38894 4676 38946
rect 4620 38892 4676 38894
rect 4396 38834 4452 38836
rect 4396 38782 4398 38834
rect 4398 38782 4450 38834
rect 4450 38782 4452 38834
rect 4396 38780 4452 38782
rect 4844 38834 4900 38836
rect 4844 38782 4846 38834
rect 4846 38782 4898 38834
rect 4898 38782 4900 38834
rect 4844 38780 4900 38782
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4620 38162 4676 38164
rect 4620 38110 4622 38162
rect 4622 38110 4674 38162
rect 4674 38110 4676 38162
rect 4620 38108 4676 38110
rect 5068 40460 5124 40516
rect 5180 40348 5236 40404
rect 6300 41692 6356 41748
rect 5740 40626 5796 40628
rect 5740 40574 5742 40626
rect 5742 40574 5794 40626
rect 5794 40574 5796 40626
rect 5740 40572 5796 40574
rect 5292 39452 5348 39508
rect 5404 38892 5460 38948
rect 4956 37996 5012 38052
rect 4284 37266 4340 37268
rect 4284 37214 4286 37266
rect 4286 37214 4338 37266
rect 4338 37214 4340 37266
rect 4284 37212 4340 37214
rect 4284 36988 4340 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4844 36428 4900 36484
rect 4284 36204 4340 36260
rect 5180 38108 5236 38164
rect 5740 38108 5796 38164
rect 5516 37772 5572 37828
rect 5068 35420 5124 35476
rect 6076 40460 6132 40516
rect 7196 40572 7252 40628
rect 6860 40514 6916 40516
rect 6860 40462 6862 40514
rect 6862 40462 6914 40514
rect 6914 40462 6916 40514
rect 6860 40460 6916 40462
rect 6188 40402 6244 40404
rect 6188 40350 6190 40402
rect 6190 40350 6242 40402
rect 6242 40350 6244 40402
rect 6188 40348 6244 40350
rect 8540 40572 8596 40628
rect 6412 38834 6468 38836
rect 6412 38782 6414 38834
rect 6414 38782 6466 38834
rect 6466 38782 6468 38834
rect 6412 38780 6468 38782
rect 5628 36428 5684 36484
rect 5852 36482 5908 36484
rect 5852 36430 5854 36482
rect 5854 36430 5906 36482
rect 5906 36430 5908 36482
rect 5852 36428 5908 36430
rect 5516 35698 5572 35700
rect 5516 35646 5518 35698
rect 5518 35646 5570 35698
rect 5570 35646 5572 35698
rect 5516 35644 5572 35646
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4284 32956 4340 33012
rect 4956 32786 5012 32788
rect 4956 32734 4958 32786
rect 4958 32734 5010 32786
rect 5010 32734 5012 32786
rect 4956 32732 5012 32734
rect 4844 32620 4900 32676
rect 4732 32508 4788 32564
rect 4620 32450 4676 32452
rect 4620 32398 4622 32450
rect 4622 32398 4674 32450
rect 4674 32398 4676 32450
rect 4620 32396 4676 32398
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4844 31948 4900 32004
rect 4396 31836 4452 31892
rect 5292 32562 5348 32564
rect 5292 32510 5294 32562
rect 5294 32510 5346 32562
rect 5346 32510 5348 32562
rect 5292 32508 5348 32510
rect 5180 31836 5236 31892
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4620 30268 4676 30324
rect 4844 30380 4900 30436
rect 4284 29986 4340 29988
rect 4284 29934 4286 29986
rect 4286 29934 4338 29986
rect 4338 29934 4340 29986
rect 4284 29932 4340 29934
rect 5964 35420 6020 35476
rect 6412 38050 6468 38052
rect 6412 37998 6414 38050
rect 6414 37998 6466 38050
rect 6466 37998 6468 38050
rect 6412 37996 6468 37998
rect 6748 38108 6804 38164
rect 6636 37996 6692 38052
rect 6636 37826 6692 37828
rect 6636 37774 6638 37826
rect 6638 37774 6690 37826
rect 6690 37774 6692 37826
rect 6636 37772 6692 37774
rect 7084 36652 7140 36708
rect 7756 38892 7812 38948
rect 7420 38556 7476 38612
rect 7644 37884 7700 37940
rect 6188 35420 6244 35476
rect 6300 36258 6356 36260
rect 6300 36206 6302 36258
rect 6302 36206 6354 36258
rect 6354 36206 6356 36258
rect 6300 36204 6356 36206
rect 6860 34524 6916 34580
rect 5740 33346 5796 33348
rect 5740 33294 5742 33346
rect 5742 33294 5794 33346
rect 5794 33294 5796 33346
rect 5740 33292 5796 33294
rect 6300 33068 6356 33124
rect 5516 32732 5572 32788
rect 5852 32674 5908 32676
rect 5852 32622 5854 32674
rect 5854 32622 5906 32674
rect 5906 32622 5908 32674
rect 5852 32620 5908 32622
rect 5628 32284 5684 32340
rect 6524 32284 6580 32340
rect 5740 31836 5796 31892
rect 6412 31500 6468 31556
rect 5404 30492 5460 30548
rect 6188 30492 6244 30548
rect 5964 30380 6020 30436
rect 3948 28700 4004 28756
rect 4172 28642 4228 28644
rect 4172 28590 4174 28642
rect 4174 28590 4226 28642
rect 4226 28590 4228 28642
rect 4172 28588 4228 28590
rect 2380 27580 2436 27636
rect 2492 26012 2548 26068
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4844 28924 4900 28980
rect 4396 28700 4452 28756
rect 4732 28700 4788 28756
rect 4508 28588 4564 28644
rect 5740 28812 5796 28868
rect 6076 29036 6132 29092
rect 5852 28700 5908 28756
rect 5964 28812 6020 28868
rect 5740 28588 5796 28644
rect 5852 27858 5908 27860
rect 5852 27806 5854 27858
rect 5854 27806 5906 27858
rect 5906 27806 5908 27858
rect 5852 27804 5908 27806
rect 5628 27692 5684 27748
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 6300 30268 6356 30324
rect 4844 26290 4900 26292
rect 4844 26238 4846 26290
rect 4846 26238 4898 26290
rect 4898 26238 4900 26290
rect 4844 26236 4900 26238
rect 4732 26066 4788 26068
rect 4732 26014 4734 26066
rect 4734 26014 4786 26066
rect 4786 26014 4788 26066
rect 4732 26012 4788 26014
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 8204 38892 8260 38948
rect 7980 38834 8036 38836
rect 7980 38782 7982 38834
rect 7982 38782 8034 38834
rect 8034 38782 8036 38834
rect 7980 38780 8036 38782
rect 7868 38722 7924 38724
rect 7868 38670 7870 38722
rect 7870 38670 7922 38722
rect 7922 38670 7924 38722
rect 7868 38668 7924 38670
rect 8316 38780 8372 38836
rect 8876 43372 8932 43428
rect 8988 42028 9044 42084
rect 8988 40572 9044 40628
rect 10332 43426 10388 43428
rect 10332 43374 10334 43426
rect 10334 43374 10386 43426
rect 10386 43374 10388 43426
rect 10332 43372 10388 43374
rect 10556 42140 10612 42196
rect 11900 43484 11956 43540
rect 11116 42082 11172 42084
rect 11116 42030 11118 42082
rect 11118 42030 11170 42082
rect 11170 42030 11172 42082
rect 11116 42028 11172 42030
rect 10108 40684 10164 40740
rect 9884 40402 9940 40404
rect 9884 40350 9886 40402
rect 9886 40350 9938 40402
rect 9938 40350 9940 40402
rect 9884 40348 9940 40350
rect 10668 40684 10724 40740
rect 10220 40626 10276 40628
rect 10220 40574 10222 40626
rect 10222 40574 10274 40626
rect 10274 40574 10276 40626
rect 10220 40572 10276 40574
rect 8988 38556 9044 38612
rect 8652 38050 8708 38052
rect 8652 37998 8654 38050
rect 8654 37998 8706 38050
rect 8706 37998 8708 38050
rect 8652 37996 8708 37998
rect 8988 36652 9044 36708
rect 7868 36482 7924 36484
rect 7868 36430 7870 36482
rect 7870 36430 7922 36482
rect 7922 36430 7924 36482
rect 7868 36428 7924 36430
rect 7532 36316 7588 36372
rect 8428 36370 8484 36372
rect 8428 36318 8430 36370
rect 8430 36318 8482 36370
rect 8482 36318 8484 36370
rect 8428 36316 8484 36318
rect 8652 36258 8708 36260
rect 8652 36206 8654 36258
rect 8654 36206 8706 36258
rect 8706 36206 8708 36258
rect 8652 36204 8708 36206
rect 7756 35308 7812 35364
rect 7420 34524 7476 34580
rect 8316 35644 8372 35700
rect 8540 35308 8596 35364
rect 8428 34524 8484 34580
rect 7420 33458 7476 33460
rect 7420 33406 7422 33458
rect 7422 33406 7474 33458
rect 7474 33406 7476 33458
rect 7420 33404 7476 33406
rect 7196 33180 7252 33236
rect 7308 33122 7364 33124
rect 7308 33070 7310 33122
rect 7310 33070 7362 33122
rect 7362 33070 7364 33122
rect 7308 33068 7364 33070
rect 8204 33234 8260 33236
rect 8204 33182 8206 33234
rect 8206 33182 8258 33234
rect 8258 33182 8260 33234
rect 8204 33180 8260 33182
rect 8428 33404 8484 33460
rect 7756 31836 7812 31892
rect 6636 30716 6692 30772
rect 7196 30380 7252 30436
rect 6636 29036 6692 29092
rect 10108 39340 10164 39396
rect 9548 38946 9604 38948
rect 9548 38894 9550 38946
rect 9550 38894 9602 38946
rect 9602 38894 9604 38946
rect 9548 38892 9604 38894
rect 9212 38668 9268 38724
rect 9660 38556 9716 38612
rect 9660 37884 9716 37940
rect 9660 37212 9716 37268
rect 8764 33516 8820 33572
rect 9212 33628 9268 33684
rect 8764 33346 8820 33348
rect 8764 33294 8766 33346
rect 8766 33294 8818 33346
rect 8818 33294 8820 33346
rect 8764 33292 8820 33294
rect 9212 33292 9268 33348
rect 8652 32562 8708 32564
rect 8652 32510 8654 32562
rect 8654 32510 8706 32562
rect 8706 32510 8708 32562
rect 8652 32508 8708 32510
rect 8428 31836 8484 31892
rect 8204 31052 8260 31108
rect 7532 30380 7588 30436
rect 7644 30268 7700 30324
rect 8092 29260 8148 29316
rect 6636 28140 6692 28196
rect 7644 28364 7700 28420
rect 5740 25452 5796 25508
rect 4620 25228 4676 25284
rect 4284 24668 4340 24724
rect 4172 24444 4228 24500
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 2044 23884 2100 23940
rect 1708 22876 1764 22932
rect 1708 22204 1764 22260
rect 5068 23938 5124 23940
rect 5068 23886 5070 23938
rect 5070 23886 5122 23938
rect 5122 23886 5124 23938
rect 5068 23884 5124 23886
rect 4620 23548 4676 23604
rect 5292 23548 5348 23604
rect 3612 23378 3668 23380
rect 3612 23326 3614 23378
rect 3614 23326 3666 23378
rect 3666 23326 3668 23378
rect 3612 23324 3668 23326
rect 2940 23100 2996 23156
rect 3164 23042 3220 23044
rect 3164 22990 3166 23042
rect 3166 22990 3218 23042
rect 3218 22990 3220 23042
rect 3164 22988 3220 22990
rect 2492 22876 2548 22932
rect 2044 21644 2100 21700
rect 2380 22204 2436 22260
rect 1932 21474 1988 21476
rect 1932 21422 1934 21474
rect 1934 21422 1986 21474
rect 1986 21422 1988 21474
rect 1932 21420 1988 21422
rect 2044 20972 2100 21028
rect 2492 21868 2548 21924
rect 3276 20860 3332 20916
rect 2828 19292 2884 19348
rect 4620 23042 4676 23044
rect 4620 22990 4622 23042
rect 4622 22990 4674 23042
rect 4674 22990 4676 23042
rect 4620 22988 4676 22990
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4620 22204 4676 22260
rect 5068 22146 5124 22148
rect 5068 22094 5070 22146
rect 5070 22094 5122 22146
rect 5122 22094 5124 22146
rect 5068 22092 5124 22094
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 4956 21308 5012 21364
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4620 21026 4676 21028
rect 4620 20974 4622 21026
rect 4622 20974 4674 21026
rect 4674 20974 4676 21026
rect 4620 20972 4676 20974
rect 3724 20076 3780 20132
rect 3612 19292 3668 19348
rect 4844 20076 4900 20132
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 7756 27804 7812 27860
rect 7756 27020 7812 27076
rect 6076 26236 6132 26292
rect 7084 26236 7140 26292
rect 6636 25452 6692 25508
rect 9100 32338 9156 32340
rect 9100 32286 9102 32338
rect 9102 32286 9154 32338
rect 9154 32286 9156 32338
rect 9100 32284 9156 32286
rect 9100 31554 9156 31556
rect 9100 31502 9102 31554
rect 9102 31502 9154 31554
rect 9154 31502 9156 31554
rect 9100 31500 9156 31502
rect 8764 31106 8820 31108
rect 8764 31054 8766 31106
rect 8766 31054 8818 31106
rect 8818 31054 8820 31106
rect 8764 31052 8820 31054
rect 8876 29372 8932 29428
rect 10556 39618 10612 39620
rect 10556 39566 10558 39618
rect 10558 39566 10610 39618
rect 10610 39566 10612 39618
rect 10556 39564 10612 39566
rect 11228 40514 11284 40516
rect 11228 40462 11230 40514
rect 11230 40462 11282 40514
rect 11282 40462 11284 40514
rect 11228 40460 11284 40462
rect 11004 40402 11060 40404
rect 11004 40350 11006 40402
rect 11006 40350 11058 40402
rect 11058 40350 11060 40402
rect 11004 40348 11060 40350
rect 11228 40012 11284 40068
rect 11004 39340 11060 39396
rect 11116 38834 11172 38836
rect 11116 38782 11118 38834
rect 11118 38782 11170 38834
rect 11170 38782 11172 38834
rect 11116 38780 11172 38782
rect 11900 42252 11956 42308
rect 11452 42140 11508 42196
rect 12572 45666 12628 45668
rect 12572 45614 12574 45666
rect 12574 45614 12626 45666
rect 12626 45614 12628 45666
rect 12572 45612 12628 45614
rect 13468 45612 13524 45668
rect 11676 40012 11732 40068
rect 11676 39618 11732 39620
rect 11676 39566 11678 39618
rect 11678 39566 11730 39618
rect 11730 39566 11732 39618
rect 11676 39564 11732 39566
rect 11452 39394 11508 39396
rect 11452 39342 11454 39394
rect 11454 39342 11506 39394
rect 11506 39342 11508 39394
rect 11452 39340 11508 39342
rect 11340 38668 11396 38724
rect 11452 38780 11508 38836
rect 10556 38108 10612 38164
rect 10220 37884 10276 37940
rect 10108 37212 10164 37268
rect 9772 35084 9828 35140
rect 10108 34300 10164 34356
rect 10444 36428 10500 36484
rect 10780 37212 10836 37268
rect 10892 36706 10948 36708
rect 10892 36654 10894 36706
rect 10894 36654 10946 36706
rect 10946 36654 10948 36706
rect 10892 36652 10948 36654
rect 10556 35084 10612 35140
rect 10332 34860 10388 34916
rect 9996 33628 10052 33684
rect 9884 33292 9940 33348
rect 9996 33068 10052 33124
rect 9884 32786 9940 32788
rect 9884 32734 9886 32786
rect 9886 32734 9938 32786
rect 9938 32734 9940 32786
rect 9884 32732 9940 32734
rect 9996 32620 10052 32676
rect 10556 34242 10612 34244
rect 10556 34190 10558 34242
rect 10558 34190 10610 34242
rect 10610 34190 10612 34242
rect 10556 34188 10612 34190
rect 11676 38668 11732 38724
rect 12460 38668 12516 38724
rect 11788 37378 11844 37380
rect 11788 37326 11790 37378
rect 11790 37326 11842 37378
rect 11842 37326 11844 37378
rect 11788 37324 11844 37326
rect 11564 36204 11620 36260
rect 10780 35138 10836 35140
rect 10780 35086 10782 35138
rect 10782 35086 10834 35138
rect 10834 35086 10836 35138
rect 10780 35084 10836 35086
rect 10892 34972 10948 35028
rect 10668 34076 10724 34132
rect 10780 34300 10836 34356
rect 11116 35868 11172 35924
rect 11452 35868 11508 35924
rect 11340 35698 11396 35700
rect 11340 35646 11342 35698
rect 11342 35646 11394 35698
rect 11394 35646 11396 35698
rect 11340 35644 11396 35646
rect 11788 35922 11844 35924
rect 11788 35870 11790 35922
rect 11790 35870 11842 35922
rect 11842 35870 11844 35922
rect 11788 35868 11844 35870
rect 12012 38162 12068 38164
rect 12012 38110 12014 38162
rect 12014 38110 12066 38162
rect 12066 38110 12068 38162
rect 12012 38108 12068 38110
rect 12908 39506 12964 39508
rect 12908 39454 12910 39506
rect 12910 39454 12962 39506
rect 12962 39454 12964 39506
rect 12908 39452 12964 39454
rect 13132 37490 13188 37492
rect 13132 37438 13134 37490
rect 13134 37438 13186 37490
rect 13186 37438 13188 37490
rect 13132 37436 13188 37438
rect 13020 37378 13076 37380
rect 13020 37326 13022 37378
rect 13022 37326 13074 37378
rect 13074 37326 13076 37378
rect 13020 37324 13076 37326
rect 13356 37266 13412 37268
rect 13356 37214 13358 37266
rect 13358 37214 13410 37266
rect 13410 37214 13412 37266
rect 13356 37212 13412 37214
rect 12908 36652 12964 36708
rect 14252 45052 14308 45108
rect 16156 46060 16212 46116
rect 14924 45052 14980 45108
rect 13804 42140 13860 42196
rect 14700 42140 14756 42196
rect 13580 41916 13636 41972
rect 13580 40012 13636 40068
rect 13580 39676 13636 39732
rect 13916 39506 13972 39508
rect 13916 39454 13918 39506
rect 13918 39454 13970 39506
rect 13970 39454 13972 39506
rect 13916 39452 13972 39454
rect 13804 39394 13860 39396
rect 13804 39342 13806 39394
rect 13806 39342 13858 39394
rect 13858 39342 13860 39394
rect 13804 39340 13860 39342
rect 14252 37378 14308 37380
rect 14252 37326 14254 37378
rect 14254 37326 14306 37378
rect 14306 37326 14308 37378
rect 14252 37324 14308 37326
rect 14140 37212 14196 37268
rect 14028 37100 14084 37156
rect 13692 36540 13748 36596
rect 11788 34914 11844 34916
rect 11788 34862 11790 34914
rect 11790 34862 11842 34914
rect 11842 34862 11844 34914
rect 11788 34860 11844 34862
rect 13244 35644 13300 35700
rect 11004 34524 11060 34580
rect 13020 34860 13076 34916
rect 12236 34690 12292 34692
rect 12236 34638 12238 34690
rect 12238 34638 12290 34690
rect 12290 34638 12292 34690
rect 12236 34636 12292 34638
rect 12908 34636 12964 34692
rect 12572 34188 12628 34244
rect 11228 33458 11284 33460
rect 11228 33406 11230 33458
rect 11230 33406 11282 33458
rect 11282 33406 11284 33458
rect 11228 33404 11284 33406
rect 12348 33404 12404 33460
rect 10444 33180 10500 33236
rect 10892 33122 10948 33124
rect 10892 33070 10894 33122
rect 10894 33070 10946 33122
rect 10946 33070 10948 33122
rect 10892 33068 10948 33070
rect 11004 32786 11060 32788
rect 11004 32734 11006 32786
rect 11006 32734 11058 32786
rect 11058 32734 11060 32786
rect 11004 32732 11060 32734
rect 10780 32674 10836 32676
rect 10780 32622 10782 32674
rect 10782 32622 10834 32674
rect 10834 32622 10836 32674
rect 10780 32620 10836 32622
rect 11116 32450 11172 32452
rect 11116 32398 11118 32450
rect 11118 32398 11170 32450
rect 11170 32398 11172 32450
rect 11116 32396 11172 32398
rect 11228 32284 11284 32340
rect 11116 31890 11172 31892
rect 11116 31838 11118 31890
rect 11118 31838 11170 31890
rect 11170 31838 11172 31890
rect 11116 31836 11172 31838
rect 10556 31778 10612 31780
rect 10556 31726 10558 31778
rect 10558 31726 10610 31778
rect 10610 31726 10612 31778
rect 10556 31724 10612 31726
rect 9436 29260 9492 29316
rect 9660 28924 9716 28980
rect 9772 28754 9828 28756
rect 9772 28702 9774 28754
rect 9774 28702 9826 28754
rect 9826 28702 9828 28754
rect 9772 28700 9828 28702
rect 9660 28642 9716 28644
rect 9660 28590 9662 28642
rect 9662 28590 9714 28642
rect 9714 28590 9716 28642
rect 9660 28588 9716 28590
rect 9884 28252 9940 28308
rect 9996 28588 10052 28644
rect 9772 27970 9828 27972
rect 9772 27918 9774 27970
rect 9774 27918 9826 27970
rect 9826 27918 9828 27970
rect 9772 27916 9828 27918
rect 8764 27746 8820 27748
rect 8764 27694 8766 27746
rect 8766 27694 8818 27746
rect 8818 27694 8820 27746
rect 8764 27692 8820 27694
rect 9548 27692 9604 27748
rect 9100 27186 9156 27188
rect 9100 27134 9102 27186
rect 9102 27134 9154 27186
rect 9154 27134 9156 27186
rect 9100 27132 9156 27134
rect 9884 27858 9940 27860
rect 9884 27806 9886 27858
rect 9886 27806 9938 27858
rect 9938 27806 9940 27858
rect 9884 27804 9940 27806
rect 10220 29426 10276 29428
rect 10220 29374 10222 29426
rect 10222 29374 10274 29426
rect 10274 29374 10276 29426
rect 10220 29372 10276 29374
rect 10444 29426 10500 29428
rect 10444 29374 10446 29426
rect 10446 29374 10498 29426
rect 10498 29374 10500 29426
rect 10444 29372 10500 29374
rect 11900 31724 11956 31780
rect 12908 33180 12964 33236
rect 12908 32956 12964 33012
rect 12460 31388 12516 31444
rect 12684 31612 12740 31668
rect 14588 37100 14644 37156
rect 14476 36988 14532 37044
rect 14140 36652 14196 36708
rect 14924 43596 14980 43652
rect 14924 42252 14980 42308
rect 14812 40348 14868 40404
rect 16268 45330 16324 45332
rect 16268 45278 16270 45330
rect 16270 45278 16322 45330
rect 16322 45278 16324 45330
rect 16268 45276 16324 45278
rect 15260 42252 15316 42308
rect 15484 42082 15540 42084
rect 15484 42030 15486 42082
rect 15486 42030 15538 42082
rect 15538 42030 15540 42082
rect 15484 42028 15540 42030
rect 15372 41970 15428 41972
rect 15372 41918 15374 41970
rect 15374 41918 15426 41970
rect 15426 41918 15428 41970
rect 15372 41916 15428 41918
rect 16268 41858 16324 41860
rect 16268 41806 16270 41858
rect 16270 41806 16322 41858
rect 16322 41806 16324 41858
rect 16268 41804 16324 41806
rect 14812 36482 14868 36484
rect 14812 36430 14814 36482
rect 14814 36430 14866 36482
rect 14866 36430 14868 36482
rect 14812 36428 14868 36430
rect 14924 37100 14980 37156
rect 17948 46114 18004 46116
rect 17948 46062 17950 46114
rect 17950 46062 18002 46114
rect 18002 46062 18004 46114
rect 17948 46060 18004 46062
rect 16828 45276 16884 45332
rect 17388 45106 17444 45108
rect 17388 45054 17390 45106
rect 17390 45054 17442 45106
rect 17442 45054 17444 45106
rect 17388 45052 17444 45054
rect 17052 44434 17108 44436
rect 17052 44382 17054 44434
rect 17054 44382 17106 44434
rect 17106 44382 17108 44434
rect 17052 44380 17108 44382
rect 17500 43650 17556 43652
rect 17500 43598 17502 43650
rect 17502 43598 17554 43650
rect 17554 43598 17556 43650
rect 17500 43596 17556 43598
rect 16716 43538 16772 43540
rect 16716 43486 16718 43538
rect 16718 43486 16770 43538
rect 16770 43486 16772 43538
rect 16716 43484 16772 43486
rect 16828 43426 16884 43428
rect 16828 43374 16830 43426
rect 16830 43374 16882 43426
rect 16882 43374 16884 43426
rect 16828 43372 16884 43374
rect 17612 43538 17668 43540
rect 17612 43486 17614 43538
rect 17614 43486 17666 43538
rect 17666 43486 17668 43538
rect 17612 43484 17668 43486
rect 17388 42812 17444 42868
rect 17724 43372 17780 43428
rect 17388 41692 17444 41748
rect 16380 40572 16436 40628
rect 17388 40572 17444 40628
rect 16044 40348 16100 40404
rect 17724 40290 17780 40292
rect 17724 40238 17726 40290
rect 17726 40238 17778 40290
rect 17778 40238 17780 40290
rect 17724 40236 17780 40238
rect 18844 45612 18900 45668
rect 18732 44156 18788 44212
rect 18508 44044 18564 44100
rect 18284 43426 18340 43428
rect 18284 43374 18286 43426
rect 18286 43374 18338 43426
rect 18338 43374 18340 43426
rect 18284 43372 18340 43374
rect 15932 39340 15988 39396
rect 18956 45276 19012 45332
rect 19852 45666 19908 45668
rect 19852 45614 19854 45666
rect 19854 45614 19906 45666
rect 19906 45614 19908 45666
rect 19852 45612 19908 45614
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 20524 45276 20580 45332
rect 19852 45164 19908 45220
rect 19516 44380 19572 44436
rect 19404 44210 19460 44212
rect 19404 44158 19406 44210
rect 19406 44158 19458 44210
rect 19458 44158 19460 44210
rect 19404 44156 19460 44158
rect 19516 43820 19572 43876
rect 19292 43484 19348 43540
rect 20188 45052 20244 45108
rect 20076 44322 20132 44324
rect 20076 44270 20078 44322
rect 20078 44270 20130 44322
rect 20130 44270 20132 44322
rect 20076 44268 20132 44270
rect 19852 44044 19908 44100
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19740 43708 19796 43764
rect 19628 43372 19684 43428
rect 19852 43314 19908 43316
rect 19852 43262 19854 43314
rect 19854 43262 19906 43314
rect 19906 43262 19908 43314
rect 19852 43260 19908 43262
rect 19516 42866 19572 42868
rect 19516 42814 19518 42866
rect 19518 42814 19570 42866
rect 19570 42814 19572 42866
rect 19516 42812 19572 42814
rect 20076 42754 20132 42756
rect 20076 42702 20078 42754
rect 20078 42702 20130 42754
rect 20130 42702 20132 42754
rect 20076 42700 20132 42702
rect 19516 42140 19572 42196
rect 18956 41298 19012 41300
rect 18956 41246 18958 41298
rect 18958 41246 19010 41298
rect 19010 41246 19012 41298
rect 18956 41244 19012 41246
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 20524 44322 20580 44324
rect 20524 44270 20526 44322
rect 20526 44270 20578 44322
rect 20578 44270 20580 44322
rect 20524 44268 20580 44270
rect 20188 42140 20244 42196
rect 19964 42028 20020 42084
rect 23548 46060 23604 46116
rect 20972 45276 21028 45332
rect 20748 45164 20804 45220
rect 20860 45052 20916 45108
rect 21420 43596 21476 43652
rect 20300 42028 20356 42084
rect 19628 41916 19684 41972
rect 20412 42700 20468 42756
rect 22764 45778 22820 45780
rect 22764 45726 22766 45778
rect 22766 45726 22818 45778
rect 22818 45726 22820 45778
rect 22764 45724 22820 45726
rect 23772 45724 23828 45780
rect 21644 43538 21700 43540
rect 21644 43486 21646 43538
rect 21646 43486 21698 43538
rect 21698 43486 21700 43538
rect 21644 43484 21700 43486
rect 25564 46114 25620 46116
rect 25564 46062 25566 46114
rect 25566 46062 25618 46114
rect 25618 46062 25620 46114
rect 25564 46060 25620 46062
rect 23436 44210 23492 44212
rect 23436 44158 23438 44210
rect 23438 44158 23490 44210
rect 23490 44158 23492 44210
rect 23436 44156 23492 44158
rect 24108 44156 24164 44212
rect 21868 43650 21924 43652
rect 21868 43598 21870 43650
rect 21870 43598 21922 43650
rect 21922 43598 21924 43650
rect 21868 43596 21924 43598
rect 21756 43260 21812 43316
rect 22092 43426 22148 43428
rect 22092 43374 22094 43426
rect 22094 43374 22146 43426
rect 22146 43374 22148 43426
rect 22092 43372 22148 43374
rect 21644 42140 21700 42196
rect 20636 41970 20692 41972
rect 20636 41918 20638 41970
rect 20638 41918 20690 41970
rect 20690 41918 20692 41970
rect 20636 41916 20692 41918
rect 19628 41244 19684 41300
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 18732 40290 18788 40292
rect 18732 40238 18734 40290
rect 18734 40238 18786 40290
rect 18786 40238 18788 40290
rect 18732 40236 18788 40238
rect 18060 39564 18116 39620
rect 18396 39676 18452 39732
rect 18172 39506 18228 39508
rect 18172 39454 18174 39506
rect 18174 39454 18226 39506
rect 18226 39454 18228 39506
rect 18172 39452 18228 39454
rect 18060 39394 18116 39396
rect 18060 39342 18062 39394
rect 18062 39342 18114 39394
rect 18114 39342 18116 39394
rect 18060 39340 18116 39342
rect 15708 37378 15764 37380
rect 15708 37326 15710 37378
rect 15710 37326 15762 37378
rect 15762 37326 15764 37378
rect 15708 37324 15764 37326
rect 19180 39618 19236 39620
rect 19180 39566 19182 39618
rect 19182 39566 19234 39618
rect 19234 39566 19236 39618
rect 19180 39564 19236 39566
rect 15820 36988 15876 37044
rect 15372 36428 15428 36484
rect 13580 35532 13636 35588
rect 13468 35084 13524 35140
rect 15036 35196 15092 35252
rect 13692 34690 13748 34692
rect 13692 34638 13694 34690
rect 13694 34638 13746 34690
rect 13746 34638 13748 34690
rect 13692 34636 13748 34638
rect 13692 34130 13748 34132
rect 13692 34078 13694 34130
rect 13694 34078 13746 34130
rect 13746 34078 13748 34130
rect 13692 34076 13748 34078
rect 13692 33346 13748 33348
rect 13692 33294 13694 33346
rect 13694 33294 13746 33346
rect 13746 33294 13748 33346
rect 13692 33292 13748 33294
rect 12684 31052 12740 31108
rect 13692 32396 13748 32452
rect 13692 31778 13748 31780
rect 13692 31726 13694 31778
rect 13694 31726 13746 31778
rect 13746 31726 13748 31778
rect 13692 31724 13748 31726
rect 15932 36540 15988 36596
rect 16828 36316 16884 36372
rect 16156 35308 16212 35364
rect 15484 35196 15540 35252
rect 16044 34914 16100 34916
rect 16044 34862 16046 34914
rect 16046 34862 16098 34914
rect 16098 34862 16100 34914
rect 16044 34860 16100 34862
rect 15260 34748 15316 34804
rect 15148 34636 15204 34692
rect 14700 33404 14756 33460
rect 13916 33234 13972 33236
rect 13916 33182 13918 33234
rect 13918 33182 13970 33234
rect 13970 33182 13972 33234
rect 13916 33180 13972 33182
rect 14028 31836 14084 31892
rect 14364 31778 14420 31780
rect 14364 31726 14366 31778
rect 14366 31726 14418 31778
rect 14418 31726 14420 31778
rect 14364 31724 14420 31726
rect 13804 31612 13860 31668
rect 13916 31500 13972 31556
rect 13692 31276 13748 31332
rect 13804 31388 13860 31444
rect 12684 30380 12740 30436
rect 13468 30380 13524 30436
rect 10668 29314 10724 29316
rect 10668 29262 10670 29314
rect 10670 29262 10722 29314
rect 10722 29262 10724 29314
rect 10668 29260 10724 29262
rect 10220 28700 10276 28756
rect 10780 28252 10836 28308
rect 10444 27858 10500 27860
rect 10444 27806 10446 27858
rect 10446 27806 10498 27858
rect 10498 27806 10500 27858
rect 10444 27804 10500 27806
rect 10108 27074 10164 27076
rect 10108 27022 10110 27074
rect 10110 27022 10162 27074
rect 10162 27022 10164 27074
rect 10108 27020 10164 27022
rect 8092 26124 8148 26180
rect 8652 26178 8708 26180
rect 8652 26126 8654 26178
rect 8654 26126 8706 26178
rect 8706 26126 8708 26178
rect 8652 26124 8708 26126
rect 6300 25282 6356 25284
rect 6300 25230 6302 25282
rect 6302 25230 6354 25282
rect 6354 25230 6356 25282
rect 6300 25228 6356 25230
rect 5852 23938 5908 23940
rect 5852 23886 5854 23938
rect 5854 23886 5906 23938
rect 5906 23886 5908 23938
rect 5852 23884 5908 23886
rect 5740 23826 5796 23828
rect 5740 23774 5742 23826
rect 5742 23774 5794 23826
rect 5794 23774 5796 23826
rect 5740 23772 5796 23774
rect 9212 26962 9268 26964
rect 9212 26910 9214 26962
rect 9214 26910 9266 26962
rect 9266 26910 9268 26962
rect 9212 26908 9268 26910
rect 10780 27580 10836 27636
rect 11452 29372 11508 29428
rect 12572 29372 12628 29428
rect 11900 29314 11956 29316
rect 11900 29262 11902 29314
rect 11902 29262 11954 29314
rect 11954 29262 11956 29314
rect 11900 29260 11956 29262
rect 11676 28140 11732 28196
rect 11900 28140 11956 28196
rect 11228 27804 11284 27860
rect 11788 27692 11844 27748
rect 11676 27634 11732 27636
rect 11676 27582 11678 27634
rect 11678 27582 11730 27634
rect 11730 27582 11732 27634
rect 11676 27580 11732 27582
rect 11004 27132 11060 27188
rect 11116 27020 11172 27076
rect 8988 25452 9044 25508
rect 9548 26124 9604 26180
rect 6972 23938 7028 23940
rect 6972 23886 6974 23938
rect 6974 23886 7026 23938
rect 7026 23886 7028 23938
rect 6972 23884 7028 23886
rect 6748 23772 6804 23828
rect 6412 23548 6468 23604
rect 10332 23884 10388 23940
rect 8316 23826 8372 23828
rect 8316 23774 8318 23826
rect 8318 23774 8370 23826
rect 8370 23774 8372 23826
rect 8316 23772 8372 23774
rect 7196 23436 7252 23492
rect 8204 23436 8260 23492
rect 9324 23212 9380 23268
rect 6524 22930 6580 22932
rect 6524 22878 6526 22930
rect 6526 22878 6578 22930
rect 6578 22878 6580 22930
rect 6524 22876 6580 22878
rect 8540 22930 8596 22932
rect 8540 22878 8542 22930
rect 8542 22878 8594 22930
rect 8594 22878 8596 22930
rect 8540 22876 8596 22878
rect 6188 22258 6244 22260
rect 6188 22206 6190 22258
rect 6190 22206 6242 22258
rect 6242 22206 6244 22258
rect 6188 22204 6244 22206
rect 7196 22204 7252 22260
rect 5404 21362 5460 21364
rect 5404 21310 5406 21362
rect 5406 21310 5458 21362
rect 5458 21310 5460 21362
rect 5404 21308 5460 21310
rect 4956 19180 5012 19236
rect 1820 18396 1876 18452
rect 2828 18450 2884 18452
rect 2828 18398 2830 18450
rect 2830 18398 2882 18450
rect 2882 18398 2884 18450
rect 2828 18396 2884 18398
rect 5068 18396 5124 18452
rect 1932 18172 1988 18228
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 1932 17500 1988 17556
rect 2492 16770 2548 16772
rect 2492 16718 2494 16770
rect 2494 16718 2546 16770
rect 2546 16718 2548 16770
rect 2492 16716 2548 16718
rect 3388 16604 3444 16660
rect 2940 15820 2996 15876
rect 3276 15372 3332 15428
rect 5516 20860 5572 20916
rect 5740 20130 5796 20132
rect 5740 20078 5742 20130
rect 5742 20078 5794 20130
rect 5794 20078 5796 20130
rect 5740 20076 5796 20078
rect 5628 19964 5684 20020
rect 6748 21868 6804 21924
rect 8204 22092 8260 22148
rect 8428 22204 8484 22260
rect 6300 20636 6356 20692
rect 6524 21362 6580 21364
rect 6524 21310 6526 21362
rect 6526 21310 6578 21362
rect 6578 21310 6580 21362
rect 6524 21308 6580 21310
rect 6748 20972 6804 21028
rect 6188 20130 6244 20132
rect 6188 20078 6190 20130
rect 6190 20078 6242 20130
rect 6242 20078 6244 20130
rect 6188 20076 6244 20078
rect 6748 20130 6804 20132
rect 6748 20078 6750 20130
rect 6750 20078 6802 20130
rect 6802 20078 6804 20130
rect 6748 20076 6804 20078
rect 8428 21586 8484 21588
rect 8428 21534 8430 21586
rect 8430 21534 8482 21586
rect 8482 21534 8484 21586
rect 8428 21532 8484 21534
rect 7980 20860 8036 20916
rect 7532 20076 7588 20132
rect 5964 19964 6020 20020
rect 5628 19234 5684 19236
rect 5628 19182 5630 19234
rect 5630 19182 5682 19234
rect 5682 19182 5684 19234
rect 5628 19180 5684 19182
rect 5964 18844 6020 18900
rect 7532 19740 7588 19796
rect 8540 20690 8596 20692
rect 8540 20638 8542 20690
rect 8542 20638 8594 20690
rect 8594 20638 8596 20690
rect 8540 20636 8596 20638
rect 8876 22204 8932 22260
rect 8988 21420 9044 21476
rect 10220 22428 10276 22484
rect 10332 21810 10388 21812
rect 10332 21758 10334 21810
rect 10334 21758 10386 21810
rect 10386 21758 10388 21810
rect 10332 21756 10388 21758
rect 8652 20130 8708 20132
rect 8652 20078 8654 20130
rect 8654 20078 8706 20130
rect 8706 20078 8708 20130
rect 8652 20076 8708 20078
rect 8428 19852 8484 19908
rect 6524 19180 6580 19236
rect 8876 20018 8932 20020
rect 8876 19966 8878 20018
rect 8878 19966 8930 20018
rect 8930 19966 8932 20018
rect 8876 19964 8932 19966
rect 9100 19740 9156 19796
rect 9212 19458 9268 19460
rect 9212 19406 9214 19458
rect 9214 19406 9266 19458
rect 9266 19406 9268 19458
rect 9212 19404 9268 19406
rect 5516 18396 5572 18452
rect 5628 18338 5684 18340
rect 5628 18286 5630 18338
rect 5630 18286 5682 18338
rect 5682 18286 5684 18338
rect 5628 18284 5684 18286
rect 6188 18284 6244 18340
rect 4844 17388 4900 17444
rect 5740 17836 5796 17892
rect 4620 16828 4676 16884
rect 4060 16268 4116 16324
rect 2492 14364 2548 14420
rect 2492 12012 2548 12068
rect 1820 11394 1876 11396
rect 1820 11342 1822 11394
rect 1822 11342 1874 11394
rect 1874 11342 1876 11394
rect 1820 11340 1876 11342
rect 4172 15708 4228 15764
rect 3836 15426 3892 15428
rect 3836 15374 3838 15426
rect 3838 15374 3890 15426
rect 3890 15374 3892 15426
rect 3836 15372 3892 15374
rect 3948 14924 4004 14980
rect 3612 14418 3668 14420
rect 3612 14366 3614 14418
rect 3614 14366 3666 14418
rect 3666 14366 3668 14418
rect 3612 14364 3668 14366
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 6188 17612 6244 17668
rect 6412 17724 6468 17780
rect 5852 17442 5908 17444
rect 5852 17390 5854 17442
rect 5854 17390 5906 17442
rect 5906 17390 5908 17442
rect 5852 17388 5908 17390
rect 5180 16828 5236 16884
rect 5068 16770 5124 16772
rect 5068 16718 5070 16770
rect 5070 16718 5122 16770
rect 5122 16718 5124 16770
rect 5068 16716 5124 16718
rect 4956 16658 5012 16660
rect 4956 16606 4958 16658
rect 4958 16606 5010 16658
rect 5010 16606 5012 16658
rect 4956 16604 5012 16606
rect 6972 18844 7028 18900
rect 7084 18674 7140 18676
rect 7084 18622 7086 18674
rect 7086 18622 7138 18674
rect 7138 18622 7140 18674
rect 7084 18620 7140 18622
rect 6972 18172 7028 18228
rect 6972 17666 7028 17668
rect 6972 17614 6974 17666
rect 6974 17614 7026 17666
rect 7026 17614 7028 17666
rect 6972 17612 7028 17614
rect 5180 16380 5236 16436
rect 5180 15426 5236 15428
rect 5180 15374 5182 15426
rect 5182 15374 5234 15426
rect 5234 15374 5236 15426
rect 5180 15372 5236 15374
rect 6412 16268 6468 16324
rect 6188 15986 6244 15988
rect 6188 15934 6190 15986
rect 6190 15934 6242 15986
rect 6242 15934 6244 15986
rect 6188 15932 6244 15934
rect 5292 15708 5348 15764
rect 5964 15820 6020 15876
rect 4396 15314 4452 15316
rect 4396 15262 4398 15314
rect 4398 15262 4450 15314
rect 4450 15262 4452 15314
rect 4396 15260 4452 15262
rect 6188 15708 6244 15764
rect 5516 15314 5572 15316
rect 5516 15262 5518 15314
rect 5518 15262 5570 15314
rect 5570 15262 5572 15314
rect 5516 15260 5572 15262
rect 4396 15036 4452 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 3724 13356 3780 13412
rect 3836 13692 3892 13748
rect 3948 12684 4004 12740
rect 3948 9212 4004 9268
rect 1708 8146 1764 8148
rect 1708 8094 1710 8146
rect 1710 8094 1762 8146
rect 1762 8094 1764 8146
rect 1708 8092 1764 8094
rect 2044 8146 2100 8148
rect 2044 8094 2046 8146
rect 2046 8094 2098 8146
rect 2098 8094 2100 8146
rect 2044 8092 2100 8094
rect 2492 8034 2548 8036
rect 2492 7982 2494 8034
rect 2494 7982 2546 8034
rect 2546 7982 2548 8034
rect 2492 7980 2548 7982
rect 5068 14530 5124 14532
rect 5068 14478 5070 14530
rect 5070 14478 5122 14530
rect 5122 14478 5124 14530
rect 5068 14476 5124 14478
rect 4956 14418 5012 14420
rect 4956 14366 4958 14418
rect 4958 14366 5010 14418
rect 5010 14366 5012 14418
rect 4956 14364 5012 14366
rect 4284 13692 4340 13748
rect 5628 14418 5684 14420
rect 5628 14366 5630 14418
rect 5630 14366 5682 14418
rect 5682 14366 5684 14418
rect 5628 14364 5684 14366
rect 6076 15372 6132 15428
rect 7308 18450 7364 18452
rect 7308 18398 7310 18450
rect 7310 18398 7362 18450
rect 7362 18398 7364 18450
rect 7308 18396 7364 18398
rect 7868 18450 7924 18452
rect 7868 18398 7870 18450
rect 7870 18398 7922 18450
rect 7922 18398 7924 18450
rect 7868 18396 7924 18398
rect 7196 17724 7252 17780
rect 6748 16044 6804 16100
rect 4508 13468 4564 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4732 12850 4788 12852
rect 4732 12798 4734 12850
rect 4734 12798 4786 12850
rect 4786 12798 4788 12850
rect 4732 12796 4788 12798
rect 4844 12124 4900 12180
rect 4732 12066 4788 12068
rect 4732 12014 4734 12066
rect 4734 12014 4786 12066
rect 4786 12014 4788 12066
rect 4732 12012 4788 12014
rect 4844 11900 4900 11956
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4732 11564 4788 11620
rect 6300 14364 6356 14420
rect 8652 18674 8708 18676
rect 8652 18622 8654 18674
rect 8654 18622 8706 18674
rect 8706 18622 8708 18674
rect 8652 18620 8708 18622
rect 9884 20130 9940 20132
rect 9884 20078 9886 20130
rect 9886 20078 9938 20130
rect 9938 20078 9940 20130
rect 9884 20076 9940 20078
rect 9660 19794 9716 19796
rect 9660 19742 9662 19794
rect 9662 19742 9714 19794
rect 9714 19742 9716 19794
rect 9660 19740 9716 19742
rect 9660 18732 9716 18788
rect 8428 18396 8484 18452
rect 8540 18172 8596 18228
rect 8876 18284 8932 18340
rect 7868 15820 7924 15876
rect 8204 16658 8260 16660
rect 8204 16606 8206 16658
rect 8206 16606 8258 16658
rect 8258 16606 8260 16658
rect 8204 16604 8260 16606
rect 7756 15426 7812 15428
rect 7756 15374 7758 15426
rect 7758 15374 7810 15426
rect 7810 15374 7812 15426
rect 7756 15372 7812 15374
rect 7196 15036 7252 15092
rect 7084 14700 7140 14756
rect 7420 13970 7476 13972
rect 7420 13918 7422 13970
rect 7422 13918 7474 13970
rect 7474 13918 7476 13970
rect 7420 13916 7476 13918
rect 6748 13692 6804 13748
rect 5292 12796 5348 12852
rect 5292 11788 5348 11844
rect 5740 12124 5796 12180
rect 5068 11340 5124 11396
rect 4284 10444 4340 10500
rect 5068 10444 5124 10500
rect 6636 13356 6692 13412
rect 5964 12684 6020 12740
rect 6412 12236 6468 12292
rect 6636 12348 6692 12404
rect 6524 12012 6580 12068
rect 6748 11954 6804 11956
rect 6748 11902 6750 11954
rect 6750 11902 6802 11954
rect 6802 11902 6804 11954
rect 6748 11900 6804 11902
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 7196 13804 7252 13860
rect 7756 13804 7812 13860
rect 7308 13746 7364 13748
rect 7308 13694 7310 13746
rect 7310 13694 7362 13746
rect 7362 13694 7364 13746
rect 7308 13692 7364 13694
rect 7532 13746 7588 13748
rect 7532 13694 7534 13746
rect 7534 13694 7586 13746
rect 7586 13694 7588 13746
rect 7532 13692 7588 13694
rect 7420 12012 7476 12068
rect 8204 16210 8260 16212
rect 8204 16158 8206 16210
rect 8206 16158 8258 16210
rect 8258 16158 8260 16210
rect 8204 16156 8260 16158
rect 8092 16098 8148 16100
rect 8092 16046 8094 16098
rect 8094 16046 8146 16098
rect 8146 16046 8148 16098
rect 8092 16044 8148 16046
rect 8428 15708 8484 15764
rect 8764 16098 8820 16100
rect 8764 16046 8766 16098
rect 8766 16046 8818 16098
rect 8818 16046 8820 16098
rect 8764 16044 8820 16046
rect 8204 15372 8260 15428
rect 9660 15708 9716 15764
rect 9100 15372 9156 15428
rect 8428 15260 8484 15316
rect 7980 13692 8036 13748
rect 8204 15036 8260 15092
rect 8316 13746 8372 13748
rect 8316 13694 8318 13746
rect 8318 13694 8370 13746
rect 8370 13694 8372 13746
rect 8316 13692 8372 13694
rect 8204 13580 8260 13636
rect 7756 12402 7812 12404
rect 7756 12350 7758 12402
rect 7758 12350 7810 12402
rect 7810 12350 7812 12402
rect 7756 12348 7812 12350
rect 8988 15314 9044 15316
rect 8988 15262 8990 15314
rect 8990 15262 9042 15314
rect 9042 15262 9044 15314
rect 8988 15260 9044 15262
rect 9772 15260 9828 15316
rect 10332 20018 10388 20020
rect 10332 19966 10334 20018
rect 10334 19966 10386 20018
rect 10386 19966 10388 20018
rect 10332 19964 10388 19966
rect 10556 25116 10612 25172
rect 11788 26908 11844 26964
rect 11340 25900 11396 25956
rect 11564 25506 11620 25508
rect 11564 25454 11566 25506
rect 11566 25454 11618 25506
rect 11618 25454 11620 25506
rect 11564 25452 11620 25454
rect 12348 28812 12404 28868
rect 13580 29820 13636 29876
rect 13804 30828 13860 30884
rect 13804 30268 13860 30324
rect 14476 31500 14532 31556
rect 14588 31164 14644 31220
rect 14812 33292 14868 33348
rect 14924 32956 14980 33012
rect 14476 30882 14532 30884
rect 14476 30830 14478 30882
rect 14478 30830 14530 30882
rect 14530 30830 14532 30882
rect 14476 30828 14532 30830
rect 15036 31724 15092 31780
rect 14924 31612 14980 31668
rect 14252 30268 14308 30324
rect 13580 28866 13636 28868
rect 13580 28814 13582 28866
rect 13582 28814 13634 28866
rect 13634 28814 13636 28866
rect 13580 28812 13636 28814
rect 12460 27746 12516 27748
rect 12460 27694 12462 27746
rect 12462 27694 12514 27746
rect 12514 27694 12516 27746
rect 12460 27692 12516 27694
rect 13580 27020 13636 27076
rect 12908 26908 12964 26964
rect 12124 26124 12180 26180
rect 11900 25900 11956 25956
rect 11228 25116 11284 25172
rect 10556 23772 10612 23828
rect 10556 23042 10612 23044
rect 10556 22990 10558 23042
rect 10558 22990 10610 23042
rect 10610 22990 10612 23042
rect 10556 22988 10612 22990
rect 10556 22092 10612 22148
rect 10668 21586 10724 21588
rect 10668 21534 10670 21586
rect 10670 21534 10722 21586
rect 10722 21534 10724 21586
rect 10668 21532 10724 21534
rect 12012 23212 12068 23268
rect 11116 22482 11172 22484
rect 11116 22430 11118 22482
rect 11118 22430 11170 22482
rect 11170 22430 11172 22482
rect 11116 22428 11172 22430
rect 10892 21532 10948 21588
rect 11116 21532 11172 21588
rect 10668 19292 10724 19348
rect 10780 19180 10836 19236
rect 9996 18956 10052 19012
rect 9996 18450 10052 18452
rect 9996 18398 9998 18450
rect 9998 18398 10050 18450
rect 10050 18398 10052 18450
rect 9996 18396 10052 18398
rect 10332 18620 10388 18676
rect 10556 18956 10612 19012
rect 11004 19852 11060 19908
rect 11004 19458 11060 19460
rect 11004 19406 11006 19458
rect 11006 19406 11058 19458
rect 11058 19406 11060 19458
rect 11004 19404 11060 19406
rect 12348 22428 12404 22484
rect 12572 24444 12628 24500
rect 13692 26908 13748 26964
rect 13692 26684 13748 26740
rect 13468 25564 13524 25620
rect 11676 21756 11732 21812
rect 11676 21586 11732 21588
rect 11676 21534 11678 21586
rect 11678 21534 11730 21586
rect 11730 21534 11732 21586
rect 11676 21532 11732 21534
rect 11788 21420 11844 21476
rect 12572 21698 12628 21700
rect 12572 21646 12574 21698
rect 12574 21646 12626 21698
rect 12626 21646 12628 21698
rect 12572 21644 12628 21646
rect 12908 22258 12964 22260
rect 12908 22206 12910 22258
rect 12910 22206 12962 22258
rect 12962 22206 12964 22258
rect 12908 22204 12964 22206
rect 12684 21532 12740 21588
rect 12124 21196 12180 21252
rect 12908 20636 12964 20692
rect 12124 20018 12180 20020
rect 12124 19966 12126 20018
rect 12126 19966 12178 20018
rect 12178 19966 12180 20018
rect 12124 19964 12180 19966
rect 11004 18450 11060 18452
rect 11004 18398 11006 18450
rect 11006 18398 11058 18450
rect 11058 18398 11060 18450
rect 11004 18396 11060 18398
rect 10892 17666 10948 17668
rect 10892 17614 10894 17666
rect 10894 17614 10946 17666
rect 10946 17614 10948 17666
rect 10892 17612 10948 17614
rect 10220 16268 10276 16324
rect 9996 16044 10052 16100
rect 9996 15708 10052 15764
rect 10780 16770 10836 16772
rect 10780 16718 10782 16770
rect 10782 16718 10834 16770
rect 10834 16718 10836 16770
rect 10780 16716 10836 16718
rect 10892 16604 10948 16660
rect 10556 16156 10612 16212
rect 10444 16044 10500 16100
rect 10220 15932 10276 15988
rect 10220 15314 10276 15316
rect 10220 15262 10222 15314
rect 10222 15262 10274 15314
rect 10274 15262 10276 15314
rect 10220 15260 10276 15262
rect 8764 14530 8820 14532
rect 8764 14478 8766 14530
rect 8766 14478 8818 14530
rect 8818 14478 8820 14530
rect 8764 14476 8820 14478
rect 9324 14418 9380 14420
rect 9324 14366 9326 14418
rect 9326 14366 9378 14418
rect 9378 14366 9380 14418
rect 9324 14364 9380 14366
rect 9660 13916 9716 13972
rect 8652 13858 8708 13860
rect 8652 13806 8654 13858
rect 8654 13806 8706 13858
rect 8706 13806 8708 13858
rect 8652 13804 8708 13806
rect 9884 13858 9940 13860
rect 9884 13806 9886 13858
rect 9886 13806 9938 13858
rect 9938 13806 9940 13858
rect 9884 13804 9940 13806
rect 9548 13634 9604 13636
rect 9548 13582 9550 13634
rect 9550 13582 9602 13634
rect 9602 13582 9604 13634
rect 9548 13580 9604 13582
rect 9884 13468 9940 13524
rect 8540 13020 8596 13076
rect 9212 13132 9268 13188
rect 8876 12684 8932 12740
rect 8764 12572 8820 12628
rect 8652 12290 8708 12292
rect 8652 12238 8654 12290
rect 8654 12238 8706 12290
rect 8706 12238 8708 12290
rect 8652 12236 8708 12238
rect 8428 12012 8484 12068
rect 7532 10498 7588 10500
rect 7532 10446 7534 10498
rect 7534 10446 7586 10498
rect 7586 10446 7588 10498
rect 7532 10444 7588 10446
rect 7196 9266 7252 9268
rect 7196 9214 7198 9266
rect 7198 9214 7250 9266
rect 7250 9214 7252 9266
rect 7196 9212 7252 9214
rect 5740 8316 5796 8372
rect 6860 8146 6916 8148
rect 6860 8094 6862 8146
rect 6862 8094 6914 8146
rect 6914 8094 6916 8146
rect 6860 8092 6916 8094
rect 4172 7644 4228 7700
rect 6188 7980 6244 8036
rect 7532 9548 7588 9604
rect 9324 12572 9380 12628
rect 9772 12738 9828 12740
rect 9772 12686 9774 12738
rect 9774 12686 9826 12738
rect 9826 12686 9828 12738
rect 9772 12684 9828 12686
rect 7980 11340 8036 11396
rect 9212 11282 9268 11284
rect 9212 11230 9214 11282
rect 9214 11230 9266 11282
rect 9266 11230 9268 11282
rect 9212 11228 9268 11230
rect 9996 13132 10052 13188
rect 10108 13020 10164 13076
rect 10444 15036 10500 15092
rect 10332 14588 10388 14644
rect 11676 19122 11732 19124
rect 11676 19070 11678 19122
rect 11678 19070 11730 19122
rect 11730 19070 11732 19122
rect 11676 19068 11732 19070
rect 11340 19010 11396 19012
rect 11340 18958 11342 19010
rect 11342 18958 11394 19010
rect 11394 18958 11396 19010
rect 11340 18956 11396 18958
rect 11452 18732 11508 18788
rect 11228 16268 11284 16324
rect 11116 14754 11172 14756
rect 11116 14702 11118 14754
rect 11118 14702 11170 14754
rect 11170 14702 11172 14754
rect 11116 14700 11172 14702
rect 10668 14476 10724 14532
rect 10892 13916 10948 13972
rect 10556 13804 10612 13860
rect 10332 13746 10388 13748
rect 10332 13694 10334 13746
rect 10334 13694 10386 13746
rect 10386 13694 10388 13746
rect 10332 13692 10388 13694
rect 10668 13356 10724 13412
rect 10220 12796 10276 12852
rect 9772 12460 9828 12516
rect 9996 12348 10052 12404
rect 10108 11340 10164 11396
rect 10780 10668 10836 10724
rect 11116 11282 11172 11284
rect 11116 11230 11118 11282
rect 11118 11230 11170 11282
rect 11170 11230 11172 11282
rect 11116 11228 11172 11230
rect 10780 9772 10836 9828
rect 9660 9548 9716 9604
rect 7420 8034 7476 8036
rect 7420 7982 7422 8034
rect 7422 7982 7474 8034
rect 7474 7982 7476 8034
rect 7420 7980 7476 7982
rect 7308 7868 7364 7924
rect 7644 8258 7700 8260
rect 7644 8206 7646 8258
rect 7646 8206 7698 8258
rect 7698 8206 7700 8258
rect 7644 8204 7700 8206
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 6524 6412 6580 6468
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 7308 6466 7364 6468
rect 7308 6414 7310 6466
rect 7310 6414 7362 6466
rect 7362 6414 7364 6466
rect 7308 6412 7364 6414
rect 7532 6412 7588 6468
rect 7196 6076 7252 6132
rect 10556 9602 10612 9604
rect 10556 9550 10558 9602
rect 10558 9550 10610 9602
rect 10610 9550 10612 9602
rect 10556 9548 10612 9550
rect 10220 8258 10276 8260
rect 10220 8206 10222 8258
rect 10222 8206 10274 8258
rect 10274 8206 10276 8258
rect 10220 8204 10276 8206
rect 8428 8034 8484 8036
rect 8428 7982 8430 8034
rect 8430 7982 8482 8034
rect 8482 7982 8484 8034
rect 8428 7980 8484 7982
rect 8316 7868 8372 7924
rect 7756 6578 7812 6580
rect 7756 6526 7758 6578
rect 7758 6526 7810 6578
rect 7810 6526 7812 6578
rect 7756 6524 7812 6526
rect 7980 6412 8036 6468
rect 8652 7698 8708 7700
rect 8652 7646 8654 7698
rect 8654 7646 8706 7698
rect 8706 7646 8708 7698
rect 8652 7644 8708 7646
rect 8652 6748 8708 6804
rect 8204 6578 8260 6580
rect 8204 6526 8206 6578
rect 8206 6526 8258 6578
rect 8258 6526 8260 6578
rect 8204 6524 8260 6526
rect 8428 6300 8484 6356
rect 8428 6130 8484 6132
rect 8428 6078 8430 6130
rect 8430 6078 8482 6130
rect 8482 6078 8484 6130
rect 8428 6076 8484 6078
rect 8652 5740 8708 5796
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 6860 3554 6916 3556
rect 6860 3502 6862 3554
rect 6862 3502 6914 3554
rect 6914 3502 6916 3554
rect 6860 3500 6916 3502
rect 6412 3442 6468 3444
rect 6412 3390 6414 3442
rect 6414 3390 6466 3442
rect 6466 3390 6468 3442
rect 6412 3388 6468 3390
rect 7308 3388 7364 3444
rect 7980 4844 8036 4900
rect 7756 4226 7812 4228
rect 7756 4174 7758 4226
rect 7758 4174 7810 4226
rect 7810 4174 7812 4226
rect 7756 4172 7812 4174
rect 8428 3554 8484 3556
rect 8428 3502 8430 3554
rect 8430 3502 8482 3554
rect 8482 3502 8484 3554
rect 8428 3500 8484 3502
rect 9772 7980 9828 8036
rect 9100 6300 9156 6356
rect 11004 8034 11060 8036
rect 11004 7982 11006 8034
rect 11006 7982 11058 8034
rect 11058 7982 11060 8034
rect 11004 7980 11060 7982
rect 10108 6748 10164 6804
rect 9996 6300 10052 6356
rect 9548 6018 9604 6020
rect 9548 5966 9550 6018
rect 9550 5966 9602 6018
rect 9602 5966 9604 6018
rect 9548 5964 9604 5966
rect 9660 5794 9716 5796
rect 9660 5742 9662 5794
rect 9662 5742 9714 5794
rect 9714 5742 9716 5794
rect 9660 5740 9716 5742
rect 10892 6860 10948 6916
rect 12124 19346 12180 19348
rect 12124 19294 12126 19346
rect 12126 19294 12178 19346
rect 12178 19294 12180 19346
rect 12124 19292 12180 19294
rect 12236 19234 12292 19236
rect 12236 19182 12238 19234
rect 12238 19182 12290 19234
rect 12290 19182 12292 19234
rect 12236 19180 12292 19182
rect 11788 17388 11844 17444
rect 11900 18396 11956 18452
rect 11788 16604 11844 16660
rect 11676 15484 11732 15540
rect 11676 15314 11732 15316
rect 11676 15262 11678 15314
rect 11678 15262 11730 15314
rect 11730 15262 11732 15314
rect 11676 15260 11732 15262
rect 11452 15036 11508 15092
rect 11564 14754 11620 14756
rect 11564 14702 11566 14754
rect 11566 14702 11618 14754
rect 11618 14702 11620 14754
rect 11564 14700 11620 14702
rect 11452 14364 11508 14420
rect 11340 13804 11396 13860
rect 13132 21756 13188 21812
rect 13132 21474 13188 21476
rect 13132 21422 13134 21474
rect 13134 21422 13186 21474
rect 13186 21422 13188 21474
rect 13132 21420 13188 21422
rect 13580 23660 13636 23716
rect 13580 23042 13636 23044
rect 13580 22990 13582 23042
rect 13582 22990 13634 23042
rect 13634 22990 13636 23042
rect 13580 22988 13636 22990
rect 13580 22428 13636 22484
rect 13804 25900 13860 25956
rect 14028 28082 14084 28084
rect 14028 28030 14030 28082
rect 14030 28030 14082 28082
rect 14082 28030 14084 28082
rect 14028 28028 14084 28030
rect 14364 28476 14420 28532
rect 14924 29820 14980 29876
rect 14588 28812 14644 28868
rect 14700 29148 14756 29204
rect 13916 25788 13972 25844
rect 14140 25228 14196 25284
rect 14028 24444 14084 24500
rect 13916 22988 13972 23044
rect 13916 22258 13972 22260
rect 13916 22206 13918 22258
rect 13918 22206 13970 22258
rect 13970 22206 13972 22258
rect 13916 22204 13972 22206
rect 13804 21420 13860 21476
rect 14924 28866 14980 28868
rect 14924 28814 14926 28866
rect 14926 28814 14978 28866
rect 14978 28814 14980 28866
rect 14924 28812 14980 28814
rect 15036 29148 15092 29204
rect 17500 35586 17556 35588
rect 17500 35534 17502 35586
rect 17502 35534 17554 35586
rect 17554 35534 17556 35586
rect 17500 35532 17556 35534
rect 16044 32732 16100 32788
rect 15596 32620 15652 32676
rect 15372 31554 15428 31556
rect 15372 31502 15374 31554
rect 15374 31502 15426 31554
rect 15426 31502 15428 31554
rect 15372 31500 15428 31502
rect 15708 31276 15764 31332
rect 15372 31218 15428 31220
rect 15372 31166 15374 31218
rect 15374 31166 15426 31218
rect 15426 31166 15428 31218
rect 15372 31164 15428 31166
rect 15484 31106 15540 31108
rect 15484 31054 15486 31106
rect 15486 31054 15538 31106
rect 15538 31054 15540 31106
rect 15484 31052 15540 31054
rect 15932 31052 15988 31108
rect 16156 31724 16212 31780
rect 15596 30156 15652 30212
rect 15260 30044 15316 30100
rect 16156 30716 16212 30772
rect 15932 30044 15988 30100
rect 16156 30156 16212 30212
rect 17164 33458 17220 33460
rect 17164 33406 17166 33458
rect 17166 33406 17218 33458
rect 17218 33406 17220 33458
rect 17164 33404 17220 33406
rect 18172 37436 18228 37492
rect 17836 37378 17892 37380
rect 17836 37326 17838 37378
rect 17838 37326 17890 37378
rect 17890 37326 17892 37378
rect 17836 37324 17892 37326
rect 18172 36594 18228 36596
rect 18172 36542 18174 36594
rect 18174 36542 18226 36594
rect 18226 36542 18228 36594
rect 18172 36540 18228 36542
rect 17948 35308 18004 35364
rect 18060 33740 18116 33796
rect 18284 34636 18340 34692
rect 17612 32732 17668 32788
rect 16604 32674 16660 32676
rect 16604 32622 16606 32674
rect 16606 32622 16658 32674
rect 16658 32622 16660 32674
rect 16604 32620 16660 32622
rect 17388 32674 17444 32676
rect 17388 32622 17390 32674
rect 17390 32622 17442 32674
rect 17442 32622 17444 32674
rect 17388 32620 17444 32622
rect 16492 32508 16548 32564
rect 16604 31276 16660 31332
rect 16268 29820 16324 29876
rect 16044 29596 16100 29652
rect 15260 29148 15316 29204
rect 16156 29538 16212 29540
rect 16156 29486 16158 29538
rect 16158 29486 16210 29538
rect 16210 29486 16212 29538
rect 16156 29484 16212 29486
rect 15372 28588 15428 28644
rect 15260 28476 15316 28532
rect 14812 27074 14868 27076
rect 14812 27022 14814 27074
rect 14814 27022 14866 27074
rect 14866 27022 14868 27074
rect 14812 27020 14868 27022
rect 14924 25506 14980 25508
rect 14924 25454 14926 25506
rect 14926 25454 14978 25506
rect 14978 25454 14980 25506
rect 14924 25452 14980 25454
rect 14364 24444 14420 24500
rect 14700 25228 14756 25284
rect 15372 27580 15428 27636
rect 15372 26962 15428 26964
rect 15372 26910 15374 26962
rect 15374 26910 15426 26962
rect 15426 26910 15428 26962
rect 15372 26908 15428 26910
rect 16492 29148 16548 29204
rect 16940 30210 16996 30212
rect 16940 30158 16942 30210
rect 16942 30158 16994 30210
rect 16994 30158 16996 30210
rect 16940 30156 16996 30158
rect 16828 30044 16884 30100
rect 16044 28252 16100 28308
rect 15596 28028 15652 28084
rect 17612 32562 17668 32564
rect 17612 32510 17614 32562
rect 17614 32510 17666 32562
rect 17666 32510 17668 32562
rect 17612 32508 17668 32510
rect 18844 37490 18900 37492
rect 18844 37438 18846 37490
rect 18846 37438 18898 37490
rect 18898 37438 18900 37490
rect 18844 37436 18900 37438
rect 18732 35196 18788 35252
rect 18956 37324 19012 37380
rect 18508 34860 18564 34916
rect 18844 34636 18900 34692
rect 18508 33740 18564 33796
rect 18284 33068 18340 33124
rect 17948 32508 18004 32564
rect 18172 32450 18228 32452
rect 18172 32398 18174 32450
rect 18174 32398 18226 32450
rect 18226 32398 18228 32450
rect 18172 32396 18228 32398
rect 18172 31778 18228 31780
rect 18172 31726 18174 31778
rect 18174 31726 18226 31778
rect 18226 31726 18228 31778
rect 18172 31724 18228 31726
rect 18060 31052 18116 31108
rect 17612 30268 17668 30324
rect 18060 30268 18116 30324
rect 17948 30098 18004 30100
rect 17948 30046 17950 30098
rect 17950 30046 18002 30098
rect 18002 30046 18004 30098
rect 17948 30044 18004 30046
rect 16940 29484 16996 29540
rect 16380 28140 16436 28196
rect 16604 28252 16660 28308
rect 15820 27970 15876 27972
rect 15820 27918 15822 27970
rect 15822 27918 15874 27970
rect 15874 27918 15876 27970
rect 15820 27916 15876 27918
rect 16268 27916 16324 27972
rect 15932 27746 15988 27748
rect 15932 27694 15934 27746
rect 15934 27694 15986 27746
rect 15986 27694 15988 27746
rect 15932 27692 15988 27694
rect 15820 27580 15876 27636
rect 15372 26012 15428 26068
rect 15260 25900 15316 25956
rect 15148 25282 15204 25284
rect 15148 25230 15150 25282
rect 15150 25230 15202 25282
rect 15202 25230 15204 25282
rect 15148 25228 15204 25230
rect 14924 23660 14980 23716
rect 14476 22482 14532 22484
rect 14476 22430 14478 22482
rect 14478 22430 14530 22482
rect 14530 22430 14532 22482
rect 14476 22428 14532 22430
rect 14812 21362 14868 21364
rect 14812 21310 14814 21362
rect 14814 21310 14866 21362
rect 14866 21310 14868 21362
rect 14812 21308 14868 21310
rect 14364 21026 14420 21028
rect 14364 20974 14366 21026
rect 14366 20974 14418 21026
rect 14418 20974 14420 21026
rect 14364 20972 14420 20974
rect 14028 19292 14084 19348
rect 13804 19234 13860 19236
rect 13804 19182 13806 19234
rect 13806 19182 13858 19234
rect 13858 19182 13860 19234
rect 13804 19180 13860 19182
rect 13468 18396 13524 18452
rect 14252 20690 14308 20692
rect 14252 20638 14254 20690
rect 14254 20638 14306 20690
rect 14306 20638 14308 20690
rect 14252 20636 14308 20638
rect 13692 17836 13748 17892
rect 13020 17724 13076 17780
rect 13580 17666 13636 17668
rect 13580 17614 13582 17666
rect 13582 17614 13634 17666
rect 13634 17614 13636 17666
rect 13580 17612 13636 17614
rect 12236 16098 12292 16100
rect 12236 16046 12238 16098
rect 12238 16046 12290 16098
rect 12290 16046 12292 16098
rect 12236 16044 12292 16046
rect 12012 14812 12068 14868
rect 11676 13020 11732 13076
rect 11788 11788 11844 11844
rect 11340 11170 11396 11172
rect 11340 11118 11342 11170
rect 11342 11118 11394 11170
rect 11394 11118 11396 11170
rect 11340 11116 11396 11118
rect 11788 11116 11844 11172
rect 11900 10722 11956 10724
rect 11900 10670 11902 10722
rect 11902 10670 11954 10722
rect 11954 10670 11956 10722
rect 11900 10668 11956 10670
rect 12348 14700 12404 14756
rect 13468 16716 13524 16772
rect 13804 16210 13860 16212
rect 13804 16158 13806 16210
rect 13806 16158 13858 16210
rect 13858 16158 13860 16210
rect 13804 16156 13860 16158
rect 12796 16044 12852 16100
rect 13020 15932 13076 15988
rect 13580 15932 13636 15988
rect 13468 15820 13524 15876
rect 12684 15538 12740 15540
rect 12684 15486 12686 15538
rect 12686 15486 12738 15538
rect 12738 15486 12740 15538
rect 12684 15484 12740 15486
rect 12572 14418 12628 14420
rect 12572 14366 12574 14418
rect 12574 14366 12626 14418
rect 12626 14366 12628 14418
rect 12572 14364 12628 14366
rect 12684 14252 12740 14308
rect 12348 13692 12404 13748
rect 12236 13132 12292 13188
rect 12684 13132 12740 13188
rect 12124 13020 12180 13076
rect 12684 12796 12740 12852
rect 12572 11788 12628 11844
rect 11900 9772 11956 9828
rect 12124 9772 12180 9828
rect 12460 11282 12516 11284
rect 12460 11230 12462 11282
rect 12462 11230 12514 11282
rect 12514 11230 12516 11282
rect 12460 11228 12516 11230
rect 12348 11170 12404 11172
rect 12348 11118 12350 11170
rect 12350 11118 12402 11170
rect 12402 11118 12404 11170
rect 12348 11116 12404 11118
rect 12572 11004 12628 11060
rect 11564 9660 11620 9716
rect 11228 7644 11284 7700
rect 11228 6860 11284 6916
rect 10668 6130 10724 6132
rect 10668 6078 10670 6130
rect 10670 6078 10722 6130
rect 10722 6078 10724 6130
rect 10668 6076 10724 6078
rect 10332 5964 10388 6020
rect 11116 6466 11172 6468
rect 11116 6414 11118 6466
rect 11118 6414 11170 6466
rect 11170 6414 11172 6466
rect 11116 6412 11172 6414
rect 11452 6748 11508 6804
rect 11788 7980 11844 8036
rect 11900 7698 11956 7700
rect 11900 7646 11902 7698
rect 11902 7646 11954 7698
rect 11954 7646 11956 7698
rect 11900 7644 11956 7646
rect 11340 6412 11396 6468
rect 11788 6466 11844 6468
rect 11788 6414 11790 6466
rect 11790 6414 11842 6466
rect 11842 6414 11844 6466
rect 11788 6412 11844 6414
rect 11004 5964 11060 6020
rect 11004 5628 11060 5684
rect 10220 4956 10276 5012
rect 10780 4898 10836 4900
rect 10780 4846 10782 4898
rect 10782 4846 10834 4898
rect 10834 4846 10836 4898
rect 10780 4844 10836 4846
rect 9100 4450 9156 4452
rect 9100 4398 9102 4450
rect 9102 4398 9154 4450
rect 9154 4398 9156 4450
rect 9100 4396 9156 4398
rect 9996 4450 10052 4452
rect 9996 4398 9998 4450
rect 9998 4398 10050 4450
rect 10050 4398 10052 4450
rect 9996 4396 10052 4398
rect 9660 4338 9716 4340
rect 9660 4286 9662 4338
rect 9662 4286 9714 4338
rect 9714 4286 9716 4338
rect 9660 4284 9716 4286
rect 9324 4172 9380 4228
rect 9324 3388 9380 3444
rect 9436 3500 9492 3556
rect 10556 4338 10612 4340
rect 10556 4286 10558 4338
rect 10558 4286 10610 4338
rect 10610 4286 10612 4338
rect 10556 4284 10612 4286
rect 10780 4226 10836 4228
rect 10780 4174 10782 4226
rect 10782 4174 10834 4226
rect 10834 4174 10836 4226
rect 10780 4172 10836 4174
rect 11564 6076 11620 6132
rect 11228 5068 11284 5124
rect 11004 4844 11060 4900
rect 11340 4956 11396 5012
rect 12012 5682 12068 5684
rect 12012 5630 12014 5682
rect 12014 5630 12066 5682
rect 12066 5630 12068 5682
rect 12012 5628 12068 5630
rect 11900 4956 11956 5012
rect 11452 3388 11508 3444
rect 12572 9772 12628 9828
rect 13020 14252 13076 14308
rect 12908 13858 12964 13860
rect 12908 13806 12910 13858
rect 12910 13806 12962 13858
rect 12962 13806 12964 13858
rect 12908 13804 12964 13806
rect 13804 15932 13860 15988
rect 13804 15314 13860 15316
rect 13804 15262 13806 15314
rect 13806 15262 13858 15314
rect 13858 15262 13860 15314
rect 13804 15260 13860 15262
rect 14140 18226 14196 18228
rect 14140 18174 14142 18226
rect 14142 18174 14194 18226
rect 14194 18174 14196 18226
rect 14140 18172 14196 18174
rect 14028 17666 14084 17668
rect 14028 17614 14030 17666
rect 14030 17614 14082 17666
rect 14082 17614 14084 17666
rect 14028 17612 14084 17614
rect 14140 16716 14196 16772
rect 14700 20914 14756 20916
rect 14700 20862 14702 20914
rect 14702 20862 14754 20914
rect 14754 20862 14756 20914
rect 14700 20860 14756 20862
rect 16156 25900 16212 25956
rect 15932 25788 15988 25844
rect 15708 25506 15764 25508
rect 15708 25454 15710 25506
rect 15710 25454 15762 25506
rect 15762 25454 15764 25506
rect 15708 25452 15764 25454
rect 15148 20802 15204 20804
rect 15148 20750 15150 20802
rect 15150 20750 15202 20802
rect 15202 20750 15204 20802
rect 15148 20748 15204 20750
rect 14700 19292 14756 19348
rect 15148 19346 15204 19348
rect 15148 19294 15150 19346
rect 15150 19294 15202 19346
rect 15202 19294 15204 19346
rect 15148 19292 15204 19294
rect 14700 18450 14756 18452
rect 14700 18398 14702 18450
rect 14702 18398 14754 18450
rect 14754 18398 14756 18450
rect 14700 18396 14756 18398
rect 14028 15932 14084 15988
rect 14252 15986 14308 15988
rect 14252 15934 14254 15986
rect 14254 15934 14306 15986
rect 14306 15934 14308 15986
rect 14252 15932 14308 15934
rect 13804 14306 13860 14308
rect 13804 14254 13806 14306
rect 13806 14254 13858 14306
rect 13858 14254 13860 14306
rect 13804 14252 13860 14254
rect 13580 13468 13636 13524
rect 13244 13356 13300 13412
rect 13580 13244 13636 13300
rect 13468 13186 13524 13188
rect 13468 13134 13470 13186
rect 13470 13134 13522 13186
rect 13522 13134 13524 13186
rect 13468 13132 13524 13134
rect 13356 12796 13412 12852
rect 13916 13804 13972 13860
rect 13468 12348 13524 12404
rect 12908 12124 12964 12180
rect 13020 12012 13076 12068
rect 13692 12178 13748 12180
rect 13692 12126 13694 12178
rect 13694 12126 13746 12178
rect 13746 12126 13748 12178
rect 13692 12124 13748 12126
rect 14476 16658 14532 16660
rect 14476 16606 14478 16658
rect 14478 16606 14530 16658
rect 14530 16606 14532 16658
rect 14476 16604 14532 16606
rect 14700 16380 14756 16436
rect 15036 16716 15092 16772
rect 15372 21308 15428 21364
rect 15372 20636 15428 20692
rect 16716 26290 16772 26292
rect 16716 26238 16718 26290
rect 16718 26238 16770 26290
rect 16770 26238 16772 26290
rect 16716 26236 16772 26238
rect 17500 29538 17556 29540
rect 17500 29486 17502 29538
rect 17502 29486 17554 29538
rect 17554 29486 17556 29538
rect 17500 29484 17556 29486
rect 17388 29202 17444 29204
rect 17388 29150 17390 29202
rect 17390 29150 17442 29202
rect 17442 29150 17444 29202
rect 17388 29148 17444 29150
rect 18620 32562 18676 32564
rect 18620 32510 18622 32562
rect 18622 32510 18674 32562
rect 18674 32510 18676 32562
rect 18620 32508 18676 32510
rect 20412 40348 20468 40404
rect 19628 39452 19684 39508
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 20300 38834 20356 38836
rect 20300 38782 20302 38834
rect 20302 38782 20354 38834
rect 20354 38782 20356 38834
rect 20300 38780 20356 38782
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19964 36764 20020 36820
rect 19740 36652 19796 36708
rect 21420 41970 21476 41972
rect 21420 41918 21422 41970
rect 21422 41918 21474 41970
rect 21474 41918 21476 41970
rect 21420 41916 21476 41918
rect 22876 43260 22932 43316
rect 22764 43148 22820 43204
rect 23996 43932 24052 43988
rect 23324 43148 23380 43204
rect 23436 43372 23492 43428
rect 23660 42700 23716 42756
rect 23212 42194 23268 42196
rect 23212 42142 23214 42194
rect 23214 42142 23266 42194
rect 23266 42142 23268 42194
rect 23212 42140 23268 42142
rect 22428 42028 22484 42084
rect 21868 41410 21924 41412
rect 21868 41358 21870 41410
rect 21870 41358 21922 41410
rect 21922 41358 21924 41410
rect 21868 41356 21924 41358
rect 22204 41692 22260 41748
rect 22316 41186 22372 41188
rect 22316 41134 22318 41186
rect 22318 41134 22370 41186
rect 22370 41134 22372 41186
rect 22316 41132 22372 41134
rect 23212 41356 23268 41412
rect 23548 41074 23604 41076
rect 23548 41022 23550 41074
rect 23550 41022 23602 41074
rect 23602 41022 23604 41074
rect 23548 41020 23604 41022
rect 23436 40908 23492 40964
rect 22988 40626 23044 40628
rect 22988 40574 22990 40626
rect 22990 40574 23042 40626
rect 23042 40574 23044 40626
rect 22988 40572 23044 40574
rect 22316 40290 22372 40292
rect 22316 40238 22318 40290
rect 22318 40238 22370 40290
rect 22370 40238 22372 40290
rect 22316 40236 22372 40238
rect 21196 37436 21252 37492
rect 22316 37772 22372 37828
rect 20748 36652 20804 36708
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19852 35420 19908 35476
rect 21196 35756 21252 35812
rect 22540 35810 22596 35812
rect 22540 35758 22542 35810
rect 22542 35758 22594 35810
rect 22594 35758 22596 35810
rect 22540 35756 22596 35758
rect 21644 35474 21700 35476
rect 21644 35422 21646 35474
rect 21646 35422 21698 35474
rect 21698 35422 21700 35474
rect 21644 35420 21700 35422
rect 21980 35474 22036 35476
rect 21980 35422 21982 35474
rect 21982 35422 22034 35474
rect 22034 35422 22036 35474
rect 21980 35420 22036 35422
rect 20524 35308 20580 35364
rect 20300 34860 20356 34916
rect 19404 33628 19460 33684
rect 19180 32620 19236 32676
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 20188 33628 20244 33684
rect 20076 33404 20132 33460
rect 19628 33234 19684 33236
rect 19628 33182 19630 33234
rect 19630 33182 19682 33234
rect 19682 33182 19684 33234
rect 19628 33180 19684 33182
rect 18620 31948 18676 32004
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19628 32620 19684 32676
rect 19068 31666 19124 31668
rect 19068 31614 19070 31666
rect 19070 31614 19122 31666
rect 19122 31614 19124 31666
rect 19068 31612 19124 31614
rect 19740 32284 19796 32340
rect 19068 30268 19124 30324
rect 20412 33628 20468 33684
rect 22764 36092 22820 36148
rect 23884 42140 23940 42196
rect 23884 40962 23940 40964
rect 23884 40910 23886 40962
rect 23886 40910 23938 40962
rect 23938 40910 23940 40962
rect 23884 40908 23940 40910
rect 24332 43314 24388 43316
rect 24332 43262 24334 43314
rect 24334 43262 24386 43314
rect 24386 43262 24388 43314
rect 24332 43260 24388 43262
rect 25340 45106 25396 45108
rect 25340 45054 25342 45106
rect 25342 45054 25394 45106
rect 25394 45054 25396 45106
rect 25340 45052 25396 45054
rect 25004 43932 25060 43988
rect 26796 44940 26852 44996
rect 24668 43538 24724 43540
rect 24668 43486 24670 43538
rect 24670 43486 24722 43538
rect 24722 43486 24724 43538
rect 24668 43484 24724 43486
rect 25564 43484 25620 43540
rect 28140 44994 28196 44996
rect 28140 44942 28142 44994
rect 28142 44942 28194 44994
rect 28194 44942 28196 44994
rect 28140 44940 28196 44942
rect 28924 46060 28980 46116
rect 30044 46114 30100 46116
rect 30044 46062 30046 46114
rect 30046 46062 30098 46114
rect 30098 46062 30100 46114
rect 30044 46060 30100 46062
rect 28588 45276 28644 45332
rect 25676 43372 25732 43428
rect 25116 42754 25172 42756
rect 25116 42702 25118 42754
rect 25118 42702 25170 42754
rect 25170 42702 25172 42754
rect 25116 42700 25172 42702
rect 24556 41020 24612 41076
rect 24220 40962 24276 40964
rect 24220 40910 24222 40962
rect 24222 40910 24274 40962
rect 24274 40910 24276 40962
rect 24220 40908 24276 40910
rect 23660 40402 23716 40404
rect 23660 40350 23662 40402
rect 23662 40350 23714 40402
rect 23714 40350 23716 40402
rect 23660 40348 23716 40350
rect 23772 40290 23828 40292
rect 23772 40238 23774 40290
rect 23774 40238 23826 40290
rect 23826 40238 23828 40290
rect 23772 40236 23828 40238
rect 24220 40402 24276 40404
rect 24220 40350 24222 40402
rect 24222 40350 24274 40402
rect 24274 40350 24276 40402
rect 24220 40348 24276 40350
rect 23884 39394 23940 39396
rect 23884 39342 23886 39394
rect 23886 39342 23938 39394
rect 23938 39342 23940 39394
rect 23884 39340 23940 39342
rect 23436 37826 23492 37828
rect 23436 37774 23438 37826
rect 23438 37774 23490 37826
rect 23490 37774 23492 37826
rect 23436 37772 23492 37774
rect 23548 38220 23604 38276
rect 23212 36428 23268 36484
rect 22652 35868 22708 35924
rect 23212 35980 23268 36036
rect 23436 35980 23492 36036
rect 23324 35474 23380 35476
rect 23324 35422 23326 35474
rect 23326 35422 23378 35474
rect 23378 35422 23380 35474
rect 23324 35420 23380 35422
rect 23100 34748 23156 34804
rect 20748 34690 20804 34692
rect 20748 34638 20750 34690
rect 20750 34638 20802 34690
rect 20802 34638 20804 34690
rect 20748 34636 20804 34638
rect 22428 34524 22484 34580
rect 20412 33458 20468 33460
rect 20412 33406 20414 33458
rect 20414 33406 20466 33458
rect 20466 33406 20468 33458
rect 20412 33404 20468 33406
rect 22204 33180 22260 33236
rect 22988 33122 23044 33124
rect 22988 33070 22990 33122
rect 22990 33070 23042 33122
rect 23042 33070 23044 33122
rect 22988 33068 23044 33070
rect 21420 32284 21476 32340
rect 21420 31948 21476 32004
rect 20972 31612 21028 31668
rect 17948 29650 18004 29652
rect 17948 29598 17950 29650
rect 17950 29598 18002 29650
rect 18002 29598 18004 29650
rect 17948 29596 18004 29598
rect 17276 28140 17332 28196
rect 16828 25788 16884 25844
rect 16940 27692 16996 27748
rect 17612 27074 17668 27076
rect 17612 27022 17614 27074
rect 17614 27022 17666 27074
rect 17666 27022 17668 27074
rect 17612 27020 17668 27022
rect 18284 29426 18340 29428
rect 18284 29374 18286 29426
rect 18286 29374 18338 29426
rect 18338 29374 18340 29426
rect 18284 29372 18340 29374
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19180 29596 19236 29652
rect 18844 29036 18900 29092
rect 18620 28140 18676 28196
rect 18508 28028 18564 28084
rect 17948 27858 18004 27860
rect 17948 27806 17950 27858
rect 17950 27806 18002 27858
rect 18002 27806 18004 27858
rect 17948 27804 18004 27806
rect 17836 26796 17892 26852
rect 17500 26012 17556 26068
rect 17388 25900 17444 25956
rect 17724 26290 17780 26292
rect 17724 26238 17726 26290
rect 17726 26238 17778 26290
rect 17778 26238 17780 26290
rect 17724 26236 17780 26238
rect 17612 25452 17668 25508
rect 18396 27074 18452 27076
rect 18396 27022 18398 27074
rect 18398 27022 18450 27074
rect 18450 27022 18452 27074
rect 18396 27020 18452 27022
rect 18284 26908 18340 26964
rect 18396 26850 18452 26852
rect 18396 26798 18398 26850
rect 18398 26798 18450 26850
rect 18450 26798 18452 26850
rect 18396 26796 18452 26798
rect 16156 25228 16212 25284
rect 18620 26796 18676 26852
rect 19292 29314 19348 29316
rect 19292 29262 19294 29314
rect 19294 29262 19346 29314
rect 19346 29262 19348 29314
rect 19292 29260 19348 29262
rect 19740 29986 19796 29988
rect 19740 29934 19742 29986
rect 19742 29934 19794 29986
rect 19794 29934 19796 29986
rect 19740 29932 19796 29934
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19516 29148 19572 29204
rect 20636 29260 20692 29316
rect 19628 29036 19684 29092
rect 19180 28924 19236 28980
rect 19068 28252 19124 28308
rect 19180 26796 19236 26852
rect 21308 31276 21364 31332
rect 22204 31836 22260 31892
rect 22092 31388 22148 31444
rect 21756 31276 21812 31332
rect 21980 31164 22036 31220
rect 20748 28924 20804 28980
rect 19404 28642 19460 28644
rect 19404 28590 19406 28642
rect 19406 28590 19458 28642
rect 19458 28590 19460 28642
rect 19404 28588 19460 28590
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19516 28028 19572 28084
rect 20076 28028 20132 28084
rect 21308 29314 21364 29316
rect 21308 29262 21310 29314
rect 21310 29262 21362 29314
rect 21362 29262 21364 29314
rect 21308 29260 21364 29262
rect 21420 29148 21476 29204
rect 21532 28700 21588 28756
rect 20860 27916 20916 27972
rect 23212 32956 23268 33012
rect 23996 38556 24052 38612
rect 23772 37772 23828 37828
rect 25452 41916 25508 41972
rect 25004 41132 25060 41188
rect 25452 41132 25508 41188
rect 25564 41356 25620 41412
rect 25228 41020 25284 41076
rect 25340 40572 25396 40628
rect 25788 41186 25844 41188
rect 25788 41134 25790 41186
rect 25790 41134 25842 41186
rect 25842 41134 25844 41186
rect 25788 41132 25844 41134
rect 25564 40348 25620 40404
rect 26908 43260 26964 43316
rect 26796 41916 26852 41972
rect 28028 43538 28084 43540
rect 28028 43486 28030 43538
rect 28030 43486 28082 43538
rect 28082 43486 28084 43538
rect 28028 43484 28084 43486
rect 27916 42812 27972 42868
rect 28028 43260 28084 43316
rect 27580 42642 27636 42644
rect 27580 42590 27582 42642
rect 27582 42590 27634 42642
rect 27634 42590 27636 42642
rect 27580 42588 27636 42590
rect 26796 41410 26852 41412
rect 26796 41358 26798 41410
rect 26798 41358 26850 41410
rect 26850 41358 26852 41410
rect 26796 41356 26852 41358
rect 26572 40908 26628 40964
rect 27356 41020 27412 41076
rect 26012 39788 26068 39844
rect 24220 39618 24276 39620
rect 24220 39566 24222 39618
rect 24222 39566 24274 39618
rect 24274 39566 24276 39618
rect 24220 39564 24276 39566
rect 27692 40962 27748 40964
rect 27692 40910 27694 40962
rect 27694 40910 27746 40962
rect 27746 40910 27748 40962
rect 27692 40908 27748 40910
rect 27020 40290 27076 40292
rect 27020 40238 27022 40290
rect 27022 40238 27074 40290
rect 27074 40238 27076 40290
rect 27020 40236 27076 40238
rect 26348 39676 26404 39732
rect 24444 38556 24500 38612
rect 24668 38780 24724 38836
rect 24444 38332 24500 38388
rect 24220 38220 24276 38276
rect 23772 35980 23828 36036
rect 23548 33292 23604 33348
rect 24444 37212 24500 37268
rect 24220 36540 24276 36596
rect 24332 36764 24388 36820
rect 24108 36482 24164 36484
rect 24108 36430 24110 36482
rect 24110 36430 24162 36482
rect 24162 36430 24164 36482
rect 24108 36428 24164 36430
rect 24220 36258 24276 36260
rect 24220 36206 24222 36258
rect 24222 36206 24274 36258
rect 24274 36206 24276 36258
rect 24220 36204 24276 36206
rect 23996 35810 24052 35812
rect 23996 35758 23998 35810
rect 23998 35758 24050 35810
rect 24050 35758 24052 35810
rect 23996 35756 24052 35758
rect 25004 38556 25060 38612
rect 23884 34748 23940 34804
rect 24668 36428 24724 36484
rect 22988 32396 23044 32452
rect 23324 31836 23380 31892
rect 23548 32956 23604 33012
rect 22652 30940 22708 30996
rect 23772 33122 23828 33124
rect 23772 33070 23774 33122
rect 23774 33070 23826 33122
rect 23826 33070 23828 33122
rect 23772 33068 23828 33070
rect 23884 31836 23940 31892
rect 23324 31164 23380 31220
rect 23436 30994 23492 30996
rect 23436 30942 23438 30994
rect 23438 30942 23490 30994
rect 23490 30942 23492 30994
rect 23436 30940 23492 30942
rect 22204 30156 22260 30212
rect 23660 29596 23716 29652
rect 24332 35644 24388 35700
rect 24668 35644 24724 35700
rect 25564 38050 25620 38052
rect 25564 37998 25566 38050
rect 25566 37998 25618 38050
rect 25618 37998 25620 38050
rect 25564 37996 25620 37998
rect 25340 37490 25396 37492
rect 25340 37438 25342 37490
rect 25342 37438 25394 37490
rect 25394 37438 25396 37490
rect 25340 37436 25396 37438
rect 26012 37436 26068 37492
rect 25900 37378 25956 37380
rect 25900 37326 25902 37378
rect 25902 37326 25954 37378
rect 25954 37326 25956 37378
rect 25900 37324 25956 37326
rect 25676 37266 25732 37268
rect 25676 37214 25678 37266
rect 25678 37214 25730 37266
rect 25730 37214 25732 37266
rect 25676 37212 25732 37214
rect 26572 39788 26628 39844
rect 26908 39730 26964 39732
rect 26908 39678 26910 39730
rect 26910 39678 26962 39730
rect 26962 39678 26964 39730
rect 26908 39676 26964 39678
rect 27692 39676 27748 39732
rect 27020 39340 27076 39396
rect 28812 43538 28868 43540
rect 28812 43486 28814 43538
rect 28814 43486 28866 43538
rect 28866 43486 28868 43538
rect 28812 43484 28868 43486
rect 28364 43372 28420 43428
rect 28252 41020 28308 41076
rect 28700 42700 28756 42756
rect 29148 42588 29204 42644
rect 29708 45330 29764 45332
rect 29708 45278 29710 45330
rect 29710 45278 29762 45330
rect 29762 45278 29764 45330
rect 29708 45276 29764 45278
rect 29372 45106 29428 45108
rect 29372 45054 29374 45106
rect 29374 45054 29426 45106
rect 29426 45054 29428 45106
rect 29372 45052 29428 45054
rect 30380 44098 30436 44100
rect 30380 44046 30382 44098
rect 30382 44046 30434 44098
rect 30434 44046 30436 44098
rect 30380 44044 30436 44046
rect 30604 44940 30660 44996
rect 29932 43708 29988 43764
rect 28700 40236 28756 40292
rect 27804 38108 27860 38164
rect 27692 37378 27748 37380
rect 27692 37326 27694 37378
rect 27694 37326 27746 37378
rect 27746 37326 27748 37378
rect 27692 37324 27748 37326
rect 24892 36316 24948 36372
rect 24892 35756 24948 35812
rect 25788 35868 25844 35924
rect 25564 35698 25620 35700
rect 25564 35646 25566 35698
rect 25566 35646 25618 35698
rect 25618 35646 25620 35698
rect 25564 35644 25620 35646
rect 27020 35922 27076 35924
rect 27020 35870 27022 35922
rect 27022 35870 27074 35922
rect 27074 35870 27076 35922
rect 27020 35868 27076 35870
rect 26124 35756 26180 35812
rect 24220 34524 24276 34580
rect 24108 33346 24164 33348
rect 24108 33294 24110 33346
rect 24110 33294 24162 33346
rect 24162 33294 24164 33346
rect 24108 33292 24164 33294
rect 24332 32396 24388 32452
rect 25900 35196 25956 35252
rect 25116 33404 25172 33460
rect 25900 33458 25956 33460
rect 25900 33406 25902 33458
rect 25902 33406 25954 33458
rect 25954 33406 25956 33458
rect 25900 33404 25956 33406
rect 25004 33234 25060 33236
rect 25004 33182 25006 33234
rect 25006 33182 25058 33234
rect 25058 33182 25060 33234
rect 25004 33180 25060 33182
rect 25228 33068 25284 33124
rect 25452 32450 25508 32452
rect 25452 32398 25454 32450
rect 25454 32398 25506 32450
rect 25506 32398 25508 32450
rect 25452 32396 25508 32398
rect 24668 32338 24724 32340
rect 24668 32286 24670 32338
rect 24670 32286 24722 32338
rect 24722 32286 24724 32338
rect 24668 32284 24724 32286
rect 25340 32284 25396 32340
rect 24780 32060 24836 32116
rect 24556 31218 24612 31220
rect 24556 31166 24558 31218
rect 24558 31166 24610 31218
rect 24610 31166 24612 31218
rect 24556 31164 24612 31166
rect 22092 28754 22148 28756
rect 22092 28702 22094 28754
rect 22094 28702 22146 28754
rect 22146 28702 22148 28754
rect 22092 28700 22148 28702
rect 24220 30156 24276 30212
rect 21644 27804 21700 27860
rect 20636 27020 20692 27076
rect 20412 26908 20468 26964
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 15596 23714 15652 23716
rect 15596 23662 15598 23714
rect 15598 23662 15650 23714
rect 15650 23662 15652 23714
rect 15596 23660 15652 23662
rect 18396 23714 18452 23716
rect 18396 23662 18398 23714
rect 18398 23662 18450 23714
rect 18450 23662 18452 23714
rect 18396 23660 18452 23662
rect 15820 22988 15876 23044
rect 16828 23042 16884 23044
rect 16828 22990 16830 23042
rect 16830 22990 16882 23042
rect 16882 22990 16884 23042
rect 16828 22988 16884 22990
rect 17612 23212 17668 23268
rect 18060 23378 18116 23380
rect 18060 23326 18062 23378
rect 18062 23326 18114 23378
rect 18114 23326 18116 23378
rect 18060 23324 18116 23326
rect 18844 23378 18900 23380
rect 18844 23326 18846 23378
rect 18846 23326 18898 23378
rect 18898 23326 18900 23378
rect 18844 23324 18900 23326
rect 15708 20914 15764 20916
rect 15708 20862 15710 20914
rect 15710 20862 15762 20914
rect 15762 20862 15764 20914
rect 15708 20860 15764 20862
rect 16156 20802 16212 20804
rect 16156 20750 16158 20802
rect 16158 20750 16210 20802
rect 16210 20750 16212 20802
rect 16156 20748 16212 20750
rect 16604 20748 16660 20804
rect 15260 16716 15316 16772
rect 15484 20018 15540 20020
rect 15484 19966 15486 20018
rect 15486 19966 15538 20018
rect 15538 19966 15540 20018
rect 15484 19964 15540 19966
rect 16716 20690 16772 20692
rect 16716 20638 16718 20690
rect 16718 20638 16770 20690
rect 16770 20638 16772 20690
rect 16716 20636 16772 20638
rect 17836 20802 17892 20804
rect 17836 20750 17838 20802
rect 17838 20750 17890 20802
rect 17890 20750 17892 20802
rect 17836 20748 17892 20750
rect 15820 19292 15876 19348
rect 16828 18396 16884 18452
rect 15484 16770 15540 16772
rect 15484 16718 15486 16770
rect 15486 16718 15538 16770
rect 15538 16718 15540 16770
rect 15484 16716 15540 16718
rect 15372 16098 15428 16100
rect 15372 16046 15374 16098
rect 15374 16046 15426 16098
rect 15426 16046 15428 16098
rect 15372 16044 15428 16046
rect 15260 15932 15316 15988
rect 14476 15820 14532 15876
rect 14812 15596 14868 15652
rect 14364 14812 14420 14868
rect 14252 14588 14308 14644
rect 14476 14588 14532 14644
rect 14700 14924 14756 14980
rect 15820 16716 15876 16772
rect 15932 16994 15988 16996
rect 15932 16942 15934 16994
rect 15934 16942 15986 16994
rect 15986 16942 15988 16994
rect 15932 16940 15988 16942
rect 15596 15596 15652 15652
rect 16156 16882 16212 16884
rect 16156 16830 16158 16882
rect 16158 16830 16210 16882
rect 16210 16830 16212 16882
rect 16156 16828 16212 16830
rect 16156 16210 16212 16212
rect 16156 16158 16158 16210
rect 16158 16158 16210 16210
rect 16210 16158 16212 16210
rect 16156 16156 16212 16158
rect 17724 20076 17780 20132
rect 18508 21196 18564 21252
rect 18284 20748 18340 20804
rect 18844 21196 18900 21252
rect 17612 18956 17668 19012
rect 17388 18450 17444 18452
rect 17388 18398 17390 18450
rect 17390 18398 17442 18450
rect 17442 18398 17444 18450
rect 17388 18396 17444 18398
rect 17836 18338 17892 18340
rect 17836 18286 17838 18338
rect 17838 18286 17890 18338
rect 17890 18286 17892 18338
rect 17836 18284 17892 18286
rect 16828 17052 16884 17108
rect 17164 17052 17220 17108
rect 17276 16940 17332 16996
rect 18060 18396 18116 18452
rect 17612 16828 17668 16884
rect 17724 16770 17780 16772
rect 17724 16718 17726 16770
rect 17726 16718 17778 16770
rect 17778 16718 17780 16770
rect 17724 16716 17780 16718
rect 17500 16604 17556 16660
rect 16156 15484 16212 15540
rect 15932 15372 15988 15428
rect 15484 15314 15540 15316
rect 15484 15262 15486 15314
rect 15486 15262 15538 15314
rect 15538 15262 15540 15314
rect 15484 15260 15540 15262
rect 16156 15314 16212 15316
rect 16156 15262 16158 15314
rect 16158 15262 16210 15314
rect 16210 15262 16212 15314
rect 16156 15260 16212 15262
rect 15708 15202 15764 15204
rect 15708 15150 15710 15202
rect 15710 15150 15762 15202
rect 15762 15150 15764 15202
rect 15708 15148 15764 15150
rect 14588 13804 14644 13860
rect 16604 15372 16660 15428
rect 14812 14530 14868 14532
rect 14812 14478 14814 14530
rect 14814 14478 14866 14530
rect 14866 14478 14868 14530
rect 14812 14476 14868 14478
rect 15484 14140 15540 14196
rect 14812 13468 14868 13524
rect 14700 12962 14756 12964
rect 14700 12910 14702 12962
rect 14702 12910 14754 12962
rect 14754 12910 14756 12962
rect 14700 12908 14756 12910
rect 14364 12460 14420 12516
rect 14028 12348 14084 12404
rect 13916 12012 13972 12068
rect 14252 11394 14308 11396
rect 14252 11342 14254 11394
rect 14254 11342 14306 11394
rect 14306 11342 14308 11394
rect 14252 11340 14308 11342
rect 13804 11282 13860 11284
rect 13804 11230 13806 11282
rect 13806 11230 13858 11282
rect 13858 11230 13860 11282
rect 13804 11228 13860 11230
rect 13356 10668 13412 10724
rect 13916 11004 13972 11060
rect 12908 9826 12964 9828
rect 12908 9774 12910 9826
rect 12910 9774 12962 9826
rect 12962 9774 12964 9826
rect 12908 9772 12964 9774
rect 14700 12124 14756 12180
rect 12796 9548 12852 9604
rect 12348 7698 12404 7700
rect 12348 7646 12350 7698
rect 12350 7646 12402 7698
rect 12402 7646 12404 7698
rect 12348 7644 12404 7646
rect 13580 8370 13636 8372
rect 13580 8318 13582 8370
rect 13582 8318 13634 8370
rect 13634 8318 13636 8370
rect 13580 8316 13636 8318
rect 13020 7644 13076 7700
rect 12684 7474 12740 7476
rect 12684 7422 12686 7474
rect 12686 7422 12738 7474
rect 12738 7422 12740 7474
rect 12684 7420 12740 7422
rect 12236 6466 12292 6468
rect 12236 6414 12238 6466
rect 12238 6414 12290 6466
rect 12290 6414 12292 6466
rect 12236 6412 12292 6414
rect 13132 7474 13188 7476
rect 13132 7422 13134 7474
rect 13134 7422 13186 7474
rect 13186 7422 13188 7474
rect 13132 7420 13188 7422
rect 12908 6690 12964 6692
rect 12908 6638 12910 6690
rect 12910 6638 12962 6690
rect 12962 6638 12964 6690
rect 12908 6636 12964 6638
rect 13244 6748 13300 6804
rect 12796 6524 12852 6580
rect 12460 5122 12516 5124
rect 12460 5070 12462 5122
rect 12462 5070 12514 5122
rect 12514 5070 12516 5122
rect 12460 5068 12516 5070
rect 12572 5010 12628 5012
rect 12572 4958 12574 5010
rect 12574 4958 12626 5010
rect 12626 4958 12628 5010
rect 12572 4956 12628 4958
rect 13804 7698 13860 7700
rect 13804 7646 13806 7698
rect 13806 7646 13858 7698
rect 13858 7646 13860 7698
rect 13804 7644 13860 7646
rect 13692 7474 13748 7476
rect 13692 7422 13694 7474
rect 13694 7422 13746 7474
rect 13746 7422 13748 7474
rect 13692 7420 13748 7422
rect 13580 6690 13636 6692
rect 13580 6638 13582 6690
rect 13582 6638 13634 6690
rect 13634 6638 13636 6690
rect 13580 6636 13636 6638
rect 13468 6300 13524 6356
rect 12348 4732 12404 4788
rect 12348 4226 12404 4228
rect 12348 4174 12350 4226
rect 12350 4174 12402 4226
rect 12402 4174 12404 4226
rect 12348 4172 12404 4174
rect 14588 12012 14644 12068
rect 14924 13020 14980 13076
rect 15596 13020 15652 13076
rect 15260 12908 15316 12964
rect 14812 11676 14868 11732
rect 15708 12962 15764 12964
rect 15708 12910 15710 12962
rect 15710 12910 15762 12962
rect 15762 12910 15764 12962
rect 15708 12908 15764 12910
rect 15820 12850 15876 12852
rect 15820 12798 15822 12850
rect 15822 12798 15874 12850
rect 15874 12798 15876 12850
rect 15820 12796 15876 12798
rect 15036 12178 15092 12180
rect 15036 12126 15038 12178
rect 15038 12126 15090 12178
rect 15090 12126 15092 12178
rect 15036 12124 15092 12126
rect 15036 11394 15092 11396
rect 15036 11342 15038 11394
rect 15038 11342 15090 11394
rect 15090 11342 15092 11394
rect 15036 11340 15092 11342
rect 15596 11170 15652 11172
rect 15596 11118 15598 11170
rect 15598 11118 15650 11170
rect 15650 11118 15652 11170
rect 15596 11116 15652 11118
rect 16380 12738 16436 12740
rect 16380 12686 16382 12738
rect 16382 12686 16434 12738
rect 16434 12686 16436 12738
rect 16380 12684 16436 12686
rect 16268 12402 16324 12404
rect 16268 12350 16270 12402
rect 16270 12350 16322 12402
rect 16322 12350 16324 12402
rect 16268 12348 16324 12350
rect 15932 12236 15988 12292
rect 16380 11676 16436 11732
rect 16044 11340 16100 11396
rect 14252 9772 14308 9828
rect 14476 9826 14532 9828
rect 14476 9774 14478 9826
rect 14478 9774 14530 9826
rect 14530 9774 14532 9826
rect 14476 9772 14532 9774
rect 14028 9602 14084 9604
rect 14028 9550 14030 9602
rect 14030 9550 14082 9602
rect 14082 9550 14084 9602
rect 14028 9548 14084 9550
rect 14252 9212 14308 9268
rect 14364 9436 14420 9492
rect 15708 10668 15764 10724
rect 14924 9714 14980 9716
rect 14924 9662 14926 9714
rect 14926 9662 14978 9714
rect 14978 9662 14980 9714
rect 14924 9660 14980 9662
rect 15260 9436 15316 9492
rect 15484 9212 15540 9268
rect 14588 8316 14644 8372
rect 14588 7644 14644 7700
rect 15148 8316 15204 8372
rect 14028 7420 14084 7476
rect 15708 9436 15764 9492
rect 15820 9548 15876 9604
rect 15820 9042 15876 9044
rect 15820 8990 15822 9042
rect 15822 8990 15874 9042
rect 15874 8990 15876 9042
rect 15820 8988 15876 8990
rect 16492 11452 16548 11508
rect 14028 6748 14084 6804
rect 14924 6636 14980 6692
rect 14252 6578 14308 6580
rect 14252 6526 14254 6578
rect 14254 6526 14306 6578
rect 14306 6526 14308 6578
rect 14252 6524 14308 6526
rect 13804 4732 13860 4788
rect 14812 4898 14868 4900
rect 14812 4846 14814 4898
rect 14814 4846 14866 4898
rect 14866 4846 14868 4898
rect 14812 4844 14868 4846
rect 15932 6636 15988 6692
rect 16716 13020 16772 13076
rect 17388 15986 17444 15988
rect 17388 15934 17390 15986
rect 17390 15934 17442 15986
rect 17442 15934 17444 15986
rect 17388 15932 17444 15934
rect 18060 15986 18116 15988
rect 18060 15934 18062 15986
rect 18062 15934 18114 15986
rect 18114 15934 18116 15986
rect 18060 15932 18116 15934
rect 18508 15932 18564 15988
rect 18732 16044 18788 16100
rect 19180 26012 19236 26068
rect 19964 26066 20020 26068
rect 19964 26014 19966 26066
rect 19966 26014 20018 26066
rect 20018 26014 20020 26066
rect 19964 26012 20020 26014
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20188 24780 20244 24836
rect 19852 23938 19908 23940
rect 19852 23886 19854 23938
rect 19854 23886 19906 23938
rect 19906 23886 19908 23938
rect 19852 23884 19908 23886
rect 20412 23938 20468 23940
rect 20412 23886 20414 23938
rect 20414 23886 20466 23938
rect 20466 23886 20468 23938
rect 20412 23884 20468 23886
rect 20524 26012 20580 26068
rect 19292 23660 19348 23716
rect 19068 20860 19124 20916
rect 19628 23714 19684 23716
rect 19628 23662 19630 23714
rect 19630 23662 19682 23714
rect 19682 23662 19684 23714
rect 19628 23660 19684 23662
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19292 23378 19348 23380
rect 19292 23326 19294 23378
rect 19294 23326 19346 23378
rect 19346 23326 19348 23378
rect 19292 23324 19348 23326
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19292 21308 19348 21364
rect 19740 20860 19796 20916
rect 19628 20802 19684 20804
rect 19628 20750 19630 20802
rect 19630 20750 19682 20802
rect 19682 20750 19684 20802
rect 19628 20748 19684 20750
rect 19516 20690 19572 20692
rect 19516 20638 19518 20690
rect 19518 20638 19570 20690
rect 19570 20638 19572 20690
rect 19516 20636 19572 20638
rect 19964 20524 20020 20580
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20188 20076 20244 20132
rect 20524 23212 20580 23268
rect 20412 20524 20468 20580
rect 20524 19852 20580 19908
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19292 18450 19348 18452
rect 19292 18398 19294 18450
rect 19294 18398 19346 18450
rect 19346 18398 19348 18450
rect 19292 18396 19348 18398
rect 19068 17724 19124 17780
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19180 16716 19236 16772
rect 20076 16156 20132 16212
rect 19628 16098 19684 16100
rect 19628 16046 19630 16098
rect 19630 16046 19682 16098
rect 19682 16046 19684 16098
rect 19628 16044 19684 16046
rect 19180 15932 19236 15988
rect 18844 15036 18900 15092
rect 17388 14476 17444 14532
rect 17276 14418 17332 14420
rect 17276 14366 17278 14418
rect 17278 14366 17330 14418
rect 17330 14366 17332 14418
rect 17276 14364 17332 14366
rect 17612 13356 17668 13412
rect 17500 13244 17556 13300
rect 17500 12402 17556 12404
rect 17500 12350 17502 12402
rect 17502 12350 17554 12402
rect 17554 12350 17556 12402
rect 17500 12348 17556 12350
rect 18172 12908 18228 12964
rect 17836 12684 17892 12740
rect 18060 12572 18116 12628
rect 16828 11004 16884 11060
rect 17836 12348 17892 12404
rect 16604 8316 16660 8372
rect 17388 10668 17444 10724
rect 17276 9826 17332 9828
rect 17276 9774 17278 9826
rect 17278 9774 17330 9826
rect 17330 9774 17332 9826
rect 17276 9772 17332 9774
rect 17052 7420 17108 7476
rect 16828 6412 16884 6468
rect 16940 6636 16996 6692
rect 16268 5292 16324 5348
rect 15708 4844 15764 4900
rect 15036 4732 15092 4788
rect 17052 6578 17108 6580
rect 17052 6526 17054 6578
rect 17054 6526 17106 6578
rect 17106 6526 17108 6578
rect 17052 6524 17108 6526
rect 18396 14252 18452 14308
rect 18620 14364 18676 14420
rect 18284 12572 18340 12628
rect 18508 12684 18564 12740
rect 17948 11506 18004 11508
rect 17948 11454 17950 11506
rect 17950 11454 18002 11506
rect 18002 11454 18004 11506
rect 17948 11452 18004 11454
rect 17836 9660 17892 9716
rect 17948 9772 18004 9828
rect 17948 9100 18004 9156
rect 17836 9042 17892 9044
rect 17836 8990 17838 9042
rect 17838 8990 17890 9042
rect 17890 8990 17892 9042
rect 17836 8988 17892 8990
rect 17500 8316 17556 8372
rect 17612 8034 17668 8036
rect 17612 7982 17614 8034
rect 17614 7982 17666 8034
rect 17666 7982 17668 8034
rect 17612 7980 17668 7982
rect 17500 6690 17556 6692
rect 17500 6638 17502 6690
rect 17502 6638 17554 6690
rect 17554 6638 17556 6690
rect 17500 6636 17556 6638
rect 17500 6412 17556 6468
rect 17164 6076 17220 6132
rect 18284 10722 18340 10724
rect 18284 10670 18286 10722
rect 18286 10670 18338 10722
rect 18338 10670 18340 10722
rect 18284 10668 18340 10670
rect 18844 14306 18900 14308
rect 18844 14254 18846 14306
rect 18846 14254 18898 14306
rect 18898 14254 18900 14306
rect 18844 14252 18900 14254
rect 18732 13634 18788 13636
rect 18732 13582 18734 13634
rect 18734 13582 18786 13634
rect 18786 13582 18788 13634
rect 18732 13580 18788 13582
rect 18732 12850 18788 12852
rect 18732 12798 18734 12850
rect 18734 12798 18786 12850
rect 18786 12798 18788 12850
rect 18732 12796 18788 12798
rect 18956 12572 19012 12628
rect 18844 12124 18900 12180
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20860 24834 20916 24836
rect 20860 24782 20862 24834
rect 20862 24782 20914 24834
rect 20914 24782 20916 24834
rect 20860 24780 20916 24782
rect 22988 28028 23044 28084
rect 22204 27970 22260 27972
rect 22204 27918 22206 27970
rect 22206 27918 22258 27970
rect 22258 27918 22260 27970
rect 22204 27916 22260 27918
rect 22876 27858 22932 27860
rect 22876 27806 22878 27858
rect 22878 27806 22930 27858
rect 22930 27806 22932 27858
rect 22876 27804 22932 27806
rect 21868 27074 21924 27076
rect 21868 27022 21870 27074
rect 21870 27022 21922 27074
rect 21922 27022 21924 27074
rect 21868 27020 21924 27022
rect 22540 27074 22596 27076
rect 22540 27022 22542 27074
rect 22542 27022 22594 27074
rect 22594 27022 22596 27074
rect 22540 27020 22596 27022
rect 21196 22428 21252 22484
rect 21308 21308 21364 21364
rect 21308 21026 21364 21028
rect 21308 20974 21310 21026
rect 21310 20974 21362 21026
rect 21362 20974 21364 21026
rect 21308 20972 21364 20974
rect 21420 20690 21476 20692
rect 21420 20638 21422 20690
rect 21422 20638 21474 20690
rect 21474 20638 21476 20690
rect 21420 20636 21476 20638
rect 20972 20076 21028 20132
rect 21644 19906 21700 19908
rect 21644 19854 21646 19906
rect 21646 19854 21698 19906
rect 21698 19854 21700 19906
rect 21644 19852 21700 19854
rect 20748 17666 20804 17668
rect 20748 17614 20750 17666
rect 20750 17614 20802 17666
rect 20802 17614 20804 17666
rect 20748 17612 20804 17614
rect 22092 23212 22148 23268
rect 22092 21868 22148 21924
rect 21980 20972 22036 21028
rect 22876 24556 22932 24612
rect 23100 23884 23156 23940
rect 22652 22482 22708 22484
rect 22652 22430 22654 22482
rect 22654 22430 22706 22482
rect 22706 22430 22708 22482
rect 22652 22428 22708 22430
rect 23100 22428 23156 22484
rect 22876 22092 22932 22148
rect 23100 21980 23156 22036
rect 22092 20690 22148 20692
rect 22092 20638 22094 20690
rect 22094 20638 22146 20690
rect 22146 20638 22148 20690
rect 22092 20636 22148 20638
rect 22540 20300 22596 20356
rect 22316 20018 22372 20020
rect 22316 19966 22318 20018
rect 22318 19966 22370 20018
rect 22370 19966 22372 20018
rect 22316 19964 22372 19966
rect 22204 18060 22260 18116
rect 22876 20300 22932 20356
rect 22988 20636 23044 20692
rect 23100 20748 23156 20804
rect 22876 18060 22932 18116
rect 23100 17948 23156 18004
rect 20972 16940 21028 16996
rect 21868 16940 21924 16996
rect 20636 16716 20692 16772
rect 21756 16380 21812 16436
rect 21420 16156 21476 16212
rect 21644 16044 21700 16100
rect 20524 15932 20580 15988
rect 20188 15314 20244 15316
rect 20188 15262 20190 15314
rect 20190 15262 20242 15314
rect 20242 15262 20244 15314
rect 20188 15260 20244 15262
rect 19516 15036 19572 15092
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20972 15314 21028 15316
rect 20972 15262 20974 15314
rect 20974 15262 21026 15314
rect 21026 15262 21028 15314
rect 20972 15260 21028 15262
rect 22540 17554 22596 17556
rect 22540 17502 22542 17554
rect 22542 17502 22594 17554
rect 22594 17502 22596 17554
rect 22540 17500 22596 17502
rect 22428 16268 22484 16324
rect 23100 16268 23156 16324
rect 21980 16044 22036 16100
rect 22092 16156 22148 16212
rect 22876 16098 22932 16100
rect 22876 16046 22878 16098
rect 22878 16046 22930 16098
rect 22930 16046 22932 16098
rect 22876 16044 22932 16046
rect 21756 14812 21812 14868
rect 19628 12796 19684 12852
rect 19404 12236 19460 12292
rect 19292 12124 19348 12180
rect 18956 11282 19012 11284
rect 18956 11230 18958 11282
rect 18958 11230 19010 11282
rect 19010 11230 19012 11282
rect 18956 11228 19012 11230
rect 18396 10556 18452 10612
rect 19068 10556 19124 10612
rect 19180 9154 19236 9156
rect 19180 9102 19182 9154
rect 19182 9102 19234 9154
rect 19234 9102 19236 9154
rect 19180 9100 19236 9102
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19740 12178 19796 12180
rect 19740 12126 19742 12178
rect 19742 12126 19794 12178
rect 19794 12126 19796 12178
rect 19740 12124 19796 12126
rect 19516 11452 19572 11508
rect 19628 11116 19684 11172
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 21420 13580 21476 13636
rect 21420 12460 21476 12516
rect 21196 12066 21252 12068
rect 21196 12014 21198 12066
rect 21198 12014 21250 12066
rect 21250 12014 21252 12066
rect 21196 12012 21252 12014
rect 22092 13244 22148 13300
rect 21980 12348 22036 12404
rect 21532 12236 21588 12292
rect 22204 12684 22260 12740
rect 22428 12850 22484 12852
rect 22428 12798 22430 12850
rect 22430 12798 22482 12850
rect 22482 12798 22484 12850
rect 22428 12796 22484 12798
rect 22316 12236 22372 12292
rect 21756 11394 21812 11396
rect 21756 11342 21758 11394
rect 21758 11342 21810 11394
rect 21810 11342 21812 11394
rect 21756 11340 21812 11342
rect 22540 11340 22596 11396
rect 23436 27020 23492 27076
rect 23660 28700 23716 28756
rect 26012 33068 26068 33124
rect 25788 32060 25844 32116
rect 26236 35308 26292 35364
rect 26684 35196 26740 35252
rect 26460 33458 26516 33460
rect 26460 33406 26462 33458
rect 26462 33406 26514 33458
rect 26514 33406 26516 33458
rect 26460 33404 26516 33406
rect 27468 35196 27524 35252
rect 28364 38162 28420 38164
rect 28364 38110 28366 38162
rect 28366 38110 28418 38162
rect 28418 38110 28420 38162
rect 28364 38108 28420 38110
rect 30828 45218 30884 45220
rect 30828 45166 30830 45218
rect 30830 45166 30882 45218
rect 30882 45166 30884 45218
rect 30828 45164 30884 45166
rect 30940 44434 30996 44436
rect 30940 44382 30942 44434
rect 30942 44382 30994 44434
rect 30994 44382 30996 44434
rect 30940 44380 30996 44382
rect 31164 44098 31220 44100
rect 31164 44046 31166 44098
rect 31166 44046 31218 44098
rect 31218 44046 31220 44098
rect 31164 44044 31220 44046
rect 30828 43538 30884 43540
rect 30828 43486 30830 43538
rect 30830 43486 30882 43538
rect 30882 43486 30884 43538
rect 30828 43484 30884 43486
rect 31276 43426 31332 43428
rect 31276 43374 31278 43426
rect 31278 43374 31330 43426
rect 31330 43374 31332 43426
rect 31276 43372 31332 43374
rect 31276 42866 31332 42868
rect 31276 42814 31278 42866
rect 31278 42814 31330 42866
rect 31330 42814 31332 42866
rect 31276 42812 31332 42814
rect 30828 41916 30884 41972
rect 31836 45218 31892 45220
rect 31836 45166 31838 45218
rect 31838 45166 31890 45218
rect 31890 45166 31892 45218
rect 31836 45164 31892 45166
rect 31500 43820 31556 43876
rect 32172 45218 32228 45220
rect 32172 45166 32174 45218
rect 32174 45166 32226 45218
rect 32226 45166 32228 45218
rect 32172 45164 32228 45166
rect 32508 45666 32564 45668
rect 32508 45614 32510 45666
rect 32510 45614 32562 45666
rect 32562 45614 32564 45666
rect 32508 45612 32564 45614
rect 31836 44322 31892 44324
rect 31836 44270 31838 44322
rect 31838 44270 31890 44322
rect 31890 44270 31892 44322
rect 31836 44268 31892 44270
rect 31948 45052 32004 45108
rect 31612 43708 31668 43764
rect 31724 43538 31780 43540
rect 31724 43486 31726 43538
rect 31726 43486 31778 43538
rect 31778 43486 31780 43538
rect 31724 43484 31780 43486
rect 31500 43372 31556 43428
rect 32172 44492 32228 44548
rect 32620 44322 32676 44324
rect 32620 44270 32622 44322
rect 32622 44270 32674 44322
rect 32674 44270 32676 44322
rect 32620 44268 32676 44270
rect 32396 44044 32452 44100
rect 32284 43372 32340 43428
rect 30940 41804 30996 41860
rect 30828 41186 30884 41188
rect 30828 41134 30830 41186
rect 30830 41134 30882 41186
rect 30882 41134 30884 41186
rect 30828 41132 30884 41134
rect 29820 40908 29876 40964
rect 30604 40402 30660 40404
rect 30604 40350 30606 40402
rect 30606 40350 30658 40402
rect 30658 40350 30660 40402
rect 30604 40348 30660 40350
rect 30940 40908 30996 40964
rect 29260 40236 29316 40292
rect 29036 38108 29092 38164
rect 30268 38668 30324 38724
rect 29260 38050 29316 38052
rect 29260 37998 29262 38050
rect 29262 37998 29314 38050
rect 29314 37998 29316 38050
rect 29260 37996 29316 37998
rect 28588 36482 28644 36484
rect 28588 36430 28590 36482
rect 28590 36430 28642 36482
rect 28642 36430 28644 36482
rect 28588 36428 28644 36430
rect 29260 36428 29316 36484
rect 29820 36482 29876 36484
rect 29820 36430 29822 36482
rect 29822 36430 29874 36482
rect 29874 36430 29876 36482
rect 29820 36428 29876 36430
rect 29148 35868 29204 35924
rect 27916 33404 27972 33460
rect 28476 34636 28532 34692
rect 26348 33122 26404 33124
rect 26348 33070 26350 33122
rect 26350 33070 26402 33122
rect 26402 33070 26404 33122
rect 26348 33068 26404 33070
rect 27132 32786 27188 32788
rect 27132 32734 27134 32786
rect 27134 32734 27186 32786
rect 27186 32734 27188 32786
rect 27132 32732 27188 32734
rect 27804 32732 27860 32788
rect 30156 35868 30212 35924
rect 32508 43932 32564 43988
rect 32956 44940 33012 44996
rect 33180 43426 33236 43428
rect 33180 43374 33182 43426
rect 33182 43374 33234 43426
rect 33234 43374 33236 43426
rect 33180 43372 33236 43374
rect 32844 42700 32900 42756
rect 31948 41804 32004 41860
rect 31836 41186 31892 41188
rect 31836 41134 31838 41186
rect 31838 41134 31890 41186
rect 31890 41134 31892 41186
rect 31836 41132 31892 41134
rect 33292 42252 33348 42308
rect 33180 41858 33236 41860
rect 33180 41806 33182 41858
rect 33182 41806 33234 41858
rect 33234 41806 33236 41858
rect 33180 41804 33236 41806
rect 32508 40348 32564 40404
rect 32396 39116 32452 39172
rect 31948 39004 32004 39060
rect 32508 39058 32564 39060
rect 32508 39006 32510 39058
rect 32510 39006 32562 39058
rect 32562 39006 32564 39058
rect 32508 39004 32564 39006
rect 33180 38946 33236 38948
rect 33180 38894 33182 38946
rect 33182 38894 33234 38946
rect 33234 38894 33236 38946
rect 33180 38892 33236 38894
rect 33068 38722 33124 38724
rect 33068 38670 33070 38722
rect 33070 38670 33122 38722
rect 33122 38670 33124 38722
rect 33068 38668 33124 38670
rect 33516 44098 33572 44100
rect 33516 44046 33518 44098
rect 33518 44046 33570 44098
rect 33570 44046 33572 44098
rect 33516 44044 33572 44046
rect 33852 43932 33908 43988
rect 33628 43708 33684 43764
rect 33628 43260 33684 43316
rect 33740 43484 33796 43540
rect 33516 42642 33572 42644
rect 33516 42590 33518 42642
rect 33518 42590 33570 42642
rect 33570 42590 33572 42642
rect 33516 42588 33572 42590
rect 33852 43372 33908 43428
rect 33852 42754 33908 42756
rect 33852 42702 33854 42754
rect 33854 42702 33906 42754
rect 33906 42702 33908 42754
rect 33852 42700 33908 42702
rect 33740 42028 33796 42084
rect 33516 41804 33572 41860
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 34972 46060 35028 46116
rect 36988 46114 37044 46116
rect 36988 46062 36990 46114
rect 36990 46062 37042 46114
rect 37042 46062 37044 46114
rect 36988 46060 37044 46062
rect 40348 46060 40404 46116
rect 34076 44380 34132 44436
rect 34300 45612 34356 45668
rect 35196 45388 35252 45444
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34524 43650 34580 43652
rect 34524 43598 34526 43650
rect 34526 43598 34578 43650
rect 34578 43598 34580 43650
rect 34524 43596 34580 43598
rect 34412 43372 34468 43428
rect 34524 42028 34580 42084
rect 34300 41692 34356 41748
rect 34076 40796 34132 40852
rect 33404 39900 33460 39956
rect 33404 39340 33460 39396
rect 33516 39116 33572 39172
rect 31724 37996 31780 38052
rect 30492 35196 30548 35252
rect 32508 35586 32564 35588
rect 32508 35534 32510 35586
rect 32510 35534 32562 35586
rect 32562 35534 32564 35586
rect 32508 35532 32564 35534
rect 31724 34748 31780 34804
rect 32060 34130 32116 34132
rect 32060 34078 32062 34130
rect 32062 34078 32114 34130
rect 32114 34078 32116 34130
rect 32060 34076 32116 34078
rect 28476 32562 28532 32564
rect 28476 32510 28478 32562
rect 28478 32510 28530 32562
rect 28530 32510 28532 32562
rect 28476 32508 28532 32510
rect 29260 32620 29316 32676
rect 28812 31948 28868 32004
rect 26796 31388 26852 31444
rect 26796 30882 26852 30884
rect 26796 30830 26798 30882
rect 26798 30830 26850 30882
rect 26850 30830 26852 30882
rect 26796 30828 26852 30830
rect 25116 30210 25172 30212
rect 25116 30158 25118 30210
rect 25118 30158 25170 30210
rect 25170 30158 25172 30210
rect 25116 30156 25172 30158
rect 24892 28700 24948 28756
rect 23548 24610 23604 24612
rect 23548 24558 23550 24610
rect 23550 24558 23602 24610
rect 23602 24558 23604 24610
rect 23548 24556 23604 24558
rect 23548 23996 23604 24052
rect 24220 23884 24276 23940
rect 24332 27468 24388 27524
rect 24668 27132 24724 27188
rect 25340 28588 25396 28644
rect 25340 27468 25396 27524
rect 24668 24722 24724 24724
rect 24668 24670 24670 24722
rect 24670 24670 24722 24722
rect 24722 24670 24724 24722
rect 24668 24668 24724 24670
rect 24332 22428 24388 22484
rect 25788 27468 25844 27524
rect 26012 27298 26068 27300
rect 26012 27246 26014 27298
rect 26014 27246 26066 27298
rect 26066 27246 26068 27298
rect 26012 27244 26068 27246
rect 26796 28588 26852 28644
rect 30268 33122 30324 33124
rect 30268 33070 30270 33122
rect 30270 33070 30322 33122
rect 30322 33070 30324 33122
rect 30268 33068 30324 33070
rect 29484 31836 29540 31892
rect 29820 32508 29876 32564
rect 29708 31778 29764 31780
rect 29708 31726 29710 31778
rect 29710 31726 29762 31778
rect 29762 31726 29764 31778
rect 29708 31724 29764 31726
rect 29596 31554 29652 31556
rect 29596 31502 29598 31554
rect 29598 31502 29650 31554
rect 29650 31502 29652 31554
rect 29596 31500 29652 31502
rect 29484 31388 29540 31444
rect 29372 31276 29428 31332
rect 29260 31218 29316 31220
rect 29260 31166 29262 31218
rect 29262 31166 29314 31218
rect 29314 31166 29316 31218
rect 29260 31164 29316 31166
rect 29372 30994 29428 30996
rect 29372 30942 29374 30994
rect 29374 30942 29426 30994
rect 29426 30942 29428 30994
rect 29372 30940 29428 30942
rect 29596 29314 29652 29316
rect 29596 29262 29598 29314
rect 29598 29262 29650 29314
rect 29650 29262 29652 29314
rect 29596 29260 29652 29262
rect 29148 28642 29204 28644
rect 29148 28590 29150 28642
rect 29150 28590 29202 28642
rect 29202 28590 29204 28642
rect 29148 28588 29204 28590
rect 28924 28364 28980 28420
rect 28140 27746 28196 27748
rect 28140 27694 28142 27746
rect 28142 27694 28194 27746
rect 28194 27694 28196 27746
rect 28140 27692 28196 27694
rect 29260 27804 29316 27860
rect 28924 27692 28980 27748
rect 29148 27746 29204 27748
rect 29148 27694 29150 27746
rect 29150 27694 29202 27746
rect 29202 27694 29204 27746
rect 29148 27692 29204 27694
rect 28588 27244 28644 27300
rect 26572 26460 26628 26516
rect 25340 24780 25396 24836
rect 25228 24722 25284 24724
rect 25228 24670 25230 24722
rect 25230 24670 25282 24722
rect 25282 24670 25284 24722
rect 25228 24668 25284 24670
rect 29596 27074 29652 27076
rect 29596 27022 29598 27074
rect 29598 27022 29650 27074
rect 29650 27022 29652 27074
rect 29596 27020 29652 27022
rect 28588 25116 28644 25172
rect 23660 22146 23716 22148
rect 23660 22094 23662 22146
rect 23662 22094 23714 22146
rect 23714 22094 23716 22146
rect 23660 22092 23716 22094
rect 23548 21980 23604 22036
rect 23436 20802 23492 20804
rect 23436 20750 23438 20802
rect 23438 20750 23490 20802
rect 23490 20750 23492 20802
rect 23436 20748 23492 20750
rect 23324 20300 23380 20356
rect 23436 20412 23492 20468
rect 23884 20578 23940 20580
rect 23884 20526 23886 20578
rect 23886 20526 23938 20578
rect 23938 20526 23940 20578
rect 23884 20524 23940 20526
rect 23996 21868 24052 21924
rect 25452 23938 25508 23940
rect 25452 23886 25454 23938
rect 25454 23886 25506 23938
rect 25506 23886 25508 23938
rect 25452 23884 25508 23886
rect 25676 23938 25732 23940
rect 25676 23886 25678 23938
rect 25678 23886 25730 23938
rect 25730 23886 25732 23938
rect 25676 23884 25732 23886
rect 26684 23938 26740 23940
rect 26684 23886 26686 23938
rect 26686 23886 26738 23938
rect 26738 23886 26740 23938
rect 26684 23884 26740 23886
rect 30604 31948 30660 32004
rect 30156 31890 30212 31892
rect 30156 31838 30158 31890
rect 30158 31838 30210 31890
rect 30210 31838 30212 31890
rect 30156 31836 30212 31838
rect 30044 31554 30100 31556
rect 30044 31502 30046 31554
rect 30046 31502 30098 31554
rect 30098 31502 30100 31554
rect 30044 31500 30100 31502
rect 30268 31554 30324 31556
rect 30268 31502 30270 31554
rect 30270 31502 30322 31554
rect 30322 31502 30324 31554
rect 30268 31500 30324 31502
rect 29932 31276 29988 31332
rect 30268 31276 30324 31332
rect 30828 33234 30884 33236
rect 30828 33182 30830 33234
rect 30830 33182 30882 33234
rect 30882 33182 30884 33234
rect 30828 33180 30884 33182
rect 31164 33180 31220 33236
rect 31052 32956 31108 33012
rect 31052 32620 31108 32676
rect 30828 31388 30884 31444
rect 30156 31218 30212 31220
rect 30156 31166 30158 31218
rect 30158 31166 30210 31218
rect 30210 31166 30212 31218
rect 30156 31164 30212 31166
rect 30268 30882 30324 30884
rect 30268 30830 30270 30882
rect 30270 30830 30322 30882
rect 30322 30830 30324 30882
rect 30268 30828 30324 30830
rect 30492 30940 30548 30996
rect 30604 30828 30660 30884
rect 30268 30044 30324 30100
rect 33404 35532 33460 35588
rect 32620 34802 32676 34804
rect 32620 34750 32622 34802
rect 32622 34750 32674 34802
rect 32674 34750 32676 34802
rect 32620 34748 32676 34750
rect 33180 34636 33236 34692
rect 33180 33292 33236 33348
rect 33292 33404 33348 33460
rect 31388 32956 31444 33012
rect 32844 32956 32900 33012
rect 31612 32508 31668 32564
rect 31276 31948 31332 32004
rect 31500 32002 31556 32004
rect 31500 31950 31502 32002
rect 31502 31950 31554 32002
rect 31554 31950 31556 32002
rect 31500 31948 31556 31950
rect 31500 31724 31556 31780
rect 31164 31388 31220 31444
rect 30940 30044 30996 30100
rect 33740 39900 33796 39956
rect 34412 39676 34468 39732
rect 34188 39004 34244 39060
rect 33852 38946 33908 38948
rect 33852 38894 33854 38946
rect 33854 38894 33906 38946
rect 33906 38894 33908 38946
rect 33852 38892 33908 38894
rect 34748 42194 34804 42196
rect 34748 42142 34750 42194
rect 34750 42142 34802 42194
rect 34802 42142 34804 42194
rect 34748 42140 34804 42142
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35420 42252 35476 42308
rect 39228 45836 39284 45892
rect 38220 45724 38276 45780
rect 36428 44882 36484 44884
rect 36428 44830 36430 44882
rect 36430 44830 36482 44882
rect 36482 44830 36484 44882
rect 36428 44828 36484 44830
rect 36764 44716 36820 44772
rect 36204 42978 36260 42980
rect 36204 42926 36206 42978
rect 36206 42926 36258 42978
rect 36258 42926 36260 42978
rect 36204 42924 36260 42926
rect 35980 42140 36036 42196
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 34636 41132 34692 41188
rect 34636 39340 34692 39396
rect 33964 37938 34020 37940
rect 33964 37886 33966 37938
rect 33966 37886 34018 37938
rect 34018 37886 34020 37938
rect 33964 37884 34020 37886
rect 35084 40908 35140 40964
rect 35532 41186 35588 41188
rect 35532 41134 35534 41186
rect 35534 41134 35586 41186
rect 35586 41134 35588 41186
rect 35532 41132 35588 41134
rect 35084 40572 35140 40628
rect 35420 40402 35476 40404
rect 35420 40350 35422 40402
rect 35422 40350 35474 40402
rect 35474 40350 35476 40402
rect 35420 40348 35476 40350
rect 34860 39788 34916 39844
rect 34860 37884 34916 37940
rect 34748 35644 34804 35700
rect 34412 34802 34468 34804
rect 34412 34750 34414 34802
rect 34414 34750 34466 34802
rect 34466 34750 34468 34802
rect 34412 34748 34468 34750
rect 33628 34130 33684 34132
rect 33628 34078 33630 34130
rect 33630 34078 33682 34130
rect 33682 34078 33684 34130
rect 33628 34076 33684 34078
rect 33628 33516 33684 33572
rect 33628 33068 33684 33124
rect 33516 32844 33572 32900
rect 33292 32562 33348 32564
rect 33292 32510 33294 32562
rect 33294 32510 33346 32562
rect 33346 32510 33348 32562
rect 33292 32508 33348 32510
rect 33516 32562 33572 32564
rect 33516 32510 33518 32562
rect 33518 32510 33570 32562
rect 33570 32510 33572 32562
rect 33516 32508 33572 32510
rect 33964 31836 34020 31892
rect 33068 31778 33124 31780
rect 33068 31726 33070 31778
rect 33070 31726 33122 31778
rect 33122 31726 33124 31778
rect 33068 31724 33124 31726
rect 33292 31500 33348 31556
rect 32396 31388 32452 31444
rect 32060 31164 32116 31220
rect 31500 30828 31556 30884
rect 31500 30098 31556 30100
rect 31500 30046 31502 30098
rect 31502 30046 31554 30098
rect 31554 30046 31556 30098
rect 31500 30044 31556 30046
rect 31836 29708 31892 29764
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35644 40572 35700 40628
rect 35644 40402 35700 40404
rect 35644 40350 35646 40402
rect 35646 40350 35698 40402
rect 35698 40350 35700 40402
rect 35644 40348 35700 40350
rect 35756 40236 35812 40292
rect 36540 41858 36596 41860
rect 36540 41806 36542 41858
rect 36542 41806 36594 41858
rect 36594 41806 36596 41858
rect 36540 41804 36596 41806
rect 37772 44492 37828 44548
rect 36988 43820 37044 43876
rect 37772 44210 37828 44212
rect 37772 44158 37774 44210
rect 37774 44158 37826 44210
rect 37826 44158 37828 44210
rect 37772 44156 37828 44158
rect 37996 44268 38052 44324
rect 37436 43372 37492 43428
rect 37212 43314 37268 43316
rect 37212 43262 37214 43314
rect 37214 43262 37266 43314
rect 37266 43262 37268 43314
rect 37212 43260 37268 43262
rect 37100 43148 37156 43204
rect 37436 43148 37492 43204
rect 37772 42588 37828 42644
rect 38444 45052 38500 45108
rect 38780 44044 38836 44100
rect 38332 43596 38388 43652
rect 39788 45778 39844 45780
rect 39788 45726 39790 45778
rect 39790 45726 39842 45778
rect 39842 45726 39844 45778
rect 39788 45724 39844 45726
rect 41468 46114 41524 46116
rect 41468 46062 41470 46114
rect 41470 46062 41522 46114
rect 41522 46062 41524 46114
rect 41468 46060 41524 46062
rect 41692 46060 41748 46116
rect 41020 45276 41076 45332
rect 42252 45330 42308 45332
rect 42252 45278 42254 45330
rect 42254 45278 42306 45330
rect 42306 45278 42308 45330
rect 42252 45276 42308 45278
rect 41132 45164 41188 45220
rect 40124 44882 40180 44884
rect 40124 44830 40126 44882
rect 40126 44830 40178 44882
rect 40178 44830 40180 44882
rect 40124 44828 40180 44830
rect 42364 44940 42420 44996
rect 44044 47740 44100 47796
rect 43708 45890 43764 45892
rect 43708 45838 43710 45890
rect 43710 45838 43762 45890
rect 43762 45838 43764 45890
rect 43708 45836 43764 45838
rect 43036 44492 43092 44548
rect 43932 44380 43988 44436
rect 41692 44322 41748 44324
rect 41692 44270 41694 44322
rect 41694 44270 41746 44322
rect 41746 44270 41748 44322
rect 41692 44268 41748 44270
rect 41244 44156 41300 44212
rect 42812 44156 42868 44212
rect 38892 43596 38948 43652
rect 41244 43596 41300 43652
rect 38668 43484 38724 43540
rect 41244 43372 41300 43428
rect 40124 43036 40180 43092
rect 37100 41804 37156 41860
rect 36204 40236 36260 40292
rect 36428 41132 36484 41188
rect 36540 40348 36596 40404
rect 36988 40236 37044 40292
rect 35644 39228 35700 39284
rect 37772 41916 37828 41972
rect 37548 41804 37604 41860
rect 37436 40402 37492 40404
rect 37436 40350 37438 40402
rect 37438 40350 37490 40402
rect 37490 40350 37492 40402
rect 37436 40348 37492 40350
rect 36652 39058 36708 39060
rect 36652 39006 36654 39058
rect 36654 39006 36706 39058
rect 36706 39006 36708 39058
rect 36652 39004 36708 39006
rect 36988 38780 37044 38836
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35084 37100 35140 37156
rect 36092 38162 36148 38164
rect 36092 38110 36094 38162
rect 36094 38110 36146 38162
rect 36146 38110 36148 38162
rect 36092 38108 36148 38110
rect 36092 37490 36148 37492
rect 36092 37438 36094 37490
rect 36094 37438 36146 37490
rect 36146 37438 36148 37490
rect 36092 37436 36148 37438
rect 35420 37378 35476 37380
rect 35420 37326 35422 37378
rect 35422 37326 35474 37378
rect 35474 37326 35476 37378
rect 35420 37324 35476 37326
rect 35980 37266 36036 37268
rect 35980 37214 35982 37266
rect 35982 37214 36034 37266
rect 36034 37214 36036 37266
rect 35980 37212 36036 37214
rect 35644 37100 35700 37156
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 34972 35532 35028 35588
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 36988 38162 37044 38164
rect 36988 38110 36990 38162
rect 36990 38110 37042 38162
rect 37042 38110 37044 38162
rect 36988 38108 37044 38110
rect 37772 39788 37828 39844
rect 37324 39394 37380 39396
rect 37324 39342 37326 39394
rect 37326 39342 37378 39394
rect 37378 39342 37380 39394
rect 37324 39340 37380 39342
rect 37212 39004 37268 39060
rect 37772 39004 37828 39060
rect 38108 41692 38164 41748
rect 38668 42140 38724 42196
rect 39228 42588 39284 42644
rect 39228 42194 39284 42196
rect 39228 42142 39230 42194
rect 39230 42142 39282 42194
rect 39282 42142 39284 42194
rect 39228 42140 39284 42142
rect 39004 42082 39060 42084
rect 39004 42030 39006 42082
rect 39006 42030 39058 42082
rect 39058 42030 39060 42082
rect 39004 42028 39060 42030
rect 39116 41858 39172 41860
rect 39116 41806 39118 41858
rect 39118 41806 39170 41858
rect 39170 41806 39172 41858
rect 39116 41804 39172 41806
rect 39788 41916 39844 41972
rect 40124 42476 40180 42532
rect 41132 42252 41188 42308
rect 40348 41804 40404 41860
rect 40796 42028 40852 42084
rect 39676 41692 39732 41748
rect 39452 41468 39508 41524
rect 38780 41186 38836 41188
rect 38780 41134 38782 41186
rect 38782 41134 38834 41186
rect 38834 41134 38836 41186
rect 38780 41132 38836 41134
rect 40684 40572 40740 40628
rect 39676 40124 39732 40180
rect 40236 40348 40292 40404
rect 40012 39788 40068 39844
rect 38108 39116 38164 39172
rect 38444 39004 38500 39060
rect 37996 38946 38052 38948
rect 37996 38894 37998 38946
rect 37998 38894 38050 38946
rect 38050 38894 38052 38946
rect 37996 38892 38052 38894
rect 38332 38834 38388 38836
rect 38332 38782 38334 38834
rect 38334 38782 38386 38834
rect 38386 38782 38388 38834
rect 38332 38780 38388 38782
rect 38668 39058 38724 39060
rect 38668 39006 38670 39058
rect 38670 39006 38722 39058
rect 38722 39006 38724 39058
rect 38668 39004 38724 39006
rect 39340 39228 39396 39284
rect 37324 36876 37380 36932
rect 37100 36204 37156 36260
rect 36316 35868 36372 35924
rect 36876 35922 36932 35924
rect 36876 35870 36878 35922
rect 36878 35870 36930 35922
rect 36930 35870 36932 35922
rect 36876 35868 36932 35870
rect 36652 35810 36708 35812
rect 36652 35758 36654 35810
rect 36654 35758 36706 35810
rect 36706 35758 36708 35810
rect 36652 35756 36708 35758
rect 35644 34860 35700 34916
rect 34860 34748 34916 34804
rect 34748 34412 34804 34468
rect 36764 35586 36820 35588
rect 36764 35534 36766 35586
rect 36766 35534 36818 35586
rect 36818 35534 36820 35586
rect 36764 35532 36820 35534
rect 36652 34300 36708 34356
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 36988 34690 37044 34692
rect 36988 34638 36990 34690
rect 36990 34638 37042 34690
rect 37042 34638 37044 34690
rect 36988 34636 37044 34638
rect 36876 33740 36932 33796
rect 37436 34354 37492 34356
rect 37436 34302 37438 34354
rect 37438 34302 37490 34354
rect 37490 34302 37492 34354
rect 37436 34300 37492 34302
rect 36764 33628 36820 33684
rect 34748 33404 34804 33460
rect 34300 33234 34356 33236
rect 34300 33182 34302 33234
rect 34302 33182 34354 33234
rect 34354 33182 34356 33234
rect 34300 33180 34356 33182
rect 33740 31388 33796 31444
rect 33740 30828 33796 30884
rect 32508 30210 32564 30212
rect 32508 30158 32510 30210
rect 32510 30158 32562 30210
rect 32562 30158 32564 30210
rect 32508 30156 32564 30158
rect 32844 30044 32900 30100
rect 33068 30156 33124 30212
rect 32508 29708 32564 29764
rect 31052 29260 31108 29316
rect 33180 29314 33236 29316
rect 33180 29262 33182 29314
rect 33182 29262 33234 29314
rect 33234 29262 33236 29314
rect 33180 29260 33236 29262
rect 34972 33346 35028 33348
rect 34972 33294 34974 33346
rect 34974 33294 35026 33346
rect 35026 33294 35028 33346
rect 34972 33292 35028 33294
rect 34524 32956 34580 33012
rect 36316 33346 36372 33348
rect 36316 33294 36318 33346
rect 36318 33294 36370 33346
rect 36370 33294 36372 33346
rect 36316 33292 36372 33294
rect 35532 33234 35588 33236
rect 35532 33182 35534 33234
rect 35534 33182 35586 33234
rect 35586 33182 35588 33234
rect 35532 33180 35588 33182
rect 35756 33122 35812 33124
rect 35756 33070 35758 33122
rect 35758 33070 35810 33122
rect 35810 33070 35812 33122
rect 35756 33068 35812 33070
rect 35532 32508 35588 32564
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 36204 33234 36260 33236
rect 36204 33182 36206 33234
rect 36206 33182 36258 33234
rect 36258 33182 36260 33234
rect 36204 33180 36260 33182
rect 36988 33068 37044 33124
rect 37212 32732 37268 32788
rect 35868 31948 35924 32004
rect 35532 31836 35588 31892
rect 37100 31890 37156 31892
rect 37100 31838 37102 31890
rect 37102 31838 37154 31890
rect 37154 31838 37156 31890
rect 37100 31836 37156 31838
rect 35644 31724 35700 31780
rect 35084 31554 35140 31556
rect 35084 31502 35086 31554
rect 35086 31502 35138 31554
rect 35138 31502 35140 31554
rect 35084 31500 35140 31502
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34860 30380 34916 30436
rect 34300 29820 34356 29876
rect 35756 31106 35812 31108
rect 35756 31054 35758 31106
rect 35758 31054 35810 31106
rect 35810 31054 35812 31106
rect 35756 31052 35812 31054
rect 36092 30770 36148 30772
rect 36092 30718 36094 30770
rect 36094 30718 36146 30770
rect 36146 30718 36148 30770
rect 36092 30716 36148 30718
rect 35644 30434 35700 30436
rect 35644 30382 35646 30434
rect 35646 30382 35698 30434
rect 35698 30382 35700 30434
rect 35644 30380 35700 30382
rect 35308 30210 35364 30212
rect 35308 30158 35310 30210
rect 35310 30158 35362 30210
rect 35362 30158 35364 30210
rect 35308 30156 35364 30158
rect 35644 29538 35700 29540
rect 35644 29486 35646 29538
rect 35646 29486 35698 29538
rect 35698 29486 35700 29538
rect 35644 29484 35700 29486
rect 36092 30098 36148 30100
rect 36092 30046 36094 30098
rect 36094 30046 36146 30098
rect 36146 30046 36148 30098
rect 36092 30044 36148 30046
rect 35980 29986 36036 29988
rect 35980 29934 35982 29986
rect 35982 29934 36034 29986
rect 36034 29934 36036 29986
rect 35980 29932 36036 29934
rect 35868 29484 35924 29540
rect 36092 29426 36148 29428
rect 36092 29374 36094 29426
rect 36094 29374 36146 29426
rect 36146 29374 36148 29426
rect 36092 29372 36148 29374
rect 33740 29260 33796 29316
rect 32172 29202 32228 29204
rect 32172 29150 32174 29202
rect 32174 29150 32226 29202
rect 32226 29150 32228 29202
rect 32172 29148 32228 29150
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 30380 27746 30436 27748
rect 30380 27694 30382 27746
rect 30382 27694 30434 27746
rect 30434 27694 30436 27746
rect 30380 27692 30436 27694
rect 30828 27746 30884 27748
rect 30828 27694 30830 27746
rect 30830 27694 30882 27746
rect 30882 27694 30884 27746
rect 30828 27692 30884 27694
rect 31388 27746 31444 27748
rect 31388 27694 31390 27746
rect 31390 27694 31442 27746
rect 31442 27694 31444 27746
rect 31388 27692 31444 27694
rect 30044 27020 30100 27076
rect 30156 27468 30212 27524
rect 30492 27580 30548 27636
rect 31164 27634 31220 27636
rect 31164 27582 31166 27634
rect 31166 27582 31218 27634
rect 31218 27582 31220 27634
rect 31164 27580 31220 27582
rect 32396 27916 32452 27972
rect 33852 27970 33908 27972
rect 33852 27918 33854 27970
rect 33854 27918 33906 27970
rect 33906 27918 33908 27970
rect 33852 27916 33908 27918
rect 32172 27692 32228 27748
rect 31388 27468 31444 27524
rect 33068 27858 33124 27860
rect 33068 27806 33070 27858
rect 33070 27806 33122 27858
rect 33122 27806 33124 27858
rect 33068 27804 33124 27806
rect 32508 27580 32564 27636
rect 33180 27580 33236 27636
rect 31612 27074 31668 27076
rect 31612 27022 31614 27074
rect 31614 27022 31666 27074
rect 31666 27022 31668 27074
rect 31612 27020 31668 27022
rect 32844 27020 32900 27076
rect 32508 26348 32564 26404
rect 32172 26290 32228 26292
rect 32172 26238 32174 26290
rect 32174 26238 32226 26290
rect 32226 26238 32228 26290
rect 32172 26236 32228 26238
rect 31500 25452 31556 25508
rect 29932 24892 29988 24948
rect 30940 24892 30996 24948
rect 28588 23884 28644 23940
rect 25788 23826 25844 23828
rect 25788 23774 25790 23826
rect 25790 23774 25842 23826
rect 25842 23774 25844 23826
rect 25788 23772 25844 23774
rect 29708 23938 29764 23940
rect 29708 23886 29710 23938
rect 29710 23886 29762 23938
rect 29762 23886 29764 23938
rect 29708 23884 29764 23886
rect 29148 23826 29204 23828
rect 29148 23774 29150 23826
rect 29150 23774 29202 23826
rect 29202 23774 29204 23826
rect 29148 23772 29204 23774
rect 25004 21868 25060 21924
rect 23996 20412 24052 20468
rect 24556 20300 24612 20356
rect 24108 20018 24164 20020
rect 24108 19966 24110 20018
rect 24110 19966 24162 20018
rect 24162 19966 24164 20018
rect 24108 19964 24164 19966
rect 24332 19906 24388 19908
rect 24332 19854 24334 19906
rect 24334 19854 24386 19906
rect 24386 19854 24388 19906
rect 24332 19852 24388 19854
rect 24108 18450 24164 18452
rect 24108 18398 24110 18450
rect 24110 18398 24162 18450
rect 24162 18398 24164 18450
rect 24108 18396 24164 18398
rect 23436 17500 23492 17556
rect 23884 18172 23940 18228
rect 23772 18060 23828 18116
rect 23996 17724 24052 17780
rect 24668 18172 24724 18228
rect 25452 22428 25508 22484
rect 25116 20076 25172 20132
rect 24892 19404 24948 19460
rect 25228 20018 25284 20020
rect 25228 19966 25230 20018
rect 25230 19966 25282 20018
rect 25282 19966 25284 20018
rect 25228 19964 25284 19966
rect 25228 18396 25284 18452
rect 25452 20076 25508 20132
rect 25676 19964 25732 20020
rect 26908 19964 26964 20020
rect 25676 19458 25732 19460
rect 25676 19406 25678 19458
rect 25678 19406 25730 19458
rect 25730 19406 25732 19458
rect 25676 19404 25732 19406
rect 25452 19292 25508 19348
rect 25900 19234 25956 19236
rect 25900 19182 25902 19234
rect 25902 19182 25954 19234
rect 25954 19182 25956 19234
rect 25900 19180 25956 19182
rect 26908 19180 26964 19236
rect 27132 19852 27188 19908
rect 25340 18620 25396 18676
rect 27132 18674 27188 18676
rect 27132 18622 27134 18674
rect 27134 18622 27186 18674
rect 27186 18622 27188 18674
rect 27132 18620 27188 18622
rect 25228 18226 25284 18228
rect 25228 18174 25230 18226
rect 25230 18174 25282 18226
rect 25282 18174 25284 18226
rect 25228 18172 25284 18174
rect 26124 18172 26180 18228
rect 24780 18060 24836 18116
rect 24332 17948 24388 18004
rect 25676 17948 25732 18004
rect 23884 17666 23940 17668
rect 23884 17614 23886 17666
rect 23886 17614 23938 17666
rect 23938 17614 23940 17666
rect 23884 17612 23940 17614
rect 23548 16268 23604 16324
rect 23324 14252 23380 14308
rect 22764 12236 22820 12292
rect 23660 15372 23716 15428
rect 23884 17388 23940 17444
rect 23996 16828 24052 16884
rect 25340 17666 25396 17668
rect 25340 17614 25342 17666
rect 25342 17614 25394 17666
rect 25394 17614 25396 17666
rect 25340 17612 25396 17614
rect 25340 16828 25396 16884
rect 25228 16210 25284 16212
rect 25228 16158 25230 16210
rect 25230 16158 25282 16210
rect 25282 16158 25284 16210
rect 25228 16156 25284 16158
rect 28252 20076 28308 20132
rect 28140 18620 28196 18676
rect 27804 18508 27860 18564
rect 26572 17612 26628 17668
rect 25676 16716 25732 16772
rect 24220 15260 24276 15316
rect 23772 14476 23828 14532
rect 25228 15426 25284 15428
rect 25228 15374 25230 15426
rect 25230 15374 25282 15426
rect 25282 15374 25284 15426
rect 25228 15372 25284 15374
rect 23884 14252 23940 14308
rect 24220 14306 24276 14308
rect 24220 14254 24222 14306
rect 24222 14254 24274 14306
rect 24274 14254 24276 14306
rect 24220 14252 24276 14254
rect 23548 13356 23604 13412
rect 23436 13244 23492 13300
rect 23996 12908 24052 12964
rect 22876 12348 22932 12404
rect 23436 12684 23492 12740
rect 22652 11170 22708 11172
rect 22652 11118 22654 11170
rect 22654 11118 22706 11170
rect 22706 11118 22708 11170
rect 22652 11116 22708 11118
rect 22652 10556 22708 10612
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 18172 8370 18228 8372
rect 18172 8318 18174 8370
rect 18174 8318 18226 8370
rect 18226 8318 18228 8370
rect 18172 8316 18228 8318
rect 19516 8764 19572 8820
rect 20188 8764 20244 8820
rect 19516 7980 19572 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 21980 9826 22036 9828
rect 21980 9774 21982 9826
rect 21982 9774 22034 9826
rect 22034 9774 22036 9826
rect 21980 9772 22036 9774
rect 22428 8764 22484 8820
rect 22876 11282 22932 11284
rect 22876 11230 22878 11282
rect 22878 11230 22930 11282
rect 22930 11230 22932 11282
rect 22876 11228 22932 11230
rect 21644 8316 21700 8372
rect 22316 8370 22372 8372
rect 22316 8318 22318 8370
rect 22318 8318 22370 8370
rect 22370 8318 22372 8370
rect 22316 8316 22372 8318
rect 20636 7474 20692 7476
rect 20636 7422 20638 7474
rect 20638 7422 20690 7474
rect 20690 7422 20692 7474
rect 20636 7420 20692 7422
rect 21532 7420 21588 7476
rect 19404 6914 19460 6916
rect 19404 6862 19406 6914
rect 19406 6862 19458 6914
rect 19458 6862 19460 6914
rect 19404 6860 19460 6862
rect 18956 6076 19012 6132
rect 20636 6524 20692 6580
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20412 6300 20468 6356
rect 20044 6244 20100 6246
rect 20188 6076 20244 6132
rect 20076 5964 20132 6020
rect 18508 5292 18564 5348
rect 19404 5292 19460 5348
rect 19180 5122 19236 5124
rect 19180 5070 19182 5122
rect 19182 5070 19234 5122
rect 19234 5070 19236 5122
rect 19180 5068 19236 5070
rect 18396 4508 18452 4564
rect 20300 5852 20356 5908
rect 20748 6130 20804 6132
rect 20748 6078 20750 6130
rect 20750 6078 20802 6130
rect 20802 6078 20804 6130
rect 20748 6076 20804 6078
rect 20636 5404 20692 5460
rect 20524 5180 20580 5236
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20412 5010 20468 5012
rect 20412 4958 20414 5010
rect 20414 4958 20466 5010
rect 20466 4958 20468 5010
rect 20412 4956 20468 4958
rect 19628 4562 19684 4564
rect 19628 4510 19630 4562
rect 19630 4510 19682 4562
rect 19682 4510 19684 4562
rect 19628 4508 19684 4510
rect 19852 4450 19908 4452
rect 19852 4398 19854 4450
rect 19854 4398 19906 4450
rect 19906 4398 19908 4450
rect 19852 4396 19908 4398
rect 18172 3948 18228 4004
rect 20860 5852 20916 5908
rect 20748 5292 20804 5348
rect 20636 4450 20692 4452
rect 20636 4398 20638 4450
rect 20638 4398 20690 4450
rect 20690 4398 20692 4450
rect 20636 4396 20692 4398
rect 18844 3948 18900 4004
rect 19516 3948 19572 4004
rect 18620 3500 18676 3556
rect 18844 3612 18900 3668
rect 15484 3388 15540 3444
rect 18508 3442 18564 3444
rect 18508 3390 18510 3442
rect 18510 3390 18562 3442
rect 18562 3390 18564 3442
rect 18508 3388 18564 3390
rect 19852 3554 19908 3556
rect 19852 3502 19854 3554
rect 19854 3502 19906 3554
rect 19906 3502 19908 3554
rect 19852 3500 19908 3502
rect 22876 7420 22932 7476
rect 24780 14812 24836 14868
rect 24556 13356 24612 13412
rect 24108 12684 24164 12740
rect 24220 12572 24276 12628
rect 24556 12402 24612 12404
rect 24556 12350 24558 12402
rect 24558 12350 24610 12402
rect 24610 12350 24612 12402
rect 24556 12348 24612 12350
rect 23884 12290 23940 12292
rect 23884 12238 23886 12290
rect 23886 12238 23938 12290
rect 23938 12238 23940 12290
rect 23884 12236 23940 12238
rect 24668 12290 24724 12292
rect 24668 12238 24670 12290
rect 24670 12238 24722 12290
rect 24722 12238 24724 12290
rect 24668 12236 24724 12238
rect 23212 12012 23268 12068
rect 23324 11228 23380 11284
rect 23436 11340 23492 11396
rect 24332 11282 24388 11284
rect 24332 11230 24334 11282
rect 24334 11230 24386 11282
rect 24386 11230 24388 11282
rect 24332 11228 24388 11230
rect 23212 10556 23268 10612
rect 23660 9660 23716 9716
rect 23548 8764 23604 8820
rect 24444 9548 24500 9604
rect 24108 9154 24164 9156
rect 24108 9102 24110 9154
rect 24110 9102 24162 9154
rect 24162 9102 24164 9154
rect 24108 9100 24164 9102
rect 24220 7420 24276 7476
rect 24220 7196 24276 7252
rect 22988 6636 23044 6692
rect 24332 6748 24388 6804
rect 22988 6076 23044 6132
rect 21644 5964 21700 6020
rect 24108 5906 24164 5908
rect 24108 5854 24110 5906
rect 24110 5854 24162 5906
rect 24162 5854 24164 5906
rect 24108 5852 24164 5854
rect 21532 5068 21588 5124
rect 20972 4956 21028 5012
rect 20860 4396 20916 4452
rect 20860 4226 20916 4228
rect 20860 4174 20862 4226
rect 20862 4174 20914 4226
rect 20914 4174 20916 4226
rect 20860 4172 20916 4174
rect 21756 5404 21812 5460
rect 22316 5234 22372 5236
rect 22316 5182 22318 5234
rect 22318 5182 22370 5234
rect 22370 5182 22372 5234
rect 22316 5180 22372 5182
rect 24668 8764 24724 8820
rect 24668 7474 24724 7476
rect 24668 7422 24670 7474
rect 24670 7422 24722 7474
rect 24722 7422 24724 7474
rect 24668 7420 24724 7422
rect 25116 14252 25172 14308
rect 25788 15148 25844 15204
rect 25564 15036 25620 15092
rect 25900 14754 25956 14756
rect 25900 14702 25902 14754
rect 25902 14702 25954 14754
rect 25954 14702 25956 14754
rect 25900 14700 25956 14702
rect 25564 14418 25620 14420
rect 25564 14366 25566 14418
rect 25566 14366 25618 14418
rect 25618 14366 25620 14418
rect 25564 14364 25620 14366
rect 25564 12908 25620 12964
rect 25228 12684 25284 12740
rect 25452 12402 25508 12404
rect 25452 12350 25454 12402
rect 25454 12350 25506 12402
rect 25506 12350 25508 12402
rect 25452 12348 25508 12350
rect 25676 12236 25732 12292
rect 25564 12066 25620 12068
rect 25564 12014 25566 12066
rect 25566 12014 25618 12066
rect 25618 12014 25620 12066
rect 25564 12012 25620 12014
rect 26460 15314 26516 15316
rect 26460 15262 26462 15314
rect 26462 15262 26514 15314
rect 26514 15262 26516 15314
rect 26460 15260 26516 15262
rect 26348 14924 26404 14980
rect 26124 14812 26180 14868
rect 26236 14530 26292 14532
rect 26236 14478 26238 14530
rect 26238 14478 26290 14530
rect 26290 14478 26292 14530
rect 26236 14476 26292 14478
rect 29260 20076 29316 20132
rect 29036 19852 29092 19908
rect 28812 19794 28868 19796
rect 28812 19742 28814 19794
rect 28814 19742 28866 19794
rect 28866 19742 28868 19794
rect 28812 19740 28868 19742
rect 29372 19964 29428 20020
rect 31052 24780 31108 24836
rect 32620 26236 32676 26292
rect 32620 25730 32676 25732
rect 32620 25678 32622 25730
rect 32622 25678 32674 25730
rect 32674 25678 32676 25730
rect 32620 25676 32676 25678
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 33852 27020 33908 27076
rect 33628 26402 33684 26404
rect 33628 26350 33630 26402
rect 33630 26350 33682 26402
rect 33682 26350 33684 26402
rect 33628 26348 33684 26350
rect 33516 26290 33572 26292
rect 33516 26238 33518 26290
rect 33518 26238 33570 26290
rect 33570 26238 33572 26290
rect 33516 26236 33572 26238
rect 35868 27074 35924 27076
rect 35868 27022 35870 27074
rect 35870 27022 35922 27074
rect 35922 27022 35924 27074
rect 35868 27020 35924 27022
rect 35980 26796 36036 26852
rect 35420 26514 35476 26516
rect 35420 26462 35422 26514
rect 35422 26462 35474 26514
rect 35474 26462 35476 26514
rect 35420 26460 35476 26462
rect 31276 24498 31332 24500
rect 31276 24446 31278 24498
rect 31278 24446 31330 24498
rect 31330 24446 31332 24498
rect 31276 24444 31332 24446
rect 30268 23100 30324 23156
rect 29932 20802 29988 20804
rect 29932 20750 29934 20802
rect 29934 20750 29986 20802
rect 29986 20750 29988 20802
rect 29932 20748 29988 20750
rect 29596 19628 29652 19684
rect 30044 20018 30100 20020
rect 30044 19966 30046 20018
rect 30046 19966 30098 20018
rect 30098 19966 30100 20018
rect 30044 19964 30100 19966
rect 30492 22428 30548 22484
rect 31388 23154 31444 23156
rect 31388 23102 31390 23154
rect 31390 23102 31442 23154
rect 31442 23102 31444 23154
rect 31388 23100 31444 23102
rect 31836 24498 31892 24500
rect 31836 24446 31838 24498
rect 31838 24446 31890 24498
rect 31890 24446 31892 24498
rect 31836 24444 31892 24446
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 33740 24780 33796 24836
rect 34636 24780 34692 24836
rect 31612 22764 31668 22820
rect 30604 21644 30660 21700
rect 31388 22482 31444 22484
rect 31388 22430 31390 22482
rect 31390 22430 31442 22482
rect 31442 22430 31444 22482
rect 31388 22428 31444 22430
rect 31164 21474 31220 21476
rect 31164 21422 31166 21474
rect 31166 21422 31218 21474
rect 31218 21422 31220 21474
rect 31164 21420 31220 21422
rect 30380 20802 30436 20804
rect 30380 20750 30382 20802
rect 30382 20750 30434 20802
rect 30434 20750 30436 20802
rect 30380 20748 30436 20750
rect 30268 19740 30324 19796
rect 29708 19516 29764 19572
rect 29484 19404 29540 19460
rect 27916 17948 27972 18004
rect 27020 16156 27076 16212
rect 27692 16604 27748 16660
rect 27692 15874 27748 15876
rect 27692 15822 27694 15874
rect 27694 15822 27746 15874
rect 27746 15822 27748 15874
rect 27692 15820 27748 15822
rect 27020 15036 27076 15092
rect 26796 14700 26852 14756
rect 26236 13580 26292 13636
rect 26348 13020 26404 13076
rect 26236 12962 26292 12964
rect 26236 12910 26238 12962
rect 26238 12910 26290 12962
rect 26290 12910 26292 12962
rect 26236 12908 26292 12910
rect 26572 13468 26628 13524
rect 26460 12348 26516 12404
rect 25228 10556 25284 10612
rect 25228 9826 25284 9828
rect 25228 9774 25230 9826
rect 25230 9774 25282 9826
rect 25282 9774 25284 9826
rect 25228 9772 25284 9774
rect 25788 9884 25844 9940
rect 25788 9100 25844 9156
rect 26124 10108 26180 10164
rect 26124 7474 26180 7476
rect 26124 7422 26126 7474
rect 26126 7422 26178 7474
rect 26178 7422 26180 7474
rect 26124 7420 26180 7422
rect 26460 10556 26516 10612
rect 26684 12796 26740 12852
rect 26684 12348 26740 12404
rect 27020 13804 27076 13860
rect 27132 14476 27188 14532
rect 27692 14812 27748 14868
rect 27692 14530 27748 14532
rect 27692 14478 27694 14530
rect 27694 14478 27746 14530
rect 27746 14478 27748 14530
rect 27692 14476 27748 14478
rect 27580 14306 27636 14308
rect 27580 14254 27582 14306
rect 27582 14254 27634 14306
rect 27634 14254 27636 14306
rect 27580 14252 27636 14254
rect 26796 11340 26852 11396
rect 26796 10780 26852 10836
rect 26908 10610 26964 10612
rect 26908 10558 26910 10610
rect 26910 10558 26962 10610
rect 26962 10558 26964 10610
rect 26908 10556 26964 10558
rect 26572 10108 26628 10164
rect 26908 10332 26964 10388
rect 26796 9602 26852 9604
rect 26796 9550 26798 9602
rect 26798 9550 26850 9602
rect 26850 9550 26852 9602
rect 26796 9548 26852 9550
rect 27020 9772 27076 9828
rect 27468 13858 27524 13860
rect 27468 13806 27470 13858
rect 27470 13806 27522 13858
rect 27522 13806 27524 13858
rect 27468 13804 27524 13806
rect 27356 13746 27412 13748
rect 27356 13694 27358 13746
rect 27358 13694 27410 13746
rect 27410 13694 27412 13746
rect 27356 13692 27412 13694
rect 27244 13020 27300 13076
rect 27468 13580 27524 13636
rect 27244 12738 27300 12740
rect 27244 12686 27246 12738
rect 27246 12686 27298 12738
rect 27298 12686 27300 12738
rect 27244 12684 27300 12686
rect 27244 12178 27300 12180
rect 27244 12126 27246 12178
rect 27246 12126 27298 12178
rect 27298 12126 27300 12178
rect 27244 12124 27300 12126
rect 28028 17500 28084 17556
rect 28140 16770 28196 16772
rect 28140 16718 28142 16770
rect 28142 16718 28194 16770
rect 28194 16718 28196 16770
rect 28140 16716 28196 16718
rect 28252 16604 28308 16660
rect 27916 14924 27972 14980
rect 28252 14812 28308 14868
rect 28140 14028 28196 14084
rect 28028 13244 28084 13300
rect 28252 13692 28308 13748
rect 29260 18508 29316 18564
rect 28812 17724 28868 17780
rect 28700 17164 28756 17220
rect 28588 15986 28644 15988
rect 28588 15934 28590 15986
rect 28590 15934 28642 15986
rect 28642 15934 28644 15986
rect 28588 15932 28644 15934
rect 28924 15260 28980 15316
rect 29708 18450 29764 18452
rect 29708 18398 29710 18450
rect 29710 18398 29762 18450
rect 29762 18398 29764 18450
rect 29708 18396 29764 18398
rect 29596 18284 29652 18340
rect 29372 17666 29428 17668
rect 29372 17614 29374 17666
rect 29374 17614 29426 17666
rect 29426 17614 29428 17666
rect 29372 17612 29428 17614
rect 30380 19404 30436 19460
rect 30492 19964 30548 20020
rect 30492 19292 30548 19348
rect 29932 17948 29988 18004
rect 29596 16994 29652 16996
rect 29596 16942 29598 16994
rect 29598 16942 29650 16994
rect 29650 16942 29652 16994
rect 29596 16940 29652 16942
rect 29708 16716 29764 16772
rect 29820 16380 29876 16436
rect 29484 15932 29540 15988
rect 29484 15596 29540 15652
rect 31164 20802 31220 20804
rect 31164 20750 31166 20802
rect 31166 20750 31218 20802
rect 31218 20750 31220 20802
rect 31164 20748 31220 20750
rect 30716 20188 30772 20244
rect 30716 19628 30772 19684
rect 30716 18508 30772 18564
rect 30268 17948 30324 18004
rect 30268 17724 30324 17780
rect 30156 17612 30212 17668
rect 30716 17666 30772 17668
rect 30716 17614 30718 17666
rect 30718 17614 30770 17666
rect 30770 17614 30772 17666
rect 30716 17612 30772 17614
rect 33516 23938 33572 23940
rect 33516 23886 33518 23938
rect 33518 23886 33570 23938
rect 33570 23886 33572 23938
rect 33516 23884 33572 23886
rect 33068 22930 33124 22932
rect 33068 22878 33070 22930
rect 33070 22878 33122 22930
rect 33122 22878 33124 22930
rect 33068 22876 33124 22878
rect 33516 23436 33572 23492
rect 33404 22428 33460 22484
rect 33180 22258 33236 22260
rect 33180 22206 33182 22258
rect 33182 22206 33234 22258
rect 33234 22206 33236 22258
rect 33180 22204 33236 22206
rect 34188 23436 34244 23492
rect 33852 22540 33908 22596
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34972 23154 35028 23156
rect 34972 23102 34974 23154
rect 34974 23102 35026 23154
rect 35026 23102 35028 23154
rect 34972 23100 35028 23102
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34412 22482 34468 22484
rect 34412 22430 34414 22482
rect 34414 22430 34466 22482
rect 34466 22430 34468 22482
rect 34412 22428 34468 22430
rect 33628 22204 33684 22260
rect 34188 22092 34244 22148
rect 31948 21756 32004 21812
rect 33964 21756 34020 21812
rect 31836 21644 31892 21700
rect 32060 21586 32116 21588
rect 32060 21534 32062 21586
rect 32062 21534 32114 21586
rect 32114 21534 32116 21586
rect 32060 21532 32116 21534
rect 31836 21474 31892 21476
rect 31836 21422 31838 21474
rect 31838 21422 31890 21474
rect 31890 21422 31892 21474
rect 31836 21420 31892 21422
rect 31612 20636 31668 20692
rect 31164 20018 31220 20020
rect 31164 19966 31166 20018
rect 31166 19966 31218 20018
rect 31218 19966 31220 20018
rect 31164 19964 31220 19966
rect 31724 19852 31780 19908
rect 31052 19794 31108 19796
rect 31052 19742 31054 19794
rect 31054 19742 31106 19794
rect 31106 19742 31108 19794
rect 31052 19740 31108 19742
rect 31948 19740 32004 19796
rect 31388 19516 31444 19572
rect 31164 19234 31220 19236
rect 31164 19182 31166 19234
rect 31166 19182 31218 19234
rect 31218 19182 31220 19234
rect 31164 19180 31220 19182
rect 31164 18396 31220 18452
rect 30940 17500 30996 17556
rect 30492 17164 30548 17220
rect 30492 16940 30548 16996
rect 30044 15874 30100 15876
rect 30044 15822 30046 15874
rect 30046 15822 30098 15874
rect 30098 15822 30100 15874
rect 30044 15820 30100 15822
rect 28924 13746 28980 13748
rect 28924 13694 28926 13746
rect 28926 13694 28978 13746
rect 28978 13694 28980 13746
rect 28924 13692 28980 13694
rect 28364 12962 28420 12964
rect 28364 12910 28366 12962
rect 28366 12910 28418 12962
rect 28418 12910 28420 12962
rect 28364 12908 28420 12910
rect 27692 11788 27748 11844
rect 27580 11228 27636 11284
rect 27356 10332 27412 10388
rect 27356 9938 27412 9940
rect 27356 9886 27358 9938
rect 27358 9886 27410 9938
rect 27410 9886 27412 9938
rect 27356 9884 27412 9886
rect 27580 9884 27636 9940
rect 27244 9660 27300 9716
rect 27468 9436 27524 9492
rect 27580 9042 27636 9044
rect 27580 8990 27582 9042
rect 27582 8990 27634 9042
rect 27634 8990 27636 9042
rect 27580 8988 27636 8990
rect 27580 8540 27636 8596
rect 28028 12124 28084 12180
rect 28252 12124 28308 12180
rect 29148 12684 29204 12740
rect 29596 13132 29652 13188
rect 29932 13692 29988 13748
rect 29708 13020 29764 13076
rect 29372 12572 29428 12628
rect 29036 12290 29092 12292
rect 29036 12238 29038 12290
rect 29038 12238 29090 12290
rect 29090 12238 29092 12290
rect 29036 12236 29092 12238
rect 29596 12124 29652 12180
rect 28476 11788 28532 11844
rect 29484 11900 29540 11956
rect 27804 11340 27860 11396
rect 29932 12178 29988 12180
rect 29932 12126 29934 12178
rect 29934 12126 29986 12178
rect 29986 12126 29988 12178
rect 29932 12124 29988 12126
rect 29820 11900 29876 11956
rect 31500 18508 31556 18564
rect 35308 22540 35364 22596
rect 35084 22482 35140 22484
rect 35084 22430 35086 22482
rect 35086 22430 35138 22482
rect 35138 22430 35140 22482
rect 35084 22428 35140 22430
rect 34748 22370 34804 22372
rect 34748 22318 34750 22370
rect 34750 22318 34802 22370
rect 34802 22318 34804 22370
rect 34748 22316 34804 22318
rect 35644 22316 35700 22372
rect 35196 22146 35252 22148
rect 35196 22094 35198 22146
rect 35198 22094 35250 22146
rect 35250 22094 35252 22146
rect 35196 22092 35252 22094
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 34076 19516 34132 19572
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 33964 19180 34020 19236
rect 32060 18396 32116 18452
rect 33516 18396 33572 18452
rect 32508 18338 32564 18340
rect 32508 18286 32510 18338
rect 32510 18286 32562 18338
rect 32562 18286 32564 18338
rect 32508 18284 32564 18286
rect 33852 18284 33908 18340
rect 33516 17164 33572 17220
rect 32956 16940 33012 16996
rect 31724 16882 31780 16884
rect 31724 16830 31726 16882
rect 31726 16830 31778 16882
rect 31778 16830 31780 16882
rect 31724 16828 31780 16830
rect 31500 15372 31556 15428
rect 31276 14530 31332 14532
rect 31276 14478 31278 14530
rect 31278 14478 31330 14530
rect 31330 14478 31332 14530
rect 31276 14476 31332 14478
rect 34076 18396 34132 18452
rect 34188 17948 34244 18004
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 36540 30882 36596 30884
rect 36540 30830 36542 30882
rect 36542 30830 36594 30882
rect 36594 30830 36596 30882
rect 36540 30828 36596 30830
rect 39900 38834 39956 38836
rect 39900 38782 39902 38834
rect 39902 38782 39954 38834
rect 39954 38782 39956 38834
rect 39900 38780 39956 38782
rect 39676 38108 39732 38164
rect 40348 38722 40404 38724
rect 40348 38670 40350 38722
rect 40350 38670 40402 38722
rect 40402 38670 40404 38722
rect 40348 38668 40404 38670
rect 39788 37772 39844 37828
rect 38892 37212 38948 37268
rect 37772 35196 37828 35252
rect 38108 36876 38164 36932
rect 38332 36370 38388 36372
rect 38332 36318 38334 36370
rect 38334 36318 38386 36370
rect 38386 36318 38388 36370
rect 38332 36316 38388 36318
rect 39228 36370 39284 36372
rect 39228 36318 39230 36370
rect 39230 36318 39282 36370
rect 39282 36318 39284 36370
rect 39228 36316 39284 36318
rect 38668 35980 38724 36036
rect 37772 34636 37828 34692
rect 38220 34636 38276 34692
rect 37772 33628 37828 33684
rect 37996 33292 38052 33348
rect 39564 36258 39620 36260
rect 39564 36206 39566 36258
rect 39566 36206 39618 36258
rect 39618 36206 39620 36258
rect 39564 36204 39620 36206
rect 40572 40124 40628 40180
rect 40572 39004 40628 39060
rect 40684 40012 40740 40068
rect 41020 41970 41076 41972
rect 41020 41918 41022 41970
rect 41022 41918 41074 41970
rect 41074 41918 41076 41970
rect 41020 41916 41076 41918
rect 41132 41020 41188 41076
rect 40908 40124 40964 40180
rect 41356 41970 41412 41972
rect 41356 41918 41358 41970
rect 41358 41918 41410 41970
rect 41410 41918 41412 41970
rect 41356 41916 41412 41918
rect 42364 43426 42420 43428
rect 42364 43374 42366 43426
rect 42366 43374 42418 43426
rect 42418 43374 42420 43426
rect 42364 43372 42420 43374
rect 41916 42866 41972 42868
rect 41916 42814 41918 42866
rect 41918 42814 41970 42866
rect 41970 42814 41972 42866
rect 41916 42812 41972 42814
rect 41804 42082 41860 42084
rect 41804 42030 41806 42082
rect 41806 42030 41858 42082
rect 41858 42030 41860 42082
rect 41804 42028 41860 42030
rect 41916 41970 41972 41972
rect 41916 41918 41918 41970
rect 41918 41918 41970 41970
rect 41970 41918 41972 41970
rect 41916 41916 41972 41918
rect 41244 40572 41300 40628
rect 41692 40796 41748 40852
rect 41468 40514 41524 40516
rect 41468 40462 41470 40514
rect 41470 40462 41522 40514
rect 41522 40462 41524 40514
rect 41468 40460 41524 40462
rect 41244 40402 41300 40404
rect 41244 40350 41246 40402
rect 41246 40350 41298 40402
rect 41298 40350 41300 40402
rect 41244 40348 41300 40350
rect 40908 39228 40964 39284
rect 40908 39058 40964 39060
rect 40908 39006 40910 39058
rect 40910 39006 40962 39058
rect 40962 39006 40964 39058
rect 40908 39004 40964 39006
rect 43820 43708 43876 43764
rect 42476 42754 42532 42756
rect 42476 42702 42478 42754
rect 42478 42702 42530 42754
rect 42530 42702 42532 42754
rect 42476 42700 42532 42702
rect 42252 42642 42308 42644
rect 42252 42590 42254 42642
rect 42254 42590 42306 42642
rect 42306 42590 42308 42642
rect 42252 42588 42308 42590
rect 42364 41692 42420 41748
rect 42140 40572 42196 40628
rect 41804 40012 41860 40068
rect 42140 40290 42196 40292
rect 42140 40238 42142 40290
rect 42142 40238 42194 40290
rect 42194 40238 42196 40290
rect 42140 40236 42196 40238
rect 41132 38946 41188 38948
rect 41132 38894 41134 38946
rect 41134 38894 41186 38946
rect 41186 38894 41188 38946
rect 41132 38892 41188 38894
rect 41020 38834 41076 38836
rect 41020 38782 41022 38834
rect 41022 38782 41074 38834
rect 41074 38782 41076 38834
rect 41020 38780 41076 38782
rect 41356 38668 41412 38724
rect 40908 38108 40964 38164
rect 40572 37324 40628 37380
rect 40684 36988 40740 37044
rect 40124 35980 40180 36036
rect 41356 37938 41412 37940
rect 41356 37886 41358 37938
rect 41358 37886 41410 37938
rect 41410 37886 41412 37938
rect 41356 37884 41412 37886
rect 41916 39058 41972 39060
rect 41916 39006 41918 39058
rect 41918 39006 41970 39058
rect 41970 39006 41972 39058
rect 41916 39004 41972 39006
rect 42476 40236 42532 40292
rect 42476 39340 42532 39396
rect 42476 39116 42532 39172
rect 41692 38050 41748 38052
rect 41692 37998 41694 38050
rect 41694 37998 41746 38050
rect 41746 37998 41748 38050
rect 41692 37996 41748 37998
rect 41020 37266 41076 37268
rect 41020 37214 41022 37266
rect 41022 37214 41074 37266
rect 41074 37214 41076 37266
rect 41020 37212 41076 37214
rect 41692 37324 41748 37380
rect 41804 36204 41860 36260
rect 40124 34972 40180 35028
rect 39116 34188 39172 34244
rect 39788 34188 39844 34244
rect 39228 33346 39284 33348
rect 39228 33294 39230 33346
rect 39230 33294 39282 33346
rect 39282 33294 39284 33346
rect 39228 33292 39284 33294
rect 38892 32956 38948 33012
rect 39116 33180 39172 33236
rect 38220 32786 38276 32788
rect 38220 32734 38222 32786
rect 38222 32734 38274 32786
rect 38274 32734 38276 32786
rect 38220 32732 38276 32734
rect 38892 32786 38948 32788
rect 38892 32734 38894 32786
rect 38894 32734 38946 32786
rect 38946 32734 38948 32786
rect 38892 32732 38948 32734
rect 38556 32674 38612 32676
rect 38556 32622 38558 32674
rect 38558 32622 38610 32674
rect 38610 32622 38612 32674
rect 38556 32620 38612 32622
rect 39228 32786 39284 32788
rect 39228 32734 39230 32786
rect 39230 32734 39282 32786
rect 39282 32734 39284 32786
rect 39228 32732 39284 32734
rect 39900 32956 39956 33012
rect 40908 32956 40964 33012
rect 40460 32620 40516 32676
rect 42476 38668 42532 38724
rect 42252 37100 42308 37156
rect 41916 35868 41972 35924
rect 41804 35196 41860 35252
rect 41468 35026 41524 35028
rect 41468 34974 41470 35026
rect 41470 34974 41522 35026
rect 41522 34974 41524 35026
rect 41468 34972 41524 34974
rect 42140 35698 42196 35700
rect 42140 35646 42142 35698
rect 42142 35646 42194 35698
rect 42194 35646 42196 35698
rect 42140 35644 42196 35646
rect 43708 42866 43764 42868
rect 43708 42814 43710 42866
rect 43710 42814 43762 42866
rect 43762 42814 43764 42866
rect 43708 42812 43764 42814
rect 43484 42754 43540 42756
rect 43484 42702 43486 42754
rect 43486 42702 43538 42754
rect 43538 42702 43540 42754
rect 43484 42700 43540 42702
rect 43148 42530 43204 42532
rect 43148 42478 43150 42530
rect 43150 42478 43202 42530
rect 43202 42478 43204 42530
rect 43148 42476 43204 42478
rect 42924 41804 42980 41860
rect 44604 46114 44660 46116
rect 44604 46062 44606 46114
rect 44606 46062 44658 46114
rect 44658 46062 44660 46114
rect 44604 46060 44660 46062
rect 44380 45164 44436 45220
rect 44156 45106 44212 45108
rect 44156 45054 44158 45106
rect 44158 45054 44210 45106
rect 44210 45054 44212 45106
rect 44156 45052 44212 45054
rect 45052 44828 45108 44884
rect 45164 49084 45220 49140
rect 45164 44716 45220 44772
rect 45276 47068 45332 47124
rect 44828 43484 44884 43540
rect 44716 43260 44772 43316
rect 44044 42924 44100 42980
rect 44828 42700 44884 42756
rect 43932 42252 43988 42308
rect 44044 42364 44100 42420
rect 43036 40572 43092 40628
rect 42812 39788 42868 39844
rect 43036 40236 43092 40292
rect 42812 38946 42868 38948
rect 42812 38894 42814 38946
rect 42814 38894 42866 38946
rect 42866 38894 42868 38946
rect 42812 38892 42868 38894
rect 42700 37884 42756 37940
rect 44940 41692 44996 41748
rect 44268 39116 44324 39172
rect 43596 38274 43652 38276
rect 43596 38222 43598 38274
rect 43598 38222 43650 38274
rect 43650 38222 43652 38274
rect 43596 38220 43652 38222
rect 43372 37996 43428 38052
rect 43820 37154 43876 37156
rect 43820 37102 43822 37154
rect 43822 37102 43874 37154
rect 43874 37102 43876 37154
rect 43820 37100 43876 37102
rect 44604 38892 44660 38948
rect 45052 41132 45108 41188
rect 45388 44994 45444 44996
rect 45388 44942 45390 44994
rect 45390 44942 45442 44994
rect 45442 44942 45444 44994
rect 45388 44940 45444 44942
rect 47180 46396 47236 46452
rect 45724 44604 45780 44660
rect 45836 44546 45892 44548
rect 45836 44494 45838 44546
rect 45838 44494 45890 44546
rect 45890 44494 45892 44546
rect 45836 44492 45892 44494
rect 45276 41356 45332 41412
rect 45164 39618 45220 39620
rect 45164 39566 45166 39618
rect 45166 39566 45218 39618
rect 45218 39566 45220 39618
rect 45164 39564 45220 39566
rect 45052 39004 45108 39060
rect 44940 38668 44996 38724
rect 45388 38668 45444 38724
rect 44828 38050 44884 38052
rect 44828 37998 44830 38050
rect 44830 37998 44882 38050
rect 44882 37998 44884 38050
rect 44828 37996 44884 37998
rect 43372 36258 43428 36260
rect 43372 36206 43374 36258
rect 43374 36206 43426 36258
rect 43426 36206 43428 36258
rect 43372 36204 43428 36206
rect 42812 36092 42868 36148
rect 43484 36092 43540 36148
rect 43596 36316 43652 36372
rect 42924 35922 42980 35924
rect 42924 35870 42926 35922
rect 42926 35870 42978 35922
rect 42978 35870 42980 35922
rect 42924 35868 42980 35870
rect 43260 35922 43316 35924
rect 43260 35870 43262 35922
rect 43262 35870 43314 35922
rect 43314 35870 43316 35922
rect 43260 35868 43316 35870
rect 43820 36428 43876 36484
rect 44044 35980 44100 36036
rect 42588 35698 42644 35700
rect 42588 35646 42590 35698
rect 42590 35646 42642 35698
rect 42642 35646 42644 35698
rect 42588 35644 42644 35646
rect 42364 35532 42420 35588
rect 42700 35026 42756 35028
rect 42700 34974 42702 35026
rect 42702 34974 42754 35026
rect 42754 34974 42756 35026
rect 42700 34972 42756 34974
rect 43148 34914 43204 34916
rect 43148 34862 43150 34914
rect 43150 34862 43202 34914
rect 43202 34862 43204 34914
rect 43148 34860 43204 34862
rect 43932 34914 43988 34916
rect 43932 34862 43934 34914
rect 43934 34862 43986 34914
rect 43986 34862 43988 34914
rect 43932 34860 43988 34862
rect 41580 33180 41636 33236
rect 42140 32956 42196 33012
rect 41804 32786 41860 32788
rect 41804 32734 41806 32786
rect 41806 32734 41858 32786
rect 41858 32734 41860 32786
rect 41804 32732 41860 32734
rect 40908 32508 40964 32564
rect 41356 32562 41412 32564
rect 41356 32510 41358 32562
rect 41358 32510 41410 32562
rect 41410 32510 41412 32562
rect 41356 32508 41412 32510
rect 41916 32562 41972 32564
rect 41916 32510 41918 32562
rect 41918 32510 41970 32562
rect 41970 32510 41972 32562
rect 41916 32508 41972 32510
rect 39900 31948 39956 32004
rect 41020 31948 41076 32004
rect 42364 32562 42420 32564
rect 42364 32510 42366 32562
rect 42366 32510 42418 32562
rect 42418 32510 42420 32562
rect 42364 32508 42420 32510
rect 43484 33346 43540 33348
rect 43484 33294 43486 33346
rect 43486 33294 43538 33346
rect 43538 33294 43540 33346
rect 43484 33292 43540 33294
rect 42924 32956 42980 33012
rect 43932 33516 43988 33572
rect 43596 32844 43652 32900
rect 43260 32732 43316 32788
rect 44268 35644 44324 35700
rect 44268 34802 44324 34804
rect 44268 34750 44270 34802
rect 44270 34750 44322 34802
rect 44322 34750 44324 34802
rect 44268 34748 44324 34750
rect 44156 33740 44212 33796
rect 44268 33292 44324 33348
rect 44268 32956 44324 33012
rect 43708 32508 43764 32564
rect 42924 32396 42980 32452
rect 44156 31890 44212 31892
rect 44156 31838 44158 31890
rect 44158 31838 44210 31890
rect 44210 31838 44212 31890
rect 44156 31836 44212 31838
rect 37996 30828 38052 30884
rect 37212 30716 37268 30772
rect 37772 30770 37828 30772
rect 37772 30718 37774 30770
rect 37774 30718 37826 30770
rect 37826 30718 37828 30770
rect 37772 30716 37828 30718
rect 43820 31778 43876 31780
rect 43820 31726 43822 31778
rect 43822 31726 43874 31778
rect 43874 31726 43876 31778
rect 43820 31724 43876 31726
rect 42588 31666 42644 31668
rect 42588 31614 42590 31666
rect 42590 31614 42642 31666
rect 42642 31614 42644 31666
rect 42588 31612 42644 31614
rect 44604 36988 44660 37044
rect 44716 36092 44772 36148
rect 44940 36428 44996 36484
rect 44940 36258 44996 36260
rect 44940 36206 44942 36258
rect 44942 36206 44994 36258
rect 44994 36206 44996 36258
rect 44940 36204 44996 36206
rect 44940 35698 44996 35700
rect 44940 35646 44942 35698
rect 44942 35646 44994 35698
rect 44994 35646 44996 35698
rect 44940 35644 44996 35646
rect 44716 35196 44772 35252
rect 44604 35084 44660 35140
rect 44716 34354 44772 34356
rect 44716 34302 44718 34354
rect 44718 34302 44770 34354
rect 44770 34302 44772 34354
rect 44716 34300 44772 34302
rect 45276 37378 45332 37380
rect 45276 37326 45278 37378
rect 45278 37326 45330 37378
rect 45330 37326 45332 37378
rect 45276 37324 45332 37326
rect 45276 36370 45332 36372
rect 45276 36318 45278 36370
rect 45278 36318 45330 36370
rect 45330 36318 45332 36370
rect 45276 36316 45332 36318
rect 45164 35756 45220 35812
rect 45612 41074 45668 41076
rect 45612 41022 45614 41074
rect 45614 41022 45666 41074
rect 45666 41022 45668 41074
rect 45612 41020 45668 41022
rect 45500 35868 45556 35924
rect 45276 35084 45332 35140
rect 45948 40572 46004 40628
rect 45948 40402 46004 40404
rect 45948 40350 45950 40402
rect 45950 40350 46002 40402
rect 46002 40350 46004 40402
rect 45948 40348 46004 40350
rect 45836 38834 45892 38836
rect 45836 38782 45838 38834
rect 45838 38782 45890 38834
rect 45890 38782 45892 38834
rect 45836 38780 45892 38782
rect 46844 43596 46900 43652
rect 47180 43596 47236 43652
rect 46508 38668 46564 38724
rect 45724 36316 45780 36372
rect 45612 35532 45668 35588
rect 45388 34972 45444 35028
rect 45836 34748 45892 34804
rect 45948 37100 46004 37156
rect 47404 40460 47460 40516
rect 47180 39116 47236 39172
rect 47292 40348 47348 40404
rect 47740 44210 47796 44212
rect 47740 44158 47742 44210
rect 47742 44158 47794 44210
rect 47794 44158 47796 44210
rect 47740 44156 47796 44158
rect 47852 43596 47908 43652
rect 47628 43372 47684 43428
rect 47068 38834 47124 38836
rect 47068 38782 47070 38834
rect 47070 38782 47122 38834
rect 47122 38782 47124 38834
rect 47068 38780 47124 38782
rect 46844 37324 46900 37380
rect 47516 38946 47572 38948
rect 47516 38894 47518 38946
rect 47518 38894 47570 38946
rect 47570 38894 47572 38946
rect 47516 38892 47572 38894
rect 47180 37100 47236 37156
rect 46620 36988 46676 37044
rect 47404 36316 47460 36372
rect 47292 35980 47348 36036
rect 46060 35810 46116 35812
rect 46060 35758 46062 35810
rect 46062 35758 46114 35810
rect 46114 35758 46116 35810
rect 46060 35756 46116 35758
rect 47180 35644 47236 35700
rect 44828 34076 44884 34132
rect 44940 33740 44996 33796
rect 45388 33516 45444 33572
rect 45500 33404 45556 33460
rect 44828 33346 44884 33348
rect 44828 33294 44830 33346
rect 44830 33294 44882 33346
rect 44882 33294 44884 33346
rect 44828 33292 44884 33294
rect 45388 33180 45444 33236
rect 45164 32508 45220 32564
rect 45164 31836 45220 31892
rect 44492 31164 44548 31220
rect 44716 31724 44772 31780
rect 45724 33404 45780 33460
rect 45052 31106 45108 31108
rect 45052 31054 45054 31106
rect 45054 31054 45106 31106
rect 45106 31054 45108 31106
rect 45052 31052 45108 31054
rect 36988 29820 37044 29876
rect 37436 29986 37492 29988
rect 37436 29934 37438 29986
rect 37438 29934 37490 29986
rect 37490 29934 37492 29986
rect 37436 29932 37492 29934
rect 37324 29708 37380 29764
rect 36764 29484 36820 29540
rect 37436 29484 37492 29540
rect 37436 28812 37492 28868
rect 39452 30098 39508 30100
rect 39452 30046 39454 30098
rect 39454 30046 39506 30098
rect 39506 30046 39508 30098
rect 39452 30044 39508 30046
rect 41132 30044 41188 30100
rect 37660 28700 37716 28756
rect 37100 28364 37156 28420
rect 38220 29426 38276 29428
rect 38220 29374 38222 29426
rect 38222 29374 38274 29426
rect 38274 29374 38276 29426
rect 38220 29372 38276 29374
rect 41356 29932 41412 29988
rect 38332 28924 38388 28980
rect 37996 28642 38052 28644
rect 37996 28590 37998 28642
rect 37998 28590 38050 28642
rect 38050 28590 38052 28642
rect 37996 28588 38052 28590
rect 37436 27970 37492 27972
rect 37436 27918 37438 27970
rect 37438 27918 37490 27970
rect 37490 27918 37492 27970
rect 37436 27916 37492 27918
rect 38892 28588 38948 28644
rect 36876 27804 36932 27860
rect 38444 27804 38500 27860
rect 36876 27580 36932 27636
rect 36428 26796 36484 26852
rect 36988 26348 37044 26404
rect 36428 25452 36484 25508
rect 38668 27634 38724 27636
rect 38668 27582 38670 27634
rect 38670 27582 38722 27634
rect 38722 27582 38724 27634
rect 38668 27580 38724 27582
rect 37324 25506 37380 25508
rect 37324 25454 37326 25506
rect 37326 25454 37378 25506
rect 37378 25454 37380 25506
rect 37324 25452 37380 25454
rect 38108 25506 38164 25508
rect 38108 25454 38110 25506
rect 38110 25454 38162 25506
rect 38162 25454 38164 25506
rect 38108 25452 38164 25454
rect 38220 25228 38276 25284
rect 38108 24946 38164 24948
rect 38108 24894 38110 24946
rect 38110 24894 38162 24946
rect 38162 24894 38164 24946
rect 38108 24892 38164 24894
rect 37772 24834 37828 24836
rect 37772 24782 37774 24834
rect 37774 24782 37826 24834
rect 37826 24782 37828 24834
rect 37772 24780 37828 24782
rect 37548 24668 37604 24724
rect 39116 26796 39172 26852
rect 39004 26290 39060 26292
rect 39004 26238 39006 26290
rect 39006 26238 39058 26290
rect 39058 26238 39060 26290
rect 39004 26236 39060 26238
rect 41580 29202 41636 29204
rect 41580 29150 41582 29202
rect 41582 29150 41634 29202
rect 41634 29150 41636 29202
rect 41580 29148 41636 29150
rect 42476 30098 42532 30100
rect 42476 30046 42478 30098
rect 42478 30046 42530 30098
rect 42530 30046 42532 30098
rect 42476 30044 42532 30046
rect 44044 30044 44100 30100
rect 42140 29932 42196 29988
rect 42252 29372 42308 29428
rect 40348 28028 40404 28084
rect 40012 27970 40068 27972
rect 40012 27918 40014 27970
rect 40014 27918 40066 27970
rect 40066 27918 40068 27970
rect 40012 27916 40068 27918
rect 41468 27858 41524 27860
rect 41468 27806 41470 27858
rect 41470 27806 41522 27858
rect 41522 27806 41524 27858
rect 41468 27804 41524 27806
rect 40908 27074 40964 27076
rect 40908 27022 40910 27074
rect 40910 27022 40962 27074
rect 40962 27022 40964 27074
rect 40908 27020 40964 27022
rect 39228 25506 39284 25508
rect 39228 25454 39230 25506
rect 39230 25454 39282 25506
rect 39282 25454 39284 25506
rect 39228 25452 39284 25454
rect 38556 25340 38612 25396
rect 38444 24668 38500 24724
rect 38668 25116 38724 25172
rect 38556 23548 38612 23604
rect 38332 23378 38388 23380
rect 38332 23326 38334 23378
rect 38334 23326 38386 23378
rect 38386 23326 38388 23378
rect 38332 23324 38388 23326
rect 38108 23100 38164 23156
rect 36204 19852 36260 19908
rect 36876 22540 36932 22596
rect 37772 22258 37828 22260
rect 37772 22206 37774 22258
rect 37774 22206 37826 22258
rect 37826 22206 37828 22258
rect 37772 22204 37828 22206
rect 38444 22258 38500 22260
rect 38444 22206 38446 22258
rect 38446 22206 38498 22258
rect 38498 22206 38500 22258
rect 38444 22204 38500 22206
rect 38780 24892 38836 24948
rect 38892 25340 38948 25396
rect 39340 24834 39396 24836
rect 39340 24782 39342 24834
rect 39342 24782 39394 24834
rect 39394 24782 39396 24834
rect 39340 24780 39396 24782
rect 38780 23212 38836 23268
rect 38892 22930 38948 22932
rect 38892 22878 38894 22930
rect 38894 22878 38946 22930
rect 38946 22878 38948 22930
rect 38892 22876 38948 22878
rect 38444 21532 38500 21588
rect 38220 21084 38276 21140
rect 36876 20860 36932 20916
rect 37660 20914 37716 20916
rect 37660 20862 37662 20914
rect 37662 20862 37714 20914
rect 37714 20862 37716 20914
rect 37660 20860 37716 20862
rect 37996 20860 38052 20916
rect 37100 20802 37156 20804
rect 37100 20750 37102 20802
rect 37102 20750 37154 20802
rect 37154 20750 37156 20802
rect 37100 20748 37156 20750
rect 36988 20690 37044 20692
rect 36988 20638 36990 20690
rect 36990 20638 37042 20690
rect 37042 20638 37044 20690
rect 36988 20636 37044 20638
rect 38108 20690 38164 20692
rect 38108 20638 38110 20690
rect 38110 20638 38162 20690
rect 38162 20638 38164 20690
rect 38108 20636 38164 20638
rect 37660 20412 37716 20468
rect 36876 19292 36932 19348
rect 35868 17948 35924 18004
rect 33292 15932 33348 15988
rect 34300 16828 34356 16884
rect 34636 16882 34692 16884
rect 34636 16830 34638 16882
rect 34638 16830 34690 16882
rect 34690 16830 34692 16882
rect 34636 16828 34692 16830
rect 33404 15538 33460 15540
rect 33404 15486 33406 15538
rect 33406 15486 33458 15538
rect 33458 15486 33460 15538
rect 33404 15484 33460 15486
rect 32172 15426 32228 15428
rect 32172 15374 32174 15426
rect 32174 15374 32226 15426
rect 32226 15374 32228 15426
rect 32172 15372 32228 15374
rect 32396 15314 32452 15316
rect 32396 15262 32398 15314
rect 32398 15262 32450 15314
rect 32450 15262 32452 15314
rect 32396 15260 32452 15262
rect 31052 13858 31108 13860
rect 31052 13806 31054 13858
rect 31054 13806 31106 13858
rect 31106 13806 31108 13858
rect 31052 13804 31108 13806
rect 31500 13746 31556 13748
rect 31500 13694 31502 13746
rect 31502 13694 31554 13746
rect 31554 13694 31556 13746
rect 31500 13692 31556 13694
rect 31388 13132 31444 13188
rect 31052 12908 31108 12964
rect 31612 13132 31668 13188
rect 31388 12402 31444 12404
rect 31388 12350 31390 12402
rect 31390 12350 31442 12402
rect 31442 12350 31444 12402
rect 31388 12348 31444 12350
rect 31276 12290 31332 12292
rect 31276 12238 31278 12290
rect 31278 12238 31330 12290
rect 31330 12238 31332 12290
rect 31276 12236 31332 12238
rect 30492 11900 30548 11956
rect 27804 10668 27860 10724
rect 26908 7532 26964 7588
rect 26124 7196 26180 7252
rect 27244 7420 27300 7476
rect 26236 6802 26292 6804
rect 26236 6750 26238 6802
rect 26238 6750 26290 6802
rect 26290 6750 26292 6802
rect 26236 6748 26292 6750
rect 26796 6690 26852 6692
rect 26796 6638 26798 6690
rect 26798 6638 26850 6690
rect 26850 6638 26852 6690
rect 26796 6636 26852 6638
rect 22316 4956 22372 5012
rect 22428 4898 22484 4900
rect 22428 4846 22430 4898
rect 22430 4846 22482 4898
rect 22482 4846 22484 4898
rect 22428 4844 22484 4846
rect 22092 4226 22148 4228
rect 22092 4174 22094 4226
rect 22094 4174 22146 4226
rect 22146 4174 22148 4226
rect 22092 4172 22148 4174
rect 21868 3666 21924 3668
rect 21868 3614 21870 3666
rect 21870 3614 21922 3666
rect 21922 3614 21924 3666
rect 21868 3612 21924 3614
rect 21532 3500 21588 3556
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 23660 4844 23716 4900
rect 24332 5180 24388 5236
rect 27916 10556 27972 10612
rect 29484 11228 29540 11284
rect 28924 10722 28980 10724
rect 28924 10670 28926 10722
rect 28926 10670 28978 10722
rect 28978 10670 28980 10722
rect 28924 10668 28980 10670
rect 28364 10610 28420 10612
rect 28364 10558 28366 10610
rect 28366 10558 28418 10610
rect 28418 10558 28420 10610
rect 28364 10556 28420 10558
rect 28252 9938 28308 9940
rect 28252 9886 28254 9938
rect 28254 9886 28306 9938
rect 28306 9886 28308 9938
rect 28252 9884 28308 9886
rect 28364 9714 28420 9716
rect 28364 9662 28366 9714
rect 28366 9662 28418 9714
rect 28418 9662 28420 9714
rect 28364 9660 28420 9662
rect 28252 9324 28308 9380
rect 27916 8988 27972 9044
rect 28700 10108 28756 10164
rect 29596 9826 29652 9828
rect 29596 9774 29598 9826
rect 29598 9774 29650 9826
rect 29650 9774 29652 9826
rect 29596 9772 29652 9774
rect 30044 11394 30100 11396
rect 30044 11342 30046 11394
rect 30046 11342 30098 11394
rect 30098 11342 30100 11394
rect 30044 11340 30100 11342
rect 31836 13916 31892 13972
rect 32060 13132 32116 13188
rect 31948 12850 32004 12852
rect 31948 12798 31950 12850
rect 31950 12798 32002 12850
rect 32002 12798 32004 12850
rect 31948 12796 32004 12798
rect 31724 11900 31780 11956
rect 31836 12236 31892 12292
rect 30716 11394 30772 11396
rect 30716 11342 30718 11394
rect 30718 11342 30770 11394
rect 30770 11342 30772 11394
rect 30716 11340 30772 11342
rect 31052 11394 31108 11396
rect 31052 11342 31054 11394
rect 31054 11342 31106 11394
rect 31106 11342 31108 11394
rect 31052 11340 31108 11342
rect 31724 11394 31780 11396
rect 31724 11342 31726 11394
rect 31726 11342 31778 11394
rect 31778 11342 31780 11394
rect 31724 11340 31780 11342
rect 31164 10668 31220 10724
rect 29932 10556 29988 10612
rect 30716 10108 30772 10164
rect 30940 9826 30996 9828
rect 30940 9774 30942 9826
rect 30942 9774 30994 9826
rect 30994 9774 30996 9826
rect 30940 9772 30996 9774
rect 28028 8428 28084 8484
rect 28476 7586 28532 7588
rect 28476 7534 28478 7586
rect 28478 7534 28530 7586
rect 28530 7534 28532 7586
rect 28476 7532 28532 7534
rect 27356 6690 27412 6692
rect 27356 6638 27358 6690
rect 27358 6638 27410 6690
rect 27410 6638 27412 6690
rect 27356 6636 27412 6638
rect 26348 6188 26404 6244
rect 24780 4844 24836 4900
rect 24668 3388 24724 3444
rect 25340 5682 25396 5684
rect 25340 5630 25342 5682
rect 25342 5630 25394 5682
rect 25394 5630 25396 5682
rect 25340 5628 25396 5630
rect 25452 5234 25508 5236
rect 25452 5182 25454 5234
rect 25454 5182 25506 5234
rect 25506 5182 25508 5234
rect 25452 5180 25508 5182
rect 25452 3500 25508 3556
rect 26572 5964 26628 6020
rect 27132 6018 27188 6020
rect 27132 5966 27134 6018
rect 27134 5966 27186 6018
rect 27186 5966 27188 6018
rect 27132 5964 27188 5966
rect 26796 5068 26852 5124
rect 27244 5628 27300 5684
rect 26348 4956 26404 5012
rect 26908 4956 26964 5012
rect 25900 3388 25956 3444
rect 27804 6466 27860 6468
rect 27804 6414 27806 6466
rect 27806 6414 27858 6466
rect 27858 6414 27860 6466
rect 27804 6412 27860 6414
rect 27692 5122 27748 5124
rect 27692 5070 27694 5122
rect 27694 5070 27746 5122
rect 27746 5070 27748 5122
rect 27692 5068 27748 5070
rect 28140 6412 28196 6468
rect 28476 4956 28532 5012
rect 32956 14418 33012 14420
rect 32956 14366 32958 14418
rect 32958 14366 33010 14418
rect 33010 14366 33012 14418
rect 32956 14364 33012 14366
rect 32844 14028 32900 14084
rect 32396 13970 32452 13972
rect 32396 13918 32398 13970
rect 32398 13918 32450 13970
rect 32450 13918 32452 13970
rect 32396 13916 32452 13918
rect 32284 13020 32340 13076
rect 32732 13020 32788 13076
rect 32508 12178 32564 12180
rect 32508 12126 32510 12178
rect 32510 12126 32562 12178
rect 32562 12126 32564 12178
rect 32508 12124 32564 12126
rect 32284 11900 32340 11956
rect 32732 12348 32788 12404
rect 32620 11228 32676 11284
rect 32396 10722 32452 10724
rect 32396 10670 32398 10722
rect 32398 10670 32450 10722
rect 32450 10670 32452 10722
rect 32396 10668 32452 10670
rect 33516 13020 33572 13076
rect 33180 12796 33236 12852
rect 33516 12348 33572 12404
rect 34636 14588 34692 14644
rect 36204 17724 36260 17780
rect 35756 16604 35812 16660
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35980 16268 36036 16324
rect 36204 15820 36260 15876
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35644 14642 35700 14644
rect 35644 14590 35646 14642
rect 35646 14590 35698 14642
rect 35698 14590 35700 14642
rect 35644 14588 35700 14590
rect 34748 14476 34804 14532
rect 34412 14418 34468 14420
rect 34412 14366 34414 14418
rect 34414 14366 34466 14418
rect 34466 14366 34468 14418
rect 34412 14364 34468 14366
rect 34076 14252 34132 14308
rect 34300 14140 34356 14196
rect 33964 12236 34020 12292
rect 33740 11954 33796 11956
rect 33740 11902 33742 11954
rect 33742 11902 33794 11954
rect 33794 11902 33796 11954
rect 33740 11900 33796 11902
rect 33180 11282 33236 11284
rect 33180 11230 33182 11282
rect 33182 11230 33234 11282
rect 33234 11230 33236 11282
rect 33180 11228 33236 11230
rect 33068 10668 33124 10724
rect 32620 9714 32676 9716
rect 32620 9662 32622 9714
rect 32622 9662 32674 9714
rect 32674 9662 32676 9714
rect 32620 9660 32676 9662
rect 32284 9548 32340 9604
rect 29820 7644 29876 7700
rect 29148 7532 29204 7588
rect 29372 6466 29428 6468
rect 29372 6414 29374 6466
rect 29374 6414 29426 6466
rect 29426 6414 29428 6466
rect 29372 6412 29428 6414
rect 29260 6130 29316 6132
rect 29260 6078 29262 6130
rect 29262 6078 29314 6130
rect 29314 6078 29316 6130
rect 29260 6076 29316 6078
rect 28588 4844 28644 4900
rect 27580 3612 27636 3668
rect 29372 5628 29428 5684
rect 29596 6636 29652 6692
rect 30156 6636 30212 6692
rect 30716 6690 30772 6692
rect 30716 6638 30718 6690
rect 30718 6638 30770 6690
rect 30770 6638 30772 6690
rect 30716 6636 30772 6638
rect 31388 6690 31444 6692
rect 31388 6638 31390 6690
rect 31390 6638 31442 6690
rect 31442 6638 31444 6690
rect 31388 6636 31444 6638
rect 29932 6018 29988 6020
rect 29932 5966 29934 6018
rect 29934 5966 29986 6018
rect 29986 5966 29988 6018
rect 29932 5964 29988 5966
rect 31164 6466 31220 6468
rect 31164 6414 31166 6466
rect 31166 6414 31218 6466
rect 31218 6414 31220 6466
rect 31164 6412 31220 6414
rect 30492 5964 30548 6020
rect 29372 5122 29428 5124
rect 29372 5070 29374 5122
rect 29374 5070 29426 5122
rect 29426 5070 29428 5122
rect 29372 5068 29428 5070
rect 30716 6076 30772 6132
rect 32172 6076 32228 6132
rect 32508 7362 32564 7364
rect 32508 7310 32510 7362
rect 32510 7310 32562 7362
rect 32562 7310 32564 7362
rect 32508 7308 32564 7310
rect 33292 9772 33348 9828
rect 32844 9324 32900 9380
rect 33180 9548 33236 9604
rect 33180 9212 33236 9268
rect 35196 14364 35252 14420
rect 35532 14476 35588 14532
rect 34076 11900 34132 11956
rect 34188 12290 34244 12292
rect 34188 12238 34190 12290
rect 34190 12238 34242 12290
rect 34242 12238 34244 12290
rect 34188 12236 34244 12238
rect 34860 12290 34916 12292
rect 34860 12238 34862 12290
rect 34862 12238 34914 12290
rect 34914 12238 34916 12290
rect 34860 12236 34916 12238
rect 34412 12178 34468 12180
rect 34412 12126 34414 12178
rect 34414 12126 34466 12178
rect 34466 12126 34468 12178
rect 34412 12124 34468 12126
rect 34412 11900 34468 11956
rect 34524 10610 34580 10612
rect 34524 10558 34526 10610
rect 34526 10558 34578 10610
rect 34578 10558 34580 10610
rect 34524 10556 34580 10558
rect 33852 10108 33908 10164
rect 33628 9938 33684 9940
rect 33628 9886 33630 9938
rect 33630 9886 33682 9938
rect 33682 9886 33684 9938
rect 33628 9884 33684 9886
rect 34188 9826 34244 9828
rect 34188 9774 34190 9826
rect 34190 9774 34242 9826
rect 34242 9774 34244 9826
rect 34188 9772 34244 9774
rect 33964 9714 34020 9716
rect 33964 9662 33966 9714
rect 33966 9662 34018 9714
rect 34018 9662 34020 9714
rect 33964 9660 34020 9662
rect 33628 8764 33684 8820
rect 32732 6690 32788 6692
rect 32732 6638 32734 6690
rect 32734 6638 32786 6690
rect 32786 6638 32788 6690
rect 32732 6636 32788 6638
rect 33852 7308 33908 7364
rect 33852 6860 33908 6916
rect 34188 6860 34244 6916
rect 34412 9938 34468 9940
rect 34412 9886 34414 9938
rect 34414 9886 34466 9938
rect 34466 9886 34468 9938
rect 34412 9884 34468 9886
rect 34524 9548 34580 9604
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35868 14418 35924 14420
rect 35868 14366 35870 14418
rect 35870 14366 35922 14418
rect 35922 14366 35924 14418
rect 35868 14364 35924 14366
rect 36092 14140 36148 14196
rect 37324 19906 37380 19908
rect 37324 19854 37326 19906
rect 37326 19854 37378 19906
rect 37378 19854 37380 19906
rect 37324 19852 37380 19854
rect 38444 19010 38500 19012
rect 38444 18958 38446 19010
rect 38446 18958 38498 19010
rect 38498 18958 38500 19010
rect 38444 18956 38500 18958
rect 37660 18508 37716 18564
rect 37100 18060 37156 18116
rect 37212 16940 37268 16996
rect 36988 15820 37044 15876
rect 37100 16156 37156 16212
rect 36316 15372 36372 15428
rect 35868 13580 35924 13636
rect 35756 13020 35812 13076
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34972 11564 35028 11620
rect 34748 10722 34804 10724
rect 34748 10670 34750 10722
rect 34750 10670 34802 10722
rect 34802 10670 34804 10722
rect 34748 10668 34804 10670
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35420 9996 35476 10052
rect 34636 9324 34692 9380
rect 34524 8764 34580 8820
rect 35644 11564 35700 11620
rect 35980 12348 36036 12404
rect 39228 23324 39284 23380
rect 40572 26236 40628 26292
rect 40236 26124 40292 26180
rect 39900 25228 39956 25284
rect 39788 24892 39844 24948
rect 41132 26908 41188 26964
rect 41132 25452 41188 25508
rect 41020 24892 41076 24948
rect 39340 23212 39396 23268
rect 38780 21084 38836 21140
rect 38668 20802 38724 20804
rect 38668 20750 38670 20802
rect 38670 20750 38722 20802
rect 38722 20750 38724 20802
rect 38668 20748 38724 20750
rect 39228 21532 39284 21588
rect 41468 26962 41524 26964
rect 41468 26910 41470 26962
rect 41470 26910 41522 26962
rect 41522 26910 41524 26962
rect 41468 26908 41524 26910
rect 41356 26236 41412 26292
rect 42028 29202 42084 29204
rect 42028 29150 42030 29202
rect 42030 29150 42082 29202
rect 42082 29150 42084 29202
rect 42028 29148 42084 29150
rect 41580 25506 41636 25508
rect 41580 25454 41582 25506
rect 41582 25454 41634 25506
rect 41634 25454 41636 25506
rect 41580 25452 41636 25454
rect 41356 24946 41412 24948
rect 41356 24894 41358 24946
rect 41358 24894 41410 24946
rect 41410 24894 41412 24946
rect 41356 24892 41412 24894
rect 41804 24892 41860 24948
rect 41580 23938 41636 23940
rect 41580 23886 41582 23938
rect 41582 23886 41634 23938
rect 41634 23886 41636 23938
rect 41580 23884 41636 23886
rect 39676 23100 39732 23156
rect 39676 22092 39732 22148
rect 39004 21084 39060 21140
rect 39564 20972 39620 21028
rect 39116 20860 39172 20916
rect 38892 20300 38948 20356
rect 39004 20412 39060 20468
rect 39228 20300 39284 20356
rect 38780 19234 38836 19236
rect 38780 19182 38782 19234
rect 38782 19182 38834 19234
rect 38834 19182 38836 19234
rect 38780 19180 38836 19182
rect 38556 18396 38612 18452
rect 39228 18172 39284 18228
rect 39228 17948 39284 18004
rect 38220 16940 38276 16996
rect 40348 21756 40404 21812
rect 39788 20690 39844 20692
rect 39788 20638 39790 20690
rect 39790 20638 39842 20690
rect 39842 20638 39844 20690
rect 39788 20636 39844 20638
rect 40012 20412 40068 20468
rect 39676 19292 39732 19348
rect 40012 18956 40068 19012
rect 39676 17724 39732 17780
rect 39340 17500 39396 17556
rect 37996 16828 38052 16884
rect 39004 16882 39060 16884
rect 39004 16830 39006 16882
rect 39006 16830 39058 16882
rect 39058 16830 39060 16882
rect 39004 16828 39060 16830
rect 38108 16322 38164 16324
rect 38108 16270 38110 16322
rect 38110 16270 38162 16322
rect 38162 16270 38164 16322
rect 38108 16268 38164 16270
rect 37772 15148 37828 15204
rect 37100 15036 37156 15092
rect 36428 13970 36484 13972
rect 36428 13918 36430 13970
rect 36430 13918 36482 13970
rect 36482 13918 36484 13970
rect 36428 13916 36484 13918
rect 37100 13970 37156 13972
rect 37100 13918 37102 13970
rect 37102 13918 37154 13970
rect 37154 13918 37156 13970
rect 37100 13916 37156 13918
rect 37548 14140 37604 14196
rect 38220 14588 38276 14644
rect 38332 15260 38388 15316
rect 38556 15426 38612 15428
rect 38556 15374 38558 15426
rect 38558 15374 38610 15426
rect 38610 15374 38612 15426
rect 38556 15372 38612 15374
rect 39788 16828 39844 16884
rect 39116 16770 39172 16772
rect 39116 16718 39118 16770
rect 39118 16718 39170 16770
rect 39170 16718 39172 16770
rect 39116 16716 39172 16718
rect 39116 15314 39172 15316
rect 39116 15262 39118 15314
rect 39118 15262 39170 15314
rect 39170 15262 39172 15314
rect 39116 15260 39172 15262
rect 38668 15202 38724 15204
rect 38668 15150 38670 15202
rect 38670 15150 38722 15202
rect 38722 15150 38724 15202
rect 38668 15148 38724 15150
rect 39900 14588 39956 14644
rect 38668 14364 38724 14420
rect 37996 13804 38052 13860
rect 38892 13804 38948 13860
rect 38108 13580 38164 13636
rect 36316 13020 36372 13076
rect 37100 12348 37156 12404
rect 35868 12290 35924 12292
rect 35868 12238 35870 12290
rect 35870 12238 35922 12290
rect 35922 12238 35924 12290
rect 35868 12236 35924 12238
rect 36316 12124 36372 12180
rect 35756 9826 35812 9828
rect 35756 9774 35758 9826
rect 35758 9774 35810 9826
rect 35810 9774 35812 9826
rect 35756 9772 35812 9774
rect 35196 9266 35252 9268
rect 35196 9214 35198 9266
rect 35198 9214 35250 9266
rect 35250 9214 35252 9266
rect 35196 9212 35252 9214
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 36092 6972 36148 7028
rect 35196 6748 35252 6804
rect 34076 6466 34132 6468
rect 34076 6414 34078 6466
rect 34078 6414 34130 6466
rect 34130 6414 34132 6466
rect 34076 6412 34132 6414
rect 33292 6130 33348 6132
rect 33292 6078 33294 6130
rect 33294 6078 33346 6130
rect 33346 6078 33348 6130
rect 33292 6076 33348 6078
rect 32508 5964 32564 6020
rect 31276 5628 31332 5684
rect 30156 5010 30212 5012
rect 30156 4958 30158 5010
rect 30158 4958 30210 5010
rect 30210 4958 30212 5010
rect 30156 4956 30212 4958
rect 28700 4508 28756 4564
rect 31612 4844 31668 4900
rect 31276 4508 31332 4564
rect 30940 4284 30996 4340
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
rect 28140 3500 28196 3556
rect 28588 3554 28644 3556
rect 28588 3502 28590 3554
rect 28590 3502 28642 3554
rect 28642 3502 28644 3554
rect 28588 3500 28644 3502
rect 28924 3500 28980 3556
rect 29596 3388 29652 3444
rect 32172 4956 32228 5012
rect 32396 4338 32452 4340
rect 32396 4286 32398 4338
rect 32398 4286 32450 4338
rect 32450 4286 32452 4338
rect 32396 4284 32452 4286
rect 32956 5180 33012 5236
rect 31612 4226 31668 4228
rect 31612 4174 31614 4226
rect 31614 4174 31666 4226
rect 31666 4174 31668 4226
rect 31612 4172 31668 4174
rect 32172 4172 32228 4228
rect 31612 3554 31668 3556
rect 31612 3502 31614 3554
rect 31614 3502 31666 3554
rect 31666 3502 31668 3554
rect 31612 3500 31668 3502
rect 33740 6076 33796 6132
rect 33740 5794 33796 5796
rect 33740 5742 33742 5794
rect 33742 5742 33794 5794
rect 33794 5742 33796 5794
rect 33740 5740 33796 5742
rect 34748 6076 34804 6132
rect 34636 5906 34692 5908
rect 34636 5854 34638 5906
rect 34638 5854 34690 5906
rect 34690 5854 34692 5906
rect 34636 5852 34692 5854
rect 34300 5740 34356 5796
rect 33964 5628 34020 5684
rect 33516 5068 33572 5124
rect 33852 5122 33908 5124
rect 33852 5070 33854 5122
rect 33854 5070 33906 5122
rect 33906 5070 33908 5122
rect 33852 5068 33908 5070
rect 34748 5794 34804 5796
rect 34748 5742 34750 5794
rect 34750 5742 34802 5794
rect 34802 5742 34804 5794
rect 34748 5740 34804 5742
rect 34972 6412 35028 6468
rect 35980 6802 36036 6804
rect 35980 6750 35982 6802
rect 35982 6750 36034 6802
rect 36034 6750 36036 6802
rect 35980 6748 36036 6750
rect 35420 6466 35476 6468
rect 35420 6414 35422 6466
rect 35422 6414 35474 6466
rect 35474 6414 35476 6466
rect 35420 6412 35476 6414
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34860 5234 34916 5236
rect 34860 5182 34862 5234
rect 34862 5182 34914 5234
rect 34914 5182 34916 5234
rect 34860 5180 34916 5182
rect 34972 4956 35028 5012
rect 35868 6466 35924 6468
rect 35868 6414 35870 6466
rect 35870 6414 35922 6466
rect 35922 6414 35924 6466
rect 35868 6412 35924 6414
rect 35644 6076 35700 6132
rect 37212 12178 37268 12180
rect 37212 12126 37214 12178
rect 37214 12126 37266 12178
rect 37266 12126 37268 12178
rect 37212 12124 37268 12126
rect 36764 11900 36820 11956
rect 36428 11116 36484 11172
rect 36540 11564 36596 11620
rect 36876 11282 36932 11284
rect 36876 11230 36878 11282
rect 36878 11230 36930 11282
rect 36930 11230 36932 11282
rect 36876 11228 36932 11230
rect 37100 11170 37156 11172
rect 37100 11118 37102 11170
rect 37102 11118 37154 11170
rect 37154 11118 37156 11170
rect 37100 11116 37156 11118
rect 37996 12402 38052 12404
rect 37996 12350 37998 12402
rect 37998 12350 38050 12402
rect 38050 12350 38052 12402
rect 37996 12348 38052 12350
rect 37772 12178 37828 12180
rect 37772 12126 37774 12178
rect 37774 12126 37826 12178
rect 37826 12126 37828 12178
rect 37772 12124 37828 12126
rect 38444 12236 38500 12292
rect 37996 11900 38052 11956
rect 36652 9996 36708 10052
rect 36988 9996 37044 10052
rect 38780 12178 38836 12180
rect 38780 12126 38782 12178
rect 38782 12126 38834 12178
rect 38834 12126 38836 12178
rect 38780 12124 38836 12126
rect 38444 10834 38500 10836
rect 38444 10782 38446 10834
rect 38446 10782 38498 10834
rect 38498 10782 38500 10834
rect 38444 10780 38500 10782
rect 39788 13858 39844 13860
rect 39788 13806 39790 13858
rect 39790 13806 39842 13858
rect 39842 13806 39844 13858
rect 39788 13804 39844 13806
rect 40236 17948 40292 18004
rect 40796 21420 40852 21476
rect 40684 20748 40740 20804
rect 41020 21810 41076 21812
rect 41020 21758 41022 21810
rect 41022 21758 41074 21810
rect 41074 21758 41076 21810
rect 41020 21756 41076 21758
rect 41244 22988 41300 23044
rect 42140 28700 42196 28756
rect 42700 29426 42756 29428
rect 42700 29374 42702 29426
rect 42702 29374 42754 29426
rect 42754 29374 42756 29426
rect 42700 29372 42756 29374
rect 42588 28588 42644 28644
rect 42700 28812 42756 28868
rect 42588 27804 42644 27860
rect 42252 27132 42308 27188
rect 42364 26962 42420 26964
rect 42364 26910 42366 26962
rect 42366 26910 42418 26962
rect 42418 26910 42420 26962
rect 42364 26908 42420 26910
rect 42812 27244 42868 27300
rect 43148 29372 43204 29428
rect 42588 26290 42644 26292
rect 42588 26238 42590 26290
rect 42590 26238 42642 26290
rect 42642 26238 42644 26290
rect 42588 26236 42644 26238
rect 42476 26124 42532 26180
rect 42588 25564 42644 25620
rect 42476 25452 42532 25508
rect 42028 24946 42084 24948
rect 42028 24894 42030 24946
rect 42030 24894 42082 24946
rect 42082 24894 42084 24946
rect 42028 24892 42084 24894
rect 42028 24556 42084 24612
rect 42252 23660 42308 23716
rect 41692 22876 41748 22932
rect 40460 20578 40516 20580
rect 40460 20526 40462 20578
rect 40462 20526 40514 20578
rect 40514 20526 40516 20578
rect 40460 20524 40516 20526
rect 41916 21474 41972 21476
rect 41916 21422 41918 21474
rect 41918 21422 41970 21474
rect 41970 21422 41972 21474
rect 41916 21420 41972 21422
rect 41804 21084 41860 21140
rect 41692 20524 41748 20580
rect 40348 17836 40404 17892
rect 40124 17724 40180 17780
rect 41804 19068 41860 19124
rect 41020 18396 41076 18452
rect 42252 23436 42308 23492
rect 42252 23042 42308 23044
rect 42252 22990 42254 23042
rect 42254 22990 42306 23042
rect 42306 22990 42308 23042
rect 42252 22988 42308 22990
rect 43260 28588 43316 28644
rect 43484 28082 43540 28084
rect 43484 28030 43486 28082
rect 43486 28030 43538 28082
rect 43538 28030 43540 28082
rect 43484 28028 43540 28030
rect 45500 32396 45556 32452
rect 45948 32786 46004 32788
rect 45948 32734 45950 32786
rect 45950 32734 46002 32786
rect 46002 32734 46004 32786
rect 45948 32732 46004 32734
rect 46172 32844 46228 32900
rect 46620 34130 46676 34132
rect 46620 34078 46622 34130
rect 46622 34078 46674 34130
rect 46674 34078 46676 34130
rect 46620 34076 46676 34078
rect 46956 34300 47012 34356
rect 47068 33068 47124 33124
rect 46844 32956 46900 33012
rect 46396 32396 46452 32452
rect 46508 32562 46564 32564
rect 46508 32510 46510 32562
rect 46510 32510 46562 32562
rect 46562 32510 46564 32562
rect 46508 32508 46564 32510
rect 44940 29314 44996 29316
rect 44940 29262 44942 29314
rect 44942 29262 44994 29314
rect 44994 29262 44996 29314
rect 44940 29260 44996 29262
rect 44044 28588 44100 28644
rect 44828 28642 44884 28644
rect 44828 28590 44830 28642
rect 44830 28590 44882 28642
rect 44882 28590 44884 28642
rect 44828 28588 44884 28590
rect 45276 28642 45332 28644
rect 45276 28590 45278 28642
rect 45278 28590 45330 28642
rect 45330 28590 45332 28642
rect 45276 28588 45332 28590
rect 44268 28028 44324 28084
rect 46060 29314 46116 29316
rect 46060 29262 46062 29314
rect 46062 29262 46114 29314
rect 46114 29262 46116 29314
rect 46060 29260 46116 29262
rect 45724 28924 45780 28980
rect 44380 27746 44436 27748
rect 44380 27694 44382 27746
rect 44382 27694 44434 27746
rect 44434 27694 44436 27746
rect 44380 27692 44436 27694
rect 43596 27244 43652 27300
rect 44268 27244 44324 27300
rect 43372 27074 43428 27076
rect 43372 27022 43374 27074
rect 43374 27022 43426 27074
rect 43426 27022 43428 27074
rect 43372 27020 43428 27022
rect 43932 27074 43988 27076
rect 43932 27022 43934 27074
rect 43934 27022 43986 27074
rect 43986 27022 43988 27074
rect 43932 27020 43988 27022
rect 44828 27186 44884 27188
rect 44828 27134 44830 27186
rect 44830 27134 44882 27186
rect 44882 27134 44884 27186
rect 44828 27132 44884 27134
rect 43932 26178 43988 26180
rect 43932 26126 43934 26178
rect 43934 26126 43986 26178
rect 43986 26126 43988 26178
rect 43932 26124 43988 26126
rect 44044 25452 44100 25508
rect 42700 24556 42756 24612
rect 42476 23660 42532 23716
rect 42588 23436 42644 23492
rect 42924 23154 42980 23156
rect 42924 23102 42926 23154
rect 42926 23102 42978 23154
rect 42978 23102 42980 23154
rect 42924 23100 42980 23102
rect 43148 23100 43204 23156
rect 43036 22258 43092 22260
rect 43036 22206 43038 22258
rect 43038 22206 43090 22258
rect 43090 22206 43092 22258
rect 43036 22204 43092 22206
rect 42028 19964 42084 20020
rect 42140 20524 42196 20580
rect 42028 18956 42084 19012
rect 41916 18620 41972 18676
rect 41020 17948 41076 18004
rect 41020 16994 41076 16996
rect 41020 16942 41022 16994
rect 41022 16942 41074 16994
rect 41074 16942 41076 16994
rect 41020 16940 41076 16942
rect 42812 20802 42868 20804
rect 42812 20750 42814 20802
rect 42814 20750 42866 20802
rect 42866 20750 42868 20802
rect 42812 20748 42868 20750
rect 43596 23884 43652 23940
rect 43820 23884 43876 23940
rect 43484 23436 43540 23492
rect 43596 23154 43652 23156
rect 43596 23102 43598 23154
rect 43598 23102 43650 23154
rect 43650 23102 43652 23154
rect 43596 23100 43652 23102
rect 43596 22146 43652 22148
rect 43596 22094 43598 22146
rect 43598 22094 43650 22146
rect 43650 22094 43652 22146
rect 43596 22092 43652 22094
rect 44268 27020 44324 27076
rect 44940 27020 44996 27076
rect 46060 27746 46116 27748
rect 46060 27694 46062 27746
rect 46062 27694 46114 27746
rect 46114 27694 46116 27746
rect 46060 27692 46116 27694
rect 46060 27074 46116 27076
rect 46060 27022 46062 27074
rect 46062 27022 46114 27074
rect 46114 27022 46116 27074
rect 46060 27020 46116 27022
rect 47852 40348 47908 40404
rect 47628 38332 47684 38388
rect 47964 39676 48020 39732
rect 48188 41410 48244 41412
rect 48188 41358 48190 41410
rect 48190 41358 48242 41410
rect 48242 41358 48244 41410
rect 48188 41356 48244 41358
rect 47740 37660 47796 37716
rect 47740 35644 47796 35700
rect 47628 35084 47684 35140
rect 47964 34972 48020 35028
rect 48188 35980 48244 36036
rect 48300 35756 48356 35812
rect 48412 37772 48468 37828
rect 48188 33458 48244 33460
rect 48188 33406 48190 33458
rect 48190 33406 48242 33458
rect 48242 33406 48244 33458
rect 48188 33404 48244 33406
rect 48188 32844 48244 32900
rect 47516 31218 47572 31220
rect 47516 31166 47518 31218
rect 47518 31166 47570 31218
rect 47570 31166 47572 31218
rect 47516 31164 47572 31166
rect 47740 31052 47796 31108
rect 45612 25618 45668 25620
rect 45612 25566 45614 25618
rect 45614 25566 45666 25618
rect 45666 25566 45668 25618
rect 45612 25564 45668 25566
rect 45052 25452 45108 25508
rect 44828 24108 44884 24164
rect 44604 23436 44660 23492
rect 44492 23042 44548 23044
rect 44492 22990 44494 23042
rect 44494 22990 44546 23042
rect 44546 22990 44548 23042
rect 44492 22988 44548 22990
rect 44940 23772 44996 23828
rect 45724 25506 45780 25508
rect 45724 25454 45726 25506
rect 45726 25454 45778 25506
rect 45778 25454 45780 25506
rect 45724 25452 45780 25454
rect 45724 25228 45780 25284
rect 45612 24834 45668 24836
rect 45612 24782 45614 24834
rect 45614 24782 45666 24834
rect 45666 24782 45668 24834
rect 45612 24780 45668 24782
rect 45836 24892 45892 24948
rect 45276 23938 45332 23940
rect 45276 23886 45278 23938
rect 45278 23886 45330 23938
rect 45330 23886 45332 23938
rect 45276 23884 45332 23886
rect 46956 25394 47012 25396
rect 46956 25342 46958 25394
rect 46958 25342 47010 25394
rect 47010 25342 47012 25394
rect 46956 25340 47012 25342
rect 47516 25394 47572 25396
rect 47516 25342 47518 25394
rect 47518 25342 47570 25394
rect 47570 25342 47572 25394
rect 47516 25340 47572 25342
rect 46844 24722 46900 24724
rect 46844 24670 46846 24722
rect 46846 24670 46898 24722
rect 46898 24670 46900 24722
rect 46844 24668 46900 24670
rect 46732 24556 46788 24612
rect 47180 24946 47236 24948
rect 47180 24894 47182 24946
rect 47182 24894 47234 24946
rect 47234 24894 47236 24946
rect 47180 24892 47236 24894
rect 47292 24722 47348 24724
rect 47292 24670 47294 24722
rect 47294 24670 47346 24722
rect 47346 24670 47348 24722
rect 47292 24668 47348 24670
rect 47068 24108 47124 24164
rect 46172 23826 46228 23828
rect 46172 23774 46174 23826
rect 46174 23774 46226 23826
rect 46226 23774 46228 23826
rect 46172 23772 46228 23774
rect 45276 23660 45332 23716
rect 45500 23548 45556 23604
rect 45276 22988 45332 23044
rect 44156 22092 44212 22148
rect 43596 21084 43652 21140
rect 43260 20524 43316 20580
rect 42700 19122 42756 19124
rect 42700 19070 42702 19122
rect 42702 19070 42754 19122
rect 42754 19070 42756 19122
rect 42700 19068 42756 19070
rect 42924 18508 42980 18564
rect 42700 18396 42756 18452
rect 42588 18060 42644 18116
rect 42252 17778 42308 17780
rect 42252 17726 42254 17778
rect 42254 17726 42306 17778
rect 42306 17726 42308 17778
rect 42252 17724 42308 17726
rect 43484 19404 43540 19460
rect 43036 17724 43092 17780
rect 43148 17948 43204 18004
rect 43484 17724 43540 17780
rect 44156 20748 44212 20804
rect 43708 19292 43764 19348
rect 43932 19628 43988 19684
rect 44268 19964 44324 20020
rect 44940 19964 44996 20020
rect 44828 19852 44884 19908
rect 44716 19404 44772 19460
rect 44268 18732 44324 18788
rect 41916 16940 41972 16996
rect 40908 16882 40964 16884
rect 40908 16830 40910 16882
rect 40910 16830 40962 16882
rect 40962 16830 40964 16882
rect 40908 16828 40964 16830
rect 41020 16716 41076 16772
rect 40460 15986 40516 15988
rect 40460 15934 40462 15986
rect 40462 15934 40514 15986
rect 40514 15934 40516 15986
rect 40460 15932 40516 15934
rect 41356 16716 41412 16772
rect 42140 16716 42196 16772
rect 41916 16156 41972 16212
rect 42364 16210 42420 16212
rect 42364 16158 42366 16210
rect 42366 16158 42418 16210
rect 42418 16158 42420 16210
rect 42364 16156 42420 16158
rect 42140 16044 42196 16100
rect 42812 17052 42868 17108
rect 43036 17388 43092 17444
rect 43372 17442 43428 17444
rect 43372 17390 43374 17442
rect 43374 17390 43426 17442
rect 43426 17390 43428 17442
rect 43372 17388 43428 17390
rect 43260 17164 43316 17220
rect 43036 16770 43092 16772
rect 43036 16718 43038 16770
rect 43038 16718 43090 16770
rect 43090 16718 43092 16770
rect 43036 16716 43092 16718
rect 43260 16268 43316 16324
rect 43820 16994 43876 16996
rect 43820 16942 43822 16994
rect 43822 16942 43874 16994
rect 43874 16942 43876 16994
rect 43820 16940 43876 16942
rect 43372 16156 43428 16212
rect 43484 16604 43540 16660
rect 42812 16098 42868 16100
rect 42812 16046 42814 16098
rect 42814 16046 42866 16098
rect 42866 16046 42868 16098
rect 42812 16044 42868 16046
rect 42476 15932 42532 15988
rect 43036 15932 43092 15988
rect 41692 15260 41748 15316
rect 42364 15314 42420 15316
rect 42364 15262 42366 15314
rect 42366 15262 42418 15314
rect 42418 15262 42420 15314
rect 42364 15260 42420 15262
rect 43372 15372 43428 15428
rect 40012 14364 40068 14420
rect 40684 14364 40740 14420
rect 39900 13692 39956 13748
rect 40124 13804 40180 13860
rect 40236 13244 40292 13300
rect 40236 12962 40292 12964
rect 40236 12910 40238 12962
rect 40238 12910 40290 12962
rect 40290 12910 40292 12962
rect 40236 12908 40292 12910
rect 40236 12460 40292 12516
rect 38892 10780 38948 10836
rect 39116 12124 39172 12180
rect 40572 13692 40628 13748
rect 41468 14588 41524 14644
rect 40908 14476 40964 14532
rect 41244 14418 41300 14420
rect 41244 14366 41246 14418
rect 41246 14366 41298 14418
rect 41298 14366 41300 14418
rect 41244 14364 41300 14366
rect 41356 14306 41412 14308
rect 41356 14254 41358 14306
rect 41358 14254 41410 14306
rect 41410 14254 41412 14306
rect 41356 14252 41412 14254
rect 41580 14364 41636 14420
rect 43148 15314 43204 15316
rect 43148 15262 43150 15314
rect 43150 15262 43202 15314
rect 43202 15262 43204 15314
rect 43148 15260 43204 15262
rect 42588 14364 42644 14420
rect 41132 13858 41188 13860
rect 41132 13806 41134 13858
rect 41134 13806 41186 13858
rect 41186 13806 41188 13858
rect 41132 13804 41188 13806
rect 41244 13244 41300 13300
rect 41468 13746 41524 13748
rect 41468 13694 41470 13746
rect 41470 13694 41522 13746
rect 41522 13694 41524 13746
rect 41468 13692 41524 13694
rect 41916 13746 41972 13748
rect 41916 13694 41918 13746
rect 41918 13694 41970 13746
rect 41970 13694 41972 13746
rect 41916 13692 41972 13694
rect 42476 14252 42532 14308
rect 43260 13804 43316 13860
rect 42700 13746 42756 13748
rect 42700 13694 42702 13746
rect 42702 13694 42754 13746
rect 42754 13694 42756 13746
rect 42700 13692 42756 13694
rect 37324 10220 37380 10276
rect 37884 10220 37940 10276
rect 37772 9996 37828 10052
rect 37324 9772 37380 9828
rect 37884 9714 37940 9716
rect 37884 9662 37886 9714
rect 37886 9662 37938 9714
rect 37938 9662 37940 9714
rect 37884 9660 37940 9662
rect 36876 8930 36932 8932
rect 36876 8878 36878 8930
rect 36878 8878 36930 8930
rect 36930 8878 36932 8930
rect 36876 8876 36932 8878
rect 37996 9772 38052 9828
rect 36652 8764 36708 8820
rect 37436 8764 37492 8820
rect 38220 10108 38276 10164
rect 41356 12460 41412 12516
rect 42252 12460 42308 12516
rect 43820 16716 43876 16772
rect 44044 17724 44100 17780
rect 44268 17666 44324 17668
rect 44268 17614 44270 17666
rect 44270 17614 44322 17666
rect 44322 17614 44324 17666
rect 44268 17612 44324 17614
rect 44156 17500 44212 17556
rect 44044 17106 44100 17108
rect 44044 17054 44046 17106
rect 44046 17054 44098 17106
rect 44098 17054 44100 17106
rect 44044 17052 44100 17054
rect 44604 18562 44660 18564
rect 44604 18510 44606 18562
rect 44606 18510 44658 18562
rect 44658 18510 44660 18562
rect 44604 18508 44660 18510
rect 44940 19346 44996 19348
rect 44940 19294 44942 19346
rect 44942 19294 44994 19346
rect 44994 19294 44996 19346
rect 44940 19292 44996 19294
rect 45276 20802 45332 20804
rect 45276 20750 45278 20802
rect 45278 20750 45330 20802
rect 45330 20750 45332 20802
rect 45276 20748 45332 20750
rect 45836 22988 45892 23044
rect 45164 20188 45220 20244
rect 46060 20860 46116 20916
rect 47068 23714 47124 23716
rect 47068 23662 47070 23714
rect 47070 23662 47122 23714
rect 47122 23662 47124 23714
rect 47068 23660 47124 23662
rect 47516 23660 47572 23716
rect 45164 19740 45220 19796
rect 44828 18450 44884 18452
rect 44828 18398 44830 18450
rect 44830 18398 44882 18450
rect 44882 18398 44884 18450
rect 44828 18396 44884 18398
rect 44828 18172 44884 18228
rect 45052 17724 45108 17780
rect 45052 17388 45108 17444
rect 43932 15932 43988 15988
rect 43932 15426 43988 15428
rect 43932 15374 43934 15426
rect 43934 15374 43986 15426
rect 43986 15374 43988 15426
rect 43932 15372 43988 15374
rect 45052 16492 45108 16548
rect 44156 15260 44212 15316
rect 44380 15148 44436 15204
rect 39228 10780 39284 10836
rect 38780 10108 38836 10164
rect 39228 9996 39284 10052
rect 39340 9884 39396 9940
rect 39564 9884 39620 9940
rect 38556 9602 38612 9604
rect 38556 9550 38558 9602
rect 38558 9550 38610 9602
rect 38610 9550 38612 9602
rect 38556 9548 38612 9550
rect 43708 14700 43764 14756
rect 43596 13020 43652 13076
rect 41356 9938 41412 9940
rect 41356 9886 41358 9938
rect 41358 9886 41410 9938
rect 41410 9886 41412 9938
rect 41356 9884 41412 9886
rect 43708 12290 43764 12292
rect 43708 12238 43710 12290
rect 43710 12238 43762 12290
rect 43762 12238 43764 12290
rect 43708 12236 43764 12238
rect 45052 15148 45108 15204
rect 44268 14642 44324 14644
rect 44268 14590 44270 14642
rect 44270 14590 44322 14642
rect 44322 14590 44324 14642
rect 44268 14588 44324 14590
rect 45276 15314 45332 15316
rect 45276 15262 45278 15314
rect 45278 15262 45330 15314
rect 45330 15262 45332 15314
rect 45276 15260 45332 15262
rect 45164 14700 45220 14756
rect 44828 14418 44884 14420
rect 44828 14366 44830 14418
rect 44830 14366 44882 14418
rect 44882 14366 44884 14418
rect 44828 14364 44884 14366
rect 45948 19740 46004 19796
rect 46396 20076 46452 20132
rect 46620 20018 46676 20020
rect 46620 19966 46622 20018
rect 46622 19966 46674 20018
rect 46674 19966 46676 20018
rect 46620 19964 46676 19966
rect 46844 19964 46900 20020
rect 45612 18172 45668 18228
rect 45836 18396 45892 18452
rect 45612 16604 45668 16660
rect 45500 16044 45556 16100
rect 45836 17500 45892 17556
rect 45836 17052 45892 17108
rect 45612 15148 45668 15204
rect 47628 24556 47684 24612
rect 47628 23548 47684 23604
rect 48188 28588 48244 28644
rect 48188 27244 48244 27300
rect 48076 27020 48132 27076
rect 47852 26236 47908 26292
rect 47852 25282 47908 25284
rect 47852 25230 47854 25282
rect 47854 25230 47906 25282
rect 47906 25230 47908 25282
rect 47852 25228 47908 25230
rect 48188 24892 48244 24948
rect 48188 24610 48244 24612
rect 48188 24558 48190 24610
rect 48190 24558 48242 24610
rect 48242 24558 48244 24610
rect 48188 24556 48244 24558
rect 46844 19010 46900 19012
rect 46844 18958 46846 19010
rect 46846 18958 46898 19010
rect 46898 18958 46900 19010
rect 46844 18956 46900 18958
rect 46284 18060 46340 18116
rect 46732 18060 46788 18116
rect 46844 18172 46900 18228
rect 46620 17666 46676 17668
rect 46620 17614 46622 17666
rect 46622 17614 46674 17666
rect 46674 17614 46676 17666
rect 46620 17612 46676 17614
rect 46172 16940 46228 16996
rect 45948 14812 46004 14868
rect 46732 17052 46788 17108
rect 46956 17666 47012 17668
rect 46956 17614 46958 17666
rect 46958 17614 47010 17666
rect 47010 17614 47012 17666
rect 46956 17612 47012 17614
rect 47180 20018 47236 20020
rect 47180 19966 47182 20018
rect 47182 19966 47234 20018
rect 47234 19966 47236 20018
rect 47180 19964 47236 19966
rect 48188 23042 48244 23044
rect 48188 22990 48190 23042
rect 48190 22990 48242 23042
rect 48242 22990 48244 23042
rect 48188 22988 48244 22990
rect 47964 22876 48020 22932
rect 48188 20914 48244 20916
rect 48188 20862 48190 20914
rect 48190 20862 48242 20914
rect 48242 20862 48244 20914
rect 48188 20860 48244 20862
rect 47964 20188 48020 20244
rect 48076 20748 48132 20804
rect 47852 19852 47908 19908
rect 48076 19628 48132 19684
rect 47068 18956 47124 19012
rect 46620 16380 46676 16436
rect 45388 14028 45444 14084
rect 44380 13970 44436 13972
rect 44380 13918 44382 13970
rect 44382 13918 44434 13970
rect 44434 13918 44436 13970
rect 44380 13916 44436 13918
rect 45724 14418 45780 14420
rect 45724 14366 45726 14418
rect 45726 14366 45778 14418
rect 45778 14366 45780 14418
rect 45724 14364 45780 14366
rect 44604 13804 44660 13860
rect 45276 13580 45332 13636
rect 44156 12236 44212 12292
rect 44380 12290 44436 12292
rect 44380 12238 44382 12290
rect 44382 12238 44434 12290
rect 44434 12238 44436 12290
rect 44380 12236 44436 12238
rect 43932 10892 43988 10948
rect 44940 12402 44996 12404
rect 44940 12350 44942 12402
rect 44942 12350 44994 12402
rect 44994 12350 44996 12402
rect 44940 12348 44996 12350
rect 45052 12290 45108 12292
rect 45052 12238 45054 12290
rect 45054 12238 45106 12290
rect 45106 12238 45108 12290
rect 45052 12236 45108 12238
rect 45948 14028 46004 14084
rect 45836 13020 45892 13076
rect 46060 13020 46116 13076
rect 45836 12348 45892 12404
rect 47292 18284 47348 18340
rect 47404 18060 47460 18116
rect 47516 18396 47572 18452
rect 47628 18338 47684 18340
rect 47628 18286 47630 18338
rect 47630 18286 47682 18338
rect 47682 18286 47684 18338
rect 47628 18284 47684 18286
rect 47628 17612 47684 17668
rect 47628 17164 47684 17220
rect 46956 15314 47012 15316
rect 46956 15262 46958 15314
rect 46958 15262 47010 15314
rect 47010 15262 47012 15314
rect 46956 15260 47012 15262
rect 47852 17164 47908 17220
rect 47964 16156 48020 16212
rect 48076 16604 48132 16660
rect 48188 17500 48244 17556
rect 47964 15932 48020 15988
rect 47068 14418 47124 14420
rect 47068 14366 47070 14418
rect 47070 14366 47122 14418
rect 47122 14366 47124 14418
rect 47068 14364 47124 14366
rect 46508 13634 46564 13636
rect 46508 13582 46510 13634
rect 46510 13582 46562 13634
rect 46562 13582 46564 13634
rect 46508 13580 46564 13582
rect 46844 13692 46900 13748
rect 46956 14028 47012 14084
rect 46620 13020 46676 13076
rect 44716 10892 44772 10948
rect 44044 10498 44100 10500
rect 44044 10446 44046 10498
rect 44046 10446 44098 10498
rect 44098 10446 44100 10498
rect 44044 10444 44100 10446
rect 42588 9602 42644 9604
rect 42588 9550 42590 9602
rect 42590 9550 42642 9602
rect 42642 9550 42644 9602
rect 42588 9548 42644 9550
rect 38220 8876 38276 8932
rect 38332 7644 38388 7700
rect 38220 7420 38276 7476
rect 36316 6972 36372 7028
rect 37548 6972 37604 7028
rect 36540 6860 36596 6916
rect 42028 8540 42084 8596
rect 43148 8876 43204 8932
rect 43932 9772 43988 9828
rect 39004 8092 39060 8148
rect 38892 7698 38948 7700
rect 38892 7646 38894 7698
rect 38894 7646 38946 7698
rect 38946 7646 38948 7698
rect 38892 7644 38948 7646
rect 40348 8146 40404 8148
rect 40348 8094 40350 8146
rect 40350 8094 40402 8146
rect 40402 8094 40404 8146
rect 40348 8092 40404 8094
rect 36204 6076 36260 6132
rect 36316 5794 36372 5796
rect 36316 5742 36318 5794
rect 36318 5742 36370 5794
rect 36370 5742 36372 5794
rect 36316 5740 36372 5742
rect 38892 6130 38948 6132
rect 38892 6078 38894 6130
rect 38894 6078 38946 6130
rect 38946 6078 38948 6130
rect 38892 6076 38948 6078
rect 40348 6130 40404 6132
rect 40348 6078 40350 6130
rect 40350 6078 40402 6130
rect 40402 6078 40404 6130
rect 40348 6076 40404 6078
rect 42812 8258 42868 8260
rect 42812 8206 42814 8258
rect 42814 8206 42866 8258
rect 42866 8206 42868 8258
rect 42812 8204 42868 8206
rect 43036 8146 43092 8148
rect 43036 8094 43038 8146
rect 43038 8094 43090 8146
rect 43090 8094 43092 8146
rect 43036 8092 43092 8094
rect 42140 7980 42196 8036
rect 42924 7868 42980 7924
rect 44940 10668 44996 10724
rect 44156 9602 44212 9604
rect 44156 9550 44158 9602
rect 44158 9550 44210 9602
rect 44210 9550 44212 9602
rect 44156 9548 44212 9550
rect 44604 8930 44660 8932
rect 44604 8878 44606 8930
rect 44606 8878 44658 8930
rect 44658 8878 44660 8930
rect 44604 8876 44660 8878
rect 45164 10444 45220 10500
rect 46060 10444 46116 10500
rect 45612 9826 45668 9828
rect 45612 9774 45614 9826
rect 45614 9774 45666 9826
rect 45666 9774 45668 9826
rect 45612 9772 45668 9774
rect 45052 8204 45108 8260
rect 43820 8146 43876 8148
rect 43820 8094 43822 8146
rect 43822 8094 43874 8146
rect 43874 8094 43876 8146
rect 43820 8092 43876 8094
rect 45836 8258 45892 8260
rect 45836 8206 45838 8258
rect 45838 8206 45890 8258
rect 45890 8206 45892 8258
rect 45836 8204 45892 8206
rect 43708 8034 43764 8036
rect 43708 7982 43710 8034
rect 43710 7982 43762 8034
rect 43762 7982 43764 8034
rect 43708 7980 43764 7982
rect 42700 7474 42756 7476
rect 42700 7422 42702 7474
rect 42702 7422 42754 7474
rect 42754 7422 42756 7474
rect 42700 7420 42756 7422
rect 43596 7420 43652 7476
rect 43148 6860 43204 6916
rect 43932 6636 43988 6692
rect 41020 6076 41076 6132
rect 35532 4508 35588 4564
rect 36652 4956 36708 5012
rect 35644 4284 35700 4340
rect 33292 4226 33348 4228
rect 33292 4174 33294 4226
rect 33294 4174 33346 4226
rect 33346 4174 33348 4226
rect 33292 4172 33348 4174
rect 35084 4172 35140 4228
rect 34300 3612 34356 3668
rect 33628 3500 33684 3556
rect 33740 3442 33796 3444
rect 33740 3390 33742 3442
rect 33742 3390 33794 3442
rect 33794 3390 33796 3442
rect 33740 3388 33796 3390
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35420 3554 35476 3556
rect 35420 3502 35422 3554
rect 35422 3502 35474 3554
rect 35474 3502 35476 3554
rect 35420 3500 35476 3502
rect 37212 4562 37268 4564
rect 37212 4510 37214 4562
rect 37214 4510 37266 4562
rect 37266 4510 37268 4562
rect 37212 4508 37268 4510
rect 37436 4338 37492 4340
rect 37436 4286 37438 4338
rect 37438 4286 37490 4338
rect 37490 4286 37492 4338
rect 37436 4284 37492 4286
rect 36988 3666 37044 3668
rect 36988 3614 36990 3666
rect 36990 3614 37042 3666
rect 37042 3614 37044 3666
rect 36988 3612 37044 3614
rect 37884 3612 37940 3668
rect 37996 3500 38052 3556
rect 47404 10498 47460 10500
rect 47404 10446 47406 10498
rect 47406 10446 47458 10498
rect 47458 10446 47460 10498
rect 47404 10444 47460 10446
rect 48076 13916 48132 13972
rect 47852 13858 47908 13860
rect 47852 13806 47854 13858
rect 47854 13806 47906 13858
rect 47906 13806 47908 13858
rect 47852 13804 47908 13806
rect 46620 8258 46676 8260
rect 46620 8206 46622 8258
rect 46622 8206 46674 8258
rect 46674 8206 46676 8258
rect 46620 8204 46676 8206
rect 48188 13746 48244 13748
rect 48188 13694 48190 13746
rect 48190 13694 48242 13746
rect 48242 13694 48244 13746
rect 48188 13692 48244 13694
rect 47964 13074 48020 13076
rect 47964 13022 47966 13074
rect 47966 13022 48018 13074
rect 48018 13022 48020 13074
rect 47964 13020 48020 13022
rect 47964 12796 48020 12852
rect 48188 12124 48244 12180
rect 47964 11506 48020 11508
rect 47964 11454 47966 11506
rect 47966 11454 48018 11506
rect 48018 11454 48020 11506
rect 47964 11452 48020 11454
rect 47628 10780 47684 10836
rect 48188 10780 48244 10836
rect 47852 10722 47908 10724
rect 47852 10670 47854 10722
rect 47854 10670 47906 10722
rect 47906 10670 47908 10722
rect 47852 10668 47908 10670
rect 47964 9436 48020 9492
rect 48188 8764 48244 8820
rect 47852 8540 47908 8596
rect 47068 8258 47124 8260
rect 47068 8206 47070 8258
rect 47070 8206 47122 8258
rect 47122 8206 47124 8258
rect 47068 8204 47124 8206
rect 46172 7980 46228 8036
rect 45612 6690 45668 6692
rect 45612 6638 45614 6690
rect 45614 6638 45666 6690
rect 45666 6638 45668 6690
rect 45612 6636 45668 6638
rect 45388 6524 45444 6580
rect 47292 6076 47348 6132
rect 41468 4956 41524 5012
rect 42700 4956 42756 5012
rect 40796 3666 40852 3668
rect 40796 3614 40798 3666
rect 40798 3614 40850 3666
rect 40850 3614 40852 3666
rect 40796 3612 40852 3614
rect 38444 3500 38500 3556
rect 39788 3554 39844 3556
rect 39788 3502 39790 3554
rect 39790 3502 39842 3554
rect 39842 3502 39844 3554
rect 39788 3500 39844 3502
rect 41692 3388 41748 3444
rect 42476 3388 42532 3444
rect 42924 3388 42980 3444
<< metal3 >>
rect 49200 49812 50000 49840
rect 44706 49756 44716 49812
rect 44772 49756 50000 49812
rect 49200 49728 50000 49756
rect 49200 49140 50000 49168
rect 45154 49084 45164 49140
rect 45220 49084 50000 49140
rect 49200 49056 50000 49084
rect 49200 48468 50000 48496
rect 44482 48412 44492 48468
rect 44548 48412 50000 48468
rect 49200 48384 50000 48412
rect 49200 47796 50000 47824
rect 44034 47740 44044 47796
rect 44100 47740 50000 47796
rect 49200 47712 50000 47740
rect 49200 47124 50000 47152
rect 45266 47068 45276 47124
rect 45332 47068 50000 47124
rect 49200 47040 50000 47068
rect 49200 46452 50000 46480
rect 47170 46396 47180 46452
rect 47236 46396 50000 46452
rect 49200 46368 50000 46396
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 16146 46060 16156 46116
rect 16212 46060 17948 46116
rect 18004 46060 18014 46116
rect 23538 46060 23548 46116
rect 23604 46060 25564 46116
rect 25620 46060 25630 46116
rect 28914 46060 28924 46116
rect 28980 46060 30044 46116
rect 30100 46060 30110 46116
rect 34962 46060 34972 46116
rect 35028 46060 36988 46116
rect 37044 46060 37054 46116
rect 40338 46060 40348 46116
rect 40404 46060 41468 46116
rect 41524 46060 41534 46116
rect 41682 46060 41692 46116
rect 41748 46060 44604 46116
rect 44660 46060 44670 46116
rect 39218 45836 39228 45892
rect 39284 45836 43708 45892
rect 43764 45836 43774 45892
rect 49200 45780 50000 45808
rect 22754 45724 22764 45780
rect 22820 45724 23772 45780
rect 23828 45724 23838 45780
rect 38210 45724 38220 45780
rect 38276 45724 39788 45780
rect 39844 45724 39854 45780
rect 43698 45724 43708 45780
rect 43764 45724 50000 45780
rect 49200 45696 50000 45724
rect 12562 45612 12572 45668
rect 12628 45612 13468 45668
rect 13524 45612 13534 45668
rect 18834 45612 18844 45668
rect 18900 45612 19852 45668
rect 19908 45612 19918 45668
rect 32498 45612 32508 45668
rect 32564 45612 34300 45668
rect 34356 45612 34366 45668
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 35186 45388 35196 45444
rect 35252 45388 43708 45444
rect 43652 45332 43708 45388
rect 16258 45276 16268 45332
rect 16324 45276 16828 45332
rect 16884 45276 16894 45332
rect 18946 45276 18956 45332
rect 19012 45276 20524 45332
rect 20580 45276 20972 45332
rect 21028 45276 21038 45332
rect 28578 45276 28588 45332
rect 28644 45276 29708 45332
rect 29764 45276 29774 45332
rect 41010 45276 41020 45332
rect 41076 45276 42252 45332
rect 42308 45276 42318 45332
rect 43652 45276 45668 45332
rect 19842 45164 19852 45220
rect 19908 45164 20748 45220
rect 20804 45164 20814 45220
rect 30818 45164 30828 45220
rect 30884 45164 31836 45220
rect 31892 45164 32172 45220
rect 32228 45164 32238 45220
rect 41122 45164 41132 45220
rect 41188 45164 44380 45220
rect 44436 45164 44446 45220
rect 0 45108 800 45136
rect 45612 45108 45668 45276
rect 49200 45108 50000 45136
rect 0 45052 4172 45108
rect 4228 45052 4238 45108
rect 14242 45052 14252 45108
rect 14308 45052 14924 45108
rect 14980 45052 17388 45108
rect 17444 45052 20188 45108
rect 20244 45052 20860 45108
rect 20916 45052 20926 45108
rect 25330 45052 25340 45108
rect 25396 45052 29372 45108
rect 29428 45052 31948 45108
rect 32004 45052 32014 45108
rect 38434 45052 38444 45108
rect 38500 45052 44156 45108
rect 44212 45052 44222 45108
rect 45612 45052 50000 45108
rect 0 45024 800 45052
rect 49200 45024 50000 45052
rect 26786 44940 26796 44996
rect 26852 44940 28140 44996
rect 28196 44940 28206 44996
rect 30594 44940 30604 44996
rect 30660 44940 32956 44996
rect 33012 44940 33022 44996
rect 42354 44940 42364 44996
rect 42420 44940 45388 44996
rect 45444 44940 45454 44996
rect 36418 44828 36428 44884
rect 36484 44828 36494 44884
rect 40114 44828 40124 44884
rect 40180 44828 45052 44884
rect 45108 44828 45118 44884
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 36428 44660 36484 44828
rect 36754 44716 36764 44772
rect 36820 44716 45164 44772
rect 45220 44716 45230 44772
rect 36428 44604 45724 44660
rect 45780 44604 45790 44660
rect 32162 44492 32172 44548
rect 32228 44492 37772 44548
rect 37828 44492 37838 44548
rect 43026 44492 43036 44548
rect 43092 44492 45836 44548
rect 45892 44492 45902 44548
rect 49200 44436 50000 44464
rect 17042 44380 17052 44436
rect 17108 44380 19516 44436
rect 19572 44380 19582 44436
rect 30930 44380 30940 44436
rect 30996 44380 34076 44436
rect 34132 44380 34142 44436
rect 43922 44380 43932 44436
rect 43988 44380 50000 44436
rect 49200 44352 50000 44380
rect 20066 44268 20076 44324
rect 20132 44268 20524 44324
rect 20580 44268 20590 44324
rect 31826 44268 31836 44324
rect 31892 44268 32620 44324
rect 32676 44268 32686 44324
rect 37986 44268 37996 44324
rect 38052 44268 41692 44324
rect 41748 44268 41758 44324
rect 18722 44156 18732 44212
rect 18788 44156 19404 44212
rect 19460 44156 19470 44212
rect 23426 44156 23436 44212
rect 23492 44156 24108 44212
rect 24164 44156 24174 44212
rect 37762 44156 37772 44212
rect 37828 44156 41244 44212
rect 41300 44156 41310 44212
rect 42802 44156 42812 44212
rect 42868 44156 47740 44212
rect 47796 44156 47806 44212
rect 18498 44044 18508 44100
rect 18564 44044 19852 44100
rect 19908 44044 19918 44100
rect 30370 44044 30380 44100
rect 30436 44044 31164 44100
rect 31220 44044 32396 44100
rect 32452 44044 32462 44100
rect 33506 44044 33516 44100
rect 33572 44044 38780 44100
rect 38836 44044 38846 44100
rect 23986 43932 23996 43988
rect 24052 43932 25004 43988
rect 25060 43932 25070 43988
rect 32498 43932 32508 43988
rect 32564 43932 33852 43988
rect 33908 43932 33918 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 19506 43820 19516 43876
rect 19572 43820 19582 43876
rect 31490 43820 31500 43876
rect 31556 43820 36988 43876
rect 37044 43820 37054 43876
rect 19516 43764 19572 43820
rect 49200 43764 50000 43792
rect 19516 43708 19740 43764
rect 19796 43708 19806 43764
rect 29922 43708 29932 43764
rect 29988 43708 31612 43764
rect 31668 43708 33628 43764
rect 33684 43708 33694 43764
rect 43810 43708 43820 43764
rect 43876 43708 50000 43764
rect 49200 43680 50000 43708
rect 14914 43596 14924 43652
rect 14980 43596 17500 43652
rect 17556 43596 17566 43652
rect 21410 43596 21420 43652
rect 21476 43596 21868 43652
rect 21924 43596 21934 43652
rect 34514 43596 34524 43652
rect 34580 43596 38332 43652
rect 38388 43596 38892 43652
rect 38948 43596 38958 43652
rect 41234 43596 41244 43652
rect 41300 43596 46844 43652
rect 46900 43596 46910 43652
rect 47170 43596 47180 43652
rect 47236 43596 47852 43652
rect 47908 43596 47918 43652
rect 4834 43484 4844 43540
rect 4900 43484 8764 43540
rect 8820 43484 11900 43540
rect 11956 43484 11966 43540
rect 16706 43484 16716 43540
rect 16772 43484 17612 43540
rect 17668 43484 17678 43540
rect 19282 43484 19292 43540
rect 19348 43484 21644 43540
rect 21700 43484 21710 43540
rect 24658 43484 24668 43540
rect 24724 43484 25564 43540
rect 25620 43484 25630 43540
rect 28018 43484 28028 43540
rect 28084 43484 28812 43540
rect 28868 43484 28878 43540
rect 30818 43484 30828 43540
rect 30884 43484 31724 43540
rect 31780 43484 33740 43540
rect 33796 43484 33806 43540
rect 38658 43484 38668 43540
rect 38724 43484 44828 43540
rect 44884 43484 44894 43540
rect 8866 43372 8876 43428
rect 8932 43372 10332 43428
rect 10388 43372 10398 43428
rect 16818 43372 16828 43428
rect 16884 43372 17724 43428
rect 17780 43372 18284 43428
rect 18340 43372 18350 43428
rect 19618 43372 19628 43428
rect 19684 43372 22092 43428
rect 22148 43372 22158 43428
rect 23426 43372 23436 43428
rect 23492 43372 25676 43428
rect 25732 43372 28364 43428
rect 28420 43372 28430 43428
rect 31266 43372 31276 43428
rect 31332 43372 31500 43428
rect 31556 43372 32284 43428
rect 32340 43372 33180 43428
rect 33236 43372 33246 43428
rect 33842 43372 33852 43428
rect 33908 43372 34412 43428
rect 34468 43372 34478 43428
rect 37426 43372 37436 43428
rect 37492 43372 41244 43428
rect 41300 43372 41310 43428
rect 42354 43372 42364 43428
rect 42420 43372 47628 43428
rect 47684 43372 47694 43428
rect 28028 43316 28084 43372
rect 19618 43260 19628 43316
rect 19684 43260 19852 43316
rect 19908 43260 19918 43316
rect 21746 43260 21756 43316
rect 21812 43260 22876 43316
rect 22932 43260 22942 43316
rect 24322 43260 24332 43316
rect 24388 43260 26908 43316
rect 26964 43260 26974 43316
rect 28018 43260 28028 43316
rect 28084 43260 28094 43316
rect 33618 43260 33628 43316
rect 33684 43260 35588 43316
rect 37202 43260 37212 43316
rect 37268 43260 44716 43316
rect 44772 43260 44782 43316
rect 35532 43204 35588 43260
rect 22754 43148 22764 43204
rect 22820 43148 23324 43204
rect 23380 43148 23390 43204
rect 35532 43148 37100 43204
rect 37156 43148 37436 43204
rect 37492 43148 37502 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 49200 43092 50000 43120
rect 40114 43036 40124 43092
rect 40180 43036 50000 43092
rect 49200 43008 50000 43036
rect 36194 42924 36204 42980
rect 36260 42924 44044 42980
rect 44100 42924 44110 42980
rect 17378 42812 17388 42868
rect 17444 42812 19516 42868
rect 19572 42812 19582 42868
rect 27906 42812 27916 42868
rect 27972 42812 31276 42868
rect 31332 42812 31342 42868
rect 41906 42812 41916 42868
rect 41972 42812 43708 42868
rect 43764 42812 43774 42868
rect 20066 42700 20076 42756
rect 20132 42700 20412 42756
rect 20468 42700 20478 42756
rect 23650 42700 23660 42756
rect 23716 42700 25116 42756
rect 25172 42700 28700 42756
rect 28756 42700 28766 42756
rect 32834 42700 32844 42756
rect 32900 42700 33852 42756
rect 33908 42700 33918 42756
rect 42466 42700 42476 42756
rect 42532 42700 43484 42756
rect 43540 42700 44828 42756
rect 44884 42700 44894 42756
rect 27570 42588 27580 42644
rect 27636 42588 29148 42644
rect 29204 42588 29214 42644
rect 33506 42588 33516 42644
rect 33572 42588 37772 42644
rect 37828 42588 37838 42644
rect 39218 42588 39228 42644
rect 39284 42588 42252 42644
rect 42308 42588 42318 42644
rect 40114 42476 40124 42532
rect 40180 42476 43148 42532
rect 43204 42476 43214 42532
rect 0 42420 800 42448
rect 49200 42420 50000 42448
rect 0 42364 1932 42420
rect 1988 42364 1998 42420
rect 44034 42364 44044 42420
rect 44100 42364 50000 42420
rect 0 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 49200 42336 50000 42364
rect 11890 42252 11900 42308
rect 11956 42252 14924 42308
rect 14980 42252 15260 42308
rect 15316 42252 15326 42308
rect 33282 42252 33292 42308
rect 33348 42252 35420 42308
rect 35476 42252 35486 42308
rect 41122 42252 41132 42308
rect 41188 42252 43932 42308
rect 43988 42252 43998 42308
rect 10546 42140 10556 42196
rect 10612 42140 11452 42196
rect 11508 42140 13804 42196
rect 13860 42140 14700 42196
rect 14756 42140 14766 42196
rect 19506 42140 19516 42196
rect 19572 42140 20188 42196
rect 20244 42140 20254 42196
rect 21634 42140 21644 42196
rect 21700 42140 23212 42196
rect 23268 42140 23884 42196
rect 23940 42140 23950 42196
rect 34738 42140 34748 42196
rect 34804 42140 35980 42196
rect 36036 42140 36046 42196
rect 38658 42140 38668 42196
rect 38724 42140 39228 42196
rect 39284 42140 39294 42196
rect 6748 42028 8204 42084
rect 8260 42028 8988 42084
rect 9044 42028 9054 42084
rect 11106 42028 11116 42084
rect 11172 42028 15484 42084
rect 15540 42028 15550 42084
rect 19618 42028 19628 42084
rect 19684 42028 19964 42084
rect 20020 42028 20030 42084
rect 20290 42028 20300 42084
rect 20356 42028 22428 42084
rect 22484 42028 22494 42084
rect 33730 42028 33740 42084
rect 33796 42028 34524 42084
rect 34580 42028 34590 42084
rect 38994 42028 39004 42084
rect 39060 42028 40796 42084
rect 40852 42028 41804 42084
rect 41860 42028 41870 42084
rect 6748 41972 6804 42028
rect 21420 41972 21476 42028
rect 6178 41916 6188 41972
rect 6244 41916 6804 41972
rect 13570 41916 13580 41972
rect 13636 41916 15372 41972
rect 15428 41916 15438 41972
rect 19618 41916 19628 41972
rect 19684 41916 20636 41972
rect 20692 41916 20702 41972
rect 21410 41916 21420 41972
rect 21476 41916 21486 41972
rect 25442 41916 25452 41972
rect 25508 41916 26796 41972
rect 26852 41916 26862 41972
rect 30818 41916 30828 41972
rect 30884 41916 37772 41972
rect 37828 41916 37838 41972
rect 39778 41916 39788 41972
rect 39844 41916 41020 41972
rect 41076 41916 41086 41972
rect 41346 41916 41356 41972
rect 41412 41916 41916 41972
rect 41972 41916 41982 41972
rect 16258 41804 16268 41860
rect 16324 41804 30940 41860
rect 30996 41804 31006 41860
rect 31938 41804 31948 41860
rect 32004 41804 33180 41860
rect 33236 41804 33516 41860
rect 33572 41804 33582 41860
rect 36530 41804 36540 41860
rect 36596 41804 37100 41860
rect 37156 41804 37166 41860
rect 37538 41804 37548 41860
rect 37604 41804 39116 41860
rect 39172 41804 39182 41860
rect 40338 41804 40348 41860
rect 40404 41804 42924 41860
rect 42980 41804 42990 41860
rect 0 41748 800 41776
rect 49200 41748 50000 41776
rect 0 41692 2044 41748
rect 2100 41692 2110 41748
rect 4918 41692 4956 41748
rect 5012 41692 5022 41748
rect 5282 41692 5292 41748
rect 5348 41692 6300 41748
rect 6356 41692 6366 41748
rect 17378 41692 17388 41748
rect 17444 41692 22204 41748
rect 22260 41692 22270 41748
rect 34290 41692 34300 41748
rect 34356 41692 38108 41748
rect 38164 41692 38174 41748
rect 39666 41692 39676 41748
rect 39732 41692 42364 41748
rect 42420 41692 42430 41748
rect 44930 41692 44940 41748
rect 44996 41692 50000 41748
rect 0 41664 800 41692
rect 49200 41664 50000 41692
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 39442 41468 39452 41524
rect 39508 41468 43708 41524
rect 43764 41468 43774 41524
rect 21858 41356 21868 41412
rect 21924 41356 23212 41412
rect 23268 41356 23278 41412
rect 25554 41356 25564 41412
rect 25620 41356 26796 41412
rect 26852 41356 26862 41412
rect 45266 41356 45276 41412
rect 45332 41356 48188 41412
rect 48244 41356 48254 41412
rect 18946 41244 18956 41300
rect 19012 41244 19628 41300
rect 19684 41244 19694 41300
rect 22306 41132 22316 41188
rect 22372 41132 25004 41188
rect 25060 41132 25452 41188
rect 25508 41132 25788 41188
rect 25844 41132 25854 41188
rect 30818 41132 30828 41188
rect 30884 41132 31836 41188
rect 31892 41132 31902 41188
rect 34626 41132 34636 41188
rect 34692 41132 35532 41188
rect 35588 41132 35598 41188
rect 36418 41132 36428 41188
rect 36484 41132 38780 41188
rect 38836 41132 38846 41188
rect 45042 41132 45052 41188
rect 45108 41132 45892 41188
rect 45836 41076 45892 41132
rect 49200 41076 50000 41104
rect 23538 41020 23548 41076
rect 23604 41020 24556 41076
rect 24612 41020 25228 41076
rect 25284 41020 25294 41076
rect 27346 41020 27356 41076
rect 27412 41020 28252 41076
rect 28308 41020 28318 41076
rect 41122 41020 41132 41076
rect 41188 41020 45612 41076
rect 45668 41020 45678 41076
rect 45836 41020 50000 41076
rect 49200 40992 50000 41020
rect 1698 40908 1708 40964
rect 1764 40908 5068 40964
rect 5124 40908 5134 40964
rect 23426 40908 23436 40964
rect 23492 40908 23884 40964
rect 23940 40908 23950 40964
rect 24210 40908 24220 40964
rect 24276 40908 26572 40964
rect 26628 40908 26638 40964
rect 27682 40908 27692 40964
rect 27748 40908 29820 40964
rect 29876 40908 29886 40964
rect 30930 40908 30940 40964
rect 30996 40908 35084 40964
rect 35140 40908 35150 40964
rect 34066 40796 34076 40852
rect 34132 40796 41692 40852
rect 41748 40796 41758 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 4274 40684 4284 40740
rect 4340 40684 10108 40740
rect 10164 40684 10668 40740
rect 10724 40684 10734 40740
rect 5730 40572 5740 40628
rect 5796 40572 7196 40628
rect 7252 40572 8540 40628
rect 8596 40572 8606 40628
rect 8978 40572 8988 40628
rect 9044 40572 10220 40628
rect 10276 40572 10286 40628
rect 16370 40572 16380 40628
rect 16436 40572 17388 40628
rect 17444 40572 17454 40628
rect 22978 40572 22988 40628
rect 23044 40572 25340 40628
rect 25396 40572 25406 40628
rect 35074 40572 35084 40628
rect 35140 40572 35644 40628
rect 35700 40572 35710 40628
rect 40674 40572 40684 40628
rect 40740 40572 41244 40628
rect 41300 40572 41310 40628
rect 42130 40572 42140 40628
rect 42196 40572 43036 40628
rect 43092 40572 45948 40628
rect 46004 40572 46014 40628
rect 4274 40460 4284 40516
rect 4340 40460 5068 40516
rect 5124 40460 6076 40516
rect 6132 40460 6142 40516
rect 6850 40460 6860 40516
rect 6916 40460 11228 40516
rect 11284 40460 11294 40516
rect 41458 40460 41468 40516
rect 41524 40460 47404 40516
rect 47460 40460 47470 40516
rect 0 40404 800 40432
rect 49200 40404 50000 40432
rect 0 40348 1932 40404
rect 1988 40348 1998 40404
rect 5170 40348 5180 40404
rect 5236 40348 6188 40404
rect 6244 40348 6254 40404
rect 9874 40348 9884 40404
rect 9940 40348 11004 40404
rect 11060 40348 11070 40404
rect 14802 40348 14812 40404
rect 14868 40348 16044 40404
rect 16100 40348 16110 40404
rect 20402 40348 20412 40404
rect 20468 40348 23660 40404
rect 23716 40348 23726 40404
rect 24210 40348 24220 40404
rect 24276 40348 25564 40404
rect 25620 40348 25630 40404
rect 30268 40348 30604 40404
rect 30660 40348 30670 40404
rect 32498 40348 32508 40404
rect 32564 40348 35420 40404
rect 35476 40348 35486 40404
rect 35634 40348 35644 40404
rect 35700 40348 36540 40404
rect 36596 40348 36606 40404
rect 37426 40348 37436 40404
rect 37492 40348 40236 40404
rect 40292 40348 40302 40404
rect 41206 40348 41244 40404
rect 41300 40348 41310 40404
rect 45938 40348 45948 40404
rect 46004 40348 47292 40404
rect 47348 40348 47358 40404
rect 47842 40348 47852 40404
rect 47908 40348 50000 40404
rect 0 40320 800 40348
rect 30268 40292 30324 40348
rect 49200 40320 50000 40348
rect 17714 40236 17724 40292
rect 17780 40236 18732 40292
rect 18788 40236 18798 40292
rect 22306 40236 22316 40292
rect 22372 40236 23772 40292
rect 23828 40236 23838 40292
rect 27010 40236 27020 40292
rect 27076 40236 28700 40292
rect 28756 40236 28766 40292
rect 29250 40236 29260 40292
rect 29316 40236 30324 40292
rect 35746 40236 35756 40292
rect 35812 40236 36204 40292
rect 36260 40236 36988 40292
rect 37044 40236 37054 40292
rect 42130 40236 42140 40292
rect 42196 40236 42476 40292
rect 42532 40236 43036 40292
rect 43092 40236 43102 40292
rect 38612 40124 39676 40180
rect 39732 40124 39742 40180
rect 40562 40124 40572 40180
rect 40628 40124 40908 40180
rect 40964 40124 40974 40180
rect 11218 40012 11228 40068
rect 11284 40012 11676 40068
rect 11732 40012 13580 40068
rect 13636 40012 13646 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 33394 39900 33404 39956
rect 33460 39900 33740 39956
rect 33796 39900 33806 39956
rect 38612 39844 38668 40124
rect 40674 40012 40684 40068
rect 40740 40012 41804 40068
rect 41860 40012 41870 40068
rect 4386 39788 4396 39844
rect 4452 39788 4956 39844
rect 5012 39788 5022 39844
rect 26002 39788 26012 39844
rect 26068 39788 26572 39844
rect 26628 39788 26638 39844
rect 34850 39788 34860 39844
rect 34916 39788 37772 39844
rect 37828 39788 38668 39844
rect 40002 39788 40012 39844
rect 40068 39788 42812 39844
rect 42868 39788 42878 39844
rect 0 39732 800 39760
rect 49200 39732 50000 39760
rect 0 39676 1932 39732
rect 1988 39676 1998 39732
rect 13570 39676 13580 39732
rect 13636 39676 18396 39732
rect 18452 39676 18462 39732
rect 26338 39676 26348 39732
rect 26404 39676 26908 39732
rect 26964 39676 27692 39732
rect 27748 39676 27758 39732
rect 34402 39676 34412 39732
rect 34468 39676 43708 39732
rect 47954 39676 47964 39732
rect 48020 39676 50000 39732
rect 0 39648 800 39676
rect 43652 39620 43708 39676
rect 49200 39648 50000 39676
rect 10546 39564 10556 39620
rect 10612 39564 11676 39620
rect 11732 39564 11742 39620
rect 18050 39564 18060 39620
rect 18116 39564 18452 39620
rect 19170 39564 19180 39620
rect 19236 39564 24220 39620
rect 24276 39564 24332 39620
rect 24388 39564 24398 39620
rect 43652 39564 45164 39620
rect 45220 39564 45230 39620
rect 18396 39508 18452 39564
rect 2482 39452 2492 39508
rect 2548 39452 5292 39508
rect 5348 39452 5358 39508
rect 12898 39452 12908 39508
rect 12964 39452 13916 39508
rect 13972 39452 13982 39508
rect 15092 39452 18172 39508
rect 18228 39452 18238 39508
rect 18396 39452 19628 39508
rect 19684 39452 19694 39508
rect 15092 39396 15148 39452
rect 4050 39340 4060 39396
rect 4116 39340 10108 39396
rect 10164 39340 11004 39396
rect 11060 39340 11070 39396
rect 11442 39340 11452 39396
rect 11508 39340 13804 39396
rect 13860 39340 15148 39396
rect 15922 39340 15932 39396
rect 15988 39340 18060 39396
rect 18116 39340 18126 39396
rect 23874 39340 23884 39396
rect 23940 39340 27020 39396
rect 27076 39340 27086 39396
rect 33394 39340 33404 39396
rect 33460 39340 34636 39396
rect 34692 39340 37324 39396
rect 37380 39340 42476 39396
rect 42532 39340 42542 39396
rect 35634 39228 35644 39284
rect 35700 39228 39340 39284
rect 39396 39228 40908 39284
rect 40964 39228 40974 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 32386 39116 32396 39172
rect 32452 39116 33516 39172
rect 33572 39116 33582 39172
rect 37212 39116 38108 39172
rect 38164 39116 38174 39172
rect 42466 39116 42476 39172
rect 42532 39116 44268 39172
rect 44324 39116 47180 39172
rect 47236 39116 47246 39172
rect 37212 39060 37268 39116
rect 49200 39060 50000 39088
rect 2370 39004 2380 39060
rect 2436 39004 3164 39060
rect 3220 39004 3230 39060
rect 3714 39004 3724 39060
rect 3780 39004 4676 39060
rect 31938 39004 31948 39060
rect 32004 39004 32014 39060
rect 32498 39004 32508 39060
rect 32564 39004 34188 39060
rect 34244 39004 34254 39060
rect 36642 39004 36652 39060
rect 36708 39004 37212 39060
rect 37268 39004 37278 39060
rect 37762 39004 37772 39060
rect 37828 39004 38444 39060
rect 38500 39004 38510 39060
rect 38658 39004 38668 39060
rect 38724 39004 40572 39060
rect 40628 39004 40638 39060
rect 40898 39004 40908 39060
rect 40964 39004 41916 39060
rect 41972 39004 41982 39060
rect 45042 39004 45052 39060
rect 45108 39004 50000 39060
rect 4620 38948 4676 39004
rect 2594 38892 2604 38948
rect 2660 38892 3612 38948
rect 3668 38892 4284 38948
rect 4340 38892 4350 38948
rect 4610 38892 4620 38948
rect 4676 38892 5404 38948
rect 5460 38892 7756 38948
rect 7812 38892 7822 38948
rect 8194 38892 8204 38948
rect 8260 38892 9548 38948
rect 9604 38892 9614 38948
rect 31948 38836 32004 39004
rect 40908 38948 40964 39004
rect 49200 38976 50000 39004
rect 33170 38892 33180 38948
rect 33236 38892 33852 38948
rect 33908 38892 33918 38948
rect 37986 38892 37996 38948
rect 38052 38892 40964 38948
rect 41122 38892 41132 38948
rect 41188 38892 42812 38948
rect 42868 38892 42878 38948
rect 44594 38892 44604 38948
rect 44660 38892 47516 38948
rect 47572 38892 47582 38948
rect 2706 38780 2716 38836
rect 2772 38780 4396 38836
rect 4452 38780 4462 38836
rect 4834 38780 4844 38836
rect 4900 38780 6412 38836
rect 6468 38780 7980 38836
rect 8036 38780 8046 38836
rect 8306 38780 8316 38836
rect 8372 38780 11116 38836
rect 11172 38780 11452 38836
rect 11508 38780 11518 38836
rect 20290 38780 20300 38836
rect 20356 38780 24668 38836
rect 24724 38780 24734 38836
rect 31948 38780 36820 38836
rect 36978 38780 36988 38836
rect 37044 38780 38332 38836
rect 38388 38780 38398 38836
rect 38612 38780 39732 38836
rect 39890 38780 39900 38836
rect 39956 38780 41020 38836
rect 41076 38780 41086 38836
rect 45826 38780 45836 38836
rect 45892 38780 47068 38836
rect 47124 38780 47134 38836
rect 4844 38724 4900 38780
rect 36764 38724 36820 38780
rect 38612 38724 38668 38780
rect 3938 38668 3948 38724
rect 4004 38668 4900 38724
rect 7420 38668 7868 38724
rect 7924 38668 7934 38724
rect 9202 38668 9212 38724
rect 9268 38668 11340 38724
rect 11396 38668 11676 38724
rect 11732 38668 12460 38724
rect 12516 38668 12526 38724
rect 30258 38668 30268 38724
rect 30324 38668 33068 38724
rect 33124 38668 33134 38724
rect 36764 38668 38668 38724
rect 39676 38724 39732 38780
rect 39676 38668 40348 38724
rect 40404 38668 41356 38724
rect 41412 38668 42476 38724
rect 42532 38668 42542 38724
rect 44930 38668 44940 38724
rect 44996 38668 45388 38724
rect 45444 38668 46508 38724
rect 46564 38668 46574 38724
rect 7420 38612 7476 38668
rect 7410 38556 7420 38612
rect 7476 38556 7486 38612
rect 8978 38556 8988 38612
rect 9044 38556 9660 38612
rect 9716 38556 9726 38612
rect 23986 38556 23996 38612
rect 24052 38556 24444 38612
rect 24500 38556 25004 38612
rect 25060 38556 25070 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 49200 38388 50000 38416
rect 24322 38332 24332 38388
rect 24388 38332 24444 38388
rect 24500 38332 24510 38388
rect 47618 38332 47628 38388
rect 47684 38332 50000 38388
rect 49200 38304 50000 38332
rect 23538 38220 23548 38276
rect 23604 38220 24220 38276
rect 24276 38220 24286 38276
rect 43586 38220 43596 38276
rect 43652 38220 44492 38276
rect 44548 38220 44558 38276
rect 4610 38108 4620 38164
rect 4676 38108 5180 38164
rect 5236 38108 5740 38164
rect 5796 38108 5806 38164
rect 6738 38108 6748 38164
rect 6804 38108 10556 38164
rect 10612 38108 12012 38164
rect 12068 38108 12078 38164
rect 27794 38108 27804 38164
rect 27860 38108 28364 38164
rect 28420 38108 29036 38164
rect 29092 38108 29102 38164
rect 36082 38108 36092 38164
rect 36148 38108 36988 38164
rect 37044 38108 37054 38164
rect 39666 38108 39676 38164
rect 39732 38108 40908 38164
rect 40964 38108 40974 38164
rect 4946 37996 4956 38052
rect 5012 37996 6412 38052
rect 6468 37996 6478 38052
rect 6626 37996 6636 38052
rect 6692 37996 8652 38052
rect 8708 37996 8718 38052
rect 25554 37996 25564 38052
rect 25620 37996 29260 38052
rect 29316 37996 29326 38052
rect 31714 37996 31724 38052
rect 31780 37996 41692 38052
rect 41748 37996 41758 38052
rect 43362 37996 43372 38052
rect 43428 37996 44828 38052
rect 44884 37996 44894 38052
rect 7634 37884 7644 37940
rect 7700 37884 9660 37940
rect 9716 37884 10220 37940
rect 10276 37884 10286 37940
rect 33954 37884 33964 37940
rect 34020 37884 34860 37940
rect 34916 37884 34926 37940
rect 41346 37884 41356 37940
rect 41412 37884 42700 37940
rect 42756 37884 42766 37940
rect 5506 37772 5516 37828
rect 5572 37772 6636 37828
rect 6692 37772 6702 37828
rect 22306 37772 22316 37828
rect 22372 37772 23436 37828
rect 23492 37772 23772 37828
rect 23828 37772 23838 37828
rect 39778 37772 39788 37828
rect 39844 37772 48412 37828
rect 48468 37772 48478 37828
rect 49200 37716 50000 37744
rect 47730 37660 47740 37716
rect 47796 37660 50000 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 49200 37632 50000 37660
rect 13122 37436 13132 37492
rect 13188 37436 14308 37492
rect 18162 37436 18172 37492
rect 18228 37436 18844 37492
rect 18900 37436 21196 37492
rect 21252 37436 21262 37492
rect 25330 37436 25340 37492
rect 25396 37436 26012 37492
rect 26068 37436 26078 37492
rect 35420 37436 36092 37492
rect 36148 37436 36158 37492
rect 14252 37380 14308 37436
rect 35420 37380 35476 37436
rect 11778 37324 11788 37380
rect 11844 37324 13020 37380
rect 13076 37324 13086 37380
rect 14242 37324 14252 37380
rect 14308 37324 15708 37380
rect 15764 37324 15774 37380
rect 17826 37324 17836 37380
rect 17892 37324 18956 37380
rect 19012 37324 19022 37380
rect 25890 37324 25900 37380
rect 25956 37324 27692 37380
rect 27748 37324 27758 37380
rect 35410 37324 35420 37380
rect 35476 37324 35486 37380
rect 40562 37324 40572 37380
rect 40628 37324 41692 37380
rect 41748 37324 45276 37380
rect 45332 37324 46844 37380
rect 46900 37324 46910 37380
rect 4274 37212 4284 37268
rect 4340 37212 9660 37268
rect 9716 37212 10108 37268
rect 10164 37212 10780 37268
rect 10836 37212 10846 37268
rect 13346 37212 13356 37268
rect 13412 37212 14140 37268
rect 14196 37212 14206 37268
rect 17836 37156 17892 37324
rect 24434 37212 24444 37268
rect 24500 37212 25676 37268
rect 25732 37212 25742 37268
rect 35970 37212 35980 37268
rect 36036 37212 36652 37268
rect 36708 37212 36718 37268
rect 38882 37212 38892 37268
rect 38948 37212 41020 37268
rect 41076 37212 41086 37268
rect 14018 37100 14028 37156
rect 14084 37100 14588 37156
rect 14644 37100 14924 37156
rect 14980 37100 17892 37156
rect 35074 37100 35084 37156
rect 35140 37100 35644 37156
rect 35700 37100 35710 37156
rect 42242 37100 42252 37156
rect 42308 37100 43820 37156
rect 43876 37100 43886 37156
rect 45938 37100 45948 37156
rect 46004 37100 47180 37156
rect 47236 37100 47246 37156
rect 0 37044 800 37072
rect 49200 37044 50000 37072
rect 0 36988 1932 37044
rect 1988 36988 1998 37044
rect 3154 36988 3164 37044
rect 3220 36988 4284 37044
rect 4340 36988 4350 37044
rect 14466 36988 14476 37044
rect 14532 36988 15820 37044
rect 15876 36988 15886 37044
rect 40674 36988 40684 37044
rect 40740 36988 44604 37044
rect 44660 36988 44670 37044
rect 46610 36988 46620 37044
rect 46676 36988 50000 37044
rect 0 36960 800 36988
rect 49200 36960 50000 36988
rect 37314 36876 37324 36932
rect 37380 36876 38108 36932
rect 38164 36876 38174 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19954 36764 19964 36820
rect 20020 36764 24332 36820
rect 24388 36764 24398 36820
rect 7074 36652 7084 36708
rect 7140 36652 8988 36708
rect 9044 36652 10892 36708
rect 10948 36652 12908 36708
rect 12964 36652 12974 36708
rect 14130 36652 14140 36708
rect 14196 36652 19740 36708
rect 19796 36652 20748 36708
rect 20804 36652 20814 36708
rect 1922 36540 1932 36596
rect 1988 36540 1998 36596
rect 13682 36540 13692 36596
rect 13748 36540 15148 36596
rect 15922 36540 15932 36596
rect 15988 36540 18172 36596
rect 18228 36540 18238 36596
rect 24210 36540 24220 36596
rect 24276 36540 24332 36596
rect 24388 36540 24398 36596
rect 0 36372 800 36400
rect 1932 36372 1988 36540
rect 15092 36484 15148 36540
rect 4834 36428 4844 36484
rect 4900 36428 5628 36484
rect 5684 36428 5694 36484
rect 5842 36428 5852 36484
rect 5908 36428 7868 36484
rect 7924 36428 10444 36484
rect 10500 36428 10510 36484
rect 14802 36428 14812 36484
rect 14868 36428 14878 36484
rect 15092 36428 15372 36484
rect 15428 36428 15438 36484
rect 23202 36428 23212 36484
rect 23268 36428 23380 36484
rect 24098 36428 24108 36484
rect 24164 36428 24668 36484
rect 24724 36428 24734 36484
rect 28578 36428 28588 36484
rect 28644 36428 29260 36484
rect 29316 36428 29820 36484
rect 29876 36428 29886 36484
rect 43810 36428 43820 36484
rect 43876 36428 44940 36484
rect 44996 36428 45006 36484
rect 14812 36372 14868 36428
rect 23324 36372 23380 36428
rect 49200 36372 50000 36400
rect 0 36316 1988 36372
rect 7522 36316 7532 36372
rect 7588 36316 8428 36372
rect 8484 36316 8494 36372
rect 14812 36316 16828 36372
rect 16884 36316 16894 36372
rect 23324 36316 24892 36372
rect 24948 36316 24958 36372
rect 38322 36316 38332 36372
rect 38388 36316 39228 36372
rect 39284 36316 39294 36372
rect 39564 36316 43596 36372
rect 43652 36316 43662 36372
rect 45266 36316 45276 36372
rect 45332 36316 45724 36372
rect 45780 36316 45790 36372
rect 47394 36316 47404 36372
rect 47460 36316 50000 36372
rect 0 36288 800 36316
rect 39564 36260 39620 36316
rect 49200 36288 50000 36316
rect 4274 36204 4284 36260
rect 4340 36204 6300 36260
rect 6356 36204 6366 36260
rect 8642 36204 8652 36260
rect 8708 36204 11564 36260
rect 11620 36204 11630 36260
rect 23772 36204 24220 36260
rect 24276 36204 24286 36260
rect 37090 36204 37100 36260
rect 37156 36204 39564 36260
rect 39620 36204 39630 36260
rect 41234 36204 41244 36260
rect 41300 36204 41804 36260
rect 41860 36204 41870 36260
rect 43362 36204 43372 36260
rect 43428 36204 44940 36260
rect 44996 36204 45006 36260
rect 22754 36092 22764 36148
rect 22820 36092 23268 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 23212 36036 23268 36092
rect 23772 36036 23828 36204
rect 42802 36092 42812 36148
rect 42868 36092 43484 36148
rect 43540 36092 44716 36148
rect 44772 36092 44782 36148
rect 23202 35980 23212 36036
rect 23268 35980 23278 36036
rect 23426 35980 23436 36036
rect 23492 35980 23772 36036
rect 23828 35980 23838 36036
rect 38658 35980 38668 36036
rect 38724 35980 40124 36036
rect 40180 35980 40190 36036
rect 44034 35980 44044 36036
rect 44100 35980 47292 36036
rect 47348 35980 48188 36036
rect 48244 35980 48254 36036
rect 11106 35868 11116 35924
rect 11172 35868 11452 35924
rect 11508 35868 11788 35924
rect 11844 35868 11854 35924
rect 22642 35868 22652 35924
rect 22708 35868 25788 35924
rect 25844 35868 25854 35924
rect 27010 35868 27020 35924
rect 27076 35868 29148 35924
rect 29204 35868 30156 35924
rect 30212 35868 30222 35924
rect 36306 35868 36316 35924
rect 36372 35868 36876 35924
rect 36932 35868 36942 35924
rect 41906 35868 41916 35924
rect 41972 35868 42924 35924
rect 42980 35868 42990 35924
rect 43250 35868 43260 35924
rect 43316 35868 45500 35924
rect 45556 35868 45566 35924
rect 21186 35756 21196 35812
rect 21252 35756 22540 35812
rect 22596 35756 22606 35812
rect 23986 35756 23996 35812
rect 24052 35756 24892 35812
rect 24948 35756 26124 35812
rect 26180 35756 26190 35812
rect 36614 35756 36652 35812
rect 36708 35756 36718 35812
rect 45154 35756 45164 35812
rect 45220 35756 46060 35812
rect 46116 35756 46126 35812
rect 47180 35756 48300 35812
rect 48356 35756 48366 35812
rect 47180 35700 47236 35756
rect 49200 35700 50000 35728
rect 2482 35644 2492 35700
rect 2548 35644 5516 35700
rect 5572 35644 5582 35700
rect 8306 35644 8316 35700
rect 8372 35644 11340 35700
rect 11396 35644 13244 35700
rect 13300 35644 13310 35700
rect 24294 35644 24332 35700
rect 24388 35644 24398 35700
rect 24658 35644 24668 35700
rect 24724 35644 25564 35700
rect 25620 35644 25630 35700
rect 34738 35644 34748 35700
rect 34804 35644 38668 35700
rect 42130 35644 42140 35700
rect 42196 35644 42588 35700
rect 42644 35644 44268 35700
rect 44324 35644 44940 35700
rect 44996 35644 47180 35700
rect 47236 35644 47246 35700
rect 47730 35644 47740 35700
rect 47796 35644 50000 35700
rect 38612 35588 38668 35644
rect 49200 35616 50000 35644
rect 1810 35532 1820 35588
rect 1876 35532 3388 35588
rect 13570 35532 13580 35588
rect 13636 35532 17500 35588
rect 17556 35532 17566 35588
rect 32498 35532 32508 35588
rect 32564 35532 33404 35588
rect 33460 35532 33470 35588
rect 34962 35532 34972 35588
rect 35028 35532 36764 35588
rect 36820 35532 36830 35588
rect 38612 35532 42364 35588
rect 42420 35532 45612 35588
rect 45668 35532 45678 35588
rect 3332 35364 3388 35532
rect 3948 35420 5068 35476
rect 5124 35420 5964 35476
rect 6020 35420 6030 35476
rect 6178 35420 6188 35476
rect 6244 35420 15148 35476
rect 19842 35420 19852 35476
rect 19908 35420 21644 35476
rect 21700 35420 21710 35476
rect 21970 35420 21980 35476
rect 22036 35420 23324 35476
rect 23380 35420 23390 35476
rect 3948 35364 4004 35420
rect 15092 35364 15148 35420
rect 3332 35308 3948 35364
rect 4004 35308 4014 35364
rect 7746 35308 7756 35364
rect 7812 35308 8540 35364
rect 8596 35308 8606 35364
rect 15092 35308 16156 35364
rect 16212 35308 17948 35364
rect 18004 35308 18014 35364
rect 20514 35308 20524 35364
rect 20580 35308 26236 35364
rect 26292 35308 26302 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 15026 35196 15036 35252
rect 15092 35196 15484 35252
rect 15540 35196 15550 35252
rect 18722 35196 18732 35252
rect 18788 35196 25900 35252
rect 25956 35196 26684 35252
rect 26740 35196 27468 35252
rect 27524 35196 30492 35252
rect 30548 35196 30558 35252
rect 37762 35196 37772 35252
rect 37828 35196 40180 35252
rect 41794 35196 41804 35252
rect 41860 35196 44716 35252
rect 44772 35196 44782 35252
rect 9762 35084 9772 35140
rect 9828 35084 10556 35140
rect 10612 35084 10622 35140
rect 10770 35084 10780 35140
rect 10836 35084 13468 35140
rect 13524 35084 13534 35140
rect 10556 35028 10612 35084
rect 40124 35028 40180 35196
rect 44594 35084 44604 35140
rect 44660 35084 45276 35140
rect 45332 35084 47628 35140
rect 47684 35084 47694 35140
rect 49200 35028 50000 35056
rect 10556 34972 10892 35028
rect 10948 34972 10958 35028
rect 40114 34972 40124 35028
rect 40180 34972 41468 35028
rect 41524 34972 42700 35028
rect 42756 34972 45388 35028
rect 45444 34972 45454 35028
rect 47954 34972 47964 35028
rect 48020 34972 50000 35028
rect 49200 34944 50000 34972
rect 10322 34860 10332 34916
rect 10388 34860 11788 34916
rect 11844 34860 13020 34916
rect 13076 34860 13086 34916
rect 16034 34860 16044 34916
rect 16100 34860 18508 34916
rect 18564 34860 20300 34916
rect 20356 34860 20366 34916
rect 35634 34860 35644 34916
rect 35700 34860 43148 34916
rect 43204 34860 43932 34916
rect 43988 34860 43998 34916
rect 3332 34748 15260 34804
rect 15316 34748 15326 34804
rect 23090 34748 23100 34804
rect 23156 34748 23884 34804
rect 23940 34748 23950 34804
rect 31714 34748 31724 34804
rect 31780 34748 32620 34804
rect 32676 34748 33236 34804
rect 34402 34748 34412 34804
rect 34468 34748 34860 34804
rect 34916 34748 37044 34804
rect 44258 34748 44268 34804
rect 44324 34748 45836 34804
rect 45892 34748 45902 34804
rect 3332 34468 3388 34748
rect 33180 34692 33236 34748
rect 36988 34692 37044 34748
rect 12226 34636 12236 34692
rect 12292 34636 12908 34692
rect 12964 34636 13692 34692
rect 13748 34636 15148 34692
rect 15204 34636 15214 34692
rect 18274 34636 18284 34692
rect 18340 34636 18844 34692
rect 18900 34636 20748 34692
rect 20804 34636 28476 34692
rect 28532 34636 28542 34692
rect 33170 34636 33180 34692
rect 33236 34636 33246 34692
rect 36978 34636 36988 34692
rect 37044 34636 37772 34692
rect 37828 34636 38220 34692
rect 38276 34636 38286 34692
rect 6850 34524 6860 34580
rect 6916 34524 7420 34580
rect 7476 34524 8428 34580
rect 8484 34524 11004 34580
rect 11060 34524 11070 34580
rect 22418 34524 22428 34580
rect 22484 34524 24220 34580
rect 24276 34524 24286 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 2034 34412 2044 34468
rect 2100 34412 3388 34468
rect 34738 34412 34748 34468
rect 34804 34412 38668 34468
rect 0 34356 800 34384
rect 38612 34356 38668 34412
rect 49200 34356 50000 34384
rect 0 34300 1708 34356
rect 1764 34300 2492 34356
rect 2548 34300 2558 34356
rect 10098 34300 10108 34356
rect 10164 34300 10780 34356
rect 10836 34300 10846 34356
rect 36642 34300 36652 34356
rect 36708 34300 37436 34356
rect 37492 34300 37502 34356
rect 38612 34300 44716 34356
rect 44772 34300 44782 34356
rect 46946 34300 46956 34356
rect 47012 34300 50000 34356
rect 0 34272 800 34300
rect 37436 34244 37492 34300
rect 49200 34272 50000 34300
rect 10546 34188 10556 34244
rect 10612 34188 12572 34244
rect 12628 34188 12638 34244
rect 37436 34188 39116 34244
rect 39172 34188 39788 34244
rect 39844 34188 39854 34244
rect 10658 34076 10668 34132
rect 10724 34076 13692 34132
rect 13748 34076 13758 34132
rect 32050 34076 32060 34132
rect 32116 34076 33628 34132
rect 33684 34076 33694 34132
rect 44818 34076 44828 34132
rect 44884 34076 46620 34132
rect 46676 34076 46686 34132
rect 18050 33740 18060 33796
rect 18116 33740 18508 33796
rect 18564 33740 18574 33796
rect 36866 33740 36876 33796
rect 36932 33740 44156 33796
rect 44212 33740 44940 33796
rect 44996 33740 45006 33796
rect 0 33684 800 33712
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 0 33628 1932 33684
rect 1988 33628 1998 33684
rect 9202 33628 9212 33684
rect 9268 33628 9996 33684
rect 10052 33628 10062 33684
rect 19394 33628 19404 33684
rect 19460 33628 20188 33684
rect 20244 33628 20412 33684
rect 20468 33628 20478 33684
rect 36754 33628 36764 33684
rect 36820 33628 37772 33684
rect 37828 33628 37838 33684
rect 0 33600 800 33628
rect 36764 33572 36820 33628
rect 8726 33516 8764 33572
rect 8820 33516 8830 33572
rect 33618 33516 33628 33572
rect 33684 33516 36820 33572
rect 43922 33516 43932 33572
rect 43988 33516 45388 33572
rect 45444 33516 45454 33572
rect 7410 33404 7420 33460
rect 7476 33404 8428 33460
rect 8484 33404 8494 33460
rect 11218 33404 11228 33460
rect 11284 33404 12348 33460
rect 12404 33404 12414 33460
rect 14690 33404 14700 33460
rect 14756 33404 17164 33460
rect 17220 33404 17230 33460
rect 20066 33404 20076 33460
rect 20132 33404 20412 33460
rect 20468 33404 20478 33460
rect 25106 33404 25116 33460
rect 25172 33404 25900 33460
rect 25956 33404 25966 33460
rect 26450 33404 26460 33460
rect 26516 33404 27916 33460
rect 27972 33404 27982 33460
rect 33282 33404 33292 33460
rect 33348 33404 34748 33460
rect 34804 33404 34814 33460
rect 45490 33404 45500 33460
rect 45556 33404 45724 33460
rect 45780 33404 48188 33460
rect 48244 33404 48254 33460
rect 1810 33292 1820 33348
rect 1876 33292 3948 33348
rect 4004 33292 4014 33348
rect 5730 33292 5740 33348
rect 5796 33292 8764 33348
rect 8820 33292 8830 33348
rect 9202 33292 9212 33348
rect 9268 33292 9884 33348
rect 9940 33292 9950 33348
rect 13682 33292 13692 33348
rect 13748 33292 14812 33348
rect 14868 33292 14878 33348
rect 23538 33292 23548 33348
rect 23604 33292 24108 33348
rect 24164 33292 24174 33348
rect 33170 33292 33180 33348
rect 33236 33292 34972 33348
rect 35028 33292 36316 33348
rect 36372 33292 36382 33348
rect 37986 33292 37996 33348
rect 38052 33292 39228 33348
rect 39284 33292 39294 33348
rect 43474 33292 43484 33348
rect 43540 33292 44268 33348
rect 44324 33292 44828 33348
rect 44884 33292 44894 33348
rect 7186 33180 7196 33236
rect 7252 33180 8204 33236
rect 8260 33180 10444 33236
rect 10500 33180 10510 33236
rect 12898 33180 12908 33236
rect 12964 33180 13916 33236
rect 13972 33180 13982 33236
rect 19618 33180 19628 33236
rect 19684 33180 22204 33236
rect 22260 33180 25004 33236
rect 25060 33180 25070 33236
rect 30818 33180 30828 33236
rect 30884 33180 31164 33236
rect 31220 33180 34300 33236
rect 34356 33180 34366 33236
rect 35522 33180 35532 33236
rect 35588 33180 36204 33236
rect 36260 33180 36270 33236
rect 39106 33180 39116 33236
rect 39172 33180 41580 33236
rect 41636 33180 45388 33236
rect 45444 33180 45454 33236
rect 6290 33068 6300 33124
rect 6356 33068 7308 33124
rect 7364 33068 9996 33124
rect 10052 33068 10062 33124
rect 10882 33068 10892 33124
rect 10948 33068 18284 33124
rect 18340 33068 18350 33124
rect 22978 33068 22988 33124
rect 23044 33068 23772 33124
rect 23828 33068 25228 33124
rect 25284 33068 25294 33124
rect 26002 33068 26012 33124
rect 26068 33068 26348 33124
rect 26404 33068 26414 33124
rect 30258 33068 30268 33124
rect 30324 33068 33628 33124
rect 33684 33068 33694 33124
rect 35746 33068 35756 33124
rect 35812 33068 36988 33124
rect 37044 33068 37054 33124
rect 38612 33068 47068 33124
rect 47124 33068 47134 33124
rect 4274 32956 4284 33012
rect 4340 32956 12908 33012
rect 12964 32956 14924 33012
rect 14980 32956 15148 33012
rect 23202 32956 23212 33012
rect 23268 32956 23548 33012
rect 23604 32956 23614 33012
rect 31042 32956 31052 33012
rect 31108 32956 31388 33012
rect 31444 32956 32844 33012
rect 32900 32956 34524 33012
rect 34580 32956 34590 33012
rect 2930 32732 2940 32788
rect 2996 32732 4956 32788
rect 5012 32732 5516 32788
rect 5572 32732 5582 32788
rect 8652 32732 8764 32788
rect 8820 32732 8830 32788
rect 9874 32732 9884 32788
rect 9940 32732 11004 32788
rect 11060 32732 11070 32788
rect 4834 32620 4844 32676
rect 4900 32620 5852 32676
rect 5908 32620 5918 32676
rect 8652 32564 8708 32732
rect 9986 32620 9996 32676
rect 10052 32620 10780 32676
rect 10836 32620 10846 32676
rect 15092 32564 15148 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 38612 32900 38668 33068
rect 38882 32956 38892 33012
rect 38948 32956 39900 33012
rect 39956 32956 39966 33012
rect 40898 32956 40908 33012
rect 40964 32956 42140 33012
rect 42196 32956 42924 33012
rect 42980 32956 42990 33012
rect 44258 32956 44268 33012
rect 44324 32956 46844 33012
rect 46900 32956 46910 33012
rect 33506 32844 33516 32900
rect 33572 32844 38668 32900
rect 43586 32844 43596 32900
rect 43652 32844 46172 32900
rect 46228 32844 48188 32900
rect 48244 32844 48254 32900
rect 16034 32732 16044 32788
rect 16100 32732 17612 32788
rect 17668 32732 17678 32788
rect 27122 32732 27132 32788
rect 27188 32732 27804 32788
rect 27860 32732 27870 32788
rect 37202 32732 37212 32788
rect 37268 32732 38220 32788
rect 38276 32732 38892 32788
rect 38948 32732 38958 32788
rect 39218 32732 39228 32788
rect 39284 32732 41804 32788
rect 41860 32732 43260 32788
rect 43316 32732 45948 32788
rect 46004 32732 46014 32788
rect 15586 32620 15596 32676
rect 15652 32620 16604 32676
rect 16660 32620 17388 32676
rect 17444 32620 17454 32676
rect 19170 32620 19180 32676
rect 19236 32620 19628 32676
rect 19684 32620 19694 32676
rect 29250 32620 29260 32676
rect 29316 32620 31052 32676
rect 31108 32620 31118 32676
rect 38546 32620 38556 32676
rect 38612 32564 38668 32676
rect 40450 32620 40460 32676
rect 40516 32620 42420 32676
rect 42364 32564 42420 32620
rect 4722 32508 4732 32564
rect 4788 32508 5292 32564
rect 5348 32508 8652 32564
rect 8708 32508 8718 32564
rect 15092 32508 16492 32564
rect 16548 32508 17612 32564
rect 17668 32508 17678 32564
rect 17938 32508 17948 32564
rect 18004 32508 18620 32564
rect 18676 32508 18686 32564
rect 28466 32508 28476 32564
rect 28532 32508 29820 32564
rect 29876 32508 29886 32564
rect 31602 32508 31612 32564
rect 31668 32508 33292 32564
rect 33348 32508 33358 32564
rect 33506 32508 33516 32564
rect 33572 32508 35532 32564
rect 35588 32508 35598 32564
rect 38612 32508 40908 32564
rect 40964 32508 40974 32564
rect 41346 32508 41356 32564
rect 41412 32508 41916 32564
rect 41972 32508 41982 32564
rect 42354 32508 42364 32564
rect 42420 32508 43708 32564
rect 43764 32508 43774 32564
rect 45154 32508 45164 32564
rect 45220 32508 46508 32564
rect 46564 32508 46574 32564
rect 17612 32452 17668 32508
rect 3938 32396 3948 32452
rect 4004 32396 4620 32452
rect 4676 32396 4686 32452
rect 11106 32396 11116 32452
rect 11172 32396 13692 32452
rect 13748 32396 13758 32452
rect 17612 32396 18172 32452
rect 18228 32396 18238 32452
rect 22978 32396 22988 32452
rect 23044 32396 23054 32452
rect 24322 32396 24332 32452
rect 24388 32396 25452 32452
rect 25508 32396 25518 32452
rect 42914 32396 42924 32452
rect 42980 32396 45500 32452
rect 45556 32396 46396 32452
rect 46452 32396 46462 32452
rect 22988 32340 23044 32396
rect 3602 32284 3612 32340
rect 3668 32284 5628 32340
rect 5684 32284 6524 32340
rect 6580 32284 6590 32340
rect 9090 32284 9100 32340
rect 9156 32284 11228 32340
rect 11284 32284 11294 32340
rect 19730 32284 19740 32340
rect 19796 32284 21420 32340
rect 21476 32284 23044 32340
rect 24658 32284 24668 32340
rect 24724 32284 25340 32340
rect 25396 32284 25406 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 24770 32060 24780 32116
rect 24836 32060 25788 32116
rect 25844 32060 25854 32116
rect 4834 31948 4844 32004
rect 4900 31948 5796 32004
rect 18610 31948 18620 32004
rect 18676 31948 21420 32004
rect 21476 31948 21486 32004
rect 28802 31948 28812 32004
rect 28868 31948 30604 32004
rect 30660 31948 31276 32004
rect 31332 31948 31342 32004
rect 31490 31948 31500 32004
rect 31556 31948 35868 32004
rect 35924 31948 35934 32004
rect 39890 31948 39900 32004
rect 39956 31948 41020 32004
rect 41076 31948 41086 32004
rect 5740 31892 5796 31948
rect 3602 31836 3612 31892
rect 3668 31836 4396 31892
rect 4452 31836 5180 31892
rect 5236 31836 5246 31892
rect 5730 31836 5740 31892
rect 5796 31836 7756 31892
rect 7812 31836 8428 31892
rect 8484 31836 11116 31892
rect 11172 31836 11182 31892
rect 13682 31836 13692 31892
rect 13748 31836 14028 31892
rect 14084 31836 14094 31892
rect 22194 31836 22204 31892
rect 22260 31836 23324 31892
rect 23380 31836 23884 31892
rect 23940 31836 23950 31892
rect 29474 31836 29484 31892
rect 29540 31836 30156 31892
rect 30212 31836 30222 31892
rect 33954 31836 33964 31892
rect 34020 31836 34030 31892
rect 35522 31836 35532 31892
rect 35588 31836 37100 31892
rect 37156 31836 44156 31892
rect 44212 31836 45164 31892
rect 45220 31836 45230 31892
rect 33964 31780 34020 31836
rect 10546 31724 10556 31780
rect 10612 31724 11900 31780
rect 11956 31724 11966 31780
rect 13682 31724 13692 31780
rect 13748 31724 14196 31780
rect 14354 31724 14364 31780
rect 14420 31724 15036 31780
rect 15092 31724 15102 31780
rect 16146 31724 16156 31780
rect 16212 31724 18172 31780
rect 18228 31724 18238 31780
rect 29698 31724 29708 31780
rect 29764 31724 31500 31780
rect 31556 31724 33068 31780
rect 33124 31724 33134 31780
rect 33964 31724 35644 31780
rect 35700 31724 35710 31780
rect 43810 31724 43820 31780
rect 43876 31724 44716 31780
rect 44772 31724 44782 31780
rect 14140 31668 14196 31724
rect 12674 31612 12684 31668
rect 12740 31612 13804 31668
rect 13860 31612 13870 31668
rect 14140 31612 14924 31668
rect 14980 31612 14990 31668
rect 19058 31612 19068 31668
rect 19124 31612 20972 31668
rect 21028 31612 21038 31668
rect 26852 31612 42588 31668
rect 42644 31612 42654 31668
rect 6402 31500 6412 31556
rect 6468 31500 9100 31556
rect 9156 31500 9166 31556
rect 13906 31500 13916 31556
rect 13972 31500 14476 31556
rect 14532 31500 14542 31556
rect 15092 31500 15372 31556
rect 15428 31500 15438 31556
rect 15092 31444 15148 31500
rect 12450 31388 12460 31444
rect 12516 31388 13804 31444
rect 13860 31388 15148 31444
rect 22082 31388 22092 31444
rect 22148 31388 26796 31444
rect 26852 31388 26908 31612
rect 29586 31500 29596 31556
rect 29652 31500 30044 31556
rect 30100 31500 30110 31556
rect 30258 31500 30268 31556
rect 30324 31500 33292 31556
rect 33348 31500 35084 31556
rect 35140 31500 35150 31556
rect 29474 31388 29484 31444
rect 29540 31388 30828 31444
rect 30884 31388 31164 31444
rect 31220 31388 31230 31444
rect 32386 31388 32396 31444
rect 32452 31388 33740 31444
rect 33796 31388 33806 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 13682 31276 13692 31332
rect 13748 31276 13860 31332
rect 15698 31276 15708 31332
rect 15764 31276 16604 31332
rect 16660 31276 16670 31332
rect 21298 31276 21308 31332
rect 21364 31276 21756 31332
rect 21812 31276 21822 31332
rect 29362 31276 29372 31332
rect 29428 31276 29932 31332
rect 29988 31276 30268 31332
rect 30324 31276 30334 31332
rect 8194 31052 8204 31108
rect 8260 31052 8764 31108
rect 8820 31052 12684 31108
rect 12740 31052 12750 31108
rect 13804 30884 13860 31276
rect 14578 31164 14588 31220
rect 14644 31164 15372 31220
rect 15428 31164 15438 31220
rect 21970 31164 21980 31220
rect 22036 31164 23324 31220
rect 23380 31164 24556 31220
rect 24612 31164 24622 31220
rect 29250 31164 29260 31220
rect 29316 31164 30156 31220
rect 30212 31164 32060 31220
rect 32116 31164 32126 31220
rect 44482 31164 44492 31220
rect 44548 31164 47516 31220
rect 47572 31164 47582 31220
rect 15474 31052 15484 31108
rect 15540 31052 15932 31108
rect 15988 31052 18060 31108
rect 18116 31052 18126 31108
rect 20972 31052 35756 31108
rect 35812 31052 35822 31108
rect 45042 31052 45052 31108
rect 45108 31052 47740 31108
rect 47796 31052 47806 31108
rect 20972 30884 21028 31052
rect 22642 30940 22652 30996
rect 22708 30940 23436 30996
rect 23492 30940 23502 30996
rect 29362 30940 29372 30996
rect 29428 30940 30492 30996
rect 30548 30940 30558 30996
rect 13794 30828 13804 30884
rect 13860 30828 13870 30884
rect 14466 30828 14476 30884
rect 14532 30828 21028 30884
rect 26786 30828 26796 30884
rect 26852 30828 30268 30884
rect 30324 30828 30334 30884
rect 30594 30828 30604 30884
rect 30660 30828 31500 30884
rect 31556 30828 31566 30884
rect 33730 30828 33740 30884
rect 33796 30828 36540 30884
rect 36596 30828 37996 30884
rect 38052 30828 38062 30884
rect 2818 30716 2828 30772
rect 2884 30716 5460 30772
rect 6626 30716 6636 30772
rect 6692 30716 16156 30772
rect 16212 30716 16222 30772
rect 36082 30716 36092 30772
rect 36148 30716 37212 30772
rect 37268 30716 37772 30772
rect 37828 30716 37838 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 5404 30548 5460 30716
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 5394 30492 5404 30548
rect 5460 30492 6188 30548
rect 6244 30492 6254 30548
rect 3378 30380 3388 30436
rect 3444 30380 4844 30436
rect 4900 30380 5964 30436
rect 6020 30380 7196 30436
rect 7252 30380 7532 30436
rect 7588 30380 7598 30436
rect 12674 30380 12684 30436
rect 12740 30380 13468 30436
rect 13524 30380 13534 30436
rect 34850 30380 34860 30436
rect 34916 30380 35644 30436
rect 35700 30380 35710 30436
rect 4610 30268 4620 30324
rect 4676 30268 6300 30324
rect 6356 30268 6366 30324
rect 7634 30268 7644 30324
rect 7700 30268 13804 30324
rect 13860 30268 14252 30324
rect 14308 30268 14318 30324
rect 17602 30268 17612 30324
rect 17668 30268 18060 30324
rect 18116 30268 18126 30324
rect 19058 30268 19068 30324
rect 19124 30268 19134 30324
rect 19068 30212 19124 30268
rect 15586 30156 15596 30212
rect 15652 30156 16156 30212
rect 16212 30156 16940 30212
rect 16996 30156 19124 30212
rect 22194 30156 22204 30212
rect 22260 30156 24220 30212
rect 24276 30156 25116 30212
rect 25172 30156 25182 30212
rect 32498 30156 32508 30212
rect 32564 30156 33068 30212
rect 33124 30156 35308 30212
rect 35364 30156 35374 30212
rect 15250 30044 15260 30100
rect 15316 30044 15932 30100
rect 15988 30044 15998 30100
rect 16818 30044 16828 30100
rect 16884 30044 17948 30100
rect 18004 30044 18014 30100
rect 30258 30044 30268 30100
rect 30324 30044 30940 30100
rect 30996 30044 31500 30100
rect 31556 30044 32844 30100
rect 32900 30044 32910 30100
rect 36082 30044 36092 30100
rect 36148 30044 38668 30100
rect 39442 30044 39452 30100
rect 39508 30044 41132 30100
rect 41188 30044 41198 30100
rect 42466 30044 42476 30100
rect 42532 30044 44044 30100
rect 44100 30044 44110 30100
rect 38612 29988 38668 30044
rect 3938 29932 3948 29988
rect 4004 29932 4284 29988
rect 4340 29932 4350 29988
rect 17948 29932 19740 29988
rect 19796 29932 19806 29988
rect 35970 29932 35980 29988
rect 36036 29932 37436 29988
rect 37492 29932 37502 29988
rect 38612 29932 41356 29988
rect 41412 29932 42140 29988
rect 42196 29932 42206 29988
rect 17948 29876 18004 29932
rect 13570 29820 13580 29876
rect 13636 29820 14924 29876
rect 14980 29820 16268 29876
rect 16324 29820 18004 29876
rect 34290 29820 34300 29876
rect 34356 29820 36988 29876
rect 37044 29820 37054 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 31826 29708 31836 29764
rect 31892 29708 32508 29764
rect 32564 29708 37324 29764
rect 37380 29708 37390 29764
rect 16034 29596 16044 29652
rect 16100 29596 17948 29652
rect 18004 29596 19180 29652
rect 19236 29596 19246 29652
rect 23650 29596 23660 29652
rect 23716 29596 26908 29652
rect 26852 29540 26908 29596
rect 16118 29484 16156 29540
rect 16212 29484 16222 29540
rect 16930 29484 16940 29540
rect 16996 29484 17500 29540
rect 17556 29484 17566 29540
rect 26852 29484 35644 29540
rect 35700 29484 35710 29540
rect 35858 29484 35868 29540
rect 35924 29484 36764 29540
rect 36820 29484 37436 29540
rect 37492 29484 37502 29540
rect 8866 29372 8876 29428
rect 8932 29372 10220 29428
rect 10276 29372 10286 29428
rect 10434 29372 10444 29428
rect 10500 29372 11452 29428
rect 11508 29372 12572 29428
rect 12628 29372 18284 29428
rect 18340 29372 18350 29428
rect 36082 29372 36092 29428
rect 36148 29372 38220 29428
rect 38276 29372 38286 29428
rect 42242 29372 42252 29428
rect 42308 29372 42700 29428
rect 42756 29372 43148 29428
rect 43204 29372 43214 29428
rect 2818 29260 2828 29316
rect 2884 29260 3276 29316
rect 3332 29260 8092 29316
rect 8148 29260 8158 29316
rect 9426 29260 9436 29316
rect 9492 29260 10668 29316
rect 10724 29260 11900 29316
rect 11956 29260 11966 29316
rect 14700 29260 19292 29316
rect 19348 29260 20636 29316
rect 20692 29260 21308 29316
rect 21364 29260 21374 29316
rect 29586 29260 29596 29316
rect 29652 29260 31052 29316
rect 31108 29260 33180 29316
rect 33236 29260 33740 29316
rect 33796 29260 33806 29316
rect 44930 29260 44940 29316
rect 44996 29260 46060 29316
rect 46116 29260 46126 29316
rect 14700 29204 14756 29260
rect 14690 29148 14700 29204
rect 14756 29148 14766 29204
rect 15026 29148 15036 29204
rect 15092 29148 15260 29204
rect 15316 29148 15326 29204
rect 16482 29148 16492 29204
rect 16548 29148 17388 29204
rect 17444 29148 17454 29204
rect 19506 29148 19516 29204
rect 19572 29148 21420 29204
rect 21476 29148 32172 29204
rect 32228 29148 32238 29204
rect 41570 29148 41580 29204
rect 41636 29148 42028 29204
rect 42084 29148 42094 29204
rect 6066 29036 6076 29092
rect 6132 29036 6636 29092
rect 6692 29036 6702 29092
rect 18834 29036 18844 29092
rect 18900 29036 19628 29092
rect 19684 29036 19694 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 4834 28924 4844 28980
rect 4900 28924 9660 28980
rect 9716 28924 9726 28980
rect 19170 28924 19180 28980
rect 19236 28924 20748 28980
rect 20804 28924 20814 28980
rect 38322 28924 38332 28980
rect 38388 28924 45724 28980
rect 45780 28924 45790 28980
rect 4844 28868 4900 28924
rect 3042 28812 3052 28868
rect 3108 28812 3724 28868
rect 3780 28812 4900 28868
rect 5730 28812 5740 28868
rect 5796 28812 5964 28868
rect 6020 28812 6030 28868
rect 12338 28812 12348 28868
rect 12404 28812 13580 28868
rect 13636 28812 14588 28868
rect 14644 28812 14654 28868
rect 14914 28812 14924 28868
rect 14980 28812 15148 28868
rect 37426 28812 37436 28868
rect 37492 28812 42700 28868
rect 42756 28812 42766 28868
rect 2930 28700 2940 28756
rect 2996 28700 3948 28756
rect 4004 28700 4396 28756
rect 4452 28700 4462 28756
rect 4722 28700 4732 28756
rect 4788 28700 5852 28756
rect 5908 28700 5918 28756
rect 9762 28700 9772 28756
rect 9828 28700 10220 28756
rect 10276 28700 11732 28756
rect 4162 28588 4172 28644
rect 4228 28588 4508 28644
rect 4564 28588 5740 28644
rect 5796 28588 5806 28644
rect 9650 28588 9660 28644
rect 9716 28588 9996 28644
rect 10052 28588 10062 28644
rect 11676 28532 11732 28700
rect 14588 28644 14644 28812
rect 15092 28756 15148 28812
rect 15092 28700 19460 28756
rect 21522 28700 21532 28756
rect 21588 28700 22092 28756
rect 22148 28700 23660 28756
rect 23716 28700 24892 28756
rect 24948 28700 24958 28756
rect 37650 28700 37660 28756
rect 37716 28700 42140 28756
rect 42196 28700 42206 28756
rect 19404 28644 19460 28700
rect 14588 28588 15372 28644
rect 15428 28588 15438 28644
rect 19394 28588 19404 28644
rect 19460 28588 19470 28644
rect 25330 28588 25340 28644
rect 25396 28588 26796 28644
rect 26852 28588 29148 28644
rect 29204 28588 29214 28644
rect 37986 28588 37996 28644
rect 38052 28588 38892 28644
rect 38948 28588 38958 28644
rect 42578 28588 42588 28644
rect 42644 28588 43260 28644
rect 43316 28588 44044 28644
rect 44100 28588 44828 28644
rect 44884 28588 44894 28644
rect 45266 28588 45276 28644
rect 45332 28588 48188 28644
rect 48244 28588 48254 28644
rect 11676 28476 14364 28532
rect 14420 28476 15260 28532
rect 15316 28476 15326 28532
rect 7634 28364 7644 28420
rect 7700 28364 20188 28420
rect 20244 28364 20254 28420
rect 28914 28364 28924 28420
rect 28980 28364 37100 28420
rect 37156 28364 37166 28420
rect 9874 28252 9884 28308
rect 9940 28252 10780 28308
rect 10836 28252 10846 28308
rect 16034 28252 16044 28308
rect 16100 28252 16604 28308
rect 16660 28252 19068 28308
rect 19124 28252 19134 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 6626 28140 6636 28196
rect 6692 28140 11676 28196
rect 11732 28140 11742 28196
rect 11890 28140 11900 28196
rect 11956 28140 16380 28196
rect 16436 28140 17276 28196
rect 17332 28140 17342 28196
rect 18284 28140 18620 28196
rect 18676 28140 18686 28196
rect 18284 28084 18340 28140
rect 14018 28028 14028 28084
rect 14084 28028 15596 28084
rect 15652 28028 18340 28084
rect 18498 28028 18508 28084
rect 18564 28028 19516 28084
rect 19572 28028 20076 28084
rect 20132 28028 20142 28084
rect 22978 28028 22988 28084
rect 23044 28028 40348 28084
rect 40404 28028 43484 28084
rect 43540 28028 44268 28084
rect 44324 28028 44334 28084
rect 9762 27916 9772 27972
rect 9828 27916 15820 27972
rect 15876 27916 16156 27972
rect 16212 27916 16268 27972
rect 16324 27916 16334 27972
rect 20850 27916 20860 27972
rect 20916 27916 22204 27972
rect 22260 27916 22270 27972
rect 32386 27916 32396 27972
rect 32452 27916 33852 27972
rect 33908 27916 33918 27972
rect 34076 27916 37436 27972
rect 37492 27916 40012 27972
rect 40068 27916 40078 27972
rect 1810 27804 1820 27860
rect 1876 27804 5852 27860
rect 5908 27804 7756 27860
rect 7812 27804 7822 27860
rect 9874 27804 9884 27860
rect 9940 27804 10444 27860
rect 10500 27804 10510 27860
rect 11218 27804 11228 27860
rect 11284 27804 17948 27860
rect 18004 27804 18014 27860
rect 21634 27804 21644 27860
rect 21700 27804 22876 27860
rect 22932 27804 22942 27860
rect 29250 27804 29260 27860
rect 29316 27804 33068 27860
rect 33124 27804 33134 27860
rect 34076 27748 34132 27916
rect 36866 27804 36876 27860
rect 36932 27804 38444 27860
rect 38500 27804 38510 27860
rect 41458 27804 41468 27860
rect 41524 27804 42588 27860
rect 42644 27804 42654 27860
rect 5618 27692 5628 27748
rect 5684 27692 8764 27748
rect 8820 27692 9548 27748
rect 9604 27692 9614 27748
rect 11778 27692 11788 27748
rect 11844 27692 12460 27748
rect 12516 27692 12526 27748
rect 15922 27692 15932 27748
rect 15988 27692 16940 27748
rect 16996 27692 17006 27748
rect 28130 27692 28140 27748
rect 28196 27692 28924 27748
rect 28980 27692 28990 27748
rect 29138 27692 29148 27748
rect 29204 27692 30380 27748
rect 30436 27692 30828 27748
rect 30884 27692 30894 27748
rect 31378 27692 31388 27748
rect 31444 27692 32172 27748
rect 32228 27692 34132 27748
rect 44370 27692 44380 27748
rect 44436 27692 46060 27748
rect 46116 27692 46126 27748
rect 2370 27580 2380 27636
rect 2436 27580 9268 27636
rect 10770 27580 10780 27636
rect 10836 27580 11676 27636
rect 11732 27580 11742 27636
rect 15362 27580 15372 27636
rect 15428 27580 15820 27636
rect 15876 27580 15886 27636
rect 30482 27580 30492 27636
rect 30548 27580 31164 27636
rect 31220 27580 32508 27636
rect 32564 27580 33180 27636
rect 33236 27580 33246 27636
rect 36866 27580 36876 27636
rect 36932 27580 38668 27636
rect 38724 27580 38734 27636
rect 9212 27524 9268 27580
rect 9212 27468 24332 27524
rect 24388 27468 25340 27524
rect 25396 27468 25788 27524
rect 25844 27468 25854 27524
rect 30146 27468 30156 27524
rect 30212 27468 31388 27524
rect 31444 27468 31454 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 26002 27244 26012 27300
rect 26068 27244 28588 27300
rect 28644 27244 28654 27300
rect 42802 27244 42812 27300
rect 42868 27244 43596 27300
rect 43652 27244 44268 27300
rect 44324 27244 48188 27300
rect 48244 27244 48254 27300
rect 9090 27132 9100 27188
rect 9156 27132 11004 27188
rect 11060 27132 11070 27188
rect 20178 27132 20188 27188
rect 20244 27132 24668 27188
rect 24724 27132 24734 27188
rect 42242 27132 42252 27188
rect 42308 27132 44828 27188
rect 44884 27132 44894 27188
rect 7746 27020 7756 27076
rect 7812 27020 10108 27076
rect 10164 27020 11116 27076
rect 11172 27020 11182 27076
rect 13570 27020 13580 27076
rect 13636 27020 14812 27076
rect 14868 27020 14878 27076
rect 17602 27020 17612 27076
rect 17668 27020 18396 27076
rect 18452 27020 18462 27076
rect 20626 27020 20636 27076
rect 20692 27020 21868 27076
rect 21924 27020 22540 27076
rect 22596 27020 22606 27076
rect 23426 27020 23436 27076
rect 23492 27020 29596 27076
rect 29652 27020 30044 27076
rect 30100 27020 31612 27076
rect 31668 27020 31678 27076
rect 32834 27020 32844 27076
rect 32900 27020 33852 27076
rect 33908 27020 35868 27076
rect 35924 27020 40908 27076
rect 40964 27020 40974 27076
rect 43362 27020 43372 27076
rect 43428 27020 43932 27076
rect 43988 27020 43998 27076
rect 44258 27020 44268 27076
rect 44324 27020 44940 27076
rect 44996 27020 46060 27076
rect 46116 27020 48076 27076
rect 48132 27020 48142 27076
rect 23436 26964 23492 27020
rect 9202 26908 9212 26964
rect 9268 26908 11788 26964
rect 11844 26908 11854 26964
rect 12898 26908 12908 26964
rect 12964 26908 13692 26964
rect 13748 26908 15372 26964
rect 15428 26908 18284 26964
rect 18340 26908 18350 26964
rect 20402 26908 20412 26964
rect 20468 26908 23492 26964
rect 41122 26908 41132 26964
rect 41188 26908 41468 26964
rect 41524 26908 42364 26964
rect 42420 26908 42430 26964
rect 17826 26796 17836 26852
rect 17892 26796 18396 26852
rect 18452 26796 18620 26852
rect 18676 26796 19180 26852
rect 19236 26796 19246 26852
rect 35970 26796 35980 26852
rect 36036 26796 36428 26852
rect 36484 26796 39116 26852
rect 39172 26796 39182 26852
rect 13654 26684 13692 26740
rect 13748 26684 13758 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 26562 26460 26572 26516
rect 26628 26460 35420 26516
rect 35476 26460 35486 26516
rect 32498 26348 32508 26404
rect 32564 26348 33628 26404
rect 33684 26348 36988 26404
rect 37044 26348 37054 26404
rect 49200 26292 50000 26320
rect 4834 26236 4844 26292
rect 4900 26236 6076 26292
rect 6132 26236 7084 26292
rect 7140 26236 7150 26292
rect 16706 26236 16716 26292
rect 16772 26236 17724 26292
rect 17780 26236 17790 26292
rect 32162 26236 32172 26292
rect 32228 26236 32620 26292
rect 32676 26236 33516 26292
rect 33572 26236 33582 26292
rect 38994 26236 39004 26292
rect 39060 26236 40572 26292
rect 40628 26236 40638 26292
rect 41346 26236 41356 26292
rect 41412 26236 42588 26292
rect 42644 26236 42654 26292
rect 47842 26236 47852 26292
rect 47908 26236 50000 26292
rect 49200 26208 50000 26236
rect 8082 26124 8092 26180
rect 8148 26124 8652 26180
rect 8708 26124 9548 26180
rect 9604 26124 9614 26180
rect 12114 26124 12124 26180
rect 12180 26124 20020 26180
rect 40226 26124 40236 26180
rect 40292 26124 42476 26180
rect 42532 26124 43932 26180
rect 43988 26124 43998 26180
rect 19964 26068 20020 26124
rect 2482 26012 2492 26068
rect 2548 26012 4732 26068
rect 4788 26012 4798 26068
rect 15362 26012 15372 26068
rect 15428 26012 17500 26068
rect 17556 26012 19180 26068
rect 19236 26012 19246 26068
rect 19954 26012 19964 26068
rect 20020 26012 20524 26068
rect 20580 26012 20590 26068
rect 11330 25900 11340 25956
rect 11396 25900 11900 25956
rect 11956 25900 13804 25956
rect 13860 25900 13870 25956
rect 15250 25900 15260 25956
rect 15316 25900 16156 25956
rect 16212 25900 17388 25956
rect 17444 25900 17454 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 13906 25788 13916 25844
rect 13972 25788 13982 25844
rect 15922 25788 15932 25844
rect 15988 25788 16828 25844
rect 16884 25788 16894 25844
rect 13916 25620 13972 25788
rect 13458 25564 13468 25620
rect 13524 25564 13972 25620
rect 31892 25676 32620 25732
rect 32676 25676 32686 25732
rect 31892 25508 31948 25676
rect 42578 25564 42588 25620
rect 42644 25564 45612 25620
rect 45668 25564 45678 25620
rect 5730 25452 5740 25508
rect 5796 25452 6636 25508
rect 6692 25452 8988 25508
rect 9044 25452 11564 25508
rect 11620 25452 11630 25508
rect 14914 25452 14924 25508
rect 14980 25452 15708 25508
rect 15764 25452 17612 25508
rect 17668 25452 17678 25508
rect 31490 25452 31500 25508
rect 31556 25452 31948 25508
rect 36418 25452 36428 25508
rect 36484 25452 37324 25508
rect 37380 25452 38108 25508
rect 38164 25452 38174 25508
rect 39218 25452 39228 25508
rect 39284 25452 41132 25508
rect 41188 25452 41198 25508
rect 41570 25452 41580 25508
rect 41636 25452 42476 25508
rect 42532 25452 42542 25508
rect 44034 25452 44044 25508
rect 44100 25452 45052 25508
rect 45108 25452 45724 25508
rect 45780 25452 45790 25508
rect 38546 25340 38556 25396
rect 38612 25340 38892 25396
rect 38948 25340 38958 25396
rect 46946 25340 46956 25396
rect 47012 25340 47516 25396
rect 47572 25340 47582 25396
rect 4610 25228 4620 25284
rect 4676 25228 6300 25284
rect 6356 25228 6366 25284
rect 14130 25228 14140 25284
rect 14196 25228 14700 25284
rect 14756 25228 14766 25284
rect 15138 25228 15148 25284
rect 15204 25228 16156 25284
rect 16212 25228 16222 25284
rect 38210 25228 38220 25284
rect 38276 25228 39900 25284
rect 39956 25228 39966 25284
rect 45714 25228 45724 25284
rect 45780 25228 47852 25284
rect 47908 25228 47918 25284
rect 10546 25116 10556 25172
rect 10612 25116 11228 25172
rect 11284 25116 11294 25172
rect 28578 25116 28588 25172
rect 28644 25116 38668 25172
rect 38724 25116 41412 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 41356 24948 41412 25116
rect 49200 24948 50000 24976
rect 29922 24892 29932 24948
rect 29988 24892 30940 24948
rect 30996 24892 31006 24948
rect 38098 24892 38108 24948
rect 38164 24892 38780 24948
rect 38836 24892 38846 24948
rect 39778 24892 39788 24948
rect 39844 24892 41020 24948
rect 41076 24892 41086 24948
rect 41346 24892 41356 24948
rect 41412 24892 41422 24948
rect 41794 24892 41804 24948
rect 41860 24892 42028 24948
rect 42084 24892 42094 24948
rect 45826 24892 45836 24948
rect 45892 24892 47180 24948
rect 47236 24892 47246 24948
rect 48178 24892 48188 24948
rect 48244 24892 50000 24948
rect 48188 24836 48244 24892
rect 49200 24864 50000 24892
rect 20178 24780 20188 24836
rect 20244 24780 20860 24836
rect 20916 24780 20926 24836
rect 25330 24780 25340 24836
rect 25396 24780 31052 24836
rect 31108 24780 33740 24836
rect 33796 24780 34636 24836
rect 34692 24780 34702 24836
rect 37762 24780 37772 24836
rect 37828 24780 39340 24836
rect 39396 24780 39406 24836
rect 45602 24780 45612 24836
rect 45668 24780 48244 24836
rect 4274 24668 4284 24724
rect 4340 24668 24668 24724
rect 24724 24668 25228 24724
rect 25284 24668 25294 24724
rect 37538 24668 37548 24724
rect 37604 24668 38444 24724
rect 38500 24668 38510 24724
rect 46834 24668 46844 24724
rect 46900 24668 47292 24724
rect 47348 24668 47358 24724
rect 22866 24556 22876 24612
rect 22932 24556 23548 24612
rect 23604 24556 23614 24612
rect 42018 24556 42028 24612
rect 42084 24556 42700 24612
rect 42756 24556 42766 24612
rect 46722 24556 46732 24612
rect 46788 24556 47628 24612
rect 47684 24556 48188 24612
rect 48244 24556 48254 24612
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 4162 24444 4172 24500
rect 4228 24444 12572 24500
rect 12628 24444 14028 24500
rect 14084 24444 14364 24500
rect 14420 24444 14430 24500
rect 31266 24444 31276 24500
rect 31332 24444 31836 24500
rect 31892 24444 31902 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 1988 24276
rect 0 24192 800 24220
rect 44818 24108 44828 24164
rect 44884 24108 47068 24164
rect 47124 24108 47134 24164
rect 23538 23996 23548 24052
rect 23604 23996 25732 24052
rect 25676 23940 25732 23996
rect 2034 23884 2044 23940
rect 2100 23884 5068 23940
rect 5124 23884 5134 23940
rect 5842 23884 5852 23940
rect 5908 23884 6972 23940
rect 7028 23884 7038 23940
rect 10322 23884 10332 23940
rect 10388 23884 19852 23940
rect 19908 23884 20412 23940
rect 20468 23884 20478 23940
rect 23090 23884 23100 23940
rect 23156 23884 24220 23940
rect 24276 23884 25452 23940
rect 25508 23884 25518 23940
rect 25666 23884 25676 23940
rect 25732 23884 26684 23940
rect 26740 23884 26750 23940
rect 28578 23884 28588 23940
rect 28644 23884 29708 23940
rect 29764 23884 33516 23940
rect 33572 23884 33582 23940
rect 41570 23884 41580 23940
rect 41636 23884 43596 23940
rect 43652 23884 43662 23940
rect 43810 23884 43820 23940
rect 43876 23884 45276 23940
rect 45332 23884 45342 23940
rect 5730 23772 5740 23828
rect 5796 23772 6748 23828
rect 6804 23772 8316 23828
rect 8372 23772 10556 23828
rect 10612 23772 10622 23828
rect 25778 23772 25788 23828
rect 25844 23772 29148 23828
rect 29204 23772 29214 23828
rect 44930 23772 44940 23828
rect 44996 23772 46172 23828
rect 46228 23772 46238 23828
rect 13570 23660 13580 23716
rect 13636 23660 14924 23716
rect 14980 23660 15596 23716
rect 15652 23660 15662 23716
rect 18386 23660 18396 23716
rect 18452 23660 19292 23716
rect 19348 23660 19628 23716
rect 19684 23660 19694 23716
rect 42242 23660 42252 23716
rect 42308 23660 42476 23716
rect 42532 23660 42542 23716
rect 45266 23660 45276 23716
rect 45332 23660 47068 23716
rect 47124 23660 47134 23716
rect 47506 23660 47516 23716
rect 47572 23660 48020 23716
rect 47964 23604 48020 23660
rect 49200 23604 50000 23632
rect 4610 23548 4620 23604
rect 4676 23548 5292 23604
rect 5348 23548 6412 23604
rect 6468 23548 6478 23604
rect 38546 23548 38556 23604
rect 38612 23548 43764 23604
rect 45490 23548 45500 23604
rect 45556 23548 47628 23604
rect 47684 23548 47694 23604
rect 47964 23548 50000 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 42252 23492 42308 23548
rect 43708 23492 43764 23548
rect 49200 23520 50000 23548
rect 7186 23436 7196 23492
rect 7252 23436 8204 23492
rect 8260 23436 8270 23492
rect 20178 23436 20188 23492
rect 20244 23436 20254 23492
rect 33506 23436 33516 23492
rect 33572 23436 34188 23492
rect 34244 23436 34254 23492
rect 42242 23436 42252 23492
rect 42308 23436 42318 23492
rect 42578 23436 42588 23492
rect 42644 23436 43484 23492
rect 43540 23436 43550 23492
rect 43708 23436 44604 23492
rect 44660 23436 44670 23492
rect 20188 23380 20244 23436
rect 3332 23324 3612 23380
rect 3668 23324 18060 23380
rect 18116 23324 18126 23380
rect 18834 23324 18844 23380
rect 18900 23324 19292 23380
rect 19348 23324 20244 23380
rect 38322 23324 38332 23380
rect 38388 23324 39228 23380
rect 39284 23324 39294 23380
rect 3332 23156 3388 23324
rect 9314 23212 9324 23268
rect 9380 23212 12012 23268
rect 12068 23212 12078 23268
rect 17602 23212 17612 23268
rect 17668 23212 20524 23268
rect 20580 23212 22092 23268
rect 22148 23212 22158 23268
rect 38770 23212 38780 23268
rect 38836 23212 39340 23268
rect 39396 23212 39406 23268
rect 2930 23100 2940 23156
rect 2996 23100 3388 23156
rect 30258 23100 30268 23156
rect 30324 23100 31388 23156
rect 31444 23100 31454 23156
rect 34962 23100 34972 23156
rect 35028 23100 38108 23156
rect 38164 23100 39676 23156
rect 39732 23100 39742 23156
rect 42914 23100 42924 23156
rect 42980 23100 43148 23156
rect 43204 23100 43596 23156
rect 43652 23100 43662 23156
rect 3154 22988 3164 23044
rect 3220 22988 4620 23044
rect 4676 22988 4686 23044
rect 10546 22988 10556 23044
rect 10612 22988 13580 23044
rect 13636 22988 13916 23044
rect 13972 22988 13982 23044
rect 15810 22988 15820 23044
rect 15876 22988 16828 23044
rect 16884 22988 16894 23044
rect 41234 22988 41244 23044
rect 41300 22988 42252 23044
rect 42308 22988 42318 23044
rect 44482 22988 44492 23044
rect 44548 22988 45276 23044
rect 45332 22988 45342 23044
rect 45826 22988 45836 23044
rect 45892 22988 48188 23044
rect 48244 22988 48254 23044
rect 0 22932 800 22960
rect 49200 22932 50000 22960
rect 0 22876 1708 22932
rect 1764 22876 2492 22932
rect 2548 22876 2558 22932
rect 6514 22876 6524 22932
rect 6580 22876 8540 22932
rect 8596 22876 8606 22932
rect 31892 22876 33068 22932
rect 33124 22876 33134 22932
rect 38882 22876 38892 22932
rect 38948 22876 41692 22932
rect 41748 22876 41758 22932
rect 47954 22876 47964 22932
rect 48020 22876 50000 22932
rect 0 22848 800 22876
rect 31892 22820 31948 22876
rect 49200 22848 50000 22876
rect 31602 22764 31612 22820
rect 31668 22764 31948 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 33842 22540 33852 22596
rect 33908 22540 35308 22596
rect 35364 22540 36876 22596
rect 36932 22540 36942 22596
rect 10210 22428 10220 22484
rect 10276 22428 11116 22484
rect 11172 22428 11182 22484
rect 12338 22428 12348 22484
rect 12404 22428 13580 22484
rect 13636 22428 14476 22484
rect 14532 22428 14542 22484
rect 21186 22428 21196 22484
rect 21252 22428 22652 22484
rect 22708 22428 22718 22484
rect 23090 22428 23100 22484
rect 23156 22428 24332 22484
rect 24388 22428 25452 22484
rect 25508 22428 25518 22484
rect 30482 22428 30492 22484
rect 30548 22428 31388 22484
rect 31444 22428 33404 22484
rect 33460 22428 33470 22484
rect 34402 22428 34412 22484
rect 34468 22428 35084 22484
rect 35140 22428 35150 22484
rect 34738 22316 34748 22372
rect 34804 22316 35644 22372
rect 35700 22316 35710 22372
rect 0 22260 800 22288
rect 0 22204 1708 22260
rect 1764 22204 2380 22260
rect 2436 22204 2446 22260
rect 4610 22204 4620 22260
rect 4676 22204 6188 22260
rect 6244 22204 7196 22260
rect 7252 22204 7262 22260
rect 8418 22204 8428 22260
rect 8484 22204 8876 22260
rect 8932 22204 8942 22260
rect 12898 22204 12908 22260
rect 12964 22204 13916 22260
rect 13972 22204 13982 22260
rect 33170 22204 33180 22260
rect 33236 22204 33628 22260
rect 33684 22204 37772 22260
rect 37828 22204 38444 22260
rect 38500 22204 38510 22260
rect 42998 22204 43036 22260
rect 43092 22204 43102 22260
rect 0 22176 800 22204
rect 5058 22092 5068 22148
rect 5124 22092 8204 22148
rect 8260 22092 10556 22148
rect 10612 22092 10622 22148
rect 22866 22092 22876 22148
rect 22932 22092 23660 22148
rect 23716 22092 23726 22148
rect 34178 22092 34188 22148
rect 34244 22092 35196 22148
rect 35252 22092 35262 22148
rect 39666 22092 39676 22148
rect 39732 22092 43596 22148
rect 43652 22092 44156 22148
rect 44212 22092 44222 22148
rect 23090 21980 23100 22036
rect 23156 21980 23548 22036
rect 23604 21980 23614 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 2482 21868 2492 21924
rect 2548 21868 6748 21924
rect 6804 21868 6814 21924
rect 22082 21868 22092 21924
rect 22148 21868 23996 21924
rect 24052 21868 25004 21924
rect 25060 21868 25070 21924
rect 10322 21756 10332 21812
rect 10388 21756 11676 21812
rect 11732 21756 13132 21812
rect 13188 21756 13198 21812
rect 31938 21756 31948 21812
rect 32004 21756 33964 21812
rect 34020 21756 34030 21812
rect 40338 21756 40348 21812
rect 40404 21756 41020 21812
rect 41076 21756 41086 21812
rect 2034 21644 2044 21700
rect 2100 21644 12572 21700
rect 12628 21644 12638 21700
rect 30594 21644 30604 21700
rect 30660 21644 31836 21700
rect 0 21588 800 21616
rect 31892 21588 31948 21700
rect 0 21532 1988 21588
rect 4274 21532 4284 21588
rect 4340 21532 8428 21588
rect 8484 21532 10668 21588
rect 10724 21532 10892 21588
rect 10948 21532 10958 21588
rect 11106 21532 11116 21588
rect 11172 21532 11676 21588
rect 11732 21532 12684 21588
rect 12740 21532 12750 21588
rect 31892 21532 32060 21588
rect 32116 21532 32126 21588
rect 38434 21532 38444 21588
rect 38500 21532 39228 21588
rect 39284 21532 39294 21588
rect 0 21504 800 21532
rect 1932 21476 1988 21532
rect 1922 21420 1932 21476
rect 1988 21420 1998 21476
rect 3332 21420 6356 21476
rect 8978 21420 8988 21476
rect 9044 21420 11788 21476
rect 11844 21420 11854 21476
rect 13122 21420 13132 21476
rect 13188 21420 13580 21476
rect 13636 21420 13804 21476
rect 13860 21420 13870 21476
rect 31154 21420 31164 21476
rect 31220 21420 31836 21476
rect 31892 21420 31902 21476
rect 40786 21420 40796 21476
rect 40852 21420 41916 21476
rect 41972 21420 41982 21476
rect 3332 21028 3388 21420
rect 4946 21308 4956 21364
rect 5012 21308 5404 21364
rect 5460 21308 5470 21364
rect 6300 21252 6356 21420
rect 6514 21308 6524 21364
rect 6580 21308 14812 21364
rect 14868 21308 15372 21364
rect 15428 21308 15438 21364
rect 19282 21308 19292 21364
rect 19348 21308 21308 21364
rect 21364 21308 21374 21364
rect 6300 21196 12124 21252
rect 12180 21196 12190 21252
rect 14364 21196 18508 21252
rect 18564 21196 18844 21252
rect 18900 21196 18910 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 14364 21028 14420 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 38210 21084 38220 21140
rect 38276 21084 38780 21140
rect 38836 21084 39004 21140
rect 39060 21084 39070 21140
rect 41794 21084 41804 21140
rect 41860 21084 43596 21140
rect 43652 21084 43662 21140
rect 2034 20972 2044 21028
rect 2100 20972 3388 21028
rect 4610 20972 4620 21028
rect 4676 20972 6748 21028
rect 6804 20972 14364 21028
rect 14420 20972 14430 21028
rect 21298 20972 21308 21028
rect 21364 20972 21980 21028
rect 22036 20972 22046 21028
rect 37660 20972 39564 21028
rect 39620 20972 39630 21028
rect 37660 20916 37716 20972
rect 49200 20916 50000 20944
rect 3266 20860 3276 20916
rect 3332 20860 5516 20916
rect 5572 20860 7980 20916
rect 8036 20860 8046 20916
rect 14690 20860 14700 20916
rect 14756 20860 15708 20916
rect 15764 20860 18340 20916
rect 19058 20860 19068 20916
rect 19124 20860 19740 20916
rect 19796 20860 19806 20916
rect 36866 20860 36876 20916
rect 36932 20860 37660 20916
rect 37716 20860 37726 20916
rect 37986 20860 37996 20916
rect 38052 20860 39116 20916
rect 39172 20860 39182 20916
rect 46050 20860 46060 20916
rect 46116 20860 48188 20916
rect 48244 20860 48254 20916
rect 48412 20860 50000 20916
rect 18284 20804 18340 20860
rect 48412 20804 48468 20860
rect 49200 20832 50000 20860
rect 15138 20748 15148 20804
rect 15204 20748 16156 20804
rect 16212 20748 16222 20804
rect 16594 20748 16604 20804
rect 16660 20748 17836 20804
rect 17892 20748 17902 20804
rect 18274 20748 18284 20804
rect 18340 20748 19628 20804
rect 19684 20748 19694 20804
rect 23090 20748 23100 20804
rect 23156 20748 23436 20804
rect 23492 20748 23502 20804
rect 29922 20748 29932 20804
rect 29988 20748 30380 20804
rect 30436 20748 31164 20804
rect 31220 20748 31230 20804
rect 37090 20748 37100 20804
rect 37156 20748 38668 20804
rect 38724 20748 38734 20804
rect 40674 20748 40684 20804
rect 40740 20748 42812 20804
rect 42868 20748 42878 20804
rect 44146 20748 44156 20804
rect 44212 20748 45276 20804
rect 45332 20748 45342 20804
rect 48066 20748 48076 20804
rect 48132 20748 48468 20804
rect 6290 20636 6300 20692
rect 6356 20636 8540 20692
rect 8596 20636 8606 20692
rect 12898 20636 12908 20692
rect 12964 20636 14252 20692
rect 14308 20636 14318 20692
rect 15362 20636 15372 20692
rect 15428 20636 16716 20692
rect 16772 20636 16782 20692
rect 17836 20580 17892 20748
rect 19506 20636 19516 20692
rect 19572 20636 21420 20692
rect 21476 20636 22092 20692
rect 22148 20636 22988 20692
rect 23044 20636 23054 20692
rect 31602 20636 31612 20692
rect 31668 20636 36988 20692
rect 37044 20636 37054 20692
rect 38098 20636 38108 20692
rect 38164 20636 39788 20692
rect 39844 20636 39854 20692
rect 17836 20524 19964 20580
rect 20020 20524 20412 20580
rect 20468 20524 20478 20580
rect 23874 20524 23884 20580
rect 23940 20524 23996 20580
rect 24052 20524 24062 20580
rect 38612 20524 40460 20580
rect 40516 20524 40526 20580
rect 41682 20524 41692 20580
rect 41748 20524 42140 20580
rect 42196 20524 42206 20580
rect 43222 20524 43260 20580
rect 43316 20524 43326 20580
rect 38612 20468 38668 20524
rect 23426 20412 23436 20468
rect 23492 20412 23996 20468
rect 24052 20412 24062 20468
rect 37650 20412 37660 20468
rect 37716 20412 38668 20468
rect 38994 20412 39004 20468
rect 39060 20412 40012 20468
rect 40068 20412 40078 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 22530 20300 22540 20356
rect 22596 20300 22876 20356
rect 22932 20300 23324 20356
rect 23380 20300 24556 20356
rect 24612 20300 24622 20356
rect 38882 20300 38892 20356
rect 38948 20300 39228 20356
rect 39284 20300 39294 20356
rect 49200 20244 50000 20272
rect 30706 20188 30716 20244
rect 30772 20188 30782 20244
rect 45154 20188 45164 20244
rect 45220 20188 45556 20244
rect 47954 20188 47964 20244
rect 48020 20188 50000 20244
rect 3714 20076 3724 20132
rect 3780 20076 4844 20132
rect 4900 20076 5740 20132
rect 5796 20076 6188 20132
rect 6244 20076 6254 20132
rect 6738 20076 6748 20132
rect 6804 20076 7532 20132
rect 7588 20076 7598 20132
rect 8642 20076 8652 20132
rect 8708 20076 9884 20132
rect 9940 20076 9950 20132
rect 17714 20076 17724 20132
rect 17780 20076 20188 20132
rect 20244 20076 20972 20132
rect 21028 20076 21038 20132
rect 25106 20076 25116 20132
rect 25172 20076 25452 20132
rect 25508 20076 25518 20132
rect 28242 20076 28252 20132
rect 28308 20076 29260 20132
rect 29316 20076 29326 20132
rect 30716 20020 30772 20188
rect 45500 20132 45556 20188
rect 49200 20160 50000 20188
rect 45500 20076 46396 20132
rect 46452 20076 46462 20132
rect 5618 19964 5628 20020
rect 5684 19964 5964 20020
rect 6020 19964 6030 20020
rect 8866 19964 8876 20020
rect 8932 19964 10332 20020
rect 10388 19964 10398 20020
rect 12114 19964 12124 20020
rect 12180 19964 15484 20020
rect 15540 19964 15550 20020
rect 22306 19964 22316 20020
rect 22372 19964 24108 20020
rect 24164 19964 24174 20020
rect 25218 19964 25228 20020
rect 25284 19964 25676 20020
rect 25732 19964 25742 20020
rect 26898 19964 26908 20020
rect 26964 19964 29372 20020
rect 29428 19964 30044 20020
rect 30100 19964 30110 20020
rect 30482 19964 30492 20020
rect 30548 19964 31164 20020
rect 31220 19964 31230 20020
rect 42018 19964 42028 20020
rect 42084 19964 44268 20020
rect 44324 19964 44334 20020
rect 44930 19964 44940 20020
rect 44996 19964 46620 20020
rect 46676 19964 46686 20020
rect 46834 19964 46844 20020
rect 46900 19964 47180 20020
rect 47236 19964 47246 20020
rect 8418 19852 8428 19908
rect 8484 19852 11004 19908
rect 11060 19852 11070 19908
rect 20514 19852 20524 19908
rect 20580 19852 21644 19908
rect 21700 19852 21710 19908
rect 24322 19852 24332 19908
rect 24388 19852 27132 19908
rect 27188 19852 29036 19908
rect 29092 19852 29102 19908
rect 30268 19852 31724 19908
rect 31780 19852 31790 19908
rect 36194 19852 36204 19908
rect 36260 19852 37324 19908
rect 37380 19852 37390 19908
rect 44818 19852 44828 19908
rect 44884 19852 47852 19908
rect 47908 19852 47918 19908
rect 30268 19796 30324 19852
rect 7522 19740 7532 19796
rect 7588 19740 9100 19796
rect 9156 19740 9660 19796
rect 9716 19740 9726 19796
rect 28802 19740 28812 19796
rect 28868 19740 30268 19796
rect 30324 19740 30334 19796
rect 31042 19740 31052 19796
rect 31108 19740 31948 19796
rect 32004 19740 32014 19796
rect 45154 19740 45164 19796
rect 45220 19740 45948 19796
rect 46004 19740 46014 19796
rect 29586 19628 29596 19684
rect 29652 19628 30716 19684
rect 30772 19628 30782 19684
rect 43922 19628 43932 19684
rect 43988 19628 48076 19684
rect 48132 19628 48142 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 29698 19516 29708 19572
rect 29764 19516 31388 19572
rect 31444 19516 34076 19572
rect 34132 19516 34142 19572
rect 9202 19404 9212 19460
rect 9268 19404 11004 19460
rect 11060 19404 11070 19460
rect 24882 19404 24892 19460
rect 24948 19404 25676 19460
rect 25732 19404 25742 19460
rect 29474 19404 29484 19460
rect 29540 19404 30380 19460
rect 30436 19404 30446 19460
rect 43474 19404 43484 19460
rect 43540 19404 44716 19460
rect 44772 19404 44782 19460
rect 2818 19292 2828 19348
rect 2884 19292 3612 19348
rect 3668 19292 3678 19348
rect 10658 19292 10668 19348
rect 10724 19292 12124 19348
rect 12180 19292 12190 19348
rect 14018 19292 14028 19348
rect 14084 19292 14700 19348
rect 14756 19292 14766 19348
rect 15138 19292 15148 19348
rect 15204 19292 15820 19348
rect 15876 19292 15886 19348
rect 25442 19292 25452 19348
rect 25508 19292 30492 19348
rect 30548 19292 30558 19348
rect 36866 19292 36876 19348
rect 36932 19292 39676 19348
rect 39732 19292 39742 19348
rect 43698 19292 43708 19348
rect 43764 19292 44940 19348
rect 44996 19292 45006 19348
rect 4946 19180 4956 19236
rect 5012 19180 5628 19236
rect 5684 19180 6524 19236
rect 6580 19180 6590 19236
rect 10770 19180 10780 19236
rect 10836 19180 12236 19236
rect 12292 19180 13804 19236
rect 13860 19180 13870 19236
rect 25890 19180 25900 19236
rect 25956 19180 26908 19236
rect 26964 19180 26974 19236
rect 31154 19180 31164 19236
rect 31220 19180 33964 19236
rect 34020 19180 34030 19236
rect 38612 19180 38780 19236
rect 38836 19180 38846 19236
rect 10556 19068 11676 19124
rect 11732 19068 11742 19124
rect 10556 19012 10612 19068
rect 38612 19012 38668 19180
rect 41794 19068 41804 19124
rect 41860 19068 42700 19124
rect 42756 19068 42766 19124
rect 9986 18956 9996 19012
rect 10052 18956 10556 19012
rect 10612 18956 10622 19012
rect 11330 18956 11340 19012
rect 11396 18956 17612 19012
rect 17668 18956 17678 19012
rect 38434 18956 38444 19012
rect 38500 18956 38668 19012
rect 40002 18956 40012 19012
rect 40068 18956 42028 19012
rect 42084 18956 42094 19012
rect 46834 18956 46844 19012
rect 46900 18956 47068 19012
rect 47124 18956 47134 19012
rect 5954 18844 5964 18900
rect 6020 18844 6972 18900
rect 7028 18844 7038 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 9650 18732 9660 18788
rect 9716 18732 11452 18788
rect 11508 18732 11518 18788
rect 44230 18732 44268 18788
rect 44324 18732 44334 18788
rect 7074 18620 7084 18676
rect 7140 18620 8652 18676
rect 8708 18620 8718 18676
rect 10322 18620 10332 18676
rect 10388 18620 10398 18676
rect 25330 18620 25340 18676
rect 25396 18620 27132 18676
rect 27188 18620 28140 18676
rect 28196 18620 28206 18676
rect 38612 18620 41916 18676
rect 41972 18620 41982 18676
rect 1810 18396 1820 18452
rect 1876 18396 2828 18452
rect 2884 18396 5068 18452
rect 5124 18396 5134 18452
rect 5506 18396 5516 18452
rect 5572 18396 7308 18452
rect 7364 18396 7868 18452
rect 7924 18396 7934 18452
rect 8418 18396 8428 18452
rect 8484 18396 9996 18452
rect 10052 18396 10062 18452
rect 10332 18340 10388 18620
rect 38612 18564 38668 18620
rect 27794 18508 27804 18564
rect 27860 18508 29260 18564
rect 29316 18508 29326 18564
rect 30706 18508 30716 18564
rect 30772 18508 31500 18564
rect 31556 18508 31566 18564
rect 37650 18508 37660 18564
rect 37716 18508 38668 18564
rect 39900 18508 40404 18564
rect 42914 18508 42924 18564
rect 42980 18508 44604 18564
rect 44660 18508 44670 18564
rect 39900 18452 39956 18508
rect 10994 18396 11004 18452
rect 11060 18396 11900 18452
rect 11956 18396 11966 18452
rect 13458 18396 13468 18452
rect 13524 18396 14700 18452
rect 14756 18396 14766 18452
rect 16818 18396 16828 18452
rect 16884 18396 17388 18452
rect 17444 18396 17454 18452
rect 18050 18396 18060 18452
rect 18116 18396 19292 18452
rect 19348 18396 19358 18452
rect 24070 18396 24108 18452
rect 24164 18396 24174 18452
rect 25218 18396 25228 18452
rect 25284 18396 29708 18452
rect 29764 18396 31164 18452
rect 31220 18396 31230 18452
rect 32050 18396 32060 18452
rect 32116 18396 33516 18452
rect 33572 18396 34076 18452
rect 34132 18396 34142 18452
rect 38546 18396 38556 18452
rect 38612 18396 39956 18452
rect 40348 18452 40404 18508
rect 40348 18396 41020 18452
rect 41076 18396 42700 18452
rect 42756 18396 42766 18452
rect 44790 18396 44828 18452
rect 44884 18396 44894 18452
rect 45826 18396 45836 18452
rect 45892 18396 47516 18452
rect 47572 18396 47582 18452
rect 5618 18284 5628 18340
rect 5684 18284 6188 18340
rect 6244 18284 6254 18340
rect 8866 18284 8876 18340
rect 8932 18284 10388 18340
rect 17826 18284 17836 18340
rect 17892 18284 29596 18340
rect 29652 18284 29662 18340
rect 32498 18284 32508 18340
rect 32564 18284 33852 18340
rect 33908 18284 33918 18340
rect 44828 18284 47292 18340
rect 47348 18284 47628 18340
rect 47684 18284 47694 18340
rect 0 18228 800 18256
rect 44828 18228 44884 18284
rect 49200 18228 50000 18256
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 6962 18172 6972 18228
rect 7028 18172 8540 18228
rect 8596 18172 8606 18228
rect 14102 18172 14140 18228
rect 14196 18172 14206 18228
rect 23846 18172 23884 18228
rect 23940 18172 23950 18228
rect 24658 18172 24668 18228
rect 24724 18172 25228 18228
rect 25284 18172 26124 18228
rect 26180 18172 26190 18228
rect 39218 18172 39228 18228
rect 39284 18172 44828 18228
rect 44884 18172 44894 18228
rect 45602 18172 45612 18228
rect 45668 18172 46844 18228
rect 46900 18172 50000 18228
rect 0 18144 800 18172
rect 49200 18144 50000 18172
rect 22194 18060 22204 18116
rect 22260 18060 22876 18116
rect 22932 18060 23772 18116
rect 23828 18060 24780 18116
rect 24836 18060 24846 18116
rect 35644 18060 37100 18116
rect 37156 18060 37166 18116
rect 42578 18060 42588 18116
rect 42644 18060 46284 18116
rect 46340 18060 46732 18116
rect 46788 18060 47404 18116
rect 47460 18060 47470 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 23090 17948 23100 18004
rect 23156 17948 24332 18004
rect 24388 17948 25676 18004
rect 25732 17948 25742 18004
rect 27906 17948 27916 18004
rect 27972 17948 29932 18004
rect 29988 17948 29998 18004
rect 30258 17948 30268 18004
rect 30324 17948 34188 18004
rect 34244 17948 34254 18004
rect 35644 17892 35700 18060
rect 35858 17948 35868 18004
rect 35924 17948 35934 18004
rect 39218 17948 39228 18004
rect 39284 17948 40236 18004
rect 40292 17948 41020 18004
rect 41076 17948 43148 18004
rect 43204 17948 43214 18004
rect 5730 17836 5740 17892
rect 5796 17836 13076 17892
rect 13682 17836 13692 17892
rect 13748 17836 35700 17892
rect 13020 17780 13076 17836
rect 6402 17724 6412 17780
rect 6468 17724 7196 17780
rect 7252 17724 7262 17780
rect 13010 17724 13020 17780
rect 13076 17724 19068 17780
rect 19124 17724 19134 17780
rect 23958 17724 23996 17780
rect 24052 17724 24062 17780
rect 28802 17724 28812 17780
rect 28868 17724 30268 17780
rect 30324 17724 30334 17780
rect 6178 17612 6188 17668
rect 6244 17612 6972 17668
rect 7028 17612 7038 17668
rect 10882 17612 10892 17668
rect 10948 17612 13580 17668
rect 13636 17612 14028 17668
rect 14084 17612 20748 17668
rect 20804 17612 20814 17668
rect 23874 17612 23884 17668
rect 23940 17612 25340 17668
rect 25396 17612 25406 17668
rect 26562 17612 26572 17668
rect 26628 17612 29372 17668
rect 29428 17612 29438 17668
rect 30146 17612 30156 17668
rect 30212 17612 30716 17668
rect 30772 17612 30782 17668
rect 0 17556 800 17584
rect 35868 17556 35924 17948
rect 38612 17836 40348 17892
rect 40404 17836 40414 17892
rect 38612 17780 38668 17836
rect 36194 17724 36204 17780
rect 36260 17724 38668 17780
rect 39666 17724 39676 17780
rect 39732 17724 40124 17780
rect 40180 17724 42252 17780
rect 42308 17724 43036 17780
rect 43092 17724 43102 17780
rect 43474 17724 43484 17780
rect 43540 17724 44044 17780
rect 44100 17724 45052 17780
rect 45108 17724 45118 17780
rect 44258 17612 44268 17668
rect 44324 17612 46620 17668
rect 46676 17612 46686 17668
rect 46946 17612 46956 17668
rect 47012 17612 47628 17668
rect 47684 17612 47694 17668
rect 49200 17556 50000 17584
rect 0 17500 1932 17556
rect 1988 17500 1998 17556
rect 22530 17500 22540 17556
rect 22596 17500 23436 17556
rect 23492 17500 28028 17556
rect 28084 17500 28094 17556
rect 30930 17500 30940 17556
rect 30996 17500 35924 17556
rect 39330 17500 39340 17556
rect 39396 17500 44156 17556
rect 44212 17500 45836 17556
rect 45892 17500 45902 17556
rect 48178 17500 48188 17556
rect 48244 17500 50000 17556
rect 0 17472 800 17500
rect 43036 17444 43092 17500
rect 49200 17472 50000 17500
rect 4834 17388 4844 17444
rect 4900 17388 5852 17444
rect 5908 17388 11788 17444
rect 11844 17388 11854 17444
rect 23846 17388 23884 17444
rect 23940 17388 23950 17444
rect 43026 17388 43036 17444
rect 43092 17388 43102 17444
rect 43362 17388 43372 17444
rect 43428 17388 45052 17444
rect 45108 17388 45118 17444
rect 44818 17276 44828 17332
rect 44884 17276 44894 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 44828 17220 44884 17276
rect 28690 17164 28700 17220
rect 28756 17164 30492 17220
rect 30548 17164 33516 17220
rect 33572 17164 33582 17220
rect 43250 17164 43260 17220
rect 43316 17164 44884 17220
rect 47618 17164 47628 17220
rect 47684 17164 47852 17220
rect 47908 17164 47918 17220
rect 16818 17052 16828 17108
rect 16884 17052 17164 17108
rect 17220 17052 17230 17108
rect 42802 17052 42812 17108
rect 42868 17052 44044 17108
rect 44100 17052 44110 17108
rect 45826 17052 45836 17108
rect 45892 17052 46732 17108
rect 46788 17052 46798 17108
rect 15922 16940 15932 16996
rect 15988 16940 17276 16996
rect 17332 16940 17342 16996
rect 20962 16940 20972 16996
rect 21028 16940 21868 16996
rect 21924 16940 29596 16996
rect 29652 16940 30492 16996
rect 30548 16940 32956 16996
rect 33012 16940 37212 16996
rect 37268 16940 38220 16996
rect 38276 16940 38286 16996
rect 41010 16940 41020 16996
rect 41076 16940 41636 16996
rect 41906 16940 41916 16996
rect 41972 16940 43820 16996
rect 43876 16940 43886 16996
rect 46162 16940 46172 16996
rect 46228 16940 46238 16996
rect 41580 16884 41636 16940
rect 4610 16828 4620 16884
rect 4676 16828 5180 16884
rect 5236 16828 5246 16884
rect 16146 16828 16156 16884
rect 16212 16828 17612 16884
rect 17668 16828 17678 16884
rect 23986 16828 23996 16884
rect 24052 16828 25340 16884
rect 25396 16828 25406 16884
rect 31714 16828 31724 16884
rect 31780 16828 34300 16884
rect 34356 16828 34636 16884
rect 34692 16828 34702 16884
rect 37986 16828 37996 16884
rect 38052 16828 39004 16884
rect 39060 16828 39070 16884
rect 39778 16828 39788 16884
rect 39844 16828 40908 16884
rect 40964 16828 40974 16884
rect 41580 16828 43876 16884
rect 43820 16772 43876 16828
rect 2482 16716 2492 16772
rect 2548 16716 5068 16772
rect 5124 16716 5134 16772
rect 10770 16716 10780 16772
rect 10836 16716 13468 16772
rect 13524 16716 13534 16772
rect 14130 16716 14140 16772
rect 14196 16716 15036 16772
rect 15092 16716 15102 16772
rect 15250 16716 15260 16772
rect 15316 16716 15484 16772
rect 15540 16716 15550 16772
rect 15810 16716 15820 16772
rect 15876 16716 17724 16772
rect 17780 16716 17790 16772
rect 19170 16716 19180 16772
rect 19236 16716 20636 16772
rect 20692 16716 20702 16772
rect 24098 16716 24108 16772
rect 24164 16716 25676 16772
rect 25732 16716 25742 16772
rect 28130 16716 28140 16772
rect 28196 16716 29708 16772
rect 29764 16716 29774 16772
rect 39106 16716 39116 16772
rect 39172 16716 41020 16772
rect 41076 16716 41086 16772
rect 41346 16716 41356 16772
rect 41412 16716 42140 16772
rect 42196 16716 43036 16772
rect 43092 16716 43102 16772
rect 43810 16716 43820 16772
rect 43876 16716 43886 16772
rect 46172 16660 46228 16940
rect 3378 16604 3388 16660
rect 3444 16604 4956 16660
rect 5012 16604 5022 16660
rect 8194 16604 8204 16660
rect 8260 16604 10892 16660
rect 10948 16604 11788 16660
rect 11844 16604 11854 16660
rect 14466 16604 14476 16660
rect 14532 16604 17500 16660
rect 17556 16604 17566 16660
rect 27682 16604 27692 16660
rect 27748 16604 28252 16660
rect 28308 16604 28318 16660
rect 31892 16604 35756 16660
rect 35812 16604 35822 16660
rect 43474 16604 43484 16660
rect 43540 16604 45612 16660
rect 45668 16604 48076 16660
rect 48132 16604 48142 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 31892 16436 31948 16604
rect 44258 16492 44268 16548
rect 44324 16492 45052 16548
rect 45108 16492 45118 16548
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 5170 16380 5180 16436
rect 5236 16380 14700 16436
rect 14756 16380 14766 16436
rect 21746 16380 21756 16436
rect 21812 16380 29820 16436
rect 29876 16380 31948 16436
rect 43026 16380 43036 16436
rect 43092 16380 46620 16436
rect 46676 16380 46686 16436
rect 4050 16268 4060 16324
rect 4116 16268 6412 16324
rect 6468 16268 6478 16324
rect 10210 16268 10220 16324
rect 10276 16268 11228 16324
rect 11284 16268 11294 16324
rect 22418 16268 22428 16324
rect 22484 16268 23100 16324
rect 23156 16268 23548 16324
rect 23604 16268 23614 16324
rect 23772 16268 27300 16324
rect 35970 16268 35980 16324
rect 36036 16268 38108 16324
rect 38164 16268 43260 16324
rect 43316 16268 43326 16324
rect 8194 16156 8204 16212
rect 8260 16156 10556 16212
rect 10612 16156 10622 16212
rect 13794 16156 13804 16212
rect 13860 16156 16156 16212
rect 16212 16156 16222 16212
rect 20066 16156 20076 16212
rect 20132 16156 21420 16212
rect 21476 16156 22092 16212
rect 22148 16156 22158 16212
rect 6738 16044 6748 16100
rect 6804 16044 8092 16100
rect 8148 16044 8764 16100
rect 8820 16044 8830 16100
rect 9986 16044 9996 16100
rect 10052 16044 10444 16100
rect 10500 16044 12236 16100
rect 12292 16044 12302 16100
rect 12786 16044 12796 16100
rect 12852 16044 15372 16100
rect 15428 16044 15438 16100
rect 18722 16044 18732 16100
rect 18788 16044 19628 16100
rect 19684 16044 19694 16100
rect 21634 16044 21644 16100
rect 21700 16044 21980 16100
rect 22036 16044 22876 16100
rect 22932 16044 22942 16100
rect 23772 15988 23828 16268
rect 27244 16212 27300 16268
rect 49200 16212 50000 16240
rect 25218 16156 25228 16212
rect 25284 16156 27020 16212
rect 27076 16156 27086 16212
rect 27244 16156 37100 16212
rect 37156 16156 37166 16212
rect 41906 16156 41916 16212
rect 41972 16156 42364 16212
rect 42420 16156 42430 16212
rect 43334 16156 43372 16212
rect 43428 16156 43438 16212
rect 47954 16156 47964 16212
rect 48020 16156 50000 16212
rect 49200 16128 50000 16156
rect 42130 16044 42140 16100
rect 42196 16044 42812 16100
rect 42868 16044 45500 16100
rect 45556 16044 45566 16100
rect 3332 15932 6188 15988
rect 6244 15932 10220 15988
rect 10276 15932 10286 15988
rect 13010 15932 13020 15988
rect 13076 15932 13580 15988
rect 13636 15932 13646 15988
rect 13794 15932 13804 15988
rect 13860 15932 14028 15988
rect 14084 15932 14094 15988
rect 14242 15932 14252 15988
rect 14308 15932 15260 15988
rect 15316 15932 15326 15988
rect 17378 15932 17388 15988
rect 17444 15932 18060 15988
rect 18116 15932 18508 15988
rect 18564 15932 19180 15988
rect 19236 15932 19246 15988
rect 20514 15932 20524 15988
rect 20580 15932 23828 15988
rect 28578 15932 28588 15988
rect 28644 15932 29484 15988
rect 29540 15932 29550 15988
rect 33282 15932 33292 15988
rect 33348 15932 40460 15988
rect 40516 15932 40526 15988
rect 42466 15932 42476 15988
rect 42532 15932 43036 15988
rect 43092 15932 43102 15988
rect 43922 15932 43932 15988
rect 43988 15932 47964 15988
rect 48020 15932 48030 15988
rect 3332 15876 3388 15932
rect 2930 15820 2940 15876
rect 2996 15820 3388 15876
rect 5954 15820 5964 15876
rect 6020 15820 7868 15876
rect 7924 15820 7934 15876
rect 13458 15820 13468 15876
rect 13524 15820 14476 15876
rect 14532 15820 14542 15876
rect 27682 15820 27692 15876
rect 27748 15820 30044 15876
rect 30100 15820 30110 15876
rect 36194 15820 36204 15876
rect 36260 15820 36988 15876
rect 37044 15820 37054 15876
rect 4162 15708 4172 15764
rect 4228 15708 5292 15764
rect 5348 15708 6188 15764
rect 6244 15708 8428 15764
rect 8484 15708 8494 15764
rect 9650 15708 9660 15764
rect 9716 15708 9996 15764
rect 10052 15708 10062 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 29484 15652 29540 15820
rect 14802 15596 14812 15652
rect 14868 15596 15596 15652
rect 15652 15596 15662 15652
rect 29474 15596 29484 15652
rect 29540 15596 29550 15652
rect 11666 15484 11676 15540
rect 11732 15484 12684 15540
rect 12740 15484 12750 15540
rect 16146 15484 16156 15540
rect 16212 15484 33404 15540
rect 33460 15484 33470 15540
rect 3266 15372 3276 15428
rect 3332 15372 3836 15428
rect 3892 15372 5180 15428
rect 5236 15372 5246 15428
rect 6066 15372 6076 15428
rect 6132 15372 7756 15428
rect 7812 15372 8204 15428
rect 8260 15372 9100 15428
rect 9156 15372 9166 15428
rect 15922 15372 15932 15428
rect 15988 15372 16604 15428
rect 16660 15372 16670 15428
rect 23650 15372 23660 15428
rect 23716 15372 25228 15428
rect 25284 15372 25294 15428
rect 31490 15372 31500 15428
rect 31556 15372 32172 15428
rect 32228 15372 32238 15428
rect 36306 15372 36316 15428
rect 36372 15372 38556 15428
rect 38612 15372 38622 15428
rect 43362 15372 43372 15428
rect 43428 15372 43932 15428
rect 43988 15372 43998 15428
rect 4386 15260 4396 15316
rect 4452 15260 5516 15316
rect 5572 15260 5582 15316
rect 8418 15260 8428 15316
rect 8484 15260 8988 15316
rect 9044 15260 9772 15316
rect 9828 15260 9838 15316
rect 10210 15260 10220 15316
rect 10276 15260 11676 15316
rect 11732 15260 11742 15316
rect 13794 15260 13804 15316
rect 13860 15260 15148 15316
rect 15474 15260 15484 15316
rect 15540 15260 16156 15316
rect 16212 15260 16222 15316
rect 20178 15260 20188 15316
rect 20244 15260 20972 15316
rect 21028 15260 21038 15316
rect 24210 15260 24220 15316
rect 24276 15260 26460 15316
rect 26516 15260 26526 15316
rect 28914 15260 28924 15316
rect 28980 15260 32396 15316
rect 32452 15260 32462 15316
rect 38322 15260 38332 15316
rect 38388 15260 39116 15316
rect 39172 15260 39182 15316
rect 41682 15260 41692 15316
rect 41748 15260 42364 15316
rect 42420 15260 43148 15316
rect 43204 15260 43214 15316
rect 44146 15260 44156 15316
rect 44212 15260 45276 15316
rect 45332 15260 46956 15316
rect 47012 15260 47022 15316
rect 15092 15204 15148 15260
rect 15092 15148 15708 15204
rect 15764 15148 15774 15204
rect 25554 15148 25564 15204
rect 25620 15148 25788 15204
rect 25844 15148 25854 15204
rect 37762 15148 37772 15204
rect 37828 15148 38668 15204
rect 38724 15148 38734 15204
rect 44370 15148 44380 15204
rect 44436 15148 45052 15204
rect 45108 15148 45612 15204
rect 45668 15148 45678 15204
rect 3948 15036 4396 15092
rect 4452 15036 4462 15092
rect 7186 15036 7196 15092
rect 7252 15036 8204 15092
rect 8260 15036 8270 15092
rect 10434 15036 10444 15092
rect 10500 15036 11452 15092
rect 11508 15036 11518 15092
rect 18834 15036 18844 15092
rect 18900 15036 19516 15092
rect 19572 15036 19582 15092
rect 25554 15036 25564 15092
rect 25620 15036 27020 15092
rect 27076 15036 27086 15092
rect 37090 15036 37100 15092
rect 37156 15036 43372 15092
rect 43428 15036 43438 15092
rect 3948 14980 4004 15036
rect 3938 14924 3948 14980
rect 4004 14924 4014 14980
rect 14690 14924 14700 14980
rect 14756 14924 14766 14980
rect 26338 14924 26348 14980
rect 26404 14924 27916 14980
rect 27972 14924 27982 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 12002 14812 12012 14868
rect 12068 14812 14364 14868
rect 14420 14812 14430 14868
rect 7074 14700 7084 14756
rect 7140 14700 11116 14756
rect 11172 14700 11182 14756
rect 11554 14700 11564 14756
rect 11620 14700 12348 14756
rect 12404 14700 12414 14756
rect 14700 14644 14756 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 21746 14812 21756 14868
rect 21812 14812 24780 14868
rect 24836 14812 26124 14868
rect 26180 14812 26190 14868
rect 27682 14812 27692 14868
rect 27748 14812 28252 14868
rect 28308 14812 28318 14868
rect 45938 14812 45948 14868
rect 46004 14812 46014 14868
rect 25890 14700 25900 14756
rect 25956 14700 26796 14756
rect 26852 14700 26862 14756
rect 43698 14700 43708 14756
rect 43764 14700 45164 14756
rect 45220 14700 45230 14756
rect 10322 14588 10332 14644
rect 10388 14588 14252 14644
rect 14308 14588 14318 14644
rect 14466 14588 14476 14644
rect 14532 14588 17668 14644
rect 34626 14588 34636 14644
rect 34692 14588 35644 14644
rect 35700 14588 35710 14644
rect 38210 14588 38220 14644
rect 38276 14588 39900 14644
rect 39956 14588 39966 14644
rect 41458 14588 41468 14644
rect 41524 14588 44268 14644
rect 44324 14588 44334 14644
rect 5058 14476 5068 14532
rect 5124 14476 8764 14532
rect 8820 14476 10668 14532
rect 10724 14476 11284 14532
rect 2482 14364 2492 14420
rect 2548 14364 3612 14420
rect 3668 14364 3678 14420
rect 4946 14364 4956 14420
rect 5012 14364 5628 14420
rect 5684 14364 5694 14420
rect 6290 14364 6300 14420
rect 6356 14364 9324 14420
rect 9380 14364 9390 14420
rect 11228 14308 11284 14476
rect 11442 14364 11452 14420
rect 11508 14364 12572 14420
rect 12628 14364 12638 14420
rect 11228 14252 12684 14308
rect 12740 14252 12750 14308
rect 13010 14252 13020 14308
rect 13076 14252 13804 14308
rect 13860 14252 13870 14308
rect 14252 14196 14308 14588
rect 14802 14476 14812 14532
rect 14868 14476 17388 14532
rect 17444 14476 17454 14532
rect 17612 14420 17668 14588
rect 23762 14476 23772 14532
rect 23828 14476 26236 14532
rect 26292 14476 26302 14532
rect 27122 14476 27132 14532
rect 27188 14476 27692 14532
rect 27748 14476 27758 14532
rect 31266 14476 31276 14532
rect 31332 14476 34748 14532
rect 34804 14476 35532 14532
rect 35588 14476 35598 14532
rect 40898 14476 40908 14532
rect 40964 14476 41636 14532
rect 41580 14420 41636 14476
rect 45948 14420 46004 14812
rect 17266 14364 17276 14420
rect 17332 14364 18620 14420
rect 18676 14364 18686 14420
rect 25526 14364 25564 14420
rect 25620 14364 25630 14420
rect 32946 14364 32956 14420
rect 33012 14364 34412 14420
rect 34468 14364 34478 14420
rect 35186 14364 35196 14420
rect 35252 14364 35868 14420
rect 35924 14364 35934 14420
rect 38658 14364 38668 14420
rect 38724 14364 40012 14420
rect 40068 14364 40078 14420
rect 40674 14364 40684 14420
rect 40740 14364 41244 14420
rect 41300 14364 41310 14420
rect 41570 14364 41580 14420
rect 41636 14364 42588 14420
rect 42644 14364 44828 14420
rect 44884 14364 44894 14420
rect 45714 14364 45724 14420
rect 45780 14364 47068 14420
rect 47124 14364 47134 14420
rect 18386 14252 18396 14308
rect 18452 14252 18844 14308
rect 18900 14252 18910 14308
rect 23314 14252 23324 14308
rect 23380 14252 23884 14308
rect 23940 14252 24220 14308
rect 24276 14252 25116 14308
rect 25172 14252 25182 14308
rect 27570 14252 27580 14308
rect 27636 14252 34076 14308
rect 34132 14252 34142 14308
rect 41346 14252 41356 14308
rect 41412 14252 42476 14308
rect 42532 14252 42542 14308
rect 14252 14140 15484 14196
rect 15540 14140 15550 14196
rect 34290 14140 34300 14196
rect 34356 14140 36092 14196
rect 36148 14140 37548 14196
rect 37604 14140 37614 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 28130 14028 28140 14084
rect 28196 14028 32844 14084
rect 32900 14028 32910 14084
rect 45378 14028 45388 14084
rect 45444 14028 45948 14084
rect 46004 14028 46956 14084
rect 47012 14028 47022 14084
rect 7410 13916 7420 13972
rect 7476 13916 9660 13972
rect 9716 13916 9726 13972
rect 10882 13916 10892 13972
rect 10948 13916 12964 13972
rect 12908 13860 12964 13916
rect 26852 13916 31108 13972
rect 31826 13916 31836 13972
rect 31892 13916 32396 13972
rect 32452 13916 36428 13972
rect 36484 13916 37100 13972
rect 37156 13916 37166 13972
rect 44370 13916 44380 13972
rect 44436 13916 48076 13972
rect 48132 13916 48142 13972
rect 26852 13860 26908 13916
rect 31052 13860 31108 13916
rect 7186 13804 7196 13860
rect 7252 13804 7756 13860
rect 7812 13804 8652 13860
rect 8708 13804 8718 13860
rect 9874 13804 9884 13860
rect 9940 13804 10556 13860
rect 10612 13804 11340 13860
rect 11396 13804 11406 13860
rect 12898 13804 12908 13860
rect 12964 13804 13916 13860
rect 13972 13804 13982 13860
rect 14578 13804 14588 13860
rect 14644 13804 26908 13860
rect 27010 13804 27020 13860
rect 27076 13804 27468 13860
rect 27524 13804 27534 13860
rect 31042 13804 31052 13860
rect 31108 13804 31118 13860
rect 37986 13804 37996 13860
rect 38052 13804 38892 13860
rect 38948 13804 39788 13860
rect 39844 13804 39854 13860
rect 40114 13804 40124 13860
rect 40180 13804 41132 13860
rect 41188 13804 43260 13860
rect 43316 13804 43326 13860
rect 44594 13804 44604 13860
rect 44660 13804 47852 13860
rect 47908 13804 47918 13860
rect 3826 13692 3836 13748
rect 3892 13692 4284 13748
rect 4340 13692 6748 13748
rect 6804 13692 7308 13748
rect 7364 13692 7374 13748
rect 7522 13692 7532 13748
rect 7588 13692 7980 13748
rect 8036 13692 8316 13748
rect 8372 13692 8382 13748
rect 10322 13692 10332 13748
rect 10388 13692 12348 13748
rect 12404 13692 12414 13748
rect 27346 13692 27356 13748
rect 27412 13692 28252 13748
rect 28308 13692 28318 13748
rect 28914 13692 28924 13748
rect 28980 13692 28990 13748
rect 29922 13692 29932 13748
rect 29988 13692 31500 13748
rect 31556 13692 31566 13748
rect 39890 13692 39900 13748
rect 39956 13692 40572 13748
rect 40628 13692 41468 13748
rect 41524 13692 41534 13748
rect 41906 13692 41916 13748
rect 41972 13692 42700 13748
rect 42756 13692 43260 13748
rect 43316 13692 43326 13748
rect 46834 13692 46844 13748
rect 46900 13692 48188 13748
rect 48244 13692 48254 13748
rect 8194 13580 8204 13636
rect 8260 13580 9548 13636
rect 9604 13580 9614 13636
rect 18722 13580 18732 13636
rect 18788 13580 21420 13636
rect 21476 13580 21486 13636
rect 26226 13580 26236 13636
rect 26292 13580 27468 13636
rect 27524 13580 27534 13636
rect 28924 13524 28980 13692
rect 35858 13580 35868 13636
rect 35924 13580 38108 13636
rect 38164 13580 38174 13636
rect 45266 13580 45276 13636
rect 45332 13580 46508 13636
rect 46564 13580 46574 13636
rect 4284 13468 4508 13524
rect 4564 13468 4900 13524
rect 9874 13468 9884 13524
rect 9940 13468 13580 13524
rect 13636 13468 13646 13524
rect 13804 13468 14812 13524
rect 14868 13468 14878 13524
rect 26562 13468 26572 13524
rect 26628 13468 28980 13524
rect 4284 13412 4340 13468
rect 3714 13356 3724 13412
rect 3780 13356 4340 13412
rect 4844 13412 4900 13468
rect 4844 13356 6636 13412
rect 6692 13356 6702 13412
rect 10658 13356 10668 13412
rect 10724 13356 13244 13412
rect 13300 13356 13310 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 13804 13300 13860 13468
rect 17602 13356 17612 13412
rect 17668 13356 23548 13412
rect 23604 13356 24556 13412
rect 24612 13356 24622 13412
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 13570 13244 13580 13300
rect 13636 13244 13860 13300
rect 17490 13244 17500 13300
rect 17556 13244 22092 13300
rect 22148 13244 23436 13300
rect 23492 13244 28028 13300
rect 28084 13244 28094 13300
rect 40226 13244 40236 13300
rect 40292 13244 41244 13300
rect 41300 13244 41310 13300
rect 9202 13132 9212 13188
rect 9268 13132 9996 13188
rect 10052 13132 10062 13188
rect 12226 13132 12236 13188
rect 12292 13132 12684 13188
rect 12740 13132 13468 13188
rect 13524 13132 13534 13188
rect 29586 13132 29596 13188
rect 29652 13132 31388 13188
rect 31444 13132 31454 13188
rect 31602 13132 31612 13188
rect 31668 13132 32060 13188
rect 32116 13132 32126 13188
rect 8530 13020 8540 13076
rect 8596 13020 10108 13076
rect 10164 13020 10174 13076
rect 11666 13020 11676 13076
rect 11732 13020 12124 13076
rect 12180 13020 12190 13076
rect 14914 13020 14924 13076
rect 14980 13020 15596 13076
rect 15652 13020 16716 13076
rect 16772 13020 16782 13076
rect 26338 13020 26348 13076
rect 26404 13020 27244 13076
rect 27300 13020 27310 13076
rect 29698 13020 29708 13076
rect 29764 13020 32284 13076
rect 32340 13020 32732 13076
rect 32788 13020 33516 13076
rect 33572 13020 33582 13076
rect 35746 13020 35756 13076
rect 35812 13020 36316 13076
rect 36372 13020 38668 13076
rect 43586 13020 43596 13076
rect 43652 13020 45836 13076
rect 45892 13020 45902 13076
rect 46050 13020 46060 13076
rect 46116 13020 46620 13076
rect 46676 13020 47964 13076
rect 48020 13020 48030 13076
rect 38612 12964 38668 13020
rect 9772 12908 14700 12964
rect 14756 12908 15148 12964
rect 15250 12908 15260 12964
rect 15316 12908 15708 12964
rect 15764 12908 18172 12964
rect 18228 12908 18238 12964
rect 23986 12908 23996 12964
rect 24052 12908 25564 12964
rect 25620 12908 26236 12964
rect 26292 12908 26302 12964
rect 28354 12908 28364 12964
rect 28420 12908 31052 12964
rect 31108 12908 31118 12964
rect 38612 12908 40236 12964
rect 40292 12908 40302 12964
rect 4722 12796 4732 12852
rect 4788 12796 5292 12852
rect 5348 12796 5358 12852
rect 9772 12740 9828 12908
rect 15092 12852 15148 12908
rect 49200 12852 50000 12880
rect 10210 12796 10220 12852
rect 10276 12796 12684 12852
rect 12740 12796 13356 12852
rect 13412 12796 13422 12852
rect 15092 12796 15820 12852
rect 15876 12796 15886 12852
rect 18722 12796 18732 12852
rect 18788 12796 19628 12852
rect 19684 12796 19694 12852
rect 22418 12796 22428 12852
rect 22484 12796 22494 12852
rect 26674 12796 26684 12852
rect 26740 12796 26908 12852
rect 31938 12796 31948 12852
rect 32004 12796 33180 12852
rect 33236 12796 33246 12852
rect 47954 12796 47964 12852
rect 48020 12796 50000 12852
rect 3938 12684 3948 12740
rect 4004 12684 5964 12740
rect 6020 12684 6030 12740
rect 8866 12684 8876 12740
rect 8932 12684 9772 12740
rect 9828 12684 9838 12740
rect 10220 12628 10276 12796
rect 22428 12740 22484 12796
rect 26852 12740 26908 12796
rect 49200 12768 50000 12796
rect 16370 12684 16380 12740
rect 16436 12684 17836 12740
rect 17892 12684 18508 12740
rect 18564 12684 18574 12740
rect 22194 12684 22204 12740
rect 22260 12684 23436 12740
rect 23492 12684 24108 12740
rect 24164 12684 25228 12740
rect 25284 12684 25294 12740
rect 26852 12684 27244 12740
rect 27300 12684 29148 12740
rect 29204 12684 29214 12740
rect 8754 12572 8764 12628
rect 8820 12572 9324 12628
rect 9380 12572 10276 12628
rect 18050 12572 18060 12628
rect 18116 12572 18284 12628
rect 18340 12572 18956 12628
rect 19012 12572 19022 12628
rect 24210 12572 24220 12628
rect 24276 12572 29372 12628
rect 29428 12572 29438 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 9762 12460 9772 12516
rect 9828 12460 14364 12516
rect 14420 12460 14430 12516
rect 21410 12460 21420 12516
rect 21476 12460 40236 12516
rect 40292 12460 41356 12516
rect 41412 12460 42252 12516
rect 42308 12460 42318 12516
rect 6626 12348 6636 12404
rect 6692 12348 7756 12404
rect 7812 12348 9996 12404
rect 10052 12348 10062 12404
rect 13458 12348 13468 12404
rect 13524 12348 14028 12404
rect 14084 12348 14094 12404
rect 16258 12348 16268 12404
rect 16324 12348 17500 12404
rect 17556 12348 17836 12404
rect 17892 12348 17902 12404
rect 21970 12348 21980 12404
rect 22036 12348 22876 12404
rect 22932 12348 22942 12404
rect 24546 12348 24556 12404
rect 24612 12348 25452 12404
rect 25508 12348 25518 12404
rect 26450 12348 26460 12404
rect 26516 12348 26684 12404
rect 26740 12348 26750 12404
rect 31378 12348 31388 12404
rect 31444 12348 32732 12404
rect 32788 12348 32798 12404
rect 33506 12348 33516 12404
rect 33572 12348 35980 12404
rect 36036 12348 36046 12404
rect 37090 12348 37100 12404
rect 37156 12348 37996 12404
rect 38052 12348 38062 12404
rect 44930 12348 44940 12404
rect 44996 12348 45836 12404
rect 45892 12348 45902 12404
rect 6402 12236 6412 12292
rect 6468 12236 8652 12292
rect 8708 12236 15932 12292
rect 15988 12236 15998 12292
rect 16268 12180 16324 12348
rect 19394 12236 19404 12292
rect 19460 12236 21532 12292
rect 21588 12236 21598 12292
rect 22306 12236 22316 12292
rect 22372 12236 22382 12292
rect 22754 12236 22764 12292
rect 22820 12236 23884 12292
rect 23940 12236 23950 12292
rect 24658 12236 24668 12292
rect 24724 12236 25676 12292
rect 25732 12236 25742 12292
rect 26852 12236 29036 12292
rect 29092 12236 29102 12292
rect 31266 12236 31276 12292
rect 31332 12236 31836 12292
rect 31892 12236 33964 12292
rect 34020 12236 34030 12292
rect 34178 12236 34188 12292
rect 34244 12236 34860 12292
rect 34916 12236 34926 12292
rect 35858 12236 35868 12292
rect 35924 12236 38444 12292
rect 38500 12236 39172 12292
rect 43698 12236 43708 12292
rect 43764 12236 44156 12292
rect 44212 12236 44222 12292
rect 44370 12236 44380 12292
rect 44436 12236 45052 12292
rect 45108 12236 45118 12292
rect 4834 12124 4844 12180
rect 4900 12124 5740 12180
rect 5796 12124 5806 12180
rect 12898 12124 12908 12180
rect 12964 12124 13692 12180
rect 13748 12124 14700 12180
rect 14756 12124 14766 12180
rect 15026 12124 15036 12180
rect 15092 12124 16324 12180
rect 18834 12124 18844 12180
rect 18900 12124 19292 12180
rect 19348 12124 19740 12180
rect 19796 12124 19806 12180
rect 22316 12068 22372 12236
rect 26852 12068 26908 12236
rect 39116 12180 39172 12236
rect 49200 12180 50000 12208
rect 27234 12124 27244 12180
rect 27300 12124 28028 12180
rect 28084 12124 28094 12180
rect 28242 12124 28252 12180
rect 28308 12124 29596 12180
rect 29652 12124 29932 12180
rect 29988 12124 29998 12180
rect 32498 12124 32508 12180
rect 32564 12124 34412 12180
rect 34468 12124 34478 12180
rect 36306 12124 36316 12180
rect 36372 12124 37212 12180
rect 37268 12124 37772 12180
rect 37828 12124 37838 12180
rect 38770 12124 38780 12180
rect 38836 12124 38846 12180
rect 39106 12124 39116 12180
rect 39172 12124 39182 12180
rect 48178 12124 48188 12180
rect 48244 12124 50000 12180
rect 2482 12012 2492 12068
rect 2548 12012 4732 12068
rect 4788 12012 4798 12068
rect 6514 12012 6524 12068
rect 6580 12012 7420 12068
rect 7476 12012 8428 12068
rect 8484 12012 13020 12068
rect 13076 12012 13086 12068
rect 13906 12012 13916 12068
rect 13972 12012 14588 12068
rect 14644 12012 14654 12068
rect 21186 12012 21196 12068
rect 21252 12012 23212 12068
rect 23268 12012 23278 12068
rect 25554 12012 25564 12068
rect 25620 12012 26908 12068
rect 38780 11956 38836 12124
rect 49200 12096 50000 12124
rect 4834 11900 4844 11956
rect 4900 11900 6748 11956
rect 6804 11900 6814 11956
rect 29474 11900 29484 11956
rect 29540 11900 29820 11956
rect 29876 11900 30492 11956
rect 30548 11900 30558 11956
rect 31714 11900 31724 11956
rect 31780 11900 32284 11956
rect 32340 11900 33740 11956
rect 33796 11900 34076 11956
rect 34132 11900 34142 11956
rect 34402 11900 34412 11956
rect 34468 11900 36764 11956
rect 36820 11900 36830 11956
rect 37986 11900 37996 11956
rect 38052 11900 38836 11956
rect 4844 11788 5292 11844
rect 5348 11788 5358 11844
rect 11778 11788 11788 11844
rect 11844 11788 12572 11844
rect 12628 11788 12638 11844
rect 27682 11788 27692 11844
rect 27748 11788 28476 11844
rect 28532 11788 28542 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 4844 11620 4900 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 14802 11676 14812 11732
rect 14868 11676 16380 11732
rect 16436 11676 16446 11732
rect 4722 11564 4732 11620
rect 4788 11564 4900 11620
rect 34962 11564 34972 11620
rect 35028 11564 35644 11620
rect 35700 11564 36540 11620
rect 36596 11564 36606 11620
rect 49200 11508 50000 11536
rect 16482 11452 16492 11508
rect 16548 11452 17948 11508
rect 18004 11452 19516 11508
rect 19572 11452 19582 11508
rect 47954 11452 47964 11508
rect 48020 11452 50000 11508
rect 1810 11340 1820 11396
rect 1876 11340 5068 11396
rect 5124 11340 5134 11396
rect 7970 11340 7980 11396
rect 8036 11340 10108 11396
rect 10164 11340 10174 11396
rect 14242 11340 14252 11396
rect 14308 11340 14318 11396
rect 15026 11340 15036 11396
rect 15092 11340 16044 11396
rect 16100 11340 16110 11396
rect 9202 11228 9212 11284
rect 9268 11228 11116 11284
rect 11172 11228 11182 11284
rect 12450 11228 12460 11284
rect 12516 11228 13804 11284
rect 13860 11228 13870 11284
rect 14252 11172 14308 11340
rect 18956 11284 19012 11452
rect 49200 11424 50000 11452
rect 21746 11340 21756 11396
rect 21812 11340 22540 11396
rect 22596 11340 23436 11396
rect 23492 11340 23502 11396
rect 26786 11340 26796 11396
rect 26852 11340 27804 11396
rect 27860 11340 27870 11396
rect 30034 11340 30044 11396
rect 30100 11340 30716 11396
rect 30772 11340 30782 11396
rect 31042 11340 31052 11396
rect 31108 11340 31724 11396
rect 31780 11340 31790 11396
rect 18946 11228 18956 11284
rect 19012 11228 19022 11284
rect 22866 11228 22876 11284
rect 22932 11228 23324 11284
rect 23380 11228 24332 11284
rect 24388 11228 24398 11284
rect 27570 11228 27580 11284
rect 27636 11228 29484 11284
rect 29540 11228 29550 11284
rect 32610 11228 32620 11284
rect 32676 11228 33180 11284
rect 33236 11228 36876 11284
rect 36932 11228 36942 11284
rect 11330 11116 11340 11172
rect 11396 11116 11788 11172
rect 11844 11116 12348 11172
rect 12404 11116 12414 11172
rect 14252 11116 15596 11172
rect 15652 11116 15662 11172
rect 19618 11116 19628 11172
rect 19684 11116 22652 11172
rect 22708 11116 22718 11172
rect 36418 11116 36428 11172
rect 36484 11116 37100 11172
rect 37156 11116 37166 11172
rect 12562 11004 12572 11060
rect 12628 11004 13916 11060
rect 13972 11004 16828 11060
rect 16884 11004 16894 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 43922 10892 43932 10948
rect 43988 10892 44716 10948
rect 44772 10892 44782 10948
rect 49200 10836 50000 10864
rect 26786 10780 26796 10836
rect 26852 10780 29988 10836
rect 38434 10780 38444 10836
rect 38500 10780 38892 10836
rect 38948 10780 39228 10836
rect 39284 10780 39294 10836
rect 47618 10780 47628 10836
rect 47684 10780 48188 10836
rect 48244 10780 50000 10836
rect 10770 10668 10780 10724
rect 10836 10668 11900 10724
rect 11956 10668 13356 10724
rect 13412 10668 13422 10724
rect 15698 10668 15708 10724
rect 15764 10668 17388 10724
rect 17444 10668 18284 10724
rect 18340 10668 18350 10724
rect 27794 10668 27804 10724
rect 27860 10668 28924 10724
rect 28980 10668 28990 10724
rect 29932 10612 29988 10780
rect 49200 10752 50000 10780
rect 31154 10668 31164 10724
rect 31220 10668 32396 10724
rect 32452 10668 33068 10724
rect 33124 10668 34748 10724
rect 34804 10668 34814 10724
rect 44930 10668 44940 10724
rect 44996 10668 47852 10724
rect 47908 10668 47918 10724
rect 18386 10556 18396 10612
rect 18452 10556 19068 10612
rect 19124 10556 19134 10612
rect 22642 10556 22652 10612
rect 22708 10556 23212 10612
rect 23268 10556 23278 10612
rect 25218 10556 25228 10612
rect 25284 10556 26460 10612
rect 26516 10556 26908 10612
rect 26964 10556 26974 10612
rect 27906 10556 27916 10612
rect 27972 10556 28364 10612
rect 28420 10556 28430 10612
rect 29922 10556 29932 10612
rect 29988 10556 34524 10612
rect 34580 10556 34590 10612
rect 4274 10444 4284 10500
rect 4340 10444 5068 10500
rect 5124 10444 7532 10500
rect 7588 10444 7598 10500
rect 44034 10444 44044 10500
rect 44100 10444 45164 10500
rect 45220 10444 45230 10500
rect 46050 10444 46060 10500
rect 46116 10444 47404 10500
rect 47460 10444 47470 10500
rect 26898 10332 26908 10388
rect 26964 10332 27356 10388
rect 27412 10332 27422 10388
rect 37314 10220 37324 10276
rect 37380 10220 37884 10276
rect 37940 10220 37950 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 26114 10108 26124 10164
rect 26180 10108 26572 10164
rect 26628 10108 26638 10164
rect 28690 10108 28700 10164
rect 28756 10108 30716 10164
rect 30772 10108 30782 10164
rect 33842 10108 33852 10164
rect 33908 10108 35028 10164
rect 38210 10108 38220 10164
rect 38276 10108 38780 10164
rect 38836 10108 38846 10164
rect 34972 10052 35028 10108
rect 34972 9996 35420 10052
rect 35476 9996 36652 10052
rect 36708 9996 36988 10052
rect 37044 9996 37054 10052
rect 37762 9996 37772 10052
rect 37828 9996 39228 10052
rect 39284 9996 39294 10052
rect 25778 9884 25788 9940
rect 25844 9884 27356 9940
rect 27412 9884 27422 9940
rect 27570 9884 27580 9940
rect 27636 9884 28252 9940
rect 28308 9884 28318 9940
rect 33618 9884 33628 9940
rect 33684 9884 34412 9940
rect 34468 9884 34478 9940
rect 38556 9884 39340 9940
rect 39396 9884 39406 9940
rect 39554 9884 39564 9940
rect 39620 9884 41356 9940
rect 41412 9884 41422 9940
rect 10770 9772 10780 9828
rect 10836 9772 11900 9828
rect 11956 9772 11966 9828
rect 12114 9772 12124 9828
rect 12180 9772 12572 9828
rect 12628 9772 12908 9828
rect 12964 9772 12974 9828
rect 14242 9772 14252 9828
rect 14308 9772 14318 9828
rect 14466 9772 14476 9828
rect 14532 9772 17276 9828
rect 17332 9772 17948 9828
rect 18004 9772 18014 9828
rect 21970 9772 21980 9828
rect 22036 9772 25228 9828
rect 25284 9772 25294 9828
rect 27010 9772 27020 9828
rect 27076 9772 29596 9828
rect 29652 9772 30940 9828
rect 30996 9772 31006 9828
rect 33282 9772 33292 9828
rect 33348 9772 34188 9828
rect 34244 9772 34254 9828
rect 12124 9716 12180 9772
rect 11554 9660 11564 9716
rect 11620 9660 12180 9716
rect 14252 9716 14308 9772
rect 34412 9716 34468 9884
rect 35746 9772 35756 9828
rect 35812 9772 37324 9828
rect 37380 9772 37996 9828
rect 38052 9772 38062 9828
rect 14252 9660 14924 9716
rect 14980 9660 17836 9716
rect 17892 9660 17902 9716
rect 23650 9660 23660 9716
rect 23716 9660 27244 9716
rect 27300 9660 28364 9716
rect 28420 9660 28430 9716
rect 32610 9660 32620 9716
rect 32676 9660 33964 9716
rect 34020 9660 34030 9716
rect 34412 9660 37884 9716
rect 37940 9660 37950 9716
rect 38556 9604 38612 9884
rect 43922 9772 43932 9828
rect 43988 9772 45612 9828
rect 45668 9772 45678 9828
rect 7522 9548 7532 9604
rect 7588 9548 9660 9604
rect 9716 9548 10556 9604
rect 10612 9548 12796 9604
rect 12852 9548 12862 9604
rect 14018 9548 14028 9604
rect 14084 9548 15820 9604
rect 15876 9548 15886 9604
rect 24434 9548 24444 9604
rect 24500 9548 26796 9604
rect 26852 9548 32284 9604
rect 32340 9548 33180 9604
rect 33236 9548 33246 9604
rect 34514 9548 34524 9604
rect 34580 9548 38556 9604
rect 38612 9548 38622 9604
rect 42578 9548 42588 9604
rect 42644 9548 44156 9604
rect 44212 9548 44222 9604
rect 49200 9492 50000 9520
rect 14130 9436 14140 9492
rect 14196 9436 14364 9492
rect 14420 9436 14430 9492
rect 15250 9436 15260 9492
rect 15316 9436 15708 9492
rect 15764 9436 15774 9492
rect 27458 9436 27468 9492
rect 27524 9436 28308 9492
rect 47954 9436 47964 9492
rect 48020 9436 50000 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 28252 9380 28308 9436
rect 49200 9408 50000 9436
rect 28242 9324 28252 9380
rect 28308 9324 28318 9380
rect 32834 9324 32844 9380
rect 32900 9324 34636 9380
rect 34692 9324 34702 9380
rect 3938 9212 3948 9268
rect 4004 9212 7196 9268
rect 7252 9212 7262 9268
rect 14242 9212 14252 9268
rect 14308 9212 15484 9268
rect 15540 9212 15550 9268
rect 33170 9212 33180 9268
rect 33236 9212 35196 9268
rect 35252 9212 35262 9268
rect 17938 9100 17948 9156
rect 18004 9100 19180 9156
rect 19236 9100 19246 9156
rect 24098 9100 24108 9156
rect 24164 9100 25788 9156
rect 25844 9100 25854 9156
rect 15810 8988 15820 9044
rect 15876 8988 17836 9044
rect 17892 8988 17902 9044
rect 27570 8988 27580 9044
rect 27636 8988 27916 9044
rect 27972 8988 27982 9044
rect 36866 8876 36876 8932
rect 36932 8876 38220 8932
rect 38276 8876 38286 8932
rect 43138 8876 43148 8932
rect 43204 8876 44604 8932
rect 44660 8876 44670 8932
rect 49200 8820 50000 8848
rect 19506 8764 19516 8820
rect 19572 8764 20188 8820
rect 20244 8764 22428 8820
rect 22484 8764 23548 8820
rect 23604 8764 24668 8820
rect 24724 8764 33628 8820
rect 33684 8764 34524 8820
rect 34580 8764 34590 8820
rect 36642 8764 36652 8820
rect 36708 8764 37436 8820
rect 37492 8764 37502 8820
rect 48178 8764 48188 8820
rect 48244 8764 50000 8820
rect 49200 8736 50000 8764
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 27570 8540 27580 8596
rect 27636 8540 28084 8596
rect 42018 8540 42028 8596
rect 42084 8540 47852 8596
rect 47908 8540 47918 8596
rect 28028 8484 28084 8540
rect 28018 8428 28028 8484
rect 28084 8428 28094 8484
rect 5730 8316 5740 8372
rect 5796 8316 10500 8372
rect 13542 8316 13580 8372
rect 13636 8316 13646 8372
rect 14578 8316 14588 8372
rect 14644 8316 15148 8372
rect 15204 8316 16604 8372
rect 16660 8316 16670 8372
rect 17490 8316 17500 8372
rect 17556 8316 18172 8372
rect 18228 8316 21644 8372
rect 21700 8316 22316 8372
rect 22372 8316 22382 8372
rect 10444 8260 10500 8316
rect 17500 8260 17556 8316
rect 7634 8204 7644 8260
rect 7700 8204 10220 8260
rect 10276 8204 10286 8260
rect 10444 8204 17556 8260
rect 42802 8204 42812 8260
rect 42868 8204 45052 8260
rect 45108 8204 45118 8260
rect 45826 8204 45836 8260
rect 45892 8204 46620 8260
rect 46676 8204 47068 8260
rect 47124 8204 47134 8260
rect 0 8148 800 8176
rect 0 8092 1708 8148
rect 1764 8092 1774 8148
rect 2034 8092 2044 8148
rect 2100 8092 6860 8148
rect 6916 8092 6926 8148
rect 38994 8092 39004 8148
rect 39060 8092 40348 8148
rect 40404 8092 40414 8148
rect 0 8064 800 8092
rect 1708 8036 1764 8092
rect 42812 8036 42868 8204
rect 43026 8092 43036 8148
rect 43092 8092 43820 8148
rect 43876 8092 43886 8148
rect 1708 7980 2492 8036
rect 2548 7980 2558 8036
rect 6178 7980 6188 8036
rect 6244 7980 7420 8036
rect 7476 7980 7486 8036
rect 8418 7980 8428 8036
rect 8484 7980 9772 8036
rect 9828 7980 11004 8036
rect 11060 7980 11788 8036
rect 11844 7980 11854 8036
rect 17602 7980 17612 8036
rect 17668 7980 19516 8036
rect 19572 7980 19582 8036
rect 42130 7980 42140 8036
rect 42196 7980 42868 8036
rect 42924 7980 43708 8036
rect 43764 7980 46172 8036
rect 46228 7980 46238 8036
rect 42924 7924 42980 7980
rect 7298 7868 7308 7924
rect 7364 7868 8316 7924
rect 8372 7868 8382 7924
rect 42914 7868 42924 7924
rect 42980 7868 42990 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4162 7644 4172 7700
rect 4228 7644 8652 7700
rect 8708 7644 8718 7700
rect 11218 7644 11228 7700
rect 11284 7644 11900 7700
rect 11956 7644 11966 7700
rect 12338 7644 12348 7700
rect 12404 7644 13020 7700
rect 13076 7644 13086 7700
rect 13794 7644 13804 7700
rect 13860 7644 14588 7700
rect 14644 7644 14654 7700
rect 29810 7644 29820 7700
rect 29876 7644 38332 7700
rect 38388 7644 38892 7700
rect 38948 7644 38958 7700
rect 11900 7588 11956 7644
rect 11900 7532 12740 7588
rect 26898 7532 26908 7588
rect 26964 7532 28476 7588
rect 28532 7532 29148 7588
rect 29204 7532 29214 7588
rect 12684 7476 12740 7532
rect 12674 7420 12684 7476
rect 12740 7420 12750 7476
rect 13122 7420 13132 7476
rect 13188 7420 13692 7476
rect 13748 7420 13758 7476
rect 14018 7420 14028 7476
rect 14084 7420 17052 7476
rect 17108 7420 17118 7476
rect 20626 7420 20636 7476
rect 20692 7420 21532 7476
rect 21588 7420 22876 7476
rect 22932 7420 24220 7476
rect 24276 7420 24286 7476
rect 24658 7420 24668 7476
rect 24724 7420 26124 7476
rect 26180 7420 27244 7476
rect 27300 7420 27310 7476
rect 38210 7420 38220 7476
rect 38276 7420 42700 7476
rect 42756 7420 43596 7476
rect 43652 7420 43662 7476
rect 32498 7308 32508 7364
rect 32564 7308 33852 7364
rect 33908 7308 33918 7364
rect 24210 7196 24220 7252
rect 24276 7196 26124 7252
rect 26180 7196 26190 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 36082 6972 36092 7028
rect 36148 6972 36316 7028
rect 36372 6972 37548 7028
rect 37604 6972 37614 7028
rect 10882 6860 10892 6916
rect 10948 6860 11228 6916
rect 11284 6860 19404 6916
rect 19460 6860 19470 6916
rect 33842 6860 33852 6916
rect 33908 6860 34188 6916
rect 34244 6860 36540 6916
rect 36596 6860 43148 6916
rect 43204 6860 43214 6916
rect 8642 6748 8652 6804
rect 8708 6748 10108 6804
rect 10164 6748 11452 6804
rect 11508 6748 11518 6804
rect 13234 6748 13244 6804
rect 13300 6748 14028 6804
rect 14084 6748 14094 6804
rect 24322 6748 24332 6804
rect 24388 6748 26236 6804
rect 26292 6748 26302 6804
rect 35186 6748 35196 6804
rect 35252 6748 35980 6804
rect 36036 6748 36046 6804
rect 12898 6636 12908 6692
rect 12964 6636 13580 6692
rect 13636 6636 14924 6692
rect 14980 6636 14990 6692
rect 15922 6636 15932 6692
rect 15988 6636 16940 6692
rect 16996 6636 17006 6692
rect 17490 6636 17500 6692
rect 17556 6636 22988 6692
rect 23044 6636 23054 6692
rect 26786 6636 26796 6692
rect 26852 6636 27356 6692
rect 27412 6636 29596 6692
rect 29652 6636 30156 6692
rect 30212 6636 30716 6692
rect 30772 6636 30782 6692
rect 31378 6636 31388 6692
rect 31444 6636 32732 6692
rect 32788 6636 32798 6692
rect 43922 6636 43932 6692
rect 43988 6636 45612 6692
rect 45668 6636 45678 6692
rect 7746 6524 7756 6580
rect 7812 6524 8204 6580
rect 8260 6524 8270 6580
rect 12786 6524 12796 6580
rect 12852 6524 14252 6580
rect 14308 6524 14318 6580
rect 17042 6524 17052 6580
rect 17108 6524 20636 6580
rect 20692 6524 20702 6580
rect 26852 6524 45388 6580
rect 45444 6524 45454 6580
rect 6514 6412 6524 6468
rect 6580 6412 7308 6468
rect 7364 6412 7374 6468
rect 7522 6412 7532 6468
rect 7588 6412 7980 6468
rect 8036 6412 11116 6468
rect 11172 6412 11340 6468
rect 11396 6412 11406 6468
rect 11778 6412 11788 6468
rect 11844 6412 12236 6468
rect 12292 6412 16828 6468
rect 16884 6412 17500 6468
rect 17556 6412 17566 6468
rect 26852 6356 26908 6524
rect 27794 6412 27804 6468
rect 27860 6412 28140 6468
rect 28196 6412 29372 6468
rect 29428 6412 31164 6468
rect 31220 6412 34076 6468
rect 34132 6412 34142 6468
rect 34962 6412 34972 6468
rect 35028 6412 35420 6468
rect 35476 6412 35486 6468
rect 35858 6412 35868 6468
rect 35924 6412 35934 6468
rect 8418 6300 8428 6356
rect 8484 6300 9100 6356
rect 9156 6300 9996 6356
rect 10052 6300 13468 6356
rect 13524 6300 13534 6356
rect 20402 6300 20412 6356
rect 20468 6300 26908 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 35868 6244 35924 6412
rect 26338 6188 26348 6244
rect 26404 6188 35924 6244
rect 49200 6132 50000 6160
rect 7186 6076 7196 6132
rect 7252 6076 8428 6132
rect 8484 6076 10668 6132
rect 10724 6076 11564 6132
rect 11620 6076 11630 6132
rect 17154 6076 17164 6132
rect 17220 6076 18956 6132
rect 19012 6076 20188 6132
rect 20244 6076 20748 6132
rect 20804 6076 20814 6132
rect 22978 6076 22988 6132
rect 23044 6076 29092 6132
rect 29250 6076 29260 6132
rect 29316 6076 30716 6132
rect 30772 6076 32172 6132
rect 32228 6076 33292 6132
rect 33348 6076 33740 6132
rect 33796 6076 34748 6132
rect 34804 6076 34814 6132
rect 35634 6076 35644 6132
rect 35700 6076 36204 6132
rect 36260 6076 38892 6132
rect 38948 6076 40348 6132
rect 40404 6076 41020 6132
rect 41076 6076 41086 6132
rect 47282 6076 47292 6132
rect 47348 6076 50000 6132
rect 29036 6020 29092 6076
rect 49200 6048 50000 6076
rect 9538 5964 9548 6020
rect 9604 5964 10332 6020
rect 10388 5964 11004 6020
rect 11060 5964 11070 6020
rect 20066 5964 20076 6020
rect 20132 5964 21644 6020
rect 21700 5964 26572 6020
rect 26628 5964 27132 6020
rect 27188 5964 27198 6020
rect 29036 5964 29932 6020
rect 29988 5964 30492 6020
rect 30548 5964 32508 6020
rect 32564 5964 32574 6020
rect 20290 5852 20300 5908
rect 20356 5852 20860 5908
rect 20916 5852 24108 5908
rect 24164 5852 34636 5908
rect 34692 5852 34702 5908
rect 8642 5740 8652 5796
rect 8708 5740 9660 5796
rect 9716 5740 9726 5796
rect 33730 5740 33740 5796
rect 33796 5740 34300 5796
rect 34356 5740 34366 5796
rect 34738 5740 34748 5796
rect 34804 5740 36316 5796
rect 36372 5740 36382 5796
rect 10994 5628 11004 5684
rect 11060 5628 12012 5684
rect 12068 5628 12078 5684
rect 25330 5628 25340 5684
rect 25396 5628 27244 5684
rect 27300 5628 27310 5684
rect 29362 5628 29372 5684
rect 29428 5628 31276 5684
rect 31332 5628 33964 5684
rect 34020 5628 34030 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 20626 5404 20636 5460
rect 20692 5404 21756 5460
rect 21812 5404 21822 5460
rect 16258 5292 16268 5348
rect 16324 5292 18508 5348
rect 18564 5292 19404 5348
rect 19460 5292 20748 5348
rect 20804 5292 20814 5348
rect 20514 5180 20524 5236
rect 20580 5180 22316 5236
rect 22372 5180 22382 5236
rect 24322 5180 24332 5236
rect 24388 5180 25452 5236
rect 25508 5180 25518 5236
rect 32946 5180 32956 5236
rect 33012 5180 34860 5236
rect 34916 5180 34926 5236
rect 11218 5068 11228 5124
rect 11284 5068 12460 5124
rect 12516 5068 12526 5124
rect 19170 5068 19180 5124
rect 19236 5068 21532 5124
rect 21588 5068 21598 5124
rect 26786 5068 26796 5124
rect 26852 5068 27692 5124
rect 27748 5068 29372 5124
rect 29428 5068 29438 5124
rect 33506 5068 33516 5124
rect 33572 5068 33852 5124
rect 33908 5068 33918 5124
rect 10210 4956 10220 5012
rect 10276 4956 11340 5012
rect 11396 4956 11406 5012
rect 11890 4956 11900 5012
rect 11956 4956 12572 5012
rect 12628 4956 12638 5012
rect 20402 4956 20412 5012
rect 20468 4956 20972 5012
rect 21028 4956 22316 5012
rect 22372 4956 26348 5012
rect 26404 4956 26414 5012
rect 26898 4956 26908 5012
rect 26964 4956 28476 5012
rect 28532 4956 28542 5012
rect 30146 4956 30156 5012
rect 30212 4956 32172 5012
rect 32228 4956 32238 5012
rect 34962 4956 34972 5012
rect 35028 4956 36652 5012
rect 36708 4956 36718 5012
rect 41458 4956 41468 5012
rect 41524 4956 42700 5012
rect 42756 4956 42766 5012
rect 7970 4844 7980 4900
rect 8036 4844 10780 4900
rect 10836 4844 11004 4900
rect 11060 4844 11070 4900
rect 14802 4844 14812 4900
rect 14868 4844 15708 4900
rect 15764 4844 15774 4900
rect 22418 4844 22428 4900
rect 22484 4844 23660 4900
rect 23716 4844 24780 4900
rect 24836 4844 24846 4900
rect 28578 4844 28588 4900
rect 28644 4844 31612 4900
rect 31668 4844 31678 4900
rect 12338 4732 12348 4788
rect 12404 4732 13804 4788
rect 13860 4732 15036 4788
rect 15092 4732 15102 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 18386 4508 18396 4564
rect 18452 4508 19628 4564
rect 19684 4508 19694 4564
rect 28690 4508 28700 4564
rect 28756 4508 31276 4564
rect 31332 4508 31342 4564
rect 35522 4508 35532 4564
rect 35588 4508 37212 4564
rect 37268 4508 37278 4564
rect 9090 4396 9100 4452
rect 9156 4396 9996 4452
rect 10052 4396 10062 4452
rect 19842 4396 19852 4452
rect 19908 4396 20636 4452
rect 20692 4396 20860 4452
rect 20916 4396 20926 4452
rect 9650 4284 9660 4340
rect 9716 4284 10556 4340
rect 10612 4284 10622 4340
rect 30930 4284 30940 4340
rect 30996 4284 32396 4340
rect 32452 4284 32462 4340
rect 35634 4284 35644 4340
rect 35700 4284 37436 4340
rect 37492 4284 37502 4340
rect 7746 4172 7756 4228
rect 7812 4172 9324 4228
rect 9380 4172 9390 4228
rect 10770 4172 10780 4228
rect 10836 4172 12348 4228
rect 12404 4172 12414 4228
rect 20850 4172 20860 4228
rect 20916 4172 22092 4228
rect 22148 4172 22158 4228
rect 31602 4172 31612 4228
rect 31668 4172 32172 4228
rect 32228 4172 32238 4228
rect 33282 4172 33292 4228
rect 33348 4172 35084 4228
rect 35140 4172 35150 4228
rect 18162 3948 18172 4004
rect 18228 3948 18844 4004
rect 18900 3948 19516 4004
rect 19572 3948 19582 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 18834 3612 18844 3668
rect 18900 3612 21868 3668
rect 21924 3612 21934 3668
rect 27570 3612 27580 3668
rect 27636 3612 29372 3668
rect 29428 3612 29438 3668
rect 34290 3612 34300 3668
rect 34356 3612 36988 3668
rect 37044 3612 37054 3668
rect 37874 3612 37884 3668
rect 37940 3612 40796 3668
rect 40852 3612 40862 3668
rect 6850 3500 6860 3556
rect 6916 3500 8428 3556
rect 8484 3500 9436 3556
rect 9492 3500 9502 3556
rect 18610 3500 18620 3556
rect 18676 3500 19852 3556
rect 19908 3500 21532 3556
rect 21588 3500 21598 3556
rect 25442 3500 25452 3556
rect 25508 3500 28140 3556
rect 28196 3500 28588 3556
rect 28644 3500 28654 3556
rect 28914 3500 28924 3556
rect 28980 3500 31612 3556
rect 31668 3500 31678 3556
rect 33618 3500 33628 3556
rect 33684 3500 35420 3556
rect 35476 3500 37996 3556
rect 38052 3500 38062 3556
rect 38434 3500 38444 3556
rect 38500 3500 39788 3556
rect 39844 3500 39854 3556
rect 6402 3388 6412 3444
rect 6468 3388 7308 3444
rect 7364 3388 7374 3444
rect 9314 3388 9324 3444
rect 9380 3388 11452 3444
rect 11508 3388 11518 3444
rect 15474 3388 15484 3444
rect 15540 3388 18508 3444
rect 18564 3388 18574 3444
rect 24658 3388 24668 3444
rect 24724 3388 25900 3444
rect 25956 3388 25966 3444
rect 29586 3388 29596 3444
rect 29652 3388 33740 3444
rect 33796 3388 33806 3444
rect 41682 3388 41692 3444
rect 41748 3388 42476 3444
rect 42532 3388 42924 3444
rect 42980 3388 42990 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 44492 48412 44548 48468
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 43708 45724 43764 45780
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 19628 43260 19684 43316
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 19628 42028 19684 42084
rect 4956 41692 5012 41748
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 43708 41468 43764 41524
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 41244 40348 41300 40404
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 4956 39788 5012 39844
rect 24332 39564 24388 39620
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 24332 38332 24388 38388
rect 44492 38220 44548 38276
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 36652 37212 36708 37268
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 24332 36540 24388 36596
rect 41244 36204 41300 36260
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 36652 35756 36708 35812
rect 24332 35644 24388 35700
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 8764 33516 8820 33572
rect 8764 32732 8820 32788
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 13692 31836 13748 31892
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 16156 29484 16212 29540
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 20188 28364 20244 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 16156 27916 16212 27972
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 20188 27132 20244 27188
rect 13692 26684 13748 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 20188 23436 20244 23492
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 43036 22204 43092 22260
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 13580 21420 13636 21476
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 23996 20524 24052 20580
rect 43260 20524 43316 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 44268 18732 44324 18788
rect 24108 18396 24164 18452
rect 44828 18396 44884 18452
rect 14140 18172 14196 18228
rect 23884 18172 23940 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 23996 17724 24052 17780
rect 23884 17388 23940 17444
rect 44828 17276 44884 17332
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 24108 16716 24164 16772
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 44268 16492 44324 16548
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 43036 16380 43092 16436
rect 43372 16156 43428 16212
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 25564 15148 25620 15204
rect 43372 15036 43428 15092
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 44268 14588 44324 14644
rect 25564 14364 25620 14420
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 43260 13692 43316 13748
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 14140 9436 14196 9492
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 13580 8316 13636 8372
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 44492 48468 44548 48478
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 19628 43316 19684 43326
rect 19628 42084 19684 43260
rect 19628 42018 19684 42028
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4956 41748 5012 41758
rect 4956 39844 5012 41692
rect 4956 39778 5012 39788
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 19808 39228 20128 40740
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 43708 45780 43764 45790
rect 43708 41524 43764 45724
rect 43708 41458 43764 41468
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 24332 39620 24388 39630
rect 24332 38388 24388 39564
rect 24332 38322 24388 38332
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 35168 36876 35488 38388
rect 41244 40404 41300 40414
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 24332 36596 24388 36606
rect 24332 35700 24388 36540
rect 24332 35634 24388 35644
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 8764 33572 8820 33582
rect 8764 32788 8820 33516
rect 8764 32722 8820 32732
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 13692 31892 13748 31902
rect 13692 26740 13748 31836
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 16156 29540 16212 29550
rect 16156 27972 16212 29484
rect 16156 27906 16212 27916
rect 19808 28252 20128 29764
rect 35168 35308 35488 36820
rect 36652 37268 36708 37278
rect 36652 35812 36708 37212
rect 41244 36260 41300 40348
rect 44492 38276 44548 48412
rect 44492 38210 44548 38220
rect 41244 36194 41300 36204
rect 36652 35746 36708 35756
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 13692 26674 13748 26684
rect 19808 26684 20128 28196
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 20188 28420 20244 28430
rect 20188 27188 20244 28364
rect 20188 23492 20244 27132
rect 20188 23426 20244 23436
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 13580 21476 13636 21486
rect 13580 8372 13636 21420
rect 19808 20412 20128 21924
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 14140 18228 14196 18238
rect 14140 9492 14196 18172
rect 14140 9426 14196 9436
rect 19808 17276 20128 18788
rect 23996 20580 24052 20590
rect 23884 18228 23940 18238
rect 23884 17444 23940 18172
rect 23996 17780 24052 20524
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 23996 17714 24052 17724
rect 24108 18452 24164 18462
rect 23884 17378 23940 17388
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 24108 16772 24164 18396
rect 24108 16706 24164 16716
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 25564 15204 25620 15214
rect 25564 14420 25620 15148
rect 25564 14354 25620 14364
rect 35168 14924 35488 16436
rect 43036 22260 43092 22270
rect 43036 16436 43092 22204
rect 43036 16370 43092 16380
rect 43260 20580 43316 20590
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 13580 8306 13636 8316
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 13356 35488 14868
rect 43260 13748 43316 20524
rect 44268 18788 44324 18798
rect 44268 16548 44324 18732
rect 44828 18452 44884 18462
rect 44828 17332 44884 18396
rect 44828 17266 44884 17276
rect 43372 16212 43428 16222
rect 43372 15092 43428 16156
rect 43372 15026 43428 15036
rect 44268 14644 44324 16492
rect 44268 14578 44324 14588
rect 43260 13682 43316 13692
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0895_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24864 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0896_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0897_
timestamp 1698431365
transform 1 0 22960 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0898_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23072 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0899_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23408 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0900_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23520 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0901_
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0902_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45360 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0903_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47152 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0904_
timestamp 1698431365
transform 1 0 47712 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0905_
timestamp 1698431365
transform 1 0 42672 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0906_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44800 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0907_
timestamp 1698431365
transform -1 0 42560 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0908_
timestamp 1698431365
transform 1 0 42784 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0909_
timestamp 1698431365
transform -1 0 45360 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0910_
timestamp 1698431365
transform -1 0 42560 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0911_
timestamp 1698431365
transform 1 0 40880 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0912_
timestamp 1698431365
transform 1 0 42672 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0913_
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0914_
timestamp 1698431365
transform -1 0 43904 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0915_
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0916_
timestamp 1698431365
transform 1 0 42112 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0917_
timestamp 1698431365
transform 1 0 47600 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0918_
timestamp 1698431365
transform -1 0 34832 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0919_
timestamp 1698431365
transform 1 0 34272 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0920_
timestamp 1698431365
transform -1 0 26656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0921_
timestamp 1698431365
transform 1 0 26656 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0922_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33600 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0923_
timestamp 1698431365
transform -1 0 32256 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0924_
timestamp 1698431365
transform -1 0 33376 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0925_
timestamp 1698431365
transform -1 0 32704 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0926_
timestamp 1698431365
transform -1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0927_
timestamp 1698431365
transform -1 0 33152 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0928_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34048 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0929_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 33264 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0930_
timestamp 1698431365
transform -1 0 43904 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0931_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43344 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0932_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44464 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0933_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45584 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0934_
timestamp 1698431365
transform -1 0 44016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _0935_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43792 0 1 25088
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0936_
timestamp 1698431365
transform -1 0 44464 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0937_
timestamp 1698431365
transform 1 0 45472 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0938_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46480 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0939_
timestamp 1698431365
transform -1 0 47264 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0940_
timestamp 1698431365
transform -1 0 44352 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0941_
timestamp 1698431365
transform -1 0 42112 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0942_
timestamp 1698431365
transform -1 0 41664 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0943_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42560 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0944_
timestamp 1698431365
transform 1 0 38192 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0945_
timestamp 1698431365
transform 1 0 41552 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0946_
timestamp 1698431365
transform -1 0 43680 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0947_
timestamp 1698431365
transform -1 0 45472 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0948_
timestamp 1698431365
transform 1 0 44464 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0949_
timestamp 1698431365
transform -1 0 45024 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0950_
timestamp 1698431365
transform 1 0 45696 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0951_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45472 0 -1 21952
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0952_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43344 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0953_
timestamp 1698431365
transform -1 0 43232 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0954_
timestamp 1698431365
transform 1 0 41776 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0955_
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0956_
timestamp 1698431365
transform -1 0 40992 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0957_
timestamp 1698431365
transform 1 0 9856 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0958_
timestamp 1698431365
transform -1 0 14000 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0959_
timestamp 1698431365
transform -1 0 7952 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0960_
timestamp 1698431365
transform -1 0 10640 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0961_
timestamp 1698431365
transform 1 0 11424 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0962_
timestamp 1698431365
transform -1 0 9856 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0963_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8288 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0964_
timestamp 1698431365
transform 1 0 7168 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0965_
timestamp 1698431365
transform 1 0 8176 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0966_
timestamp 1698431365
transform 1 0 10640 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0967_
timestamp 1698431365
transform -1 0 9184 0 -1 36064
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0968_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11200 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0969_
timestamp 1698431365
transform 1 0 17808 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0970_
timestamp 1698431365
transform 1 0 18144 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _0971_
timestamp 1698431365
transform -1 0 21168 0 -1 31360
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _0972_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0973_
timestamp 1698431365
transform -1 0 17696 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0974_
timestamp 1698431365
transform -1 0 19824 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0975_
timestamp 1698431365
transform -1 0 15232 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  _0976_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 28224
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0977_
timestamp 1698431365
transform -1 0 18256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0978_
timestamp 1698431365
transform -1 0 13888 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0979_
timestamp 1698431365
transform 1 0 14336 0 1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0980_
timestamp 1698431365
transform -1 0 14000 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0981_
timestamp 1698431365
transform 1 0 13552 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0982_
timestamp 1698431365
transform -1 0 14224 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0983_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14224 0 1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0984_
timestamp 1698431365
transform -1 0 13104 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0985_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11984 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0986_
timestamp 1698431365
transform -1 0 17920 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0987_
timestamp 1698431365
transform -1 0 17808 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0988_
timestamp 1698431365
transform -1 0 16912 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0989_
timestamp 1698431365
transform -1 0 16352 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0990_
timestamp 1698431365
transform 1 0 14896 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0991_
timestamp 1698431365
transform -1 0 15680 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0992_
timestamp 1698431365
transform 1 0 15344 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0993_
timestamp 1698431365
transform -1 0 15680 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0994_
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0995_
timestamp 1698431365
transform -1 0 16128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0996_
timestamp 1698431365
transform 1 0 14672 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0997_
timestamp 1698431365
transform 1 0 13664 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0998_
timestamp 1698431365
transform 1 0 14224 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0999_
timestamp 1698431365
transform 1 0 6272 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1000_
timestamp 1698431365
transform 1 0 6832 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1001_
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1002_
timestamp 1698431365
transform 1 0 7056 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1003_
timestamp 1698431365
transform 1 0 7392 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1004_
timestamp 1698431365
transform 1 0 7056 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1005_
timestamp 1698431365
transform 1 0 7056 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1006_
timestamp 1698431365
transform -1 0 4928 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1007_
timestamp 1698431365
transform 1 0 6944 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1008_
timestamp 1698431365
transform 1 0 6832 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1009_
timestamp 1698431365
transform 1 0 10528 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1010_
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1011_
timestamp 1698431365
transform 1 0 6048 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1012_
timestamp 1698431365
transform -1 0 6720 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1013_
timestamp 1698431365
transform -1 0 12880 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1014_
timestamp 1698431365
transform 1 0 9856 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1015_
timestamp 1698431365
transform 1 0 12432 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1016_
timestamp 1698431365
transform 1 0 10080 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1017_
timestamp 1698431365
transform -1 0 9408 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1018_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1019_
timestamp 1698431365
transform 1 0 11200 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1020_
timestamp 1698431365
transform -1 0 12880 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1021_
timestamp 1698431365
transform -1 0 13776 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1022_
timestamp 1698431365
transform -1 0 12096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1023_
timestamp 1698431365
transform 1 0 10976 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1024_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12096 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1025_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10752 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1026_
timestamp 1698431365
transform -1 0 14448 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1027_
timestamp 1698431365
transform 1 0 11312 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1028_
timestamp 1698431365
transform -1 0 9520 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1029_
timestamp 1698431365
transform -1 0 10080 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1030_
timestamp 1698431365
transform -1 0 8848 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1031_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1032_
timestamp 1698431365
transform -1 0 10640 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1033_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14224 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1034_
timestamp 1698431365
transform -1 0 15680 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1035_
timestamp 1698431365
transform 1 0 14112 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1036_
timestamp 1698431365
transform -1 0 47600 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1037_
timestamp 1698431365
transform 1 0 44688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1038_
timestamp 1698431365
transform 1 0 42112 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1039_
timestamp 1698431365
transform 1 0 43680 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1040_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44464 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1041_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40992 0 1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1042_
timestamp 1698431365
transform 1 0 41552 0 -1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1043_
timestamp 1698431365
transform -1 0 33488 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1044_
timestamp 1698431365
transform 1 0 34720 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1045_
timestamp 1698431365
transform -1 0 33376 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1046_
timestamp 1698431365
transform -1 0 37744 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1047_
timestamp 1698431365
transform -1 0 34608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1048_
timestamp 1698431365
transform 1 0 34720 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1049_
timestamp 1698431365
transform 1 0 36400 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1050_
timestamp 1698431365
transform -1 0 38080 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1051_
timestamp 1698431365
transform -1 0 38304 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1052_
timestamp 1698431365
transform 1 0 36736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1053_
timestamp 1698431365
transform 1 0 36624 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1054_
timestamp 1698431365
transform -1 0 37408 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1055_
timestamp 1698431365
transform 1 0 31808 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1056_
timestamp 1698431365
transform -1 0 28224 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1057_
timestamp 1698431365
transform 1 0 27440 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1058_
timestamp 1698431365
transform -1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1059_
timestamp 1698431365
transform -1 0 27216 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1060_
timestamp 1698431365
transform 1 0 26544 0 -1 10976
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1061_
timestamp 1698431365
transform -1 0 28112 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1062_
timestamp 1698431365
transform -1 0 26544 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1063_
timestamp 1698431365
transform 1 0 26656 0 -1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1064_
timestamp 1698431365
transform -1 0 33712 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1065_
timestamp 1698431365
transform -1 0 32144 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1066_
timestamp 1698431365
transform -1 0 31024 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1067_
timestamp 1698431365
transform 1 0 30912 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1068_
timestamp 1698431365
transform -1 0 24864 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1069_
timestamp 1698431365
transform -1 0 22960 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1070_
timestamp 1698431365
transform -1 0 18704 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1071_
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1072_
timestamp 1698431365
transform -1 0 29008 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1073_
timestamp 1698431365
transform -1 0 31248 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1074_
timestamp 1698431365
transform 1 0 23744 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1075_
timestamp 1698431365
transform 1 0 24976 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1076_
timestamp 1698431365
transform -1 0 19600 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1077_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24752 0 1 12544
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1078_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28896 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1079_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29232 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1080_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32032 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1081_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1082_
timestamp 1698431365
transform 1 0 38640 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1083_
timestamp 1698431365
transform 1 0 35728 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1084_
timestamp 1698431365
transform 1 0 31920 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1085_
timestamp 1698431365
transform 1 0 28672 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1086_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29344 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1087_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1088_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28784 0 -1 12544
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1089_
timestamp 1698431365
transform 1 0 30352 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1090_
timestamp 1698431365
transform 1 0 31584 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1091_
timestamp 1698431365
transform 1 0 35840 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1092_
timestamp 1698431365
transform 1 0 37072 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1093_
timestamp 1698431365
transform -1 0 7616 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1094_
timestamp 1698431365
transform 1 0 10640 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1095_
timestamp 1698431365
transform 1 0 10864 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1096_
timestamp 1698431365
transform 1 0 11312 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1097_
timestamp 1698431365
transform -1 0 5488 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1098_
timestamp 1698431365
transform 1 0 8960 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1099_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9968 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1100_
timestamp 1698431365
transform 1 0 11088 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1101_
timestamp 1698431365
transform 1 0 11536 0 -1 32928
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1102_
timestamp 1698431365
transform -1 0 14560 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1103_
timestamp 1698431365
transform 1 0 35840 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1104_
timestamp 1698431365
transform 1 0 37632 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1105_
timestamp 1698431365
transform -1 0 37520 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1106_
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1107_
timestamp 1698431365
transform -1 0 33600 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1108_
timestamp 1698431365
transform -1 0 30464 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1109_
timestamp 1698431365
transform 1 0 10192 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1110_
timestamp 1698431365
transform 1 0 10640 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1111_
timestamp 1698431365
transform -1 0 12768 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1112_
timestamp 1698431365
transform -1 0 10640 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1113_
timestamp 1698431365
transform 1 0 14224 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1114_
timestamp 1698431365
transform -1 0 27328 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1115_
timestamp 1698431365
transform -1 0 21840 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1116_
timestamp 1698431365
transform 1 0 20160 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1117_
timestamp 1698431365
transform -1 0 14224 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1118_
timestamp 1698431365
transform 1 0 12208 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1119_
timestamp 1698431365
transform -1 0 12096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1120_
timestamp 1698431365
transform 1 0 11312 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1121_
timestamp 1698431365
transform -1 0 12208 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1122_
timestamp 1698431365
transform 1 0 6608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1123_
timestamp 1698431365
transform -1 0 23968 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1124_
timestamp 1698431365
transform -1 0 11984 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1125_
timestamp 1698431365
transform 1 0 7952 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1126_
timestamp 1698431365
transform 1 0 7056 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1127_
timestamp 1698431365
transform -1 0 11312 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1128_
timestamp 1698431365
transform 1 0 6720 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1129_
timestamp 1698431365
transform 1 0 11312 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1130_
timestamp 1698431365
transform 1 0 8064 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1131_
timestamp 1698431365
transform 1 0 7168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1132_
timestamp 1698431365
transform 1 0 6720 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1133_
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1134_
timestamp 1698431365
transform 1 0 7840 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1135_
timestamp 1698431365
transform 1 0 9296 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1136_
timestamp 1698431365
transform 1 0 10640 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1137_
timestamp 1698431365
transform 1 0 9744 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1138_
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1139_
timestamp 1698431365
transform 1 0 16576 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1140_
timestamp 1698431365
transform 1 0 12208 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1141_
timestamp 1698431365
transform 1 0 10528 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1142_
timestamp 1698431365
transform 1 0 12096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1143_
timestamp 1698431365
transform 1 0 13440 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1144_
timestamp 1698431365
transform 1 0 12544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1145_
timestamp 1698431365
transform -1 0 27664 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1146_
timestamp 1698431365
transform 1 0 19824 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1147_
timestamp 1698431365
transform -1 0 19824 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1148_
timestamp 1698431365
transform -1 0 21840 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1149_
timestamp 1698431365
transform 1 0 20048 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1150_
timestamp 1698431365
transform 1 0 19376 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1151_
timestamp 1698431365
transform -1 0 21616 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1152_
timestamp 1698431365
transform -1 0 24304 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1153_
timestamp 1698431365
transform -1 0 22624 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1154_
timestamp 1698431365
transform -1 0 21168 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1155_
timestamp 1698431365
transform 1 0 23184 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1156_
timestamp 1698431365
transform -1 0 24864 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1157_
timestamp 1698431365
transform -1 0 30688 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1158_
timestamp 1698431365
transform 1 0 25984 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1159_
timestamp 1698431365
transform 1 0 23632 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1160_
timestamp 1698431365
transform 1 0 26320 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1161_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1162_
timestamp 1698431365
transform 1 0 27664 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1163_
timestamp 1698431365
transform -1 0 28224 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1164_
timestamp 1698431365
transform 1 0 27216 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1165_
timestamp 1698431365
transform 1 0 28560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1166_
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1167_
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1168_
timestamp 1698431365
transform 1 0 30016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1169_
timestamp 1698431365
transform -1 0 31584 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1170_
timestamp 1698431365
transform 1 0 30800 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1171_
timestamp 1698431365
transform 1 0 33152 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1172_
timestamp 1698431365
transform 1 0 33712 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1173_
timestamp 1698431365
transform -1 0 34496 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1174_
timestamp 1698431365
transform 1 0 33488 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1175_
timestamp 1698431365
transform -1 0 35728 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1176_
timestamp 1698431365
transform 1 0 35728 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1177_
timestamp 1698431365
transform 1 0 34496 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1178_
timestamp 1698431365
transform 1 0 47376 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1179_
timestamp 1698431365
transform -1 0 45696 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1180_
timestamp 1698431365
transform 1 0 41328 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1181_
timestamp 1698431365
transform 1 0 45696 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1182_
timestamp 1698431365
transform 1 0 42560 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1183_
timestamp 1698431365
transform 1 0 41776 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1184_
timestamp 1698431365
transform 1 0 41888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1185_
timestamp 1698431365
transform -1 0 44128 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1186_
timestamp 1698431365
transform 1 0 42336 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1187_
timestamp 1698431365
transform -1 0 45136 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1188_
timestamp 1698431365
transform 1 0 42784 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1189_
timestamp 1698431365
transform 1 0 44576 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1190_
timestamp 1698431365
transform 1 0 45584 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1191_
timestamp 1698431365
transform -1 0 44352 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1192_
timestamp 1698431365
transform -1 0 48160 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1193_
timestamp 1698431365
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1194_
timestamp 1698431365
transform -1 0 48048 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1195_
timestamp 1698431365
transform -1 0 48384 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1196_
timestamp 1698431365
transform -1 0 47488 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1197_
timestamp 1698431365
transform 1 0 46480 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1198_
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1199_
timestamp 1698431365
transform 1 0 46480 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1200_
timestamp 1698431365
transform 1 0 46592 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1201_
timestamp 1698431365
transform 1 0 44688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1202_
timestamp 1698431365
transform 1 0 46928 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1203_
timestamp 1698431365
transform 1 0 46032 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1204_
timestamp 1698431365
transform 1 0 45696 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1205_
timestamp 1698431365
transform -1 0 46480 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1206_
timestamp 1698431365
transform 1 0 43568 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1207_
timestamp 1698431365
transform 1 0 47040 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1208_
timestamp 1698431365
transform 1 0 46144 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1209_
timestamp 1698431365
transform 1 0 44128 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1210_
timestamp 1698431365
transform 1 0 46256 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1211_
timestamp 1698431365
transform 1 0 44576 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1212_
timestamp 1698431365
transform -1 0 28000 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1213_
timestamp 1698431365
transform -1 0 15008 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1214_
timestamp 1698431365
transform -1 0 4368 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1215_
timestamp 1698431365
transform 1 0 5600 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1216_
timestamp 1698431365
transform -1 0 5936 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1217_
timestamp 1698431365
transform -1 0 8512 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1218_
timestamp 1698431365
transform -1 0 5488 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1219_
timestamp 1698431365
transform 1 0 6944 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1220_
timestamp 1698431365
transform 1 0 6272 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1221_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6832 0 1 37632
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1222_
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1223_
timestamp 1698431365
transform -1 0 7728 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1224_
timestamp 1698431365
transform -1 0 8064 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1225_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7056 0 1 28224
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1226_
timestamp 1698431365
transform -1 0 16688 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1227_
timestamp 1698431365
transform -1 0 10416 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1228_
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1229_
timestamp 1698431365
transform -1 0 9856 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1230_
timestamp 1698431365
transform 1 0 10416 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1231_
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1232_
timestamp 1698431365
transform -1 0 6496 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1233_
timestamp 1698431365
transform 1 0 6608 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1234_
timestamp 1698431365
transform -1 0 7392 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1235_
timestamp 1698431365
transform 1 0 8400 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1236_
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1237_
timestamp 1698431365
transform -1 0 8512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1238_
timestamp 1698431365
transform -1 0 9072 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1239_
timestamp 1698431365
transform -1 0 12208 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1240_
timestamp 1698431365
transform -1 0 11984 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1241_
timestamp 1698431365
transform -1 0 14112 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1242_
timestamp 1698431365
transform 1 0 7056 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1243_
timestamp 1698431365
transform 1 0 9520 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1244_
timestamp 1698431365
transform -1 0 12432 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1245_
timestamp 1698431365
transform 1 0 8400 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1246_
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1247_
timestamp 1698431365
transform 1 0 10192 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1248_
timestamp 1698431365
transform 1 0 9632 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1249_
timestamp 1698431365
transform 1 0 7728 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1250_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9408 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1251_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9968 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1252_
timestamp 1698431365
transform 1 0 10304 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1253_
timestamp 1698431365
transform -1 0 17360 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1254_
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1255_
timestamp 1698431365
transform 1 0 16688 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1256_
timestamp 1698431365
transform 1 0 14448 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1257_
timestamp 1698431365
transform -1 0 16352 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1258_
timestamp 1698431365
transform 1 0 15456 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1259_
timestamp 1698431365
transform 1 0 17360 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1260_
timestamp 1698431365
transform 1 0 16352 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1261_
timestamp 1698431365
transform -1 0 18144 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1262_
timestamp 1698431365
transform 1 0 27776 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1263_
timestamp 1698431365
transform 1 0 26880 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1264_
timestamp 1698431365
transform -1 0 25536 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1265_
timestamp 1698431365
transform 1 0 22624 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1266_
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1267_
timestamp 1698431365
transform -1 0 23968 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1268_
timestamp 1698431365
transform 1 0 22400 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1269_
timestamp 1698431365
transform 1 0 22512 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1270_
timestamp 1698431365
transform -1 0 24416 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1271_
timestamp 1698431365
transform -1 0 26992 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1272_
timestamp 1698431365
transform -1 0 32704 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1273_
timestamp 1698431365
transform -1 0 31920 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1274_
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1275_
timestamp 1698431365
transform -1 0 28112 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1276_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1277_
timestamp 1698431365
transform -1 0 34272 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1278_
timestamp 1698431365
transform -1 0 34048 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1279_
timestamp 1698431365
transform -1 0 34944 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1280_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27888 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1281_
timestamp 1698431365
transform 1 0 29680 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1282_
timestamp 1698431365
transform 1 0 23520 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1283_
timestamp 1698431365
transform 1 0 24976 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1284_
timestamp 1698431365
transform 1 0 26880 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1285_
timestamp 1698431365
transform 1 0 27440 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1286_
timestamp 1698431365
transform 1 0 29792 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1287_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1288_
timestamp 1698431365
transform -1 0 45360 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1289_
timestamp 1698431365
transform -1 0 37520 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1290_
timestamp 1698431365
transform 1 0 37296 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1291_
timestamp 1698431365
transform -1 0 38304 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1292_
timestamp 1698431365
transform 1 0 38304 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1293_
timestamp 1698431365
transform -1 0 41776 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1294_
timestamp 1698431365
transform -1 0 36624 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1295_
timestamp 1698431365
transform -1 0 41776 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1296_
timestamp 1698431365
transform 1 0 37744 0 1 25088
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1297_
timestamp 1698431365
transform -1 0 39088 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1298_
timestamp 1698431365
transform -1 0 38528 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1299_
timestamp 1698431365
transform -1 0 40208 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1300_
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1301_
timestamp 1698431365
transform 1 0 37520 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1302_
timestamp 1698431365
transform -1 0 39536 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1303_
timestamp 1698431365
transform 1 0 38864 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1304_
timestamp 1698431365
transform 1 0 39536 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1305_
timestamp 1698431365
transform 1 0 37968 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1306_
timestamp 1698431365
transform -1 0 42672 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1307_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1308_
timestamp 1698431365
transform 1 0 37296 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1309_
timestamp 1698431365
transform 1 0 37744 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1310_
timestamp 1698431365
transform 1 0 39872 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1311_
timestamp 1698431365
transform -1 0 39760 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1312_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1313_
timestamp 1698431365
transform 1 0 39088 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1314_
timestamp 1698431365
transform -1 0 39648 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1315_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38528 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1316_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42000 0 1 26656
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1317_
timestamp 1698431365
transform -1 0 38976 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1318_
timestamp 1698431365
transform -1 0 37520 0 -1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1319_
timestamp 1698431365
transform 1 0 35168 0 -1 26656
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1320_
timestamp 1698431365
transform -1 0 26768 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1321_
timestamp 1698431365
transform 1 0 22960 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1322_
timestamp 1698431365
transform 1 0 23744 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1323_
timestamp 1698431365
transform 1 0 23968 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1324_
timestamp 1698431365
transform -1 0 25200 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1325_
timestamp 1698431365
transform 1 0 23632 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1326_
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1327_
timestamp 1698431365
transform 1 0 25536 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1328_
timestamp 1698431365
transform 1 0 24528 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1329_
timestamp 1698431365
transform 1 0 23744 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1330_
timestamp 1698431365
transform -1 0 26768 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1331_
timestamp 1698431365
transform 1 0 25536 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1332_
timestamp 1698431365
transform -1 0 24864 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1333_
timestamp 1698431365
transform -1 0 24416 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1334_
timestamp 1698431365
transform 1 0 26880 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1335_
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1336_
timestamp 1698431365
transform -1 0 27104 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1337_
timestamp 1698431365
transform -1 0 25536 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1338_
timestamp 1698431365
transform 1 0 25648 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1339_
timestamp 1698431365
transform -1 0 27440 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1340_
timestamp 1698431365
transform -1 0 24192 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1341_
timestamp 1698431365
transform 1 0 27440 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1342_
timestamp 1698431365
transform 1 0 28560 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1343_
timestamp 1698431365
transform -1 0 27776 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1344_
timestamp 1698431365
transform 1 0 26656 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1345_
timestamp 1698431365
transform 1 0 26432 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1346_
timestamp 1698431365
transform 1 0 27664 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1347_
timestamp 1698431365
transform -1 0 25312 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1348_
timestamp 1698431365
transform -1 0 23744 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1349_
timestamp 1698431365
transform -1 0 26432 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1350_
timestamp 1698431365
transform 1 0 25312 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1351_
timestamp 1698431365
transform 1 0 23744 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1352_
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1353_
timestamp 1698431365
transform -1 0 23744 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1354_
timestamp 1698431365
transform -1 0 23744 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1355_
timestamp 1698431365
transform -1 0 23632 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1356_
timestamp 1698431365
transform -1 0 23184 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1357_
timestamp 1698431365
transform 1 0 22288 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1358_
timestamp 1698431365
transform 1 0 21504 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1359_
timestamp 1698431365
transform 1 0 22624 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1360_
timestamp 1698431365
transform -1 0 19376 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1361_
timestamp 1698431365
transform 1 0 18144 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1362_
timestamp 1698431365
transform -1 0 21616 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1363_
timestamp 1698431365
transform 1 0 20272 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1364_
timestamp 1698431365
transform 1 0 19152 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1365_
timestamp 1698431365
transform -1 0 20496 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1366_
timestamp 1698431365
transform -1 0 18704 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1367_
timestamp 1698431365
transform -1 0 17024 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1368_
timestamp 1698431365
transform 1 0 19600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1369_
timestamp 1698431365
transform -1 0 20496 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1370_
timestamp 1698431365
transform 1 0 19264 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1371_
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1372_
timestamp 1698431365
transform -1 0 17920 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1373_
timestamp 1698431365
transform 1 0 20496 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1374_
timestamp 1698431365
transform -1 0 21616 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1375_
timestamp 1698431365
transform -1 0 22512 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1376_
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1377_
timestamp 1698431365
transform 1 0 18592 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1378_
timestamp 1698431365
transform -1 0 24416 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1379_
timestamp 1698431365
transform -1 0 20384 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1380_
timestamp 1698431365
transform -1 0 28000 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1381_
timestamp 1698431365
transform 1 0 25760 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1382_
timestamp 1698431365
transform 1 0 23184 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1383_
timestamp 1698431365
transform -1 0 25536 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1384_
timestamp 1698431365
transform 1 0 23632 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1385_
timestamp 1698431365
transform -1 0 23408 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1386_
timestamp 1698431365
transform 1 0 23632 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1387_
timestamp 1698431365
transform 1 0 19600 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1388_
timestamp 1698431365
transform 1 0 19936 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1389_
timestamp 1698431365
transform 1 0 25312 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1390_
timestamp 1698431365
transform 1 0 26656 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1391_
timestamp 1698431365
transform -1 0 23072 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1392_
timestamp 1698431365
transform 1 0 23072 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1393_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21392 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1394_
timestamp 1698431365
transform -1 0 20048 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1395_
timestamp 1698431365
transform -1 0 19488 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1396_
timestamp 1698431365
transform 1 0 22064 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1397_
timestamp 1698431365
transform -1 0 26096 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1398_
timestamp 1698431365
transform 1 0 21616 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1399_
timestamp 1698431365
transform 1 0 22848 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1400_
timestamp 1698431365
transform -1 0 18368 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1401_
timestamp 1698431365
transform -1 0 20048 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1402_
timestamp 1698431365
transform -1 0 20160 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1403_
timestamp 1698431365
transform 1 0 19264 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1404_
timestamp 1698431365
transform 1 0 33040 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1405_
timestamp 1698431365
transform -1 0 35056 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1406_
timestamp 1698431365
transform -1 0 42000 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1407_
timestamp 1698431365
transform -1 0 36288 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1408_
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1409_
timestamp 1698431365
transform -1 0 45360 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1410_
timestamp 1698431365
transform -1 0 42896 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1411_
timestamp 1698431365
transform -1 0 41664 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1412_
timestamp 1698431365
transform -1 0 15456 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1413_
timestamp 1698431365
transform 1 0 16128 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1414_
timestamp 1698431365
transform 1 0 15232 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1415_
timestamp 1698431365
transform -1 0 18256 0 1 25088
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1416_
timestamp 1698431365
transform -1 0 18256 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1417_
timestamp 1698431365
transform 1 0 15008 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1418_
timestamp 1698431365
transform -1 0 16128 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1419_
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1420_
timestamp 1698431365
transform -1 0 16912 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1421_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11424 0 1 34496
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1422_
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1423_
timestamp 1698431365
transform -1 0 11200 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1424_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11536 0 -1 34496
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1425_
timestamp 1698431365
transform 1 0 14896 0 -1 25088
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1426_
timestamp 1698431365
transform 1 0 15680 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1427_
timestamp 1698431365
transform -1 0 16800 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1428_
timestamp 1698431365
transform 1 0 11984 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1429_
timestamp 1698431365
transform 1 0 12544 0 -1 12544
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1430_
timestamp 1698431365
transform -1 0 15232 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1431_
timestamp 1698431365
transform 1 0 8624 0 1 15680
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1432_
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1433_
timestamp 1698431365
transform -1 0 10416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1434_
timestamp 1698431365
transform -1 0 9072 0 -1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1435_
timestamp 1698431365
transform 1 0 7504 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1436_
timestamp 1698431365
transform -1 0 11872 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1437_
timestamp 1698431365
transform 1 0 11088 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1438_
timestamp 1698431365
transform -1 0 11088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1439_
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1440_
timestamp 1698431365
transform 1 0 17360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1441_
timestamp 1698431365
transform 1 0 17584 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1442_
timestamp 1698431365
transform 1 0 14336 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1443_
timestamp 1698431365
transform 1 0 15344 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1444_
timestamp 1698431365
transform 1 0 15680 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1445_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15232 0 1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1446_
timestamp 1698431365
transform 1 0 37632 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1447_
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1448_
timestamp 1698431365
transform 1 0 34944 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1449_
timestamp 1698431365
transform 1 0 37296 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1450_
timestamp 1698431365
transform 1 0 33600 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1451_
timestamp 1698431365
transform 1 0 33712 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1452_
timestamp 1698431365
transform -1 0 35392 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1453_
timestamp 1698431365
transform 1 0 27216 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1454_
timestamp 1698431365
transform 1 0 27776 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1455_
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1456_
timestamp 1698431365
transform 1 0 24080 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1457_
timestamp 1698431365
transform 1 0 25424 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1458_
timestamp 1698431365
transform 1 0 26096 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1459_
timestamp 1698431365
transform 1 0 26992 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1460_
timestamp 1698431365
transform 1 0 32704 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1461_
timestamp 1698431365
transform -1 0 27664 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1462_
timestamp 1698431365
transform -1 0 28112 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1463_
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1464_
timestamp 1698431365
transform 1 0 26656 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1465_
timestamp 1698431365
transform 1 0 34832 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1466_
timestamp 1698431365
transform 1 0 35392 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1467_
timestamp 1698431365
transform 1 0 33936 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1468_
timestamp 1698431365
transform 1 0 33040 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1469_
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1470_
timestamp 1698431365
transform -1 0 45360 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1471_
timestamp 1698431365
transform -1 0 43904 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1472_
timestamp 1698431365
transform -1 0 43680 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1473_
timestamp 1698431365
transform 1 0 37408 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1474_
timestamp 1698431365
transform 1 0 37856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1475_
timestamp 1698431365
transform -1 0 43680 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1476_
timestamp 1698431365
transform -1 0 40320 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1477_
timestamp 1698431365
transform 1 0 38640 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1478_
timestamp 1698431365
transform -1 0 42000 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1479_
timestamp 1698431365
transform 1 0 42112 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1480_
timestamp 1698431365
transform -1 0 42560 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1481_
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1482_
timestamp 1698431365
transform 1 0 40208 0 1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1483_
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1484_
timestamp 1698431365
transform -1 0 37856 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1485_
timestamp 1698431365
transform -1 0 32032 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1486_
timestamp 1698431365
transform 1 0 33600 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1487_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32816 0 1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1488_
timestamp 1698431365
transform -1 0 31584 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1489_
timestamp 1698431365
transform -1 0 30688 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1490_
timestamp 1698431365
transform -1 0 29568 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1491_
timestamp 1698431365
transform 1 0 29568 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1492_
timestamp 1698431365
transform 1 0 26432 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1493_
timestamp 1698431365
transform -1 0 28000 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1494_
timestamp 1698431365
transform -1 0 31360 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1495_
timestamp 1698431365
transform -1 0 29904 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1496_
timestamp 1698431365
transform 1 0 29904 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1497_
timestamp 1698431365
transform 1 0 28672 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1498_
timestamp 1698431365
transform -1 0 29904 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1499_
timestamp 1698431365
transform 1 0 30464 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1500_
timestamp 1698431365
transform -1 0 32256 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1501_
timestamp 1698431365
transform -1 0 30912 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1502_
timestamp 1698431365
transform 1 0 30800 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1503_
timestamp 1698431365
transform 1 0 34160 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1504_
timestamp 1698431365
transform 1 0 33600 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1505_
timestamp 1698431365
transform 1 0 34720 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1506_
timestamp 1698431365
transform -1 0 36064 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1507_
timestamp 1698431365
transform -1 0 5152 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1508_
timestamp 1698431365
transform -1 0 24528 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1509_
timestamp 1698431365
transform -1 0 23968 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1510_
timestamp 1698431365
transform -1 0 10080 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1511_
timestamp 1698431365
transform 1 0 2240 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1512_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3360 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1513_
timestamp 1698431365
transform 1 0 4816 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1514_
timestamp 1698431365
transform 1 0 23968 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1515_
timestamp 1698431365
transform -1 0 4144 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1516_
timestamp 1698431365
transform 1 0 4144 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1517_
timestamp 1698431365
transform -1 0 3024 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1518_
timestamp 1698431365
transform 1 0 23968 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1519_
timestamp 1698431365
transform -1 0 7616 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1520_
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1521_
timestamp 1698431365
transform 1 0 4480 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1522_
timestamp 1698431365
transform 1 0 4816 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1523_
timestamp 1698431365
transform -1 0 5040 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1524_
timestamp 1698431365
transform -1 0 3808 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1525_
timestamp 1698431365
transform -1 0 3472 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1526_
timestamp 1698431365
transform -1 0 3472 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1527_
timestamp 1698431365
transform 1 0 2352 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1528_
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1529_
timestamp 1698431365
transform 1 0 4368 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1530_
timestamp 1698431365
transform 1 0 5600 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1531_
timestamp 1698431365
transform -1 0 6384 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1532_
timestamp 1698431365
transform -1 0 6160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1533_
timestamp 1698431365
transform -1 0 5488 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1534_
timestamp 1698431365
transform 1 0 6720 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1535_
timestamp 1698431365
transform 1 0 7728 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1536_
timestamp 1698431365
transform -1 0 20160 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1537_
timestamp 1698431365
transform -1 0 6048 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1538_
timestamp 1698431365
transform -1 0 5824 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1539_
timestamp 1698431365
transform -1 0 3360 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1540_
timestamp 1698431365
transform -1 0 19040 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1541_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5040 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1542_
timestamp 1698431365
transform -1 0 6048 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1543_
timestamp 1698431365
transform -1 0 6160 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1544_
timestamp 1698431365
transform -1 0 5264 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1545_
timestamp 1698431365
transform -1 0 4032 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1546_
timestamp 1698431365
transform -1 0 3248 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1547_
timestamp 1698431365
transform 1 0 6048 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1548_
timestamp 1698431365
transform 1 0 5824 0 1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1549_
timestamp 1698431365
transform 1 0 6048 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1550_
timestamp 1698431365
transform 1 0 6160 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1551_
timestamp 1698431365
transform 1 0 14672 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1552_
timestamp 1698431365
transform 1 0 15008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1553_
timestamp 1698431365
transform -1 0 15008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1554_
timestamp 1698431365
transform -1 0 18592 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1555_
timestamp 1698431365
transform 1 0 17696 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1556_
timestamp 1698431365
transform 1 0 19600 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1557_
timestamp 1698431365
transform 1 0 16016 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1558_
timestamp 1698431365
transform -1 0 21616 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1559_
timestamp 1698431365
transform -1 0 19488 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1560_
timestamp 1698431365
transform 1 0 21952 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1561_
timestamp 1698431365
transform 1 0 21840 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1562_
timestamp 1698431365
transform -1 0 23296 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1563_
timestamp 1698431365
transform 1 0 22624 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1564_
timestamp 1698431365
transform -1 0 24192 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1565_
timestamp 1698431365
transform -1 0 23632 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1566_
timestamp 1698431365
transform 1 0 22400 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1567_
timestamp 1698431365
transform -1 0 22848 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1568_
timestamp 1698431365
transform -1 0 20496 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1569_
timestamp 1698431365
transform 1 0 24640 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1570_
timestamp 1698431365
transform 1 0 24528 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1571_
timestamp 1698431365
transform 1 0 22848 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1572_
timestamp 1698431365
transform -1 0 27440 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1573_
timestamp 1698431365
transform -1 0 26096 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1574_
timestamp 1698431365
transform -1 0 27776 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1575_
timestamp 1698431365
transform -1 0 25984 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1576_
timestamp 1698431365
transform 1 0 30016 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1577_
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1578_
timestamp 1698431365
transform 1 0 30128 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1579_
timestamp 1698431365
transform 1 0 31024 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1580_
timestamp 1698431365
transform -1 0 30016 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1581_
timestamp 1698431365
transform -1 0 31808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1582_
timestamp 1698431365
transform 1 0 31584 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1583_
timestamp 1698431365
transform -1 0 30688 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1584_
timestamp 1698431365
transform 1 0 30016 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1585_
timestamp 1698431365
transform -1 0 31584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1586_
timestamp 1698431365
transform 1 0 28112 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1587_
timestamp 1698431365
transform -1 0 30352 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1588_
timestamp 1698431365
transform 1 0 25312 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1589_
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1590_
timestamp 1698431365
transform 1 0 24864 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1591_
timestamp 1698431365
transform 1 0 32928 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1592_
timestamp 1698431365
transform 1 0 33152 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1593_
timestamp 1698431365
transform 1 0 34048 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1594_
timestamp 1698431365
transform 1 0 34944 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1595_
timestamp 1698431365
transform -1 0 34048 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1596_
timestamp 1698431365
transform 1 0 31248 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1597_
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1598_
timestamp 1698431365
transform -1 0 32368 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1599_
timestamp 1698431365
transform -1 0 31920 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1600_
timestamp 1698431365
transform -1 0 31696 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1601_
timestamp 1698431365
transform 1 0 32032 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1602_
timestamp 1698431365
transform 1 0 32256 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1603_
timestamp 1698431365
transform 1 0 33152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1604_
timestamp 1698431365
transform -1 0 33264 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1605_
timestamp 1698431365
transform -1 0 34048 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1606_
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1607_
timestamp 1698431365
transform -1 0 30688 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1608_
timestamp 1698431365
transform -1 0 31584 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1609_
timestamp 1698431365
transform -1 0 30688 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1610_
timestamp 1698431365
transform -1 0 29792 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1611_
timestamp 1698431365
transform -1 0 26208 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1612_
timestamp 1698431365
transform 1 0 45360 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1613_
timestamp 1698431365
transform 1 0 36400 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1614_
timestamp 1698431365
transform 1 0 38080 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1615_
timestamp 1698431365
transform 1 0 38752 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1616_
timestamp 1698431365
transform 1 0 45808 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1617_
timestamp 1698431365
transform 1 0 45360 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1618_
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1619_
timestamp 1698431365
transform -1 0 44240 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1620_
timestamp 1698431365
transform -1 0 46144 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1621_
timestamp 1698431365
transform 1 0 46144 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1622_
timestamp 1698431365
transform -1 0 43008 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1623_
timestamp 1698431365
transform 1 0 43120 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1624_
timestamp 1698431365
transform 1 0 42000 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1625_
timestamp 1698431365
transform 1 0 40768 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1626_
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1627_
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1628_
timestamp 1698431365
transform 1 0 39872 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1629_
timestamp 1698431365
transform -1 0 37520 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1630_
timestamp 1698431365
transform 1 0 36960 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1631_
timestamp 1698431365
transform 1 0 39648 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1632_
timestamp 1698431365
transform 1 0 38192 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1633_
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1634_
timestamp 1698431365
transform -1 0 44128 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1635_
timestamp 1698431365
transform 1 0 38976 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1636_
timestamp 1698431365
transform 1 0 37632 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1637_
timestamp 1698431365
transform -1 0 35952 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1638_
timestamp 1698431365
transform 1 0 35840 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1639_
timestamp 1698431365
transform 1 0 34720 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1640_
timestamp 1698431365
transform 1 0 36512 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1641_
timestamp 1698431365
transform 1 0 34272 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1642_
timestamp 1698431365
transform 1 0 43344 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1643_
timestamp 1698431365
transform 1 0 38192 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1644_
timestamp 1698431365
transform -1 0 44464 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1645_
timestamp 1698431365
transform -1 0 45472 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1646_
timestamp 1698431365
transform 1 0 31472 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1647_
timestamp 1698431365
transform -1 0 45136 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1648_
timestamp 1698431365
transform 1 0 46816 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1649_
timestamp 1698431365
transform 1 0 47264 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1650_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1651_
timestamp 1698431365
transform 1 0 37520 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1652_
timestamp 1698431365
transform 1 0 41776 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1653_
timestamp 1698431365
transform 1 0 41552 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1654_
timestamp 1698431365
transform 1 0 36064 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1655_
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1656_
timestamp 1698431365
transform 1 0 39200 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1657_
timestamp 1698431365
transform -1 0 31696 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1658_
timestamp 1698431365
transform 1 0 41664 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1659_
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1660_
timestamp 1698431365
transform 1 0 38864 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1661_
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1662_
timestamp 1698431365
transform -1 0 35952 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1663_
timestamp 1698431365
transform -1 0 35728 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1664_
timestamp 1698431365
transform -1 0 32480 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1665_
timestamp 1698431365
transform 1 0 21280 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1666_
timestamp 1698431365
transform 1 0 18256 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1667_
timestamp 1698431365
transform -1 0 19824 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1668_
timestamp 1698431365
transform -1 0 3360 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1669_
timestamp 1698431365
transform -1 0 6832 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1670_
timestamp 1698431365
transform -1 0 6160 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1671_
timestamp 1698431365
transform 1 0 19824 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1672_
timestamp 1698431365
transform 1 0 9632 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1673_
timestamp 1698431365
transform -1 0 8960 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1674_
timestamp 1698431365
transform 1 0 8848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1675_
timestamp 1698431365
transform 1 0 7952 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1676_
timestamp 1698431365
transform 1 0 10976 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1677_
timestamp 1698431365
transform -1 0 9184 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1678_
timestamp 1698431365
transform 1 0 10080 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1679_
timestamp 1698431365
transform -1 0 12880 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1680_
timestamp 1698431365
transform -1 0 12208 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1681_
timestamp 1698431365
transform 1 0 18256 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1682_
timestamp 1698431365
transform 1 0 18256 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1683_
timestamp 1698431365
transform 1 0 18928 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1684_
timestamp 1698431365
transform 1 0 19152 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1685_
timestamp 1698431365
transform 1 0 20384 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1686_
timestamp 1698431365
transform -1 0 18928 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1687_
timestamp 1698431365
transform 1 0 18480 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1688_
timestamp 1698431365
transform 1 0 19376 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1689_
timestamp 1698431365
transform -1 0 18256 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1690_
timestamp 1698431365
transform -1 0 15904 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1691_
timestamp 1698431365
transform -1 0 15120 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1692_
timestamp 1698431365
transform -1 0 15456 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1693_
timestamp 1698431365
transform -1 0 15120 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1694_
timestamp 1698431365
transform 1 0 2240 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1695_
timestamp 1698431365
transform 1 0 4816 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1696_
timestamp 1698431365
transform -1 0 5712 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1697_
timestamp 1698431365
transform 1 0 3696 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1698_
timestamp 1698431365
transform -1 0 4368 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1699_
timestamp 1698431365
transform 1 0 21616 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1700_
timestamp 1698431365
transform -1 0 22624 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1701_
timestamp 1698431365
transform 1 0 3136 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1702_
timestamp 1698431365
transform 1 0 4480 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1703_
timestamp 1698431365
transform -1 0 10640 0 1 14112
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1704_
timestamp 1698431365
transform 1 0 15120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1705_
timestamp 1698431365
transform 1 0 5936 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1706_
timestamp 1698431365
transform 1 0 6048 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1707_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13552 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1708_
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1709_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1710_
timestamp 1698431365
transform -1 0 19376 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1711_
timestamp 1698431365
transform 1 0 17136 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1712_
timestamp 1698431365
transform 1 0 15456 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1713_
timestamp 1698431365
transform 1 0 17584 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1714_
timestamp 1698431365
transform 1 0 17808 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1715_
timestamp 1698431365
transform -1 0 18592 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1716_
timestamp 1698431365
transform -1 0 17920 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1717_
timestamp 1698431365
transform 1 0 18144 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1718_
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1719_
timestamp 1698431365
transform 1 0 18480 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1720_
timestamp 1698431365
transform 1 0 21952 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1721_
timestamp 1698431365
transform 1 0 18816 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1722_
timestamp 1698431365
transform 1 0 17920 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1723_
timestamp 1698431365
transform -1 0 22512 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1724_
timestamp 1698431365
transform 1 0 21280 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1725_
timestamp 1698431365
transform 1 0 21504 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1726_
timestamp 1698431365
transform -1 0 19712 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1727_
timestamp 1698431365
transform -1 0 23632 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1728_
timestamp 1698431365
transform -1 0 23072 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1729_
timestamp 1698431365
transform -1 0 22064 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1730_
timestamp 1698431365
transform 1 0 21280 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1731_
timestamp 1698431365
transform -1 0 22064 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1732_
timestamp 1698431365
transform 1 0 23296 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1733_
timestamp 1698431365
transform 1 0 23072 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1734_
timestamp 1698431365
transform 1 0 23744 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1735_
timestamp 1698431365
transform 1 0 21168 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1736_
timestamp 1698431365
transform 1 0 23072 0 1 10976
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1737_
timestamp 1698431365
transform 1 0 29120 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1738_
timestamp 1698431365
transform -1 0 30352 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1739_
timestamp 1698431365
transform 1 0 32144 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1740_
timestamp 1698431365
transform 1 0 32704 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1741_
timestamp 1698431365
transform 1 0 33824 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1742_
timestamp 1698431365
transform 1 0 37184 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1743_
timestamp 1698431365
transform 1 0 38528 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1744_
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1745_
timestamp 1698431365
transform 1 0 37520 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1746_
timestamp 1698431365
transform 1 0 38640 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1747_
timestamp 1698431365
transform -1 0 36176 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1748_
timestamp 1698431365
transform 1 0 35504 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1749_
timestamp 1698431365
transform 1 0 35280 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1750_
timestamp 1698431365
transform -1 0 36624 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1751_
timestamp 1698431365
transform 1 0 37968 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1752_
timestamp 1698431365
transform 1 0 38304 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1753_
timestamp 1698431365
transform 1 0 38416 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1754_
timestamp 1698431365
transform -1 0 38416 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1755_
timestamp 1698431365
transform -1 0 40768 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1756_
timestamp 1698431365
transform 1 0 39424 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1757_
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1758_
timestamp 1698431365
transform 1 0 41104 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1759_
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1760_
timestamp 1698431365
transform -1 0 42896 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1761_
timestamp 1698431365
transform 1 0 43792 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1762_
timestamp 1698431365
transform -1 0 43792 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1763_
timestamp 1698431365
transform 1 0 43680 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1764_
timestamp 1698431365
transform 1 0 43344 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1765_
timestamp 1698431365
transform 1 0 43680 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1766_
timestamp 1698431365
transform 1 0 44240 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1767_
timestamp 1698431365
transform -1 0 42672 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1768_
timestamp 1698431365
transform -1 0 43008 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1769_
timestamp 1698431365
transform -1 0 41888 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1770_
timestamp 1698431365
transform -1 0 43456 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1771_
timestamp 1698431365
transform -1 0 41440 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1772_
timestamp 1698431365
transform -1 0 14784 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1773_
timestamp 1698431365
transform -1 0 14336 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1774_
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1775_
timestamp 1698431365
transform 1 0 12768 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1776_
timestamp 1698431365
transform -1 0 15008 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1777_
timestamp 1698431365
transform -1 0 14672 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1778_
timestamp 1698431365
transform 1 0 15120 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1779_
timestamp 1698431365
transform -1 0 14224 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1780_
timestamp 1698431365
transform 1 0 9856 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1781_
timestamp 1698431365
transform -1 0 18816 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1782_
timestamp 1698431365
transform 1 0 10752 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1783_
timestamp 1698431365
transform 1 0 10080 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1784_
timestamp 1698431365
transform 1 0 9632 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1785_
timestamp 1698431365
transform -1 0 19040 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1786_
timestamp 1698431365
transform -1 0 11872 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1787_
timestamp 1698431365
transform 1 0 10976 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1788_
timestamp 1698431365
transform 1 0 11984 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1789_
timestamp 1698431365
transform -1 0 14224 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1790_
timestamp 1698431365
transform 1 0 12208 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1791_
timestamp 1698431365
transform 1 0 15008 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1792_
timestamp 1698431365
transform 1 0 17808 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1793_
timestamp 1698431365
transform 1 0 15232 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1794_
timestamp 1698431365
transform 1 0 14784 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1795_
timestamp 1698431365
transform 1 0 17920 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1796_
timestamp 1698431365
transform 1 0 15232 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1797_
timestamp 1698431365
transform -1 0 15456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1798_
timestamp 1698431365
transform 1 0 15232 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1799_
timestamp 1698431365
transform 1 0 14336 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1800_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28896 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1801_
timestamp 1698431365
transform 1 0 10976 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1802_
timestamp 1698431365
transform 1 0 8064 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1803_
timestamp 1698431365
transform -1 0 7504 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1804_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7168 0 -1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1805_
timestamp 1698431365
transform 1 0 7168 0 1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1806_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1807_
timestamp 1698431365
transform 1 0 11424 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1808_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1809_
timestamp 1698431365
transform -1 0 19376 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1810_
timestamp 1698431365
transform 1 0 21168 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1811_
timestamp 1698431365
transform 1 0 22736 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1812_
timestamp 1698431365
transform -1 0 28560 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1813_
timestamp 1698431365
transform 1 0 28560 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1814_
timestamp 1698431365
transform 1 0 30464 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1815_
timestamp 1698431365
transform 1 0 33600 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1816_
timestamp 1698431365
transform 1 0 35392 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1817_
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1818_
timestamp 1698431365
transform 1 0 41552 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1819_
timestamp 1698431365
transform 1 0 44352 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1820_
timestamp 1698431365
transform 1 0 44912 0 1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1821_
timestamp 1698431365
transform 1 0 45136 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1822_
timestamp 1698431365
transform 1 0 45136 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1823_
timestamp 1698431365
transform 1 0 44912 0 -1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1824_
timestamp 1698431365
transform 1 0 44912 0 1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1825_
timestamp 1698431365
transform 1 0 25312 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1826_
timestamp 1698431365
transform -1 0 30800 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1827_
timestamp 1698431365
transform -1 0 32256 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1828_
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1829_
timestamp 1698431365
transform 1 0 20832 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1830_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1831_
timestamp 1698431365
transform 1 0 14000 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1832_
timestamp 1698431365
transform 1 0 15904 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1833_
timestamp 1698431365
transform 1 0 19264 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1834_
timestamp 1698431365
transform 1 0 19600 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1835_
timestamp 1698431365
transform -1 0 28784 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1836_
timestamp 1698431365
transform 1 0 18144 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1837_
timestamp 1698431365
transform 1 0 21392 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1838_
timestamp 1698431365
transform 1 0 18368 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1839_
timestamp 1698431365
transform 1 0 26544 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1840_
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1841_
timestamp 1698431365
transform 1 0 29680 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1842_
timestamp 1698431365
transform -1 0 37968 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1843_
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1844_
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1845_
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1846_
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1847_
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1848_
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1849_
timestamp 1698431365
transform 1 0 5712 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1850_
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1851_
timestamp 1698431365
transform 1 0 7504 0 1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1852_
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1853_
timestamp 1698431365
transform 1 0 2576 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1854_
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1855_
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1856_
timestamp 1698431365
transform 1 0 11984 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1857_
timestamp 1698431365
transform 1 0 17360 0 1 21952
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1858_
timestamp 1698431365
transform 1 0 17920 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1859_
timestamp 1698431365
transform 1 0 21952 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1860_
timestamp 1698431365
transform 1 0 20272 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1861_
timestamp 1698431365
transform 1 0 19152 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1862_
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1863_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1864_
timestamp 1698431365
transform -1 0 32032 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1865_
timestamp 1698431365
transform 1 0 31024 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1866_
timestamp 1698431365
transform 1 0 29456 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1867_
timestamp 1698431365
transform 1 0 25536 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1868_
timestamp 1698431365
transform 1 0 34720 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1869_
timestamp 1698431365
transform 1 0 33824 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1870_
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1871_
timestamp 1698431365
transform 1 0 33376 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1872_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1873_
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1874_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1875_
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1876_
timestamp 1698431365
transform 1 0 45136 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1877_
timestamp 1698431365
transform 1 0 41216 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1878_
timestamp 1698431365
transform 1 0 38976 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1879_
timestamp 1698431365
transform 1 0 37520 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1880_
timestamp 1698431365
transform 1 0 37072 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1881_
timestamp 1698431365
transform 1 0 33040 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1882_
timestamp 1698431365
transform 1 0 33264 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1883_
timestamp 1698431365
transform 1 0 45136 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1884_
timestamp 1698431365
transform -1 0 46816 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1885_
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1886_
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1887_
timestamp 1698431365
transform 1 0 37968 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1888_
timestamp 1698431365
transform 1 0 38864 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1889_
timestamp 1698431365
transform 1 0 35616 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1890_
timestamp 1698431365
transform 1 0 31584 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1891_
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1892_
timestamp 1698431365
transform 1 0 3696 0 -1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1893_
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1894_
timestamp 1698431365
transform 1 0 9632 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1895_
timestamp 1698431365
transform 1 0 9856 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1896_
timestamp 1698431365
transform -1 0 23184 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1897_
timestamp 1698431365
transform -1 0 21840 0 -1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1898_
timestamp 1698431365
transform 1 0 13776 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1899_
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1900_
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1901_
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1902_
timestamp 1698431365
transform 1 0 4032 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1903_
timestamp 1698431365
transform 1 0 7056 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1904_
timestamp 1698431365
transform -1 0 20496 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1905_
timestamp 1698431365
transform -1 0 20496 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1906_
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1907_
timestamp 1698431365
transform 1 0 20832 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1908_
timestamp 1698431365
transform 1 0 19936 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1909_
timestamp 1698431365
transform 1 0 20496 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1910_
timestamp 1698431365
transform 1 0 23968 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1911_
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1912_
timestamp 1698431365
transform -1 0 35952 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1913_
timestamp 1698431365
transform -1 0 41328 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1914_
timestamp 1698431365
transform -1 0 42336 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1915_
timestamp 1698431365
transform 1 0 34496 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1916_
timestamp 1698431365
transform 1 0 36624 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1917_
timestamp 1698431365
transform 1 0 41104 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1918_
timestamp 1698431365
transform 1 0 41216 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1919_
timestamp 1698431365
transform 1 0 45136 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1920_
timestamp 1698431365
transform 1 0 45136 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1921_
timestamp 1698431365
transform 1 0 38528 0 1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1922_
timestamp 1698431365
transform 1 0 39536 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1923_
timestamp 1698431365
transform -1 0 12768 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1924_
timestamp 1698431365
transform -1 0 15120 0 -1 42336
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1925_
timestamp 1698431365
transform 1 0 7952 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1926_
timestamp 1698431365
transform 1 0 5936 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1927_
timestamp 1698431365
transform 1 0 11424 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1928_
timestamp 1698431365
transform 1 0 14560 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1929_
timestamp 1698431365
transform 1 0 14672 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1930_
timestamp 1698431365
transform -1 0 18144 0 1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1934_
timestamp 1698431365
transform 1 0 37520 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1935_
timestamp 1698431365
transform 1 0 39536 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1936_
timestamp 1698431365
transform -1 0 35616 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1937_
timestamp 1698431365
transform 1 0 43792 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1938_
timestamp 1698431365
transform 1 0 32032 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1939_
timestamp 1698431365
transform 1 0 31696 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1940_
timestamp 1698431365
transform 1 0 39648 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1941_
timestamp 1698431365
transform 1 0 30688 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1942_
timestamp 1698431365
transform 1 0 33040 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1943_
timestamp 1698431365
transform 1 0 35952 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1944_
timestamp 1698431365
transform 1 0 37968 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1945_
timestamp 1698431365
transform 1 0 32368 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1946_
timestamp 1698431365
transform 1 0 33040 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1947_
timestamp 1698431365
transform 1 0 40992 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1948_
timestamp 1698431365
transform 1 0 33376 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1949_
timestamp 1698431365
transform -1 0 47040 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1950_
timestamp 1698431365
transform 1 0 30016 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1951_
timestamp 1698431365
transform 1 0 33600 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1952_
timestamp 1698431365
transform 1 0 37296 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1953_
timestamp 1698431365
transform 1 0 38752 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1954_
timestamp 1698431365
transform 1 0 38192 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1955_
timestamp 1698431365
transform 1 0 32368 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1956_
timestamp 1698431365
transform -1 0 37632 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0962__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__A1
timestamp 1698431365
transform 1 0 18144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__B2
timestamp 1698431365
transform 1 0 21392 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__I
timestamp 1698431365
transform 1 0 12880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0973__I
timestamp 1698431365
transform 1 0 16912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0979__B2
timestamp 1698431365
transform 1 0 19712 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__I
timestamp 1698431365
transform -1 0 13664 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__I
timestamp 1698431365
transform 1 0 18368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1026__B
timestamp 1698431365
transform -1 0 13552 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1071__B2
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__C2
timestamp 1698431365
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__A1
timestamp 1698431365
transform -1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__B
timestamp 1698431365
transform 1 0 14672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__B
timestamp 1698431365
transform -1 0 37184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__A2
timestamp 1698431365
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__A1
timestamp 1698431365
transform -1 0 9968 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__A1
timestamp 1698431365
transform 1 0 17472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__A2
timestamp 1698431365
transform 1 0 13888 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__A2
timestamp 1698431365
transform -1 0 35840 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__A2
timestamp 1698431365
transform 1 0 34496 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__I
timestamp 1698431365
transform 1 0 22064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__A1
timestamp 1698431365
transform 1 0 13104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__B
timestamp 1698431365
transform 1 0 14448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1118__A1
timestamp 1698431365
transform 1 0 12768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A1
timestamp 1698431365
transform 1 0 10304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__B
timestamp 1698431365
transform 1 0 12320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__A1
timestamp 1698431365
transform 1 0 11088 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1123__I
timestamp 1698431365
transform 1 0 24864 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1124__I
timestamp 1698431365
transform 1 0 12208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__A1
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1126__A1
timestamp 1698431365
transform -1 0 8176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__I
timestamp 1698431365
transform 1 0 17472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__A2
timestamp 1698431365
transform 1 0 13552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1144__A2
timestamp 1698431365
transform 1 0 11872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A2
timestamp 1698431365
transform 1 0 20720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__I
timestamp 1698431365
transform -1 0 30016 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__I
timestamp 1698431365
transform 1 0 32480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1179__I
timestamp 1698431365
transform 1 0 46592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1181__I
timestamp 1698431365
transform 1 0 47040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1188__I
timestamp 1698431365
transform 1 0 42560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1190__B
timestamp 1698431365
transform -1 0 45584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__I
timestamp 1698431365
transform 1 0 47488 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1196__B
timestamp 1698431365
transform -1 0 42672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__B
timestamp 1698431365
transform 1 0 46256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1202__B
timestamp 1698431365
transform 1 0 48048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__B
timestamp 1698431365
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__B
timestamp 1698431365
transform -1 0 46256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1269__B2
timestamp 1698431365
transform -1 0 22512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A1
timestamp 1698431365
transform 1 0 27664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1331__B
timestamp 1698431365
transform 1 0 25312 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1340__I
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1381__I
timestamp 1698431365
transform 1 0 26656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1387__A1
timestamp 1698431365
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__B
timestamp 1698431365
transform -1 0 20496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1401__A1
timestamp 1698431365
transform -1 0 20496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__A3
timestamp 1698431365
transform -1 0 19264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__B
timestamp 1698431365
transform 1 0 20384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__A1
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1424__A1
timestamp 1698431365
transform 1 0 17920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1426__A1
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__A1
timestamp 1698431365
transform 1 0 16128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1444__A1
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1492__A1
timestamp 1698431365
transform 1 0 26208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__B
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1510__I
timestamp 1698431365
transform 1 0 10304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A2
timestamp 1698431365
transform -1 0 2240 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__A1
timestamp 1698431365
transform 1 0 5712 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__A1
timestamp 1698431365
transform -1 0 3360 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__I
timestamp 1698431365
transform 1 0 7616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__A1
timestamp 1698431365
transform 1 0 3248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1535__A1
timestamp 1698431365
transform 1 0 8624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1536__I
timestamp 1698431365
transform 1 0 20384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1539__A1
timestamp 1698431365
transform 1 0 3584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1540__I
timestamp 1698431365
transform 1 0 19264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A1
timestamp 1698431365
transform 1 0 3472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A1
timestamp 1698431365
transform 1 0 18368 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A2
timestamp 1698431365
transform 1 0 23520 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__C
timestamp 1698431365
transform -1 0 23744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__A1
timestamp 1698431365
transform 1 0 19600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1569__I
timestamp 1698431365
transform -1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__A1
timestamp 1698431365
transform 1 0 24416 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A2
timestamp 1698431365
transform 1 0 26656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__I
timestamp 1698431365
transform 1 0 24640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A1
timestamp 1698431365
transform 1 0 31584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__A1
timestamp 1698431365
transform 1 0 29568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__A1
timestamp 1698431365
transform 1 0 25312 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A3
timestamp 1698431365
transform -1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__B
timestamp 1698431365
transform 1 0 45136 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A2
timestamp 1698431365
transform 1 0 42112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__I
timestamp 1698431365
transform 1 0 31248 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__A2
timestamp 1698431365
transform 1 0 42560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__B
timestamp 1698431365
transform 1 0 44240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__A2
timestamp 1698431365
transform -1 0 47152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__B
timestamp 1698431365
transform -1 0 47600 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__B
timestamp 1698431365
transform 1 0 41552 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__B
timestamp 1698431365
transform 1 0 40320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__I
timestamp 1698431365
transform 1 0 30576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__B
timestamp 1698431365
transform -1 0 38640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__B
timestamp 1698431365
transform 1 0 37744 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__B
timestamp 1698431365
transform 1 0 34832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__A1
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__I
timestamp 1698431365
transform 1 0 17360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A2
timestamp 1698431365
transform 1 0 3584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A1
timestamp 1698431365
transform 1 0 6384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__A1
timestamp 1698431365
transform 1 0 9408 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A1
timestamp 1698431365
transform 1 0 11872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__A1
timestamp 1698431365
transform 1 0 12432 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A1
timestamp 1698431365
transform 1 0 21280 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A1
timestamp 1698431365
transform 1 0 20496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A2
timestamp 1698431365
transform 1 0 19152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__I
timestamp 1698431365
transform -1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A2
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__A2
timestamp 1698431365
transform 1 0 15456 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__A1
timestamp 1698431365
transform -1 0 14784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A1
timestamp 1698431365
transform 1 0 5712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__A1
timestamp 1698431365
transform 1 0 4592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__I
timestamp 1698431365
transform 1 0 22512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__I
timestamp 1698431365
transform -1 0 23072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__A1
timestamp 1698431365
transform 1 0 5712 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__A1
timestamp 1698431365
transform 1 0 7728 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__A3
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A1
timestamp 1698431365
transform 1 0 10528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__I
timestamp 1698431365
transform 1 0 19600 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__A1
timestamp 1698431365
transform 1 0 18704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__A1
timestamp 1698431365
transform 1 0 18144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__C
timestamp 1698431365
transform 1 0 20160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__A1
timestamp 1698431365
transform 1 0 22848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__A1
timestamp 1698431365
transform -1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__A1
timestamp 1698431365
transform 1 0 22288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__C
timestamp 1698431365
transform 1 0 23520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__A1
timestamp 1698431365
transform 1 0 29456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__C
timestamp 1698431365
transform 1 0 33600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A1
timestamp 1698431365
transform -1 0 38528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__C
timestamp 1698431365
transform 1 0 38528 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__A1
timestamp 1698431365
transform 1 0 35728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__C
timestamp 1698431365
transform 1 0 37072 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1757__A1
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__A1
timestamp 1698431365
transform 1 0 42000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__A1
timestamp 1698431365
transform 1 0 43456 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A1
timestamp 1698431365
transform -1 0 44240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__A1
timestamp 1698431365
transform 1 0 40320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A1
timestamp 1698431365
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__B
timestamp 1698431365
transform -1 0 14112 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__A2
timestamp 1698431365
transform 1 0 14896 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__B
timestamp 1698431365
transform 1 0 16240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__I
timestamp 1698431365
transform 1 0 19040 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__CLK
timestamp 1698431365
transform 1 0 32144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__CLK
timestamp 1698431365
transform 1 0 10528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__CLK
timestamp 1698431365
transform 1 0 8400 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__CLK
timestamp 1698431365
transform 1 0 7392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__CLK
timestamp 1698431365
transform 1 0 10640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__CLK
timestamp 1698431365
transform 1 0 12880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__CLK
timestamp 1698431365
transform 1 0 14896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__CLK
timestamp 1698431365
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__CLK
timestamp 1698431365
transform 1 0 29232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__CLK
timestamp 1698431365
transform 1 0 32032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__CLK
timestamp 1698431365
transform 1 0 33264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__CLK
timestamp 1698431365
transform 1 0 34720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__CLK
timestamp 1698431365
transform 1 0 38864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__CLK
timestamp 1698431365
transform 1 0 41328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__CLK
timestamp 1698431365
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__CLK
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__CLK
timestamp 1698431365
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__CLK
timestamp 1698431365
transform 1 0 44464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__CLK
timestamp 1698431365
transform 1 0 44688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__CLK
timestamp 1698431365
transform 1 0 29232 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__CLK
timestamp 1698431365
transform 1 0 30800 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__CLK
timestamp 1698431365
transform -1 0 29456 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__CLK
timestamp 1698431365
transform 1 0 29232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__CLK
timestamp 1698431365
transform 1 0 33152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__CLK
timestamp 1698431365
transform -1 0 38192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__CLK
timestamp 1698431365
transform 1 0 5040 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__CLK
timestamp 1698431365
transform 1 0 8960 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__CLK
timestamp 1698431365
transform 1 0 5040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__CLK
timestamp 1698431365
transform 1 0 5936 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__CLK
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__CLK
timestamp 1698431365
transform 1 0 5824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__CLK
timestamp 1698431365
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__CLK
timestamp 1698431365
transform 1 0 15456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__CLK
timestamp 1698431365
transform 1 0 32144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__CLK
timestamp 1698431365
transform -1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1879__CLK
timestamp 1698431365
transform 1 0 41440 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__CLK
timestamp 1698431365
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__CLK
timestamp 1698431365
transform 1 0 32816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__CLK
timestamp 1698431365
transform 1 0 42672 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__CLK
timestamp 1698431365
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__CLK
timestamp 1698431365
transform 1 0 36624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1886__CLK
timestamp 1698431365
transform 1 0 40992 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__CLK
timestamp 1698431365
transform 1 0 38864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__CLK
timestamp 1698431365
transform 1 0 35952 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__CLK
timestamp 1698431365
transform 1 0 44128 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__CLK
timestamp 1698431365
transform 1 0 33712 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__CLK
timestamp 1698431365
transform 1 0 4592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__CLK
timestamp 1698431365
transform 1 0 8064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1893__CLK
timestamp 1698431365
transform -1 0 8512 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__CLK
timestamp 1698431365
transform 1 0 13552 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__CLK
timestamp 1698431365
transform -1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__CLK
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__CLK
timestamp 1698431365
transform 1 0 7504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1903__CLK
timestamp 1698431365
transform 1 0 10528 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__CLK
timestamp 1698431365
transform 1 0 32480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__CLK
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__CLK
timestamp 1698431365
transform 1 0 41552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__CLK
timestamp 1698431365
transform 1 0 42560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__CLK
timestamp 1698431365
transform 1 0 34272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__CLK
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__CLK
timestamp 1698431365
transform 1 0 40880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__CLK
timestamp 1698431365
transform -1 0 41216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__CLK
timestamp 1698431365
transform 1 0 43568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__CLK
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1925__CLK
timestamp 1698431365
transform 1 0 11424 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__CLK
timestamp 1698431365
transform 1 0 9184 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1927__CLK
timestamp 1698431365
transform 1 0 12432 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1935__I
timestamp 1698431365
transform -1 0 39536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1936__I
timestamp 1698431365
transform 1 0 35280 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1937__I
timestamp 1698431365
transform 1 0 43120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1938__I
timestamp 1698431365
transform -1 0 31360 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__I
timestamp 1698431365
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__I
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__I
timestamp 1698431365
transform -1 0 38192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__I
timestamp 1698431365
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__I
timestamp 1698431365
transform -1 0 29680 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__I
timestamp 1698431365
transform 1 0 30352 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__I
timestamp 1698431365
transform 1 0 34272 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__I
timestamp 1698431365
transform 1 0 32144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_clk_I
timestamp 1698431365
transform 1 0 14000 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_clk_I
timestamp 1698431365
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_clk_I
timestamp 1698431365
transform 1 0 21840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_clk_I
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_clk_I
timestamp 1698431365
transform 1 0 12656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_clk_I
timestamp 1698431365
transform 1 0 10864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_clk_I
timestamp 1698431365
transform 1 0 20720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_clk_I
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_clk_I
timestamp 1698431365
transform 1 0 29568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_clk_I
timestamp 1698431365
transform -1 0 29680 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_clk_I
timestamp 1698431365
transform 1 0 37184 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_clk_I
timestamp 1698431365
transform 1 0 38416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_clk_I
timestamp 1698431365
transform 1 0 28448 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_clk_I
timestamp 1698431365
transform 1 0 30240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_clk_I
timestamp 1698431365
transform 1 0 37968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_clk_I
timestamp 1698431365
transform 1 0 36736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout115_I
timestamp 1698431365
transform 1 0 48160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout121_I
timestamp 1698431365
transform 1 0 29904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout123_I
timestamp 1698431365
transform -1 0 30912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout124_I
timestamp 1698431365
transform 1 0 44240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout125_I
timestamp 1698431365
transform -1 0 46704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 29680 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 28336 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 22848 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 22400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 20608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 16352 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 15904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 19152 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 30464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 24864 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 12768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 6496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 2464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 7392 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 6944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 7840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 13664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 18256 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 18704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 23408 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 25984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 13552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 31920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 32368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 37968 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 37296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 42560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 48384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 47712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 44464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 44016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 47040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 10192 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 45696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 46928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 12096 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 15456 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 14784 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform 1 0 2464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform 1 0 21840 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform 1 0 28448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform -1 0 46480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform -1 0 27328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform -1 0 31024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output63_I
timestamp 1698431365
transform -1 0 42448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output93_I
timestamp 1698431365
transform -1 0 4928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output108_I
timestamp 1698431365
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output110_I
timestamp 1698431365
transform 1 0 6272 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output111_I
timestamp 1698431365
transform 1 0 4704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14000 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1698431365
transform 1 0 10192 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1698431365
transform -1 0 21168 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1698431365
transform -1 0 12656 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1698431365
transform 1 0 9856 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1698431365
transform 1 0 17584 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1698431365
transform -1 0 19040 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1698431365
transform 1 0 29792 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1698431365
transform -1 0 33712 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1698431365
transform 1 0 38080 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1698431365
transform 1 0 38640 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1698431365
transform 1 0 29792 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1698431365
transform -1 0 34160 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1698431365
transform 1 0 39088 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1698431365
transform 1 0 37632 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout115
timestamp 1698431365
transform -1 0 48272 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout116
timestamp 1698431365
transform 1 0 47488 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout117
timestamp 1698431365
transform 1 0 37968 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout118
timestamp 1698431365
transform 1 0 34048 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout119
timestamp 1698431365
transform 1 0 32032 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout120
timestamp 1698431365
transform 1 0 32032 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout121
timestamp 1698431365
transform 1 0 31360 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout122
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout123
timestamp 1698431365
transform -1 0 32032 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout124
timestamp 1698431365
transform -1 0 45248 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout125
timestamp 1698431365
transform -1 0 47376 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout126
timestamp 1698431365
transform -1 0 31696 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout127
timestamp 1698431365
transform -1 0 40880 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout128
timestamp 1698431365
transform 1 0 44800 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout129
timestamp 1698431365
transform 1 0 18368 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout130
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  fanout131 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15456 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout132
timestamp 1698431365
transform 1 0 10080 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout133
timestamp 1698431365
transform -1 0 10864 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout134
timestamp 1698431365
transform -1 0 46032 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout135
timestamp 1698431365
transform 1 0 42896 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout136
timestamp 1698431365
transform -1 0 44128 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout137
timestamp 1698431365
transform 1 0 25424 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout138
timestamp 1698431365
transform -1 0 16576 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout139
timestamp 1698431365
transform 1 0 12208 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout140
timestamp 1698431365
transform -1 0 8848 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout141
timestamp 1698431365
transform -1 0 11648 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_46 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_334 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38752 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_338
timestamp 1698431365
transform 1 0 39200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_418
timestamp 1698431365
transform 1 0 48160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_34 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_50
timestamp 1698431365
transform 1 0 6944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_54
timestamp 1698431365
transform 1 0 7392 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_119
timestamp 1698431365
transform 1 0 14672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_123
timestamp 1698431365
transform 1 0 15120 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_146
timestamp 1698431365
transform 1 0 17696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_148
timestamp 1698431365
transform 1 0 17920 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_151
timestamp 1698431365
transform 1 0 18256 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_208
timestamp 1698431365
transform 1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_325
timestamp 1698431365
transform 1 0 37744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_329
timestamp 1698431365
transform 1 0 38192 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_345
timestamp 1698431365
transform 1 0 39984 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_354
timestamp 1698431365
transform 1 0 40992 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_359
timestamp 1698431365
transform 1 0 41552 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_363
timestamp 1698431365
transform 1 0 42000 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_365
timestamp 1698431365
transform 1 0 42224 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_368
timestamp 1698431365
transform 1 0 42560 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_400
timestamp 1698431365
transform 1 0 46144 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698431365
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_45
timestamp 1698431365
transform 1 0 6384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_47
timestamp 1698431365
transform 1 0 6608 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_95
timestamp 1698431365
transform 1 0 11984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_109
timestamp 1698431365
transform 1 0 13552 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_112
timestamp 1698431365
transform 1 0 13888 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_116
timestamp 1698431365
transform 1 0 14336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_118
timestamp 1698431365
transform 1 0 14560 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_131
timestamp 1698431365
transform 1 0 16016 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_165
timestamp 1698431365
transform 1 0 19824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_181
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_190
timestamp 1698431365
transform 1 0 22624 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_194
timestamp 1698431365
transform 1 0 23072 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_255
timestamp 1698431365
transform 1 0 29904 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_321 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_419
timestamp 1698431365
transform 1 0 48272 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_18
timestamp 1698431365
transform 1 0 3360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_55
timestamp 1698431365
transform 1 0 7504 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_61
timestamp 1698431365
transform 1 0 8176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_65
timestamp 1698431365
transform 1 0 8624 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_69
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_80
timestamp 1698431365
transform 1 0 10304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_82
timestamp 1698431365
transform 1 0 10528 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_111
timestamp 1698431365
transform 1 0 13776 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_127
timestamp 1698431365
transform 1 0 15568 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_135
timestamp 1698431365
transform 1 0 16464 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_146
timestamp 1698431365
transform 1 0 17696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_148
timestamp 1698431365
transform 1 0 17920 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_163
timestamp 1698431365
transform 1 0 19600 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_171
timestamp 1698431365
transform 1 0 20496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_175
timestamp 1698431365
transform 1 0 20944 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_191
timestamp 1698431365
transform 1 0 22736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_207
timestamp 1698431365
transform 1 0 24528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_216
timestamp 1698431365
transform 1 0 25536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_220
timestamp 1698431365
transform 1 0 25984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_222
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_241
timestamp 1698431365
transform 1 0 28336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_247
timestamp 1698431365
transform 1 0 29008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_251
timestamp 1698431365
transform 1 0 29456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_253
timestamp 1698431365
transform 1 0 29680 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_256
timestamp 1698431365
transform 1 0 30016 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_260
timestamp 1698431365
transform 1 0 30464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_262
timestamp 1698431365
transform 1 0 30688 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_271
timestamp 1698431365
transform 1 0 31696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_275
timestamp 1698431365
transform 1 0 32144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_284
timestamp 1698431365
transform 1 0 33152 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_295
timestamp 1698431365
transform 1 0 34384 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_333
timestamp 1698431365
transform 1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_337
timestamp 1698431365
transform 1 0 39088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_345
timestamp 1698431365
transform 1 0 39984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_347
timestamp 1698431365
transform 1 0 40208 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_381
timestamp 1698431365
transform 1 0 44016 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_413
timestamp 1698431365
transform 1 0 47600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_417
timestamp 1698431365
transform 1 0 48048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_419
timestamp 1698431365
transform 1 0 48272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_45
timestamp 1698431365
transform 1 0 6384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_67
timestamp 1698431365
transform 1 0 8848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_71
timestamp 1698431365
transform 1 0 9296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_95
timestamp 1698431365
transform 1 0 11984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_99
timestamp 1698431365
transform 1 0 12432 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_142
timestamp 1698431365
transform 1 0 17248 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_146
timestamp 1698431365
transform 1 0 17696 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_154
timestamp 1698431365
transform 1 0 18592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_156
timestamp 1698431365
transform 1 0 18816 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_167
timestamp 1698431365
transform 1 0 20048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_183
timestamp 1698431365
transform 1 0 21840 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_228
timestamp 1698431365
transform 1 0 26880 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_240
timestamp 1698431365
transform 1 0 28224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_255
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_270
timestamp 1698431365
transform 1 0 31584 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_276
timestamp 1698431365
transform 1 0 32256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_278
timestamp 1698431365
transform 1 0 32480 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_287
timestamp 1698431365
transform 1 0 33488 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_296
timestamp 1698431365
transform 1 0 34496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_300
timestamp 1698431365
transform 1 0 34944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_302
timestamp 1698431365
transform 1 0 35168 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_321
timestamp 1698431365
transform 1 0 37296 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_328
timestamp 1698431365
transform 1 0 38080 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_344
timestamp 1698431365
transform 1 0 39872 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_352
timestamp 1698431365
transform 1 0 40768 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_356
timestamp 1698431365
transform 1 0 41216 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_369
timestamp 1698431365
transform 1 0 42672 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_391
timestamp 1698431365
transform 1 0 45136 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_393
timestamp 1698431365
transform 1 0 45360 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_18
timestamp 1698431365
transform 1 0 3360 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_20
timestamp 1698431365
transform 1 0 3584 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_52
timestamp 1698431365
transform 1 0 7168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_56
timestamp 1698431365
transform 1 0 7616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_60
timestamp 1698431365
transform 1 0 8064 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_67
timestamp 1698431365
transform 1 0 8848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_76
timestamp 1698431365
transform 1 0 9856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_78
timestamp 1698431365
transform 1 0 10080 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_85
timestamp 1698431365
transform 1 0 10864 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_93
timestamp 1698431365
transform 1 0 11760 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_116
timestamp 1698431365
transform 1 0 14336 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_120
timestamp 1698431365
transform 1 0 14784 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_200
timestamp 1698431365
transform 1 0 23744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_214
timestamp 1698431365
transform 1 0 25312 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_223
timestamp 1698431365
transform 1 0 26320 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_231
timestamp 1698431365
transform 1 0 27216 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_240
timestamp 1698431365
transform 1 0 28224 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_247
timestamp 1698431365
transform 1 0 29008 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_263
timestamp 1698431365
transform 1 0 30800 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_271
timestamp 1698431365
transform 1 0 31696 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_275
timestamp 1698431365
transform 1 0 32144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_277
timestamp 1698431365
transform 1 0 32368 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_295
timestamp 1698431365
transform 1 0 34384 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_311
timestamp 1698431365
transform 1 0 36176 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_319
timestamp 1698431365
transform 1 0 37072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_325
timestamp 1698431365
transform 1 0 37744 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_329
timestamp 1698431365
transform 1 0 38192 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_338
timestamp 1698431365
transform 1 0 39200 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_382
timestamp 1698431365
transform 1 0 44128 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_414
timestamp 1698431365
transform 1 0 47712 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_418
timestamp 1698431365
transform 1 0 48160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_8
timestamp 1698431365
transform 1 0 2240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_12
timestamp 1698431365
transform 1 0 2688 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_28
timestamp 1698431365
transform 1 0 4480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_45
timestamp 1698431365
transform 1 0 6384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_47
timestamp 1698431365
transform 1 0 6608 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_68
timestamp 1698431365
transform 1 0 8960 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_70
timestamp 1698431365
transform 1 0 9184 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_91
timestamp 1698431365
transform 1 0 11536 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_99
timestamp 1698431365
transform 1 0 12432 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_111
timestamp 1698431365
transform 1 0 13776 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_127
timestamp 1698431365
transform 1 0 15568 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_135
timestamp 1698431365
transform 1 0 16464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_139
timestamp 1698431365
transform 1 0 16912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_141
timestamp 1698431365
transform 1 0 17136 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_148
timestamp 1698431365
transform 1 0 17920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_152
timestamp 1698431365
transform 1 0 18368 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_168
timestamp 1698431365
transform 1 0 20160 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_185
timestamp 1698431365
transform 1 0 22064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_189
timestamp 1698431365
transform 1 0 22512 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_197
timestamp 1698431365
transform 1 0 23408 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_201
timestamp 1698431365
transform 1 0 23856 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_231
timestamp 1698431365
transform 1 0 27216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_239
timestamp 1698431365
transform 1 0 28112 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_243
timestamp 1698431365
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_276
timestamp 1698431365
transform 1 0 32256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_309
timestamp 1698431365
transform 1 0 35952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_313
timestamp 1698431365
transform 1 0 36400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_327
timestamp 1698431365
transform 1 0 37968 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_357
timestamp 1698431365
transform 1 0 41328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_361
timestamp 1698431365
transform 1 0 41776 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_382
timestamp 1698431365
transform 1 0 44128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_384
timestamp 1698431365
transform 1 0 44352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_389
timestamp 1698431365
transform 1 0 44912 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_402
timestamp 1698431365
transform 1 0 46368 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_406
timestamp 1698431365
transform 1 0 46816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_410
timestamp 1698431365
transform 1 0 47264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_34
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_50
timestamp 1698431365
transform 1 0 6944 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_57
timestamp 1698431365
transform 1 0 7728 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_65
timestamp 1698431365
transform 1 0 8624 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_101
timestamp 1698431365
transform 1 0 12656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_105
timestamp 1698431365
transform 1 0 13104 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_113
timestamp 1698431365
transform 1 0 14000 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_122
timestamp 1698431365
transform 1 0 15008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_132
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_154
timestamp 1698431365
transform 1 0 18592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_166
timestamp 1698431365
transform 1 0 19936 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_170
timestamp 1698431365
transform 1 0 20384 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_186
timestamp 1698431365
transform 1 0 22176 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_194
timestamp 1698431365
transform 1 0 23072 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_220
timestamp 1698431365
transform 1 0 25984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_222
timestamp 1698431365
transform 1 0 26208 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_247
timestamp 1698431365
transform 1 0 29008 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_259
timestamp 1698431365
transform 1 0 30352 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_275
timestamp 1698431365
transform 1 0 32144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_286
timestamp 1698431365
transform 1 0 33376 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_290
timestamp 1698431365
transform 1 0 33824 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_304
timestamp 1698431365
transform 1 0 35392 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_312
timestamp 1698431365
transform 1 0 36288 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_332
timestamp 1698431365
transform 1 0 38528 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_348
timestamp 1698431365
transform 1 0 40320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_356
timestamp 1698431365
transform 1 0 41216 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_388
timestamp 1698431365
transform 1 0 44800 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_404
timestamp 1698431365
transform 1 0 46592 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_49
timestamp 1698431365
transform 1 0 6832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_80
timestamp 1698431365
transform 1 0 10304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_84
timestamp 1698431365
transform 1 0 10752 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_88
timestamp 1698431365
transform 1 0 11200 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_109
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_144
timestamp 1698431365
transform 1 0 17472 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_190
timestamp 1698431365
transform 1 0 22624 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_243
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_260
timestamp 1698431365
transform 1 0 30464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_262
timestamp 1698431365
transform 1 0 30688 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_267
timestamp 1698431365
transform 1 0 31248 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_309
timestamp 1698431365
transform 1 0 35952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_323
timestamp 1698431365
transform 1 0 37520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_330
timestamp 1698431365
transform 1 0 38304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_334
timestamp 1698431365
transform 1 0 38752 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_336
timestamp 1698431365
transform 1 0 38976 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_366
timestamp 1698431365
transform 1 0 42336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_370
timestamp 1698431365
transform 1 0 42784 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_379
timestamp 1698431365
transform 1 0 43792 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_391
timestamp 1698431365
transform 1 0 45136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_393
timestamp 1698431365
transform 1 0 45360 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_18
timestamp 1698431365
transform 1 0 3360 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_22
timestamp 1698431365
transform 1 0 3808 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_53
timestamp 1698431365
transform 1 0 7280 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_57
timestamp 1698431365
transform 1 0 7728 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_65
timestamp 1698431365
transform 1 0 8624 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_88
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_96
timestamp 1698431365
transform 1 0 12096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_98
timestamp 1698431365
transform 1 0 12320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_105
timestamp 1698431365
transform 1 0 13104 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_113
timestamp 1698431365
transform 1 0 14000 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_120
timestamp 1698431365
transform 1 0 14784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_138
timestamp 1698431365
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_163
timestamp 1698431365
transform 1 0 19600 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_195
timestamp 1698431365
transform 1 0 23184 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_201
timestamp 1698431365
transform 1 0 23856 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_224
timestamp 1698431365
transform 1 0 26432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_249
timestamp 1698431365
transform 1 0 29232 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_257
timestamp 1698431365
transform 1 0 30128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_265
timestamp 1698431365
transform 1 0 31024 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_290
timestamp 1698431365
transform 1 0 33824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_294
timestamp 1698431365
transform 1 0 34272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_311
timestamp 1698431365
transform 1 0 36176 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_322
timestamp 1698431365
transform 1 0 37408 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_343
timestamp 1698431365
transform 1 0 39760 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_347
timestamp 1698431365
transform 1 0 40208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_368
timestamp 1698431365
transform 1 0 42560 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_413
timestamp 1698431365
transform 1 0 47600 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_31
timestamp 1698431365
transform 1 0 4816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_41
timestamp 1698431365
transform 1 0 5936 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_57
timestamp 1698431365
transform 1 0 7728 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_65
timestamp 1698431365
transform 1 0 8624 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_124
timestamp 1698431365
transform 1 0 15232 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_130
timestamp 1698431365
transform 1 0 15904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_134
timestamp 1698431365
transform 1 0 16352 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_142
timestamp 1698431365
transform 1 0 17248 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_164
timestamp 1698431365
transform 1 0 19712 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_172
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_187
timestamp 1698431365
transform 1 0 22288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_231
timestamp 1698431365
transform 1 0 27216 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_239
timestamp 1698431365
transform 1 0 28112 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_249
timestamp 1698431365
transform 1 0 29232 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_258
timestamp 1698431365
transform 1 0 30240 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_269
timestamp 1698431365
transform 1 0 31472 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_297
timestamp 1698431365
transform 1 0 34608 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_322
timestamp 1698431365
transform 1 0 37408 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_330
timestamp 1698431365
transform 1 0 38304 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_346
timestamp 1698431365
transform 1 0 40096 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_350
timestamp 1698431365
transform 1 0 40544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_352
timestamp 1698431365
transform 1 0 40768 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_391
timestamp 1698431365
transform 1 0 45136 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_393
timestamp 1698431365
transform 1 0 45360 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_10
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_14
timestamp 1698431365
transform 1 0 2912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_50
timestamp 1698431365
transform 1 0 6944 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_55
timestamp 1698431365
transform 1 0 7504 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_59
timestamp 1698431365
transform 1 0 7952 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_63
timestamp 1698431365
transform 1 0 8400 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_80
timestamp 1698431365
transform 1 0 10304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_84
timestamp 1698431365
transform 1 0 10752 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_125
timestamp 1698431365
transform 1 0 15344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_127
timestamp 1698431365
transform 1 0 15568 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_137
timestamp 1698431365
transform 1 0 16688 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_139
timestamp 1698431365
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_188
timestamp 1698431365
transform 1 0 22400 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_199
timestamp 1698431365
transform 1 0 23632 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_204
timestamp 1698431365
transform 1 0 24192 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_218
timestamp 1698431365
transform 1 0 25760 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_263
timestamp 1698431365
transform 1 0 30800 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_286
timestamp 1698431365
transform 1 0 33376 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_306
timestamp 1698431365
transform 1 0 35616 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_339
timestamp 1698431365
transform 1 0 39312 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_347
timestamp 1698431365
transform 1 0 40208 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_360
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_368
timestamp 1698431365
transform 1 0 42560 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_372
timestamp 1698431365
transform 1 0 43008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_380
timestamp 1698431365
transform 1 0 43904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_18
timestamp 1698431365
transform 1 0 3360 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_49
timestamp 1698431365
transform 1 0 6832 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_65
timestamp 1698431365
transform 1 0 8624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_83
timestamp 1698431365
transform 1 0 10640 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_99
timestamp 1698431365
transform 1 0 12432 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_103
timestamp 1698431365
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_111
timestamp 1698431365
transform 1 0 13776 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_115
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_136
timestamp 1698431365
transform 1 0 16576 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_144
timestamp 1698431365
transform 1 0 17472 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_151
timestamp 1698431365
transform 1 0 18256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_163
timestamp 1698431365
transform 1 0 19600 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_234
timestamp 1698431365
transform 1 0 27552 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_257
timestamp 1698431365
transform 1 0 30128 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_265
timestamp 1698431365
transform 1 0 31024 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_269
timestamp 1698431365
transform 1 0 31472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_271
timestamp 1698431365
transform 1 0 31696 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_280
timestamp 1698431365
transform 1 0 32704 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_312
timestamp 1698431365
transform 1 0 36288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_333
timestamp 1698431365
transform 1 0 38640 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_341
timestamp 1698431365
transform 1 0 39536 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_343
timestamp 1698431365
transform 1 0 39760 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_352
timestamp 1698431365
transform 1 0 40768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_31
timestamp 1698431365
transform 1 0 4816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_35
timestamp 1698431365
transform 1 0 5264 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_43
timestamp 1698431365
transform 1 0 6160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_47
timestamp 1698431365
transform 1 0 6608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_49
timestamp 1698431365
transform 1 0 6832 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_67
timestamp 1698431365
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_83
timestamp 1698431365
transform 1 0 10640 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_91
timestamp 1698431365
transform 1 0 11536 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_115
timestamp 1698431365
transform 1 0 14224 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_131
timestamp 1698431365
transform 1 0 16016 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_144
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_153
timestamp 1698431365
transform 1 0 18480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_157
timestamp 1698431365
transform 1 0 18928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_165
timestamp 1698431365
transform 1 0 19824 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_195
timestamp 1698431365
transform 1 0 23184 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_203
timestamp 1698431365
transform 1 0 24080 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_228
timestamp 1698431365
transform 1 0 26880 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_240
timestamp 1698431365
transform 1 0 28224 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_244
timestamp 1698431365
transform 1 0 28672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_253
timestamp 1698431365
transform 1 0 29680 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_261
timestamp 1698431365
transform 1 0 30576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_263
timestamp 1698431365
transform 1 0 30800 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_274
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_286
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_288
timestamp 1698431365
transform 1 0 33600 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_304
timestamp 1698431365
transform 1 0 35392 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_316
timestamp 1698431365
transform 1 0 36736 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_320
timestamp 1698431365
transform 1 0 37184 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_327
timestamp 1698431365
transform 1 0 37968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_335
timestamp 1698431365
transform 1 0 38864 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_339
timestamp 1698431365
transform 1 0 39312 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_371
timestamp 1698431365
transform 1 0 42896 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_379
timestamp 1698431365
transform 1 0 43792 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_385
timestamp 1698431365
transform 1 0 44464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_389
timestamp 1698431365
transform 1 0 44912 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_395
timestamp 1698431365
transform 1 0 45584 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_409
timestamp 1698431365
transform 1 0 47152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_411
timestamp 1698431365
transform 1 0 47376 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_27
timestamp 1698431365
transform 1 0 4368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_43
timestamp 1698431365
transform 1 0 6160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_45
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_83
timestamp 1698431365
transform 1 0 10640 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698431365
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_131
timestamp 1698431365
transform 1 0 16016 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_139
timestamp 1698431365
transform 1 0 16912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_161
timestamp 1698431365
transform 1 0 19376 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_165
timestamp 1698431365
transform 1 0 19824 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_189
timestamp 1698431365
transform 1 0 22512 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_197
timestamp 1698431365
transform 1 0 23408 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_201
timestamp 1698431365
transform 1 0 23856 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_225
timestamp 1698431365
transform 1 0 26544 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_238
timestamp 1698431365
transform 1 0 28000 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698431365
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_256
timestamp 1698431365
transform 1 0 30016 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_273
timestamp 1698431365
transform 1 0 31920 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_277
timestamp 1698431365
transform 1 0 32368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_279
timestamp 1698431365
transform 1 0 32592 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_285
timestamp 1698431365
transform 1 0 33264 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_293
timestamp 1698431365
transform 1 0 34160 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_312
timestamp 1698431365
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_325
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_332
timestamp 1698431365
transform 1 0 38528 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_348
timestamp 1698431365
transform 1 0 40320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_352
timestamp 1698431365
transform 1 0 40768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_354
timestamp 1698431365
transform 1 0 40992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_361
timestamp 1698431365
transform 1 0 41776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_365
timestamp 1698431365
transform 1 0 42224 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_393
timestamp 1698431365
transform 1 0 45360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_403
timestamp 1698431365
transform 1 0 46480 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_413
timestamp 1698431365
transform 1 0 47600 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_6
timestamp 1698431365
transform 1 0 2016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_20
timestamp 1698431365
transform 1 0 3584 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_39
timestamp 1698431365
transform 1 0 5712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_41
timestamp 1698431365
transform 1 0 5936 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_46
timestamp 1698431365
transform 1 0 6496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_48
timestamp 1698431365
transform 1 0 6720 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_94
timestamp 1698431365
transform 1 0 11872 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_105
timestamp 1698431365
transform 1 0 13104 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_130
timestamp 1698431365
transform 1 0 15904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_134
timestamp 1698431365
transform 1 0 16352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_171
timestamp 1698431365
transform 1 0 20496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_173
timestamp 1698431365
transform 1 0 20720 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_203
timestamp 1698431365
transform 1 0 24080 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698431365
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_229
timestamp 1698431365
transform 1 0 26992 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_235
timestamp 1698431365
transform 1 0 27664 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_243
timestamp 1698431365
transform 1 0 28560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_299
timestamp 1698431365
transform 1 0 34832 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_315
timestamp 1698431365
transform 1 0 36624 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_339
timestamp 1698431365
transform 1 0 39312 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_347
timestamp 1698431365
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_368
timestamp 1698431365
transform 1 0 42560 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_398
timestamp 1698431365
transform 1 0 45920 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_400
timestamp 1698431365
transform 1 0 46144 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_403
timestamp 1698431365
transform 1 0 46480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_405
timestamp 1698431365
transform 1 0 46704 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_410
timestamp 1698431365
transform 1 0 47264 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_417
timestamp 1698431365
transform 1 0 48048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_419
timestamp 1698431365
transform 1 0 48272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_28
timestamp 1698431365
transform 1 0 4480 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_30
timestamp 1698431365
transform 1 0 4704 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_33
timestamp 1698431365
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_41
timestamp 1698431365
transform 1 0 5936 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_48
timestamp 1698431365
transform 1 0 6720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_50
timestamp 1698431365
transform 1 0 6944 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_64
timestamp 1698431365
transform 1 0 8512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_84
timestamp 1698431365
transform 1 0 10752 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_86
timestamp 1698431365
transform 1 0 10976 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_113
timestamp 1698431365
transform 1 0 14000 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_123
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_141
timestamp 1698431365
transform 1 0 17136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698431365
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_190
timestamp 1698431365
transform 1 0 22624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_194
timestamp 1698431365
transform 1 0 23072 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_210
timestamp 1698431365
transform 1 0 24864 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_219
timestamp 1698431365
transform 1 0 25872 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_227
timestamp 1698431365
transform 1 0 26768 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_231
timestamp 1698431365
transform 1 0 27216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_238
timestamp 1698431365
transform 1 0 28000 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_240
timestamp 1698431365
transform 1 0 28224 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_260
timestamp 1698431365
transform 1 0 30464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_262
timestamp 1698431365
transform 1 0 30688 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_289
timestamp 1698431365
transform 1 0 33712 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_293
timestamp 1698431365
transform 1 0 34160 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_296
timestamp 1698431365
transform 1 0 34496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_300
timestamp 1698431365
transform 1 0 34944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_302
timestamp 1698431365
transform 1 0 35168 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_325
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_334
timestamp 1698431365
transform 1 0 38752 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_342
timestamp 1698431365
transform 1 0 39648 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_346
timestamp 1698431365
transform 1 0 40096 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_372
timestamp 1698431365
transform 1 0 43008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_384
timestamp 1698431365
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_37
timestamp 1698431365
transform 1 0 5488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_41
timestamp 1698431365
transform 1 0 5936 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_43
timestamp 1698431365
transform 1 0 6160 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_76
timestamp 1698431365
transform 1 0 9856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_78
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_113
timestamp 1698431365
transform 1 0 14000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_123
timestamp 1698431365
transform 1 0 15120 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_125
timestamp 1698431365
transform 1 0 15344 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_185
timestamp 1698431365
transform 1 0 22064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_205
timestamp 1698431365
transform 1 0 24304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_233
timestamp 1698431365
transform 1 0 27440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_247
timestamp 1698431365
transform 1 0 29008 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_251
timestamp 1698431365
transform 1 0 29456 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_294
timestamp 1698431365
transform 1 0 34272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_325
timestamp 1698431365
transform 1 0 37744 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_348
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_391
timestamp 1698431365
transform 1 0 45136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_393
timestamp 1698431365
transform 1 0 45360 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698431365
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_39
timestamp 1698431365
transform 1 0 5712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_42
timestamp 1698431365
transform 1 0 6048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_44
timestamp 1698431365
transform 1 0 6272 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_54
timestamp 1698431365
transform 1 0 7392 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_70
timestamp 1698431365
transform 1 0 9184 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_78
timestamp 1698431365
transform 1 0 10080 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698431365
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_115
timestamp 1698431365
transform 1 0 14224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_117
timestamp 1698431365
transform 1 0 14448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_146
timestamp 1698431365
transform 1 0 17696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_148
timestamp 1698431365
transform 1 0 17920 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_181
timestamp 1698431365
transform 1 0 21616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_187
timestamp 1698431365
transform 1 0 22288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_192
timestamp 1698431365
transform 1 0 22848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_196
timestamp 1698431365
transform 1 0 23296 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_206
timestamp 1698431365
transform 1 0 24416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_210
timestamp 1698431365
transform 1 0 24864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_212
timestamp 1698431365
transform 1 0 25088 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_229
timestamp 1698431365
transform 1 0 26992 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_270
timestamp 1698431365
transform 1 0 31584 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_286
timestamp 1698431365
transform 1 0 33376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_300
timestamp 1698431365
transform 1 0 34944 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_304
timestamp 1698431365
transform 1 0 35392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_306
timestamp 1698431365
transform 1 0 35616 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_319
timestamp 1698431365
transform 1 0 37072 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_354
timestamp 1698431365
transform 1 0 40992 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_362
timestamp 1698431365
transform 1 0 41888 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_378
timestamp 1698431365
transform 1 0 43680 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_380
timestamp 1698431365
transform 1 0 43904 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_411
timestamp 1698431365
transform 1 0 47376 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_418
timestamp 1698431365
transform 1 0 48160 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_10
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_46
timestamp 1698431365
transform 1 0 6496 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_56
timestamp 1698431365
transform 1 0 7616 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_76
timestamp 1698431365
transform 1 0 9856 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_93
timestamp 1698431365
transform 1 0 11760 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_101
timestamp 1698431365
transform 1 0 12656 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_105
timestamp 1698431365
transform 1 0 13104 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_117
timestamp 1698431365
transform 1 0 14448 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_121
timestamp 1698431365
transform 1 0 14896 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698431365
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_158
timestamp 1698431365
transform 1 0 19040 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_188
timestamp 1698431365
transform 1 0 22400 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_196
timestamp 1698431365
transform 1 0 23296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_216
timestamp 1698431365
transform 1 0 25536 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_224
timestamp 1698431365
transform 1 0 26432 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_244
timestamp 1698431365
transform 1 0 28672 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_248
timestamp 1698431365
transform 1 0 29120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_250
timestamp 1698431365
transform 1 0 29344 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_292
timestamp 1698431365
transform 1 0 34048 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_308
timestamp 1698431365
transform 1 0 35840 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_312
timestamp 1698431365
transform 1 0 36288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_314
timestamp 1698431365
transform 1 0 36512 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_344
timestamp 1698431365
transform 1 0 39872 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_348
timestamp 1698431365
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_364
timestamp 1698431365
transform 1 0 42112 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_366
timestamp 1698431365
transform 1 0 42336 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_399
timestamp 1698431365
transform 1 0 46032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_403
timestamp 1698431365
transform 1 0 46480 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_10
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_17
timestamp 1698431365
transform 1 0 3248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_21
timestamp 1698431365
transform 1 0 3696 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_29
timestamp 1698431365
transform 1 0 4592 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_33
timestamp 1698431365
transform 1 0 5040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_43
timestamp 1698431365
transform 1 0 6160 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_59
timestamp 1698431365
transform 1 0 7952 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_72
timestamp 1698431365
transform 1 0 9408 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_79
timestamp 1698431365
transform 1 0 10192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_99
timestamp 1698431365
transform 1 0 12432 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_109
timestamp 1698431365
transform 1 0 13552 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_114
timestamp 1698431365
transform 1 0 14112 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_116
timestamp 1698431365
transform 1 0 14336 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_125
timestamp 1698431365
transform 1 0 15344 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_133
timestamp 1698431365
transform 1 0 16240 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_137
timestamp 1698431365
transform 1 0 16688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_143
timestamp 1698431365
transform 1 0 17360 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_159
timestamp 1698431365
transform 1 0 19152 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_209
timestamp 1698431365
transform 1 0 24752 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_221
timestamp 1698431365
transform 1 0 26096 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_225
timestamp 1698431365
transform 1 0 26544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_233
timestamp 1698431365
transform 1 0 27440 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_253
timestamp 1698431365
transform 1 0 29680 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_262
timestamp 1698431365
transform 1 0 30688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_264
timestamp 1698431365
transform 1 0 30912 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_294
timestamp 1698431365
transform 1 0 34272 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_310
timestamp 1698431365
transform 1 0 36064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_321
timestamp 1698431365
transform 1 0 37296 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_329
timestamp 1698431365
transform 1 0 38192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_375
timestamp 1698431365
transform 1 0 43344 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_381
timestamp 1698431365
transform 1 0 44016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_417
timestamp 1698431365
transform 1 0 48048 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_419
timestamp 1698431365
transform 1 0 48272 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_31
timestamp 1698431365
transform 1 0 4816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_35
timestamp 1698431365
transform 1 0 5264 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_50
timestamp 1698431365
transform 1 0 6944 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_58
timestamp 1698431365
transform 1 0 7840 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_92
timestamp 1698431365
transform 1 0 11648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_94
timestamp 1698431365
transform 1 0 11872 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_124
timestamp 1698431365
transform 1 0 15232 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_128
timestamp 1698431365
transform 1 0 15680 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_146
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_177
timestamp 1698431365
transform 1 0 21168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_179
timestamp 1698431365
transform 1 0 21392 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_241
timestamp 1698431365
transform 1 0 28336 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_272
timestamp 1698431365
transform 1 0 31808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_326
timestamp 1698431365
transform 1 0 37856 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_334
timestamp 1698431365
transform 1 0 38752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_341
timestamp 1698431365
transform 1 0 39536 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_356
timestamp 1698431365
transform 1 0 41216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_358
timestamp 1698431365
transform 1 0 41440 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_412
timestamp 1698431365
transform 1 0 47488 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_24
timestamp 1698431365
transform 1 0 4032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_26
timestamp 1698431365
transform 1 0 4256 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_39
timestamp 1698431365
transform 1 0 5712 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_81
timestamp 1698431365
transform 1 0 10416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_85
timestamp 1698431365
transform 1 0 10864 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_89
timestamp 1698431365
transform 1 0 11312 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698431365
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_113
timestamp 1698431365
transform 1 0 14000 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_130
timestamp 1698431365
transform 1 0 15904 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_181
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_183
timestamp 1698431365
transform 1 0 21840 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_204
timestamp 1698431365
transform 1 0 24192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_206
timestamp 1698431365
transform 1 0 24416 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_215
timestamp 1698431365
transform 1 0 25424 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_231
timestamp 1698431365
transform 1 0 27216 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_239
timestamp 1698431365
transform 1 0 28112 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_271
timestamp 1698431365
transform 1 0 31696 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_303
timestamp 1698431365
transform 1 0 35280 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_372
timestamp 1698431365
transform 1 0 43008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_374
timestamp 1698431365
transform 1 0 43232 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_383
timestamp 1698431365
transform 1 0 44240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_28
timestamp 1698431365
transform 1 0 4480 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_32
timestamp 1698431365
transform 1 0 4928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_34
timestamp 1698431365
transform 1 0 5152 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_57
timestamp 1698431365
transform 1 0 7728 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_59
timestamp 1698431365
transform 1 0 7952 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_88
timestamp 1698431365
transform 1 0 11200 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_97
timestamp 1698431365
transform 1 0 12208 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_102
timestamp 1698431365
transform 1 0 12768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_104
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_107
timestamp 1698431365
transform 1 0 13328 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_115
timestamp 1698431365
transform 1 0 14224 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_125
timestamp 1698431365
transform 1 0 15344 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_133
timestamp 1698431365
transform 1 0 16240 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698431365
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_162
timestamp 1698431365
transform 1 0 19488 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_194
timestamp 1698431365
transform 1 0 23072 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_200
timestamp 1698431365
transform 1 0 23744 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_204
timestamp 1698431365
transform 1 0 24192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_228
timestamp 1698431365
transform 1 0 26880 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_232
timestamp 1698431365
transform 1 0 27328 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_234
timestamp 1698431365
transform 1 0 27552 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_239
timestamp 1698431365
transform 1 0 28112 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_255
timestamp 1698431365
transform 1 0 29904 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_259
timestamp 1698431365
transform 1 0 30352 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_261
timestamp 1698431365
transform 1 0 30576 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_298
timestamp 1698431365
transform 1 0 34720 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_330
timestamp 1698431365
transform 1 0 38304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_342
timestamp 1698431365
transform 1 0 39648 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698431365
transform 1 0 40096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_358
timestamp 1698431365
transform 1 0 41440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_368
timestamp 1698431365
transform 1 0 42560 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_372
timestamp 1698431365
transform 1 0 43008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_374
timestamp 1698431365
transform 1 0 43232 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_31
timestamp 1698431365
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_41
timestamp 1698431365
transform 1 0 5936 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_46
timestamp 1698431365
transform 1 0 6496 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_54
timestamp 1698431365
transform 1 0 7392 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_58
timestamp 1698431365
transform 1 0 7840 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698431365
transform 1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_119
timestamp 1698431365
transform 1 0 14672 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_135
timestamp 1698431365
transform 1 0 16464 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_181
timestamp 1698431365
transform 1 0 21616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_202
timestamp 1698431365
transform 1 0 23968 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_220
timestamp 1698431365
transform 1 0 25984 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698431365
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_255
timestamp 1698431365
transform 1 0 29904 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_262
timestamp 1698431365
transform 1 0 30688 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_266
timestamp 1698431365
transform 1 0 31136 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_275
timestamp 1698431365
transform 1 0 32144 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_279
timestamp 1698431365
transform 1 0 32592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_281
timestamp 1698431365
transform 1 0 32816 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_306
timestamp 1698431365
transform 1 0 35616 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698431365
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_323
timestamp 1698431365
transform 1 0 37520 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_335
timestamp 1698431365
transform 1 0 38864 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_339
timestamp 1698431365
transform 1 0 39312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_375
timestamp 1698431365
transform 1 0 43344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_379
timestamp 1698431365
transform 1 0 43792 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_383
timestamp 1698431365
transform 1 0 44240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_393
timestamp 1698431365
transform 1 0 45360 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_18
timestamp 1698431365
transform 1 0 3360 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_22
timestamp 1698431365
transform 1 0 3808 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_26
timestamp 1698431365
transform 1 0 4256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_40
timestamp 1698431365
transform 1 0 5824 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_48
timestamp 1698431365
transform 1 0 6720 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_56
timestamp 1698431365
transform 1 0 7616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_60
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_62
timestamp 1698431365
transform 1 0 8288 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_80
timestamp 1698431365
transform 1 0 10304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_96
timestamp 1698431365
transform 1 0 12096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_100
timestamp 1698431365
transform 1 0 12544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_104
timestamp 1698431365
transform 1 0 12992 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_108
timestamp 1698431365
transform 1 0 13440 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_158
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_162
timestamp 1698431365
transform 1 0 19488 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_166
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_168
timestamp 1698431365
transform 1 0 20160 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_198
timestamp 1698431365
transform 1 0 23520 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698431365
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_241
timestamp 1698431365
transform 1 0 28336 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_249
timestamp 1698431365
transform 1 0 29232 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_253
timestamp 1698431365
transform 1 0 29680 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698431365
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_292
timestamp 1698431365
transform 1 0 34048 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_296
timestamp 1698431365
transform 1 0 34496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_342
timestamp 1698431365
transform 1 0 39648 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_360
timestamp 1698431365
transform 1 0 41664 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_380
timestamp 1698431365
transform 1 0 43904 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_384
timestamp 1698431365
transform 1 0 44352 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_42
timestamp 1698431365
transform 1 0 6048 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_46
timestamp 1698431365
transform 1 0 6496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_64
timestamp 1698431365
transform 1 0 8512 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_80
timestamp 1698431365
transform 1 0 10304 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_88
timestamp 1698431365
transform 1 0 11200 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_92
timestamp 1698431365
transform 1 0 11648 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_103
timestamp 1698431365
transform 1 0 12880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_123
timestamp 1698431365
transform 1 0 15120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_125
timestamp 1698431365
transform 1 0 15344 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_132
timestamp 1698431365
transform 1 0 16128 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_148
timestamp 1698431365
transform 1 0 17920 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_154
timestamp 1698431365
transform 1 0 18592 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_168
timestamp 1698431365
transform 1 0 20160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_181
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_183
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_213
timestamp 1698431365
transform 1 0 25200 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_224
timestamp 1698431365
transform 1 0 26432 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_228
timestamp 1698431365
transform 1 0 26880 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_236
timestamp 1698431365
transform 1 0 27776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_238
timestamp 1698431365
transform 1 0 28000 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_259
timestamp 1698431365
transform 1 0 30352 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_275
timestamp 1698431365
transform 1 0 32144 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_283
timestamp 1698431365
transform 1 0 33040 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_292
timestamp 1698431365
transform 1 0 34048 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_308
timestamp 1698431365
transform 1 0 35840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698431365
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_329
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_345
timestamp 1698431365
transform 1 0 39984 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_369
timestamp 1698431365
transform 1 0 42672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_374
timestamp 1698431365
transform 1 0 43232 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_382
timestamp 1698431365
transform 1 0 44128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_415
timestamp 1698431365
transform 1 0 47824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_419
timestamp 1698431365
transform 1 0 48272 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_28
timestamp 1698431365
transform 1 0 4480 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_32
timestamp 1698431365
transform 1 0 4928 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_65
timestamp 1698431365
transform 1 0 8624 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_78
timestamp 1698431365
transform 1 0 10080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_82
timestamp 1698431365
transform 1 0 10528 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_150
timestamp 1698431365
transform 1 0 18144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_183
timestamp 1698431365
transform 1 0 21840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_196
timestamp 1698431365
transform 1 0 23296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_200
timestamp 1698431365
transform 1 0 23744 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_262
timestamp 1698431365
transform 1 0 30688 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698431365
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_292
timestamp 1698431365
transform 1 0 34048 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_308
timestamp 1698431365
transform 1 0 35840 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_316
timestamp 1698431365
transform 1 0 36736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_320
timestamp 1698431365
transform 1 0 37184 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_345
timestamp 1698431365
transform 1 0 39984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_381
timestamp 1698431365
transform 1 0 44016 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_389
timestamp 1698431365
transform 1 0 44912 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_393
timestamp 1698431365
transform 1 0 45360 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_416
timestamp 1698431365
transform 1 0 47936 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_31
timestamp 1698431365
transform 1 0 4816 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_49
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_53
timestamp 1698431365
transform 1 0 7280 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_95
timestamp 1698431365
transform 1 0 11984 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_103
timestamp 1698431365
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_115
timestamp 1698431365
transform 1 0 14224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_119
timestamp 1698431365
transform 1 0 14672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_151
timestamp 1698431365
transform 1 0 18256 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_161
timestamp 1698431365
transform 1 0 19376 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_169
timestamp 1698431365
transform 1 0 20272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698431365
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_189
timestamp 1698431365
transform 1 0 22512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_196
timestamp 1698431365
transform 1 0 23296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_204
timestamp 1698431365
transform 1 0 24192 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_284
timestamp 1698431365
transform 1 0 33152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_323
timestamp 1698431365
transform 1 0 37520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_403
timestamp 1698431365
transform 1 0 46480 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_405
timestamp 1698431365
transform 1 0 46704 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_18
timestamp 1698431365
transform 1 0 3360 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_26
timestamp 1698431365
transform 1 0 4256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_28
timestamp 1698431365
transform 1 0 4480 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_45
timestamp 1698431365
transform 1 0 6384 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_49
timestamp 1698431365
transform 1 0 6832 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_56
timestamp 1698431365
transform 1 0 7616 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_63
timestamp 1698431365
transform 1 0 8400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_67
timestamp 1698431365
transform 1 0 8848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_104
timestamp 1698431365
transform 1 0 12992 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_120
timestamp 1698431365
transform 1 0 14784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_122
timestamp 1698431365
transform 1 0 15008 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_151
timestamp 1698431365
transform 1 0 18256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_169
timestamp 1698431365
transform 1 0 20272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_173
timestamp 1698431365
transform 1 0 20720 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_181
timestamp 1698431365
transform 1 0 21616 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_190
timestamp 1698431365
transform 1 0 22624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_194
timestamp 1698431365
transform 1 0 23072 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_226
timestamp 1698431365
transform 1 0 26656 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_258
timestamp 1698431365
transform 1 0 30240 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_292
timestamp 1698431365
transform 1 0 34048 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_300
timestamp 1698431365
transform 1 0 34944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_347
timestamp 1698431365
transform 1 0 40208 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_349
timestamp 1698431365
transform 1 0 40432 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_385
timestamp 1698431365
transform 1 0 44464 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_55
timestamp 1698431365
transform 1 0 7504 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_58
timestamp 1698431365
transform 1 0 7840 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_148
timestamp 1698431365
transform 1 0 17920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_156
timestamp 1698431365
transform 1 0 18816 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698431365
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_187
timestamp 1698431365
transform 1 0 22288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_191
timestamp 1698431365
transform 1 0 22736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_193
timestamp 1698431365
transform 1 0 22960 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_208
timestamp 1698431365
transform 1 0 24640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_212
timestamp 1698431365
transform 1 0 25088 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_222
timestamp 1698431365
transform 1 0 26208 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698431365
transform 1 0 28000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_251
timestamp 1698431365
transform 1 0 29456 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_254
timestamp 1698431365
transform 1 0 29792 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_262
timestamp 1698431365
transform 1 0 30688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_272
timestamp 1698431365
transform 1 0 31808 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_276
timestamp 1698431365
transform 1 0 32256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_278
timestamp 1698431365
transform 1 0 32480 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_285
timestamp 1698431365
transform 1 0 33264 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_301
timestamp 1698431365
transform 1 0 35056 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_305
timestamp 1698431365
transform 1 0 35504 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_325
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_393
timestamp 1698431365
transform 1 0 45360 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_31
timestamp 1698431365
transform 1 0 4816 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_89
timestamp 1698431365
transform 1 0 11312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_97
timestamp 1698431365
transform 1 0 12208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_101
timestamp 1698431365
transform 1 0 12656 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_115
timestamp 1698431365
transform 1 0 14224 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_123
timestamp 1698431365
transform 1 0 15120 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_134
timestamp 1698431365
transform 1 0 16352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_165
timestamp 1698431365
transform 1 0 19824 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_195
timestamp 1698431365
transform 1 0 23184 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_270
timestamp 1698431365
transform 1 0 31584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_311
timestamp 1698431365
transform 1 0 36176 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_319
timestamp 1698431365
transform 1 0 37072 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_354
timestamp 1698431365
transform 1 0 40992 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_360
timestamp 1698431365
transform 1 0 41664 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_390
timestamp 1698431365
transform 1 0 45024 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_48
timestamp 1698431365
transform 1 0 6720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_50
timestamp 1698431365
transform 1 0 6944 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_78
timestamp 1698431365
transform 1 0 10080 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_86
timestamp 1698431365
transform 1 0 10976 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_90
timestamp 1698431365
transform 1 0 11424 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_103
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_112
timestamp 1698431365
transform 1 0 13888 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_183
timestamp 1698431365
transform 1 0 21840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_187
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_195
timestamp 1698431365
transform 1 0 23184 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_199
timestamp 1698431365
transform 1 0 23632 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_201
timestamp 1698431365
transform 1 0 23856 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_207
timestamp 1698431365
transform 1 0 24528 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_239
timestamp 1698431365
transform 1 0 28112 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698431365
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_276
timestamp 1698431365
transform 1 0 32256 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_308
timestamp 1698431365
transform 1 0 35840 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_312
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_329
timestamp 1698431365
transform 1 0 38192 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_343
timestamp 1698431365
transform 1 0 39760 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_351
timestamp 1698431365
transform 1 0 40656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_355
timestamp 1698431365
transform 1 0 41104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_363
timestamp 1698431365
transform 1 0 42000 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_371
timestamp 1698431365
transform 1 0 42896 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_375
timestamp 1698431365
transform 1 0 43344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_377
timestamp 1698431365
transform 1 0 43568 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_403
timestamp 1698431365
transform 1 0 46480 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_419
timestamp 1698431365
transform 1 0 48272 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_6
timestamp 1698431365
transform 1 0 2016 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_8
timestamp 1698431365
transform 1 0 2240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_15
timestamp 1698431365
transform 1 0 3024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_19
timestamp 1698431365
transform 1 0 3472 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_35
timestamp 1698431365
transform 1 0 5264 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_37
timestamp 1698431365
transform 1 0 5488 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_46
timestamp 1698431365
transform 1 0 6496 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_62
timestamp 1698431365
transform 1 0 8288 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_76
timestamp 1698431365
transform 1 0 9856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_92
timestamp 1698431365
transform 1 0 11648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_96
timestamp 1698431365
transform 1 0 12096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_100
timestamp 1698431365
transform 1 0 12544 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_103
timestamp 1698431365
transform 1 0 12880 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_107
timestamp 1698431365
transform 1 0 13328 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_110
timestamp 1698431365
transform 1 0 13664 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_137
timestamp 1698431365
transform 1 0 16688 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_146
timestamp 1698431365
transform 1 0 17696 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_158
timestamp 1698431365
transform 1 0 19040 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_176
timestamp 1698431365
transform 1 0 21056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_180
timestamp 1698431365
transform 1 0 21504 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_196
timestamp 1698431365
transform 1 0 23296 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_204
timestamp 1698431365
transform 1 0 24192 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_208
timestamp 1698431365
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_224
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_254
timestamp 1698431365
transform 1 0 29792 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_270
timestamp 1698431365
transform 1 0 31584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_272
timestamp 1698431365
transform 1 0 31808 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_278
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_286
timestamp 1698431365
transform 1 0 33376 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_294
timestamp 1698431365
transform 1 0 34272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_301
timestamp 1698431365
transform 1 0 35056 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_323
timestamp 1698431365
transform 1 0 37520 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_327
timestamp 1698431365
transform 1 0 37968 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_336
timestamp 1698431365
transform 1 0 38976 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_344
timestamp 1698431365
transform 1 0 39872 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_372
timestamp 1698431365
transform 1 0 43008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_374
timestamp 1698431365
transform 1 0 43232 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_10
timestamp 1698431365
transform 1 0 2464 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_19
timestamp 1698431365
transform 1 0 3472 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_23
timestamp 1698431365
transform 1 0 3920 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_33
timestamp 1698431365
transform 1 0 5040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_43
timestamp 1698431365
transform 1 0 6160 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_59
timestamp 1698431365
transform 1 0 7952 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_67
timestamp 1698431365
transform 1 0 8848 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_71
timestamp 1698431365
transform 1 0 9296 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698431365
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_115
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_135
timestamp 1698431365
transform 1 0 16464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_156
timestamp 1698431365
transform 1 0 18816 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_162
timestamp 1698431365
transform 1 0 19488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_166
timestamp 1698431365
transform 1 0 19936 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_208
timestamp 1698431365
transform 1 0 24640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_210
timestamp 1698431365
transform 1 0 24864 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_227
timestamp 1698431365
transform 1 0 26768 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_243
timestamp 1698431365
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_255
timestamp 1698431365
transform 1 0 29904 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_262
timestamp 1698431365
transform 1 0 30688 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_266
timestamp 1698431365
transform 1 0 31136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_280
timestamp 1698431365
transform 1 0 32704 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_300
timestamp 1698431365
transform 1 0 34944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_312
timestamp 1698431365
transform 1 0 36288 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_326
timestamp 1698431365
transform 1 0 37856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_330
timestamp 1698431365
transform 1 0 38304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_369
timestamp 1698431365
transform 1 0 42672 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_377
timestamp 1698431365
transform 1 0 43568 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_383
timestamp 1698431365
transform 1 0 44240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_419
timestamp 1698431365
transform 1 0 48272 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_31
timestamp 1698431365
transform 1 0 4816 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_47
timestamp 1698431365
transform 1 0 6608 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_51
timestamp 1698431365
transform 1 0 7056 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_57
timestamp 1698431365
transform 1 0 7728 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_61
timestamp 1698431365
transform 1 0 8176 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_74
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_101
timestamp 1698431365
transform 1 0 12656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_118
timestamp 1698431365
transform 1 0 14560 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_120
timestamp 1698431365
transform 1 0 14784 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_130
timestamp 1698431365
transform 1 0 15904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_177
timestamp 1698431365
transform 1 0 21168 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_220
timestamp 1698431365
transform 1 0 25984 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_238
timestamp 1698431365
transform 1 0 28000 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_246
timestamp 1698431365
transform 1 0 28896 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_268
timestamp 1698431365
transform 1 0 31360 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_298
timestamp 1698431365
transform 1 0 34720 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_330
timestamp 1698431365
transform 1 0 38304 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698431365
transform 1 0 40096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_384
timestamp 1698431365
transform 1 0 44352 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_392
timestamp 1698431365
transform 1 0 45248 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_401
timestamp 1698431365
transform 1 0 46256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_405
timestamp 1698431365
transform 1 0 46704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_409
timestamp 1698431365
transform 1 0 47152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_413
timestamp 1698431365
transform 1 0 47600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_417
timestamp 1698431365
transform 1 0 48048 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_10
timestamp 1698431365
transform 1 0 2464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_14
timestamp 1698431365
transform 1 0 2912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_22
timestamp 1698431365
transform 1 0 3808 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_30
timestamp 1698431365
transform 1 0 4704 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_66
timestamp 1698431365
transform 1 0 8736 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_75
timestamp 1698431365
transform 1 0 9744 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_102
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_113
timestamp 1698431365
transform 1 0 14000 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_183
timestamp 1698431365
transform 1 0 21840 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_187
timestamp 1698431365
transform 1 0 22288 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_191
timestamp 1698431365
transform 1 0 22736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_193
timestamp 1698431365
transform 1 0 22960 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_203
timestamp 1698431365
transform 1 0 24080 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_235
timestamp 1698431365
transform 1 0 27664 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_243
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_285
timestamp 1698431365
transform 1 0 33264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_287
timestamp 1698431365
transform 1 0 33488 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_306
timestamp 1698431365
transform 1 0 35616 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_310
timestamp 1698431365
transform 1 0 36064 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_313
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_321
timestamp 1698431365
transform 1 0 37296 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_325
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_329
timestamp 1698431365
transform 1 0 38192 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_333
timestamp 1698431365
transform 1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_335
timestamp 1698431365
transform 1 0 38864 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_365
timestamp 1698431365
transform 1 0 42224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_367
timestamp 1698431365
transform 1 0 42448 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_376
timestamp 1698431365
transform 1 0 43456 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_10
timestamp 1698431365
transform 1 0 2464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_18
timestamp 1698431365
transform 1 0 3360 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_22
timestamp 1698431365
transform 1 0 3808 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_26
timestamp 1698431365
transform 1 0 4256 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_28
timestamp 1698431365
transform 1 0 4480 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_43
timestamp 1698431365
transform 1 0 6160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_47
timestamp 1698431365
transform 1 0 6608 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_74
timestamp 1698431365
transform 1 0 9632 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_89
timestamp 1698431365
transform 1 0 11312 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698431365
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_148
timestamp 1698431365
transform 1 0 17920 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_181
timestamp 1698431365
transform 1 0 21616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_197
timestamp 1698431365
transform 1 0 23408 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_224
timestamp 1698431365
transform 1 0 26432 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_232
timestamp 1698431365
transform 1 0 27328 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_240
timestamp 1698431365
transform 1 0 28224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_292
timestamp 1698431365
transform 1 0 34048 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_296
timestamp 1698431365
transform 1 0 34496 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_327
timestamp 1698431365
transform 1 0 37968 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_340
timestamp 1698431365
transform 1 0 39424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_372
timestamp 1698431365
transform 1 0 43008 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_376
timestamp 1698431365
transform 1 0 43456 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_383
timestamp 1698431365
transform 1 0 44240 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_411
timestamp 1698431365
transform 1 0 47376 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_418
timestamp 1698431365
transform 1 0 48160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_33
timestamp 1698431365
transform 1 0 5040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_49
timestamp 1698431365
transform 1 0 6832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_51
timestamp 1698431365
transform 1 0 7056 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_56
timestamp 1698431365
transform 1 0 7616 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_72
timestamp 1698431365
transform 1 0 9408 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_82
timestamp 1698431365
transform 1 0 10528 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_84
timestamp 1698431365
transform 1 0 10752 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_117
timestamp 1698431365
transform 1 0 14448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_150
timestamp 1698431365
transform 1 0 18144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_154
timestamp 1698431365
transform 1 0 18592 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_168
timestamp 1698431365
transform 1 0 20160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_172
timestamp 1698431365
transform 1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_185
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_189
timestamp 1698431365
transform 1 0 22512 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_238
timestamp 1698431365
transform 1 0 28000 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_242
timestamp 1698431365
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698431365
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_255
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_257
timestamp 1698431365
transform 1 0 30128 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_371
timestamp 1698431365
transform 1 0 42896 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_8
timestamp 1698431365
transform 1 0 2240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_12
timestamp 1698431365
transform 1 0 2688 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_20
timestamp 1698431365
transform 1 0 3584 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_58
timestamp 1698431365
transform 1 0 7840 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_62
timestamp 1698431365
transform 1 0 8288 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_76
timestamp 1698431365
transform 1 0 9856 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_89
timestamp 1698431365
transform 1 0 11312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_138
timestamp 1698431365
transform 1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_144
timestamp 1698431365
transform 1 0 17472 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_171
timestamp 1698431365
transform 1 0 20496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_175
timestamp 1698431365
transform 1 0 20944 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_207
timestamp 1698431365
transform 1 0 24528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_209
timestamp 1698431365
transform 1 0 24752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_244
timestamp 1698431365
transform 1 0 28672 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_260
timestamp 1698431365
transform 1 0 30464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_293
timestamp 1698431365
transform 1 0 34160 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_309
timestamp 1698431365
transform 1 0 35952 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_313
timestamp 1698431365
transform 1 0 36400 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_315
timestamp 1698431365
transform 1 0 36624 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_385
timestamp 1698431365
transform 1 0 44464 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_408
timestamp 1698431365
transform 1 0 47040 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_417
timestamp 1698431365
transform 1 0 48048 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_419
timestamp 1698431365
transform 1 0 48272 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_28
timestamp 1698431365
transform 1 0 4480 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_53
timestamp 1698431365
transform 1 0 7280 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_113
timestamp 1698431365
transform 1 0 14000 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_115
timestamp 1698431365
transform 1 0 14224 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_158
timestamp 1698431365
transform 1 0 19040 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_167
timestamp 1698431365
transform 1 0 20048 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_197
timestamp 1698431365
transform 1 0 23408 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_205
timestamp 1698431365
transform 1 0 24304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_213
timestamp 1698431365
transform 1 0 25200 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_217
timestamp 1698431365
transform 1 0 25648 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_224
timestamp 1698431365
transform 1 0 26432 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_228
timestamp 1698431365
transform 1 0 26880 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_276
timestamp 1698431365
transform 1 0 32256 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_284
timestamp 1698431365
transform 1 0 33152 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_292
timestamp 1698431365
transform 1 0 34048 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_302
timestamp 1698431365
transform 1 0 35168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_310
timestamp 1698431365
transform 1 0 36064 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_356
timestamp 1698431365
transform 1 0 41216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_360
timestamp 1698431365
transform 1 0 41664 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_364
timestamp 1698431365
transform 1 0 42112 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_367
timestamp 1698431365
transform 1 0 42448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_371
timestamp 1698431365
transform 1 0 42896 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_39
timestamp 1698431365
transform 1 0 5712 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_43
timestamp 1698431365
transform 1 0 6160 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_97
timestamp 1698431365
transform 1 0 12208 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_105
timestamp 1698431365
transform 1 0 13104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_109
timestamp 1698431365
transform 1 0 13552 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_146
timestamp 1698431365
transform 1 0 17696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_232
timestamp 1698431365
transform 1 0 27328 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_248
timestamp 1698431365
transform 1 0 29120 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_256
timestamp 1698431365
transform 1 0 30016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_284
timestamp 1698431365
transform 1 0 33152 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_322
timestamp 1698431365
transform 1 0 37408 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_338
timestamp 1698431365
transform 1 0 39200 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_354
timestamp 1698431365
transform 1 0 40992 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_357
timestamp 1698431365
transform 1 0 41328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_361
timestamp 1698431365
transform 1 0 41776 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_363
timestamp 1698431365
transform 1 0 42000 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_366
timestamp 1698431365
transform 1 0 42336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_382
timestamp 1698431365
transform 1 0 44128 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_42
timestamp 1698431365
transform 1 0 6048 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_46
timestamp 1698431365
transform 1 0 6496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_50
timestamp 1698431365
transform 1 0 6944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_60
timestamp 1698431365
transform 1 0 8064 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_66
timestamp 1698431365
transform 1 0 8736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_72
timestamp 1698431365
transform 1 0 9408 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_80
timestamp 1698431365
transform 1 0 10304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_82
timestamp 1698431365
transform 1 0 10528 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_87
timestamp 1698431365
transform 1 0 11088 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_95
timestamp 1698431365
transform 1 0 11984 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_99
timestamp 1698431365
transform 1 0 12432 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_112
timestamp 1698431365
transform 1 0 13888 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_116
timestamp 1698431365
transform 1 0 14336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_118
timestamp 1698431365
transform 1 0 14560 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_156
timestamp 1698431365
transform 1 0 18816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_162
timestamp 1698431365
transform 1 0 19488 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_185
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_194
timestamp 1698431365
transform 1 0 23072 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_209
timestamp 1698431365
transform 1 0 24752 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_213
timestamp 1698431365
transform 1 0 25200 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_215
timestamp 1698431365
transform 1 0 25424 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_251
timestamp 1698431365
transform 1 0 29456 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_282
timestamp 1698431365
transform 1 0 32928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_286
timestamp 1698431365
transform 1 0 33376 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_302
timestamp 1698431365
transform 1 0 35168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_304
timestamp 1698431365
transform 1 0 35392 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_309
timestamp 1698431365
transform 1 0 35952 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_321
timestamp 1698431365
transform 1 0 37296 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_323
timestamp 1698431365
transform 1 0 37520 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_332
timestamp 1698431365
transform 1 0 38528 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_348
timestamp 1698431365
transform 1 0 40320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_352
timestamp 1698431365
transform 1 0 40768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_356
timestamp 1698431365
transform 1 0 41216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_358
timestamp 1698431365
transform 1 0 41440 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_367
timestamp 1698431365
transform 1 0 42448 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_28
timestamp 1698431365
transform 1 0 4480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_30
timestamp 1698431365
transform 1 0 4704 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_37
timestamp 1698431365
transform 1 0 5488 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_45
timestamp 1698431365
transform 1 0 6384 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_64
timestamp 1698431365
transform 1 0 8512 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_68
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_112
timestamp 1698431365
transform 1 0 13888 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_132
timestamp 1698431365
transform 1 0 16128 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_158
timestamp 1698431365
transform 1 0 19040 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698431365
transform 1 0 19488 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_192
timestamp 1698431365
transform 1 0 22848 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_226
timestamp 1698431365
transform 1 0 26656 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698431365
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698431365
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698431365
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_306
timestamp 1698431365
transform 1 0 35616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_316
timestamp 1698431365
transform 1 0 36736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_318
timestamp 1698431365
transform 1 0 36960 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_348
timestamp 1698431365
transform 1 0 40320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_381
timestamp 1698431365
transform 1 0 44016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_385
timestamp 1698431365
transform 1 0 44464 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_31
timestamp 1698431365
transform 1 0 4816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_48
timestamp 1698431365
transform 1 0 6720 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_97
timestamp 1698431365
transform 1 0 12208 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_111
timestamp 1698431365
transform 1 0 13776 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_114
timestamp 1698431365
transform 1 0 14112 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_146
timestamp 1698431365
transform 1 0 17696 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_162
timestamp 1698431365
transform 1 0 19488 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698431365
transform 1 0 20608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698431365
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_213
timestamp 1698431365
transform 1 0 25200 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_243
timestamp 1698431365
transform 1 0 28560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_251
timestamp 1698431365
transform 1 0 29456 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_253
timestamp 1698431365
transform 1 0 29680 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_260
timestamp 1698431365
transform 1 0 30464 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_268
timestamp 1698431365
transform 1 0 31360 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_272
timestamp 1698431365
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_274
timestamp 1698431365
transform 1 0 32032 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_277
timestamp 1698431365
transform 1 0 32368 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_312
timestamp 1698431365
transform 1 0 36288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_314
timestamp 1698431365
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_321
timestamp 1698431365
transform 1 0 37296 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_325
timestamp 1698431365
transform 1 0 37744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_329
timestamp 1698431365
transform 1 0 38192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_333
timestamp 1698431365
transform 1 0 38640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_337
timestamp 1698431365
transform 1 0 39088 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_393
timestamp 1698431365
transform 1 0 45360 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_6
timestamp 1698431365
transform 1 0 2016 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_33
timestamp 1698431365
transform 1 0 5040 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_41
timestamp 1698431365
transform 1 0 5936 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_43
timestamp 1698431365
transform 1 0 6160 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_76
timestamp 1698431365
transform 1 0 9856 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_89
timestamp 1698431365
transform 1 0 11312 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_119
timestamp 1698431365
transform 1 0 14672 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_123
timestamp 1698431365
transform 1 0 15120 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_132
timestamp 1698431365
transform 1 0 16128 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_156
timestamp 1698431365
transform 1 0 18816 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_160
timestamp 1698431365
transform 1 0 19264 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_164
timestamp 1698431365
transform 1 0 19712 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_171
timestamp 1698431365
transform 1 0 20496 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_187
timestamp 1698431365
transform 1 0 22288 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_195
timestamp 1698431365
transform 1 0 23184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_197
timestamp 1698431365
transform 1 0 23408 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_204
timestamp 1698431365
transform 1 0 24192 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_208
timestamp 1698431365
transform 1 0 24640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_244
timestamp 1698431365
transform 1 0 28672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_275
timestamp 1698431365
transform 1 0 32144 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_294
timestamp 1698431365
transform 1 0 34272 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_298
timestamp 1698431365
transform 1 0 34720 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_314
timestamp 1698431365
transform 1 0 36512 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_335
timestamp 1698431365
transform 1 0 38864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_337
timestamp 1698431365
transform 1 0 39088 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_360
timestamp 1698431365
transform 1 0 41664 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_14
timestamp 1698431365
transform 1 0 2912 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_31
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_53
timestamp 1698431365
transform 1 0 7280 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_62
timestamp 1698431365
transform 1 0 8288 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_72
timestamp 1698431365
transform 1 0 9408 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_84
timestamp 1698431365
transform 1 0 10752 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_94
timestamp 1698431365
transform 1 0 11872 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_96
timestamp 1698431365
transform 1 0 12096 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_115
timestamp 1698431365
transform 1 0 14224 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_117
timestamp 1698431365
transform 1 0 14448 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_161
timestamp 1698431365
transform 1 0 19376 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_170
timestamp 1698431365
transform 1 0 20384 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698431365
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_193
timestamp 1698431365
transform 1 0 22960 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_197
timestamp 1698431365
transform 1 0 23408 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_199
timestamp 1698431365
transform 1 0 23632 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_206
timestamp 1698431365
transform 1 0 24416 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_222
timestamp 1698431365
transform 1 0 26208 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_230
timestamp 1698431365
transform 1 0 27104 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_238
timestamp 1698431365
transform 1 0 28000 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_242
timestamp 1698431365
transform 1 0 28448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_255
timestamp 1698431365
transform 1 0 29904 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_259
timestamp 1698431365
transform 1 0 30352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_263
timestamp 1698431365
transform 1 0 30800 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_275
timestamp 1698431365
transform 1 0 32144 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_291
timestamp 1698431365
transform 1 0 33936 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_293
timestamp 1698431365
transform 1 0 34160 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_296
timestamp 1698431365
transform 1 0 34496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_298
timestamp 1698431365
transform 1 0 34720 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_301
timestamp 1698431365
transform 1 0 35056 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_305
timestamp 1698431365
transform 1 0 35504 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_323
timestamp 1698431365
transform 1 0 37520 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_356
timestamp 1698431365
transform 1 0 41216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_358
timestamp 1698431365
transform 1 0 41440 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_393
timestamp 1698431365
transform 1 0 45360 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_34
timestamp 1698431365
transform 1 0 5152 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_94
timestamp 1698431365
transform 1 0 11872 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_99
timestamp 1698431365
transform 1 0 12432 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_115
timestamp 1698431365
transform 1 0 14224 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_119
timestamp 1698431365
transform 1 0 14672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_121
timestamp 1698431365
transform 1 0 14896 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_126
timestamp 1698431365
transform 1 0 15456 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_134
timestamp 1698431365
transform 1 0 16352 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_138
timestamp 1698431365
transform 1 0 16800 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_148
timestamp 1698431365
transform 1 0 17920 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_152
timestamp 1698431365
transform 1 0 18368 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_195
timestamp 1698431365
transform 1 0 23184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_197
timestamp 1698431365
transform 1 0 23408 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_218
timestamp 1698431365
transform 1 0 25760 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_227
timestamp 1698431365
transform 1 0 26768 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_271
timestamp 1698431365
transform 1 0 31696 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_286
timestamp 1698431365
transform 1 0 33376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_288
timestamp 1698431365
transform 1 0 33600 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_307
timestamp 1698431365
transform 1 0 35728 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_309
timestamp 1698431365
transform 1 0 35952 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_316
timestamp 1698431365
transform 1 0 36736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_31
timestamp 1698431365
transform 1 0 4816 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_66
timestamp 1698431365
transform 1 0 8736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_70
timestamp 1698431365
transform 1 0 9184 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_102
timestamp 1698431365
transform 1 0 12768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_104
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_115
timestamp 1698431365
transform 1 0 14224 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_119
timestamp 1698431365
transform 1 0 14672 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_123
timestamp 1698431365
transform 1 0 15120 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_127
timestamp 1698431365
transform 1 0 15568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_129
timestamp 1698431365
transform 1 0 15792 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_159
timestamp 1698431365
transform 1 0 19152 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_189
timestamp 1698431365
transform 1 0 22512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_193
timestamp 1698431365
transform 1 0 22960 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_206
timestamp 1698431365
transform 1 0 24416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_216
timestamp 1698431365
transform 1 0 25536 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_265
timestamp 1698431365
transform 1 0 31024 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_269
timestamp 1698431365
transform 1 0 31472 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_299
timestamp 1698431365
transform 1 0 34832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_28
timestamp 1698431365
transform 1 0 4480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_30
timestamp 1698431365
transform 1 0 4704 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_37
timestamp 1698431365
transform 1 0 5488 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_41
timestamp 1698431365
transform 1 0 5936 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_57
timestamp 1698431365
transform 1 0 7728 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_65
timestamp 1698431365
transform 1 0 8624 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_69
timestamp 1698431365
transform 1 0 9072 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_80
timestamp 1698431365
transform 1 0 10304 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_131
timestamp 1698431365
transform 1 0 16016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_135
timestamp 1698431365
transform 1 0 16464 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_139
timestamp 1698431365
transform 1 0 16912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_150
timestamp 1698431365
transform 1 0 18144 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_158
timestamp 1698431365
transform 1 0 19040 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_162
timestamp 1698431365
transform 1 0 19488 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_164
timestamp 1698431365
transform 1 0 19712 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_181
timestamp 1698431365
transform 1 0 21616 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_189
timestamp 1698431365
transform 1 0 22512 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_193
timestamp 1698431365
transform 1 0 22960 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_200
timestamp 1698431365
transform 1 0 23744 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_208
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_244
timestamp 1698431365
transform 1 0 28672 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_260
timestamp 1698431365
transform 1 0 30464 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_268
timestamp 1698431365
transform 1 0 31360 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_272
timestamp 1698431365
transform 1 0 31808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_274
timestamp 1698431365
transform 1 0 32032 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_277
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_286
timestamp 1698431365
transform 1 0 33376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_343
timestamp 1698431365
transform 1 0 39760 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_28
timestamp 1698431365
transform 1 0 4480 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_32
timestamp 1698431365
transform 1 0 4928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_53
timestamp 1698431365
transform 1 0 7280 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_57
timestamp 1698431365
transform 1 0 7728 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_88
timestamp 1698431365
transform 1 0 11200 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_92
timestamp 1698431365
transform 1 0 11648 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_100
timestamp 1698431365
transform 1 0 12544 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698431365
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_119
timestamp 1698431365
transform 1 0 14672 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_151
timestamp 1698431365
transform 1 0 18256 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_159
timestamp 1698431365
transform 1 0 19152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_170
timestamp 1698431365
transform 1 0 20384 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_185
timestamp 1698431365
transform 1 0 22064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_193
timestamp 1698431365
transform 1 0 22960 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_200
timestamp 1698431365
transform 1 0 23744 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_220
timestamp 1698431365
transform 1 0 25984 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_224
timestamp 1698431365
transform 1 0 26432 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_236
timestamp 1698431365
transform 1 0 27776 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_276
timestamp 1698431365
transform 1 0 32256 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_380
timestamp 1698431365
transform 1 0 43904 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_384
timestamp 1698431365
transform 1 0 44352 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_393
timestamp 1698431365
transform 1 0 45360 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_28
timestamp 1698431365
transform 1 0 4480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_32
timestamp 1698431365
transform 1 0 4928 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_64
timestamp 1698431365
transform 1 0 8512 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_68
timestamp 1698431365
transform 1 0 8960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_76
timestamp 1698431365
transform 1 0 9856 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_86
timestamp 1698431365
transform 1 0 10976 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_118
timestamp 1698431365
transform 1 0 14560 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_156
timestamp 1698431365
transform 1 0 18816 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_160
timestamp 1698431365
transform 1 0 19264 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_162
timestamp 1698431365
transform 1 0 19488 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_167
timestamp 1698431365
transform 1 0 20048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_169
timestamp 1698431365
transform 1 0 20272 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_172
timestamp 1698431365
transform 1 0 20608 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_198
timestamp 1698431365
transform 1 0 23520 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_234
timestamp 1698431365
transform 1 0 27552 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_249
timestamp 1698431365
transform 1 0 29232 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_257
timestamp 1698431365
transform 1 0 30128 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_260
timestamp 1698431365
transform 1 0 30464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_264
timestamp 1698431365
transform 1 0 30912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698431365
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_111
timestamp 1698431365
transform 1 0 13776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_142
timestamp 1698431365
transform 1 0 17248 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_146
timestamp 1698431365
transform 1 0 17696 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_155
timestamp 1698431365
transform 1 0 18704 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_181
timestamp 1698431365
transform 1 0 21616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_185
timestamp 1698431365
transform 1 0 22064 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_193
timestamp 1698431365
transform 1 0 22960 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_199
timestamp 1698431365
transform 1 0 23632 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_207
timestamp 1698431365
transform 1 0 24528 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_209
timestamp 1698431365
transform 1 0 24752 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_212
timestamp 1698431365
transform 1 0 25088 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_228
timestamp 1698431365
transform 1 0 26880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_232
timestamp 1698431365
transform 1 0 27328 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_236
timestamp 1698431365
transform 1 0 27776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_238
timestamp 1698431365
transform 1 0 28000 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_253
timestamp 1698431365
transform 1 0 29680 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_257
timestamp 1698431365
transform 1 0 30128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_261
timestamp 1698431365
transform 1 0 30576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_419
timestamp 1698431365
transform 1 0 48272 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_76
timestamp 1698431365
transform 1 0 9856 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_79
timestamp 1698431365
transform 1 0 10192 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_95
timestamp 1698431365
transform 1 0 11984 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_98
timestamp 1698431365
transform 1 0 12320 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_104
timestamp 1698431365
transform 1 0 12992 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_122
timestamp 1698431365
transform 1 0 15008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_126
timestamp 1698431365
transform 1 0 15456 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_130
timestamp 1698431365
transform 1 0 15904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_171
timestamp 1698431365
transform 1 0 20496 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_173
timestamp 1698431365
transform 1 0 20720 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_203
timestamp 1698431365
transform 1 0 24080 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_247
timestamp 1698431365
transform 1 0 29008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_251
timestamp 1698431365
transform 1 0 29456 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_255
timestamp 1698431365
transform 1 0 29904 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_295
timestamp 1698431365
transform 1 0 34384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_297
timestamp 1698431365
transform 1 0 34608 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_354
timestamp 1698431365
transform 1 0 40992 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_419
timestamp 1698431365
transform 1 0 48272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_36
timestamp 1698431365
transform 1 0 5376 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_52
timestamp 1698431365
transform 1 0 7168 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_60
timestamp 1698431365
transform 1 0 8064 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_64
timestamp 1698431365
transform 1 0 8512 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_70
timestamp 1698431365
transform 1 0 9184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_72
timestamp 1698431365
transform 1 0 9408 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_85
timestamp 1698431365
transform 1 0 10864 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_89
timestamp 1698431365
transform 1 0 11312 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_106
timestamp 1698431365
transform 1 0 13216 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_115
timestamp 1698431365
transform 1 0 14224 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_117
timestamp 1698431365
transform 1 0 14448 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_184
timestamp 1698431365
transform 1 0 21952 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_188
timestamp 1698431365
transform 1 0 22400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_418
timestamp 1698431365
transform 1 0 48160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 28896 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 28336 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 23520 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 22848 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 21280 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 17024 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 15904 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 20384 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 33040 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 24864 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 12096 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 7616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 8288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 8288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 13664 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 18704 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 19712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 24192 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 13552 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 31808 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 32704 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 37744 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform -1 0 43232 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform -1 0 48384 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform -1 0 48384 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 48384 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 48384 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 47712 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 10864 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 48384 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform -1 0 48384 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 9520 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 11424 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform -1 0 15904 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 14560 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698431365
transform -1 0 21952 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform 1 0 9856 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698431365
transform -1 0 28784 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform 1 0 45360 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform 1 0 27328 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform -1 0 34384 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output49 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48384 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output50
timestamp 1698431365
transform 1 0 34720 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output51
timestamp 1698431365
transform 1 0 45472 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output52
timestamp 1698431365
transform 1 0 33712 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output53
timestamp 1698431365
transform 1 0 37632 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output54
timestamp 1698431365
transform 1 0 40320 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output55
timestamp 1698431365
transform 1 0 41552 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output56
timestamp 1698431365
transform 1 0 37632 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output57
timestamp 1698431365
transform 1 0 38640 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output58
timestamp 1698431365
transform 1 0 44016 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output59
timestamp 1698431365
transform 1 0 32704 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output60
timestamp 1698431365
transform 1 0 45472 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output61
timestamp 1698431365
transform 1 0 38640 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output62
timestamp 1698431365
transform 1 0 41552 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output63
timestamp 1698431365
transform 1 0 45472 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output64
timestamp 1698431365
transform 1 0 45472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output65
timestamp 1698431365
transform 1 0 37632 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output66
timestamp 1698431365
transform 1 0 41552 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output67
timestamp 1698431365
transform 1 0 41104 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output68
timestamp 1698431365
transform 1 0 43456 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output69
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output70
timestamp 1698431365
transform 1 0 33712 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output71
timestamp 1698431365
transform 1 0 45472 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output72
timestamp 1698431365
transform -1 0 37632 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output73
timestamp 1698431365
transform 1 0 45472 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output74
timestamp 1698431365
transform 1 0 42560 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output75
timestamp 1698431365
transform 1 0 45472 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output76
timestamp 1698431365
transform 1 0 42560 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output77
timestamp 1698431365
transform -1 0 48384 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output78
timestamp 1698431365
transform 1 0 35840 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output79
timestamp 1698431365
transform 1 0 41552 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output80
timestamp 1698431365
transform 1 0 42560 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output81
timestamp 1698431365
transform 1 0 24416 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output82
timestamp 1698431365
transform -1 0 4480 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output83
timestamp 1698431365
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output84
timestamp 1698431365
transform -1 0 4480 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output85
timestamp 1698431365
transform 1 0 10864 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output86
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output87
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output88
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output89
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output90
timestamp 1698431365
transform 1 0 24304 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output91
timestamp 1698431365
transform -1 0 28000 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output92
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output93
timestamp 1698431365
transform -1 0 4480 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output94
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output95
timestamp 1698431365
transform 1 0 33712 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output96
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output97
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output98
timestamp 1698431365
transform 1 0 45472 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output99
timestamp 1698431365
transform 1 0 45472 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output100
timestamp 1698431365
transform 1 0 45472 0 1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output101
timestamp 1698431365
transform 1 0 45472 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output102
timestamp 1698431365
transform 1 0 45472 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output103
timestamp 1698431365
transform 1 0 45472 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output104
timestamp 1698431365
transform -1 0 4480 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output105
timestamp 1698431365
transform 1 0 45472 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output106
timestamp 1698431365
transform 1 0 45472 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output107
timestamp 1698431365
transform -1 0 4480 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output108
timestamp 1698431365
transform -1 0 4480 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output109
timestamp 1698431365
transform 1 0 16800 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output110
timestamp 1698431365
transform -1 0 4480 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output111
timestamp 1698431365
transform -1 0 4480 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output112
timestamp 1698431365
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output113
timestamp 1698431365
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output114
timestamp 1698431365
transform 1 0 28896 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_55 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_106
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_107
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_108
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_109
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simpleuart_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41552 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simpleuart_143
timestamp 1698431365
transform 1 0 46928 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  simpleuart_144 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47936 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_118
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_119
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_120
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_121
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_122
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_123
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_124
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_125
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_126
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_128
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_129
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_130
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_131
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_132
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_133
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_134
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_135
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_136
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_137
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_138
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_139
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_140
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_141
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_142
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_143
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_144
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_145
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_146
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_147
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_148
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_149
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_150
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_151
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_152
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_153
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_154
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_155
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_156
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_157
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_158
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_159
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_160
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_161
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_162
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_163
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_164
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_165
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_166
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_167
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_168
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_169
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_170
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_171
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_172
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_173
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_174
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_175
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_176
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_177
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_178
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_179
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_180
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_181
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_183
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_184
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_185
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_186
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_187
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_188
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_189
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_190
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_191
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_192
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_193
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_194
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_195
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_196
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_197
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_198
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_199
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_200
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_201
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_202
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_203
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_204
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_205
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_206
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_207
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_208
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_209
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_210
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_211
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_212
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_213
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_214
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_215
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_216
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_217
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_218
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_219
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_220
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_221
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_222
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_223
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_224
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_225
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_226
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_227
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_228
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_229
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_230
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_231
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_232
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_233
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_234
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_235
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_236
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_237
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_238
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_239
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_240
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_241
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_242
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_243
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_244
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_245
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_246
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_247
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_248
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_249
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_250
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_251
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_252
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_253
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_254
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_255
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_256
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_257
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_258
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_259
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_260
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_261
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_262
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_263
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_264
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_265
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_266
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_267
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_268
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_269
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_270
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_271
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_272
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_273
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_274
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_275
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_276
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_277
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_278
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_279
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_280
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_281
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_282
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_283
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_284
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_285
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_286
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_287
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_288
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_289
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_290
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_291
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_292
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_293
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_294
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_295
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_296
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_297
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_298
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_299
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_300
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_301
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_302
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_303
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_304
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_305
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_306
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_307
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_308
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_309
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_310
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_311
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_312
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_313
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_314
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_315
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_316
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_317
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_318
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_319
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_320
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_321
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_322
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_323
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_324
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_325
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_326
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_327
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_328
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_329
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_330
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_331
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_332
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_333
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_334
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_335
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_336
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_337
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_338
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_339
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_340
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_341
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_342
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_343
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_344
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_345
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_346
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_347
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_348
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_349
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_350
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_351
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_352
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_353
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_354
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_355
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_356
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_357
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_358
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_359
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_360
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_361
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_362
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_363
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_364
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_365
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_366
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_367
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_368
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_369
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_370
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_371
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_372
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_373
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_374
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_375
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_376
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_377
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_378
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_379
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_380
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_381
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_382
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_383
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_384
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_385
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_386
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_387
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_388
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_389
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_390
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_391
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_392
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_393
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_394
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_395
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_396
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_397
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_398
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_399
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_400
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_401
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_402
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_403
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_404
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_405
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_406
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_407
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_408
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_409
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_410
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_411
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_412
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_413
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_414
timestamp 1698431365
transform 1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_415
timestamp 1698431365
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_416
timestamp 1698431365
transform 1 0 16576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_417
timestamp 1698431365
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_418
timestamp 1698431365
transform 1 0 24192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_419
timestamp 1698431365
transform 1 0 28000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_420
timestamp 1698431365
transform 1 0 31808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_421
timestamp 1698431365
transform 1 0 35616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_422
timestamp 1698431365
transform 1 0 39424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_423
timestamp 1698431365
transform 1 0 43232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_424
timestamp 1698431365
transform 1 0 47040 0 1 45472
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 45024 800 45136 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 27552 49200 27664 50000 0 FreeSans 448 90 0 0 reg_dat_di[0]
port 1 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 reg_dat_di[10]
port 2 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 reg_dat_di[11]
port 3 nsew signal input
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 reg_dat_di[12]
port 4 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 reg_dat_di[13]
port 5 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 reg_dat_di[14]
port 6 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 reg_dat_di[15]
port 7 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 reg_dat_di[16]
port 8 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 reg_dat_di[17]
port 9 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 reg_dat_di[18]
port 10 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 reg_dat_di[19]
port 11 nsew signal input
flabel metal2 s 28224 49200 28336 50000 0 FreeSans 448 90 0 0 reg_dat_di[1]
port 12 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 reg_dat_di[20]
port 13 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 reg_dat_di[21]
port 14 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 reg_dat_di[22]
port 15 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 reg_dat_di[23]
port 16 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 reg_dat_di[24]
port 17 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 reg_dat_di[25]
port 18 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 reg_dat_di[26]
port 19 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 reg_dat_di[27]
port 20 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 reg_dat_di[28]
port 21 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 reg_dat_di[29]
port 22 nsew signal input
flabel metal2 s 24864 49200 24976 50000 0 FreeSans 448 90 0 0 reg_dat_di[2]
port 23 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 reg_dat_di[30]
port 24 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 reg_dat_di[31]
port 25 nsew signal input
flabel metal2 s 22848 49200 22960 50000 0 FreeSans 448 90 0 0 reg_dat_di[3]
port 26 nsew signal input
flabel metal2 s 18816 49200 18928 50000 0 FreeSans 448 90 0 0 reg_dat_di[4]
port 27 nsew signal input
flabel metal2 s 16800 49200 16912 50000 0 FreeSans 448 90 0 0 reg_dat_di[5]
port 28 nsew signal input
flabel metal2 s 17472 49200 17584 50000 0 FreeSans 448 90 0 0 reg_dat_di[6]
port 29 nsew signal input
flabel metal2 s 19488 49200 19600 50000 0 FreeSans 448 90 0 0 reg_dat_di[7]
port 30 nsew signal input
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 reg_dat_di[8]
port 31 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 reg_dat_di[9]
port 32 nsew signal input
flabel metal3 s 49200 34272 50000 34384 0 FreeSans 448 0 0 0 reg_dat_do[0]
port 33 nsew signal tristate
flabel metal3 s 49200 49728 50000 49840 0 FreeSans 448 0 0 0 reg_dat_do[10]
port 34 nsew signal tristate
flabel metal3 s 49200 35616 50000 35728 0 FreeSans 448 0 0 0 reg_dat_do[11]
port 35 nsew signal tristate
flabel metal3 s 49200 49056 50000 49168 0 FreeSans 448 0 0 0 reg_dat_do[12]
port 36 nsew signal tristate
flabel metal2 s 45024 49200 45136 50000 0 FreeSans 448 90 0 0 reg_dat_do[13]
port 37 nsew signal tristate
flabel metal2 s 40320 49200 40432 50000 0 FreeSans 448 90 0 0 reg_dat_do[14]
port 38 nsew signal tristate
flabel metal3 s 49200 48384 50000 48496 0 FreeSans 448 0 0 0 reg_dat_do[15]
port 39 nsew signal tristate
flabel metal3 s 49200 43008 50000 43120 0 FreeSans 448 0 0 0 reg_dat_do[16]
port 40 nsew signal tristate
flabel metal3 s 49200 44352 50000 44464 0 FreeSans 448 0 0 0 reg_dat_do[17]
port 41 nsew signal tristate
flabel metal2 s 42336 49200 42448 50000 0 FreeSans 448 90 0 0 reg_dat_do[18]
port 42 nsew signal tristate
flabel metal3 s 49200 45024 50000 45136 0 FreeSans 448 0 0 0 reg_dat_do[19]
port 43 nsew signal tristate
flabel metal3 s 49200 38304 50000 38416 0 FreeSans 448 0 0 0 reg_dat_do[1]
port 44 nsew signal tristate
flabel metal2 s 44352 49200 44464 50000 0 FreeSans 448 90 0 0 reg_dat_do[20]
port 45 nsew signal tristate
flabel metal3 s 49200 42336 50000 42448 0 FreeSans 448 0 0 0 reg_dat_do[21]
port 46 nsew signal tristate
flabel metal3 s 49200 34944 50000 35056 0 FreeSans 448 0 0 0 reg_dat_do[22]
port 47 nsew signal tristate
flabel metal3 s 49200 36288 50000 36400 0 FreeSans 448 0 0 0 reg_dat_do[23]
port 48 nsew signal tristate
flabel metal3 s 49200 45696 50000 45808 0 FreeSans 448 0 0 0 reg_dat_do[24]
port 49 nsew signal tristate
flabel metal3 s 49200 43680 50000 43792 0 FreeSans 448 0 0 0 reg_dat_do[25]
port 50 nsew signal tristate
flabel metal2 s 40992 49200 41104 50000 0 FreeSans 448 90 0 0 reg_dat_do[26]
port 51 nsew signal tristate
flabel metal2 s 41664 49200 41776 50000 0 FreeSans 448 90 0 0 reg_dat_do[27]
port 52 nsew signal tristate
flabel metal2 s 43008 49200 43120 50000 0 FreeSans 448 90 0 0 reg_dat_do[28]
port 53 nsew signal tristate
flabel metal3 s 49200 47712 50000 47824 0 FreeSans 448 0 0 0 reg_dat_do[29]
port 54 nsew signal tristate
flabel metal3 s 49200 40320 50000 40432 0 FreeSans 448 0 0 0 reg_dat_do[2]
port 55 nsew signal tristate
flabel metal2 s 45696 49200 45808 50000 0 FreeSans 448 90 0 0 reg_dat_do[30]
port 56 nsew signal tristate
flabel metal3 s 49200 37632 50000 37744 0 FreeSans 448 0 0 0 reg_dat_do[31]
port 57 nsew signal tristate
flabel metal3 s 49200 38976 50000 39088 0 FreeSans 448 0 0 0 reg_dat_do[3]
port 58 nsew signal tristate
flabel metal3 s 49200 39648 50000 39760 0 FreeSans 448 0 0 0 reg_dat_do[4]
port 59 nsew signal tristate
flabel metal3 s 49200 41664 50000 41776 0 FreeSans 448 0 0 0 reg_dat_do[5]
port 60 nsew signal tristate
flabel metal3 s 49200 36960 50000 37072 0 FreeSans 448 0 0 0 reg_dat_do[6]
port 61 nsew signal tristate
flabel metal2 s 34944 49200 35056 50000 0 FreeSans 448 90 0 0 reg_dat_do[7]
port 62 nsew signal tristate
flabel metal2 s 43680 49200 43792 50000 0 FreeSans 448 90 0 0 reg_dat_do[8]
port 63 nsew signal tristate
flabel metal3 s 49200 40992 50000 41104 0 FreeSans 448 0 0 0 reg_dat_do[9]
port 64 nsew signal tristate
flabel metal2 s 32928 49200 33040 50000 0 FreeSans 448 90 0 0 reg_dat_re
port 65 nsew signal input
flabel metal2 s 23520 49200 23632 50000 0 FreeSans 448 90 0 0 reg_dat_wait
port 66 nsew signal tristate
flabel metal2 s 24192 49200 24304 50000 0 FreeSans 448 90 0 0 reg_dat_we
port 67 nsew signal input
flabel metal2 s 12768 49200 12880 50000 0 FreeSans 448 90 0 0 reg_div_di[0]
port 68 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 reg_div_di[10]
port 69 nsew signal input
flabel metal3 s 0 8064 800 8176 0 FreeSans 448 0 0 0 reg_div_di[11]
port 70 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 reg_div_di[12]
port 71 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 reg_div_di[13]
port 72 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 reg_div_di[14]
port 73 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 reg_div_di[15]
port 74 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 reg_div_di[16]
port 75 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 reg_div_di[17]
port 76 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 reg_div_di[18]
port 77 nsew signal input
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 reg_div_di[19]
port 78 nsew signal input
flabel metal2 s 13440 49200 13552 50000 0 FreeSans 448 90 0 0 reg_div_di[1]
port 79 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 reg_div_di[20]
port 80 nsew signal input
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 reg_div_di[21]
port 81 nsew signal input
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 reg_div_di[22]
port 82 nsew signal input
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 reg_div_di[23]
port 83 nsew signal input
flabel metal2 s 41664 0 41776 800 0 FreeSans 448 90 0 0 reg_div_di[24]
port 84 nsew signal input
flabel metal3 s 49200 8736 50000 8848 0 FreeSans 448 0 0 0 reg_div_di[25]
port 85 nsew signal input
flabel metal3 s 49200 10752 50000 10864 0 FreeSans 448 0 0 0 reg_div_di[26]
port 86 nsew signal input
flabel metal3 s 49200 17472 50000 17584 0 FreeSans 448 0 0 0 reg_div_di[27]
port 87 nsew signal input
flabel metal3 s 49200 20832 50000 20944 0 FreeSans 448 0 0 0 reg_div_di[28]
port 88 nsew signal input
flabel metal3 s 49200 23520 50000 23632 0 FreeSans 448 0 0 0 reg_div_di[29]
port 89 nsew signal input
flabel metal2 s 10080 49200 10192 50000 0 FreeSans 448 90 0 0 reg_div_di[2]
port 90 nsew signal input
flabel metal3 s 49200 24864 50000 24976 0 FreeSans 448 0 0 0 reg_div_di[30]
port 91 nsew signal input
flabel metal3 s 49200 12096 50000 12208 0 FreeSans 448 0 0 0 reg_div_di[31]
port 92 nsew signal input
flabel metal2 s 9408 49200 9520 50000 0 FreeSans 448 90 0 0 reg_div_di[3]
port 93 nsew signal input
flabel metal2 s 12096 49200 12208 50000 0 FreeSans 448 90 0 0 reg_div_di[4]
port 94 nsew signal input
flabel metal2 s 15456 49200 15568 50000 0 FreeSans 448 90 0 0 reg_div_di[5]
port 95 nsew signal input
flabel metal2 s 14784 49200 14896 50000 0 FreeSans 448 90 0 0 reg_div_di[6]
port 96 nsew signal input
flabel metal3 s 0 34272 800 34384 0 FreeSans 448 0 0 0 reg_div_di[7]
port 97 nsew signal input
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 reg_div_di[8]
port 98 nsew signal input
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 reg_div_di[9]
port 99 nsew signal input
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 reg_div_do[0]
port 100 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 reg_div_do[10]
port 101 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 reg_div_do[11]
port 102 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 reg_div_do[12]
port 103 nsew signal tristate
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 reg_div_do[13]
port 104 nsew signal tristate
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 reg_div_do[14]
port 105 nsew signal tristate
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 reg_div_do[15]
port 106 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 reg_div_do[16]
port 107 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 reg_div_do[17]
port 108 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 reg_div_do[18]
port 109 nsew signal tristate
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 reg_div_do[19]
port 110 nsew signal tristate
flabel metal3 s 0 42336 800 42448 0 FreeSans 448 0 0 0 reg_div_do[1]
port 111 nsew signal tristate
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 reg_div_do[20]
port 112 nsew signal tristate
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 reg_div_do[21]
port 113 nsew signal tristate
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 reg_div_do[22]
port 114 nsew signal tristate
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 reg_div_do[23]
port 115 nsew signal tristate
flabel metal3 s 49200 6048 50000 6160 0 FreeSans 448 0 0 0 reg_div_do[24]
port 116 nsew signal tristate
flabel metal3 s 49200 9408 50000 9520 0 FreeSans 448 0 0 0 reg_div_do[25]
port 117 nsew signal tristate
flabel metal3 s 49200 11424 50000 11536 0 FreeSans 448 0 0 0 reg_div_do[26]
port 118 nsew signal tristate
flabel metal3 s 49200 16128 50000 16240 0 FreeSans 448 0 0 0 reg_div_do[27]
port 119 nsew signal tristate
flabel metal3 s 49200 20160 50000 20272 0 FreeSans 448 0 0 0 reg_div_do[28]
port 120 nsew signal tristate
flabel metal3 s 49200 22848 50000 22960 0 FreeSans 448 0 0 0 reg_div_do[29]
port 121 nsew signal tristate
flabel metal3 s 0 41664 800 41776 0 FreeSans 448 0 0 0 reg_div_do[2]
port 122 nsew signal tristate
flabel metal3 s 49200 26208 50000 26320 0 FreeSans 448 0 0 0 reg_div_do[30]
port 123 nsew signal tristate
flabel metal3 s 49200 12768 50000 12880 0 FreeSans 448 0 0 0 reg_div_do[31]
port 124 nsew signal tristate
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 reg_div_do[3]
port 125 nsew signal tristate
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 reg_div_do[4]
port 126 nsew signal tristate
flabel metal2 s 16128 49200 16240 50000 0 FreeSans 448 90 0 0 reg_div_do[5]
port 127 nsew signal tristate
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 reg_div_do[6]
port 128 nsew signal tristate
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 reg_div_do[7]
port 129 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 reg_div_do[8]
port 130 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 reg_div_do[9]
port 131 nsew signal tristate
flabel metal2 s 18144 49200 18256 50000 0 FreeSans 448 90 0 0 reg_div_we[0]
port 132 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 reg_div_we[1]
port 133 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 reg_div_we[2]
port 134 nsew signal input
flabel metal3 s 49200 18144 50000 18256 0 FreeSans 448 0 0 0 reg_div_we[3]
port 135 nsew signal input
flabel metal2 s 26880 49200 26992 50000 0 FreeSans 448 90 0 0 resetn
port 136 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 uart_in[0]
port 137 nsew signal input
flabel metal2 s 33600 49200 33712 50000 0 FreeSans 448 90 0 0 uart_in[1]
port 138 nsew signal input
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 uart_oeb[0]
port 139 nsew signal tristate
flabel metal3 s 49200 47040 50000 47152 0 FreeSans 448 0 0 0 uart_oeb[1]
port 140 nsew signal tristate
flabel metal2 s 28896 49200 29008 50000 0 FreeSans 448 90 0 0 uart_out[0]
port 141 nsew signal tristate
flabel metal3 s 49200 46368 50000 46480 0 FreeSans 448 0 0 0 uart_out[1]
port 142 nsew signal tristate
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vdd
port 143 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vdd
port 143 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vss
port 144 nsew ground bidirectional
rlabel metal1 24976 46256 24976 46256 0 vdd
rlabel metal1 24976 45472 24976 45472 0 vss
rlabel metal2 29848 38668 29848 38668 0 _0000_
rlabel metal2 12488 23520 12488 23520 0 _0001_
rlabel metal2 11872 21560 11872 21560 0 _0002_
rlabel metal2 6552 6216 6552 6216 0 _0003_
rlabel metal2 6216 7784 6216 7784 0 _0004_
rlabel metal2 8120 4760 8120 4760 0 _0005_
rlabel metal2 10024 8624 10024 8624 0 _0006_
rlabel metal3 11592 4200 11592 4200 0 _0007_
rlabel metal3 13552 6552 13552 6552 0 _0008_
rlabel metal3 19040 4536 19040 4536 0 _0009_
rlabel metal3 21504 4200 21504 4200 0 _0010_
rlabel metal2 23912 6328 23912 6328 0 _0011_
rlabel metal2 27608 4648 27608 4648 0 _0012_
rlabel metal2 29456 4424 29456 4424 0 _0013_
rlabel metal2 31304 5208 31304 5208 0 _0014_
rlabel metal2 34552 5096 34552 5096 0 _0015_
rlabel metal3 35560 5768 35560 5768 0 _0016_
rlabel metal2 41720 6216 41720 6216 0 _0017_
rlabel metal2 42560 8344 42560 8344 0 _0018_
rlabel metal2 45304 10528 45304 10528 0 _0019_
rlabel metal2 45864 16632 45864 16632 0 _0020_
rlabel metal2 46872 20440 46872 20440 0 _0021_
rlabel metal2 46088 23296 46088 23296 0 _0022_
rlabel metal2 46424 25536 46424 25536 0 _0023_
rlabel metal3 45416 12376 45416 12376 0 _0024_
rlabel metal2 26096 37128 26096 37128 0 _0025_
rlabel metal2 29848 40712 29848 40712 0 _0026_
rlabel metal3 29624 42840 29624 42840 0 _0027_
rlabel metal2 25424 43736 25424 43736 0 _0028_
rlabel metal2 22904 43344 22904 43344 0 _0029_
rlabel metal2 18424 44688 18424 44688 0 _0030_
rlabel metal2 14952 43904 14952 43904 0 _0031_
rlabel metal2 16856 41384 16856 41384 0 _0032_
rlabel metal2 20104 40040 20104 40040 0 _0033_
rlabel metal2 20496 37352 20496 37352 0 _0034_
rlabel metal2 27160 35952 27160 35952 0 _0035_
rlabel metal2 19096 36008 19096 36008 0 _0036_
rlabel metal2 22344 30352 22344 30352 0 _0037_
rlabel metal2 19320 32984 19320 32984 0 _0038_
rlabel metal2 27496 30296 27496 30296 0 _0039_
rlabel metal2 29624 34104 29624 34104 0 _0040_
rlabel metal2 30632 36120 30632 36120 0 _0041_
rlabel metal2 37016 32872 37016 32872 0 _0042_
rlabel metal2 2520 40376 2520 40376 0 _0043_
rlabel metal2 6440 41496 6440 41496 0 _0044_
rlabel metal2 2520 38192 2520 38192 0 _0045_
rlabel metal3 4032 35672 4032 35672 0 _0046_
rlabel metal2 2520 30632 2520 30632 0 _0047_
rlabel metal2 2576 27944 2576 27944 0 _0048_
rlabel metal2 6608 27944 6608 27944 0 _0049_
rlabel metal2 2520 25816 2520 25816 0 _0050_
rlabel metal2 8456 25816 8456 25816 0 _0051_
rlabel metal2 2856 23408 2856 23408 0 _0052_
rlabel metal2 3528 18592 3528 18592 0 _0053_
rlabel metal2 2744 19656 2744 19656 0 _0054_
rlabel metal2 2520 22064 2520 22064 0 _0055_
rlabel metal2 12936 20384 12936 20384 0 _0056_
rlabel metal2 18312 22680 18312 22680 0 _0057_
rlabel metal2 18816 20104 18816 20104 0 _0058_
rlabel metal2 22960 24024 22960 24024 0 _0059_
rlabel metal2 21224 22736 21224 22736 0 _0060_
rlabel metal2 20104 18592 20104 18592 0 _0061_
rlabel metal2 25928 18984 25928 18984 0 _0062_
rlabel metal2 25704 22736 25704 22736 0 _0063_
rlabel metal2 31080 16352 31080 16352 0 _0064_
rlabel metal2 31976 19544 31976 19544 0 _0065_
rlabel metal2 30744 21336 30744 21336 0 _0066_
rlabel metal2 26488 25984 26488 25984 0 _0067_
rlabel metal3 35224 22344 35224 22344 0 _0068_
rlabel metal2 34552 20748 34552 20748 0 _0069_
rlabel metal2 30968 24864 30968 24864 0 _0070_
rlabel metal2 33880 25088 33880 25088 0 _0071_
rlabel metal2 32424 28000 32424 28000 0 _0072_
rlabel metal2 29960 28224 29960 28224 0 _0073_
rlabel metal2 25928 27440 25928 27440 0 _0074_
rlabel metal2 45752 31416 45752 31416 0 _0075_
rlabel metal2 46088 33488 46088 33488 0 _0076_
rlabel metal2 42280 33712 42280 33712 0 _0077_
rlabel metal2 39928 31920 39928 31920 0 _0078_
rlabel metal2 38472 34104 38472 34104 0 _0079_
rlabel metal2 38024 36680 38024 36680 0 _0080_
rlabel metal2 35000 37688 35000 37688 0 _0081_
rlabel metal2 34552 35280 34552 35280 0 _0082_
rlabel metal3 45640 35784 45640 35784 0 _0083_
rlabel metal3 46480 38808 46480 38808 0 _0084_
rlabel metal2 41160 40824 41160 40824 0 _0085_
rlabel metal2 41776 36568 41776 36568 0 _0086_
rlabel metal2 39480 39256 39480 39256 0 _0087_
rlabel metal3 40432 41944 40432 41944 0 _0088_
rlabel metal2 37128 41552 37128 41552 0 _0089_
rlabel metal3 33992 40376 33992 40376 0 _0090_
rlabel metal2 2856 32816 2856 32816 0 _0091_
rlabel metal3 5376 32648 5376 32648 0 _0092_
rlabel metal2 6440 31584 6440 31584 0 _0093_
rlabel metal2 10360 29848 10360 29848 0 _0094_
rlabel metal2 10808 27384 10808 27384 0 _0095_
rlabel metal3 21560 27944 21560 27944 0 _0096_
rlabel metal3 20552 24808 20552 24808 0 _0097_
rlabel metal2 14448 16968 14448 16968 0 _0098_
rlabel metal3 3808 16744 3808 16744 0 _0099_
rlabel metal2 2520 14112 2520 14112 0 _0100_
rlabel metal2 2520 11760 2520 11760 0 _0101_
rlabel metal2 4928 10696 4928 10696 0 _0102_
rlabel metal2 8008 10640 8008 10640 0 _0103_
rlabel metal2 18536 14896 18536 14896 0 _0104_
rlabel metal2 19544 7784 19544 7784 0 _0105_
rlabel metal2 19992 9632 19992 9632 0 _0106_
rlabel metal2 21784 15792 21784 15792 0 _0107_
rlabel metal2 20888 12600 20888 12600 0 _0108_
rlabel metal2 21448 7952 21448 7952 0 _0109_
rlabel metal2 24920 8792 24920 8792 0 _0110_
rlabel metal2 29960 8624 29960 8624 0 _0111_
rlabel metal2 35000 8960 35000 8960 0 _0112_
rlabel metal2 39032 7728 39032 7728 0 _0113_
rlabel metal3 40488 9912 40488 9912 0 _0114_
rlabel metal2 35448 17360 35448 17360 0 _0115_
rlabel metal2 37520 18312 37520 18312 0 _0116_
rlabel metal2 42000 11480 42000 11480 0 _0117_
rlabel metal2 42168 13272 42168 13272 0 _0118_
rlabel metal3 45248 27720 45248 27720 0 _0119_
rlabel metal3 45528 29288 45528 29288 0 _0120_
rlabel metal2 41160 29792 41160 29792 0 _0121_
rlabel metal2 40936 21840 40936 21840 0 _0122_
rlabel metal3 12432 37352 12432 37352 0 _0123_
rlabel metal2 14168 42280 14168 42280 0 _0124_
rlabel metal2 8904 43120 8904 43120 0 _0125_
rlabel metal3 9072 40488 9072 40488 0 _0126_
rlabel metal2 12432 38920 12432 38920 0 _0127_
rlabel metal2 15512 39256 15512 39256 0 _0128_
rlabel metal2 15624 37016 15624 37016 0 _0129_
rlabel metal2 14728 34048 14728 34048 0 _0130_
rlabel metal2 26208 22232 26208 22232 0 _0131_
rlabel metal2 30464 20216 30464 20216 0 _0132_
rlabel metal3 30800 20776 30800 20776 0 _0133_
rlabel metal2 31360 19992 31360 19992 0 _0134_
rlabel metal3 30856 23128 30856 23128 0 _0135_
rlabel metal3 31528 21448 31528 21448 0 _0136_
rlabel metal2 29960 23688 29960 23688 0 _0137_
rlabel metal2 31416 22008 31416 22008 0 _0138_
rlabel metal2 28616 23856 28616 23856 0 _0139_
rlabel metal3 27496 23800 27496 23800 0 _0140_
rlabel metal2 26264 25200 26264 25200 0 _0141_
rlabel metal2 31080 24752 31080 24752 0 _0142_
rlabel metal3 34776 22456 34776 22456 0 _0143_
rlabel metal2 34328 23016 34328 23016 0 _0144_
rlabel metal2 34216 21840 34216 21840 0 _0145_
rlabel metal2 31640 22680 31640 22680 0 _0146_
rlabel metal2 31976 23520 31976 23520 0 _0147_
rlabel metal3 31584 24472 31584 24472 0 _0148_
rlabel metal2 31472 24696 31472 24696 0 _0149_
rlabel metal2 33376 24472 33376 24472 0 _0150_
rlabel metal2 33320 25200 33320 25200 0 _0151_
rlabel metal2 32760 27328 32760 27328 0 _0152_
rlabel metal2 33152 26488 33152 26488 0 _0153_
rlabel metal2 30296 27384 30296 27384 0 _0154_
rlabel metal3 29792 27720 29792 27720 0 _0155_
rlabel metal2 28616 27440 28616 27440 0 _0156_
rlabel metal2 45640 33656 45640 33656 0 _0157_
rlabel metal2 37240 34496 37240 34496 0 _0158_
rlabel metal2 45528 31752 45528 31752 0 _0159_
rlabel metal3 40544 32760 40544 32760 0 _0160_
rlabel metal2 46144 31080 46144 31080 0 _0161_
rlabel metal2 44912 33544 44912 33544 0 _0162_
rlabel metal2 43960 33432 43960 33432 0 _0163_
rlabel metal2 46760 34216 46760 34216 0 _0164_
rlabel metal2 42392 33768 42392 33768 0 _0165_
rlabel metal2 43064 33320 43064 33320 0 _0166_
rlabel metal2 40992 35112 40992 35112 0 _0167_
rlabel metal3 41664 32536 41664 32536 0 _0168_
rlabel metal2 40600 40600 40600 40600 0 _0169_
rlabel metal3 37632 34664 37632 34664 0 _0170_
rlabel metal2 39816 33488 39816 33488 0 _0171_
rlabel metal2 39928 32872 39928 32872 0 _0172_
rlabel metal2 37240 39928 37240 39928 0 _0173_
rlabel metal2 43624 36400 43624 36400 0 _0174_
rlabel metal3 38808 36344 38808 36344 0 _0175_
rlabel metal2 35224 40152 35224 40152 0 _0176_
rlabel metal3 35448 37408 35448 37408 0 _0177_
rlabel metal2 35000 35224 35000 35224 0 _0178_
rlabel metal2 43624 35392 43624 35392 0 _0179_
rlabel metal2 40936 40264 40936 40264 0 _0180_
rlabel metal2 44184 36624 44184 36624 0 _0181_
rlabel metal2 47208 41384 47208 41384 0 _0182_
rlabel metal3 46088 38920 46088 38920 0 _0183_
rlabel metal2 47488 45192 47488 45192 0 _0184_
rlabel metal3 40432 42056 40432 42056 0 _0185_
rlabel metal2 42168 36960 42168 36960 0 _0186_
rlabel metal2 39368 39088 39368 39088 0 _0187_
rlabel metal3 40488 38808 40488 38808 0 _0188_
rlabel metal2 39704 41832 39704 41832 0 _0189_
rlabel metal3 41664 41944 41664 41944 0 _0190_
rlabel metal2 37576 41496 37576 41496 0 _0191_
rlabel metal2 35112 40488 35112 40488 0 _0192_
rlabel metal2 21448 28840 21448 28840 0 _0193_
rlabel metal3 19936 16744 19936 16744 0 _0194_
rlabel metal2 22120 16128 22120 16128 0 _0195_
rlabel metal2 19096 16968 19096 16968 0 _0196_
rlabel metal2 5992 32760 5992 32760 0 _0197_
rlabel metal3 27272 16240 27272 16240 0 _0198_
rlabel metal2 9240 32592 9240 32592 0 _0199_
rlabel metal2 9016 32256 9016 32256 0 _0200_
rlabel metal2 11256 28616 11256 28616 0 _0201_
rlabel metal2 18368 30072 18368 30072 0 _0202_
rlabel metal3 9576 29400 9576 29400 0 _0203_
rlabel metal2 12040 28168 12040 28168 0 _0204_
rlabel metal2 19656 29232 19656 29232 0 _0205_
rlabel metal2 18928 30072 18928 30072 0 _0206_
rlabel metal2 19880 29512 19880 29512 0 _0207_
rlabel metal2 20440 29400 20440 29400 0 _0208_
rlabel metal2 19208 25816 19208 25816 0 _0209_
rlabel metal2 19376 26264 19376 26264 0 _0210_
rlabel metal2 17696 15960 17696 15960 0 _0211_
rlabel metal2 15176 15680 15176 15680 0 _0212_
rlabel metal2 3304 15344 3304 15344 0 _0213_
rlabel metal2 14952 17304 14952 17304 0 _0214_
rlabel metal2 3416 16016 3416 16016 0 _0215_
rlabel metal2 3976 13272 3976 13272 0 _0216_
rlabel metal2 3976 15148 3976 15148 0 _0217_
rlabel metal2 22736 26488 22736 26488 0 _0218_
rlabel metal2 21672 16016 21672 16016 0 _0219_
rlabel metal2 4480 12040 4480 12040 0 _0220_
rlabel metal2 15512 14336 15512 14336 0 _0221_
rlabel metal2 15960 13608 15960 13608 0 _0222_
rlabel metal2 6216 12432 6216 12432 0 _0223_
rlabel metal3 17976 14392 17976 14392 0 _0224_
rlabel metal2 9576 12096 9576 12096 0 _0225_
rlabel metal2 21448 12040 21448 12040 0 _0226_
rlabel metal2 17920 14728 17920 14728 0 _0227_
rlabel metal2 17864 12824 17864 12824 0 _0228_
rlabel metal2 19208 10612 19208 10612 0 _0229_
rlabel metal2 17752 8680 17752 8680 0 _0230_
rlabel metal2 18872 12488 18872 12488 0 _0231_
rlabel metal2 18984 9744 18984 9744 0 _0232_
rlabel metal2 19432 10864 19432 10864 0 _0233_
rlabel metal2 22456 15484 22456 15484 0 _0234_
rlabel metal3 22232 12040 22232 12040 0 _0235_
rlabel metal2 21448 15540 21448 15540 0 _0236_
rlabel metal2 21728 11592 21728 11592 0 _0237_
rlabel metal2 22680 10864 22680 10864 0 _0238_
rlabel metal2 24360 10472 24360 10472 0 _0239_
rlabel metal2 21728 11368 21728 11368 0 _0240_
rlabel metal2 21896 8680 21896 8680 0 _0241_
rlabel metal2 23912 9856 23912 9856 0 _0242_
rlabel metal2 24360 9184 24360 9184 0 _0243_
rlabel metal2 36232 17640 36232 17640 0 _0244_
rlabel metal2 26824 10976 26824 10976 0 _0245_
rlabel metal2 30184 9408 30184 9408 0 _0246_
rlabel metal3 33320 9688 33320 9688 0 _0247_
rlabel metal3 34048 9912 34048 9912 0 _0248_
rlabel metal2 38472 8232 38472 8232 0 _0249_
rlabel metal2 38808 10360 38808 10360 0 _0250_
rlabel metal2 38920 12320 38920 12320 0 _0251_
rlabel metal2 35672 10864 35672 10864 0 _0252_
rlabel metal3 37464 15400 37464 15400 0 _0253_
rlabel metal2 36456 16856 36456 16856 0 _0254_
rlabel metal2 38472 15232 38472 15232 0 _0255_
rlabel metal2 38248 15792 38248 15792 0 _0256_
rlabel metal3 38248 15176 38248 15176 0 _0257_
rlabel metal2 41160 12264 41160 12264 0 _0258_
rlabel metal2 40376 14168 40376 14168 0 _0259_
rlabel metal2 42504 14000 42504 14000 0 _0260_
rlabel metal2 43344 24920 43344 24920 0 _0261_
rlabel metal2 44072 27384 44072 27384 0 _0262_
rlabel metal2 43736 29512 43736 29512 0 _0263_
rlabel metal2 44072 29848 44072 29848 0 _0264_
rlabel metal2 44184 29120 44184 29120 0 _0265_
rlabel metal2 41496 29848 41496 29848 0 _0266_
rlabel metal2 42112 25144 42112 25144 0 _0267_
rlabel metal2 41272 22344 41272 22344 0 _0268_
rlabel metal2 15736 38080 15736 38080 0 _0269_
rlabel metal2 15512 41496 15512 41496 0 _0270_
rlabel metal2 13608 36960 13608 36960 0 _0271_
rlabel metal2 11480 41328 11480 41328 0 _0272_
rlabel metal2 14280 42728 14280 42728 0 _0273_
rlabel metal2 13608 42336 13608 42336 0 _0274_
rlabel metal2 10136 42840 10136 42840 0 _0275_
rlabel metal2 18424 39592 18424 39592 0 _0276_
rlabel metal2 11032 42392 11032 42392 0 _0277_
rlabel metal3 10472 40376 10472 40376 0 _0278_
rlabel metal2 18200 39060 18200 39060 0 _0279_
rlabel metal2 11592 40040 11592 40040 0 _0280_
rlabel metal2 12264 39872 12264 39872 0 _0281_
rlabel metal3 13440 39480 13440 39480 0 _0282_
rlabel metal2 15288 39480 15288 39480 0 _0283_
rlabel metal2 15960 39144 15960 39144 0 _0284_
rlabel metal2 15064 37184 15064 37184 0 _0285_
rlabel metal3 17080 36568 17080 36568 0 _0286_
rlabel metal2 14840 35168 14840 35168 0 _0287_
rlabel metal2 15512 35112 15512 35112 0 _0288_
rlabel metal2 23352 31136 23352 31136 0 _0289_
rlabel metal2 23408 35112 23408 35112 0 _0290_
rlabel metal2 23240 32032 23240 32032 0 _0291_
rlabel metal2 23688 30576 23688 30576 0 _0292_
rlabel metal2 23688 32872 23688 32872 0 _0293_
rlabel metal2 45192 41104 45192 41104 0 _0294_
rlabel metal2 47880 36568 47880 36568 0 _0295_
rlabel metal3 44184 36232 44184 36232 0 _0296_
rlabel metal2 41776 43288 41776 43288 0 _0297_
rlabel metal2 44856 42672 44856 42672 0 _0298_
rlabel metal3 41272 40040 41272 40040 0 _0299_
rlabel metal2 43400 38304 43400 38304 0 _0300_
rlabel metal2 40152 42224 40152 42224 0 _0301_
rlabel metal3 45304 44184 45304 44184 0 _0302_
rlabel metal2 34160 40600 34160 40600 0 _0303_
rlabel metal2 26600 33096 26600 33096 0 _0304_
rlabel metal2 30408 35840 30408 35840 0 _0305_
rlabel metal3 33544 38920 33544 38920 0 _0306_
rlabel metal2 32872 32312 32872 32312 0 _0307_
rlabel metal3 33936 30184 33936 30184 0 _0308_
rlabel metal2 29288 31416 29288 31416 0 _0309_
rlabel metal2 35560 32872 35560 32872 0 _0310_
rlabel metal3 32200 34776 32200 34776 0 _0311_
rlabel metal2 33096 32088 33096 32088 0 _0312_
rlabel metal2 32480 31528 32480 31528 0 _0313_
rlabel metal3 43288 23128 43288 23128 0 _0314_
rlabel metal2 42840 21448 42840 21448 0 _0315_
rlabel metal2 42504 25424 42504 25424 0 _0316_
rlabel metal2 44072 28560 44072 28560 0 _0317_
rlabel metal2 43680 24920 43680 24920 0 _0318_
rlabel metal2 42056 22680 42056 22680 0 _0319_
rlabel metal2 45080 20384 45080 20384 0 _0320_
rlabel metal2 45752 16576 45752 16576 0 _0321_
rlabel metal2 43904 18424 43904 18424 0 _0322_
rlabel metal3 46144 15288 46144 15288 0 _0323_
rlabel metal2 39256 17528 39256 17528 0 _0324_
rlabel metal2 41832 18760 41832 18760 0 _0325_
rlabel metal2 38528 23128 38528 23128 0 _0326_
rlabel metal2 43288 17304 43288 17304 0 _0327_
rlabel metal2 42056 19096 42056 19096 0 _0328_
rlabel metal2 42952 18480 42952 18480 0 _0329_
rlabel metal2 43400 15568 43400 15568 0 _0330_
rlabel metal2 45192 18088 45192 18088 0 _0331_
rlabel metal2 44744 18928 44744 18928 0 _0332_
rlabel metal3 44912 25480 44912 25480 0 _0333_
rlabel metal2 46648 18592 46648 18592 0 _0334_
rlabel metal2 43960 20384 43960 20384 0 _0335_
rlabel metal2 43624 21000 43624 21000 0 _0336_
rlabel metal2 42952 24472 42952 24472 0 _0337_
rlabel metal2 42392 23240 42392 23240 0 _0338_
rlabel metal2 40824 21112 40824 21112 0 _0339_
rlabel metal2 37688 20272 37688 20272 0 _0340_
rlabel metal3 11144 39592 11144 39592 0 _0341_
rlabel metal2 15176 34440 15176 34440 0 _0342_
rlabel metal3 7728 33208 7728 33208 0 _0343_
rlabel metal2 10248 32872 10248 32872 0 _0344_
rlabel via2 12376 33432 12376 33432 0 _0345_
rlabel metal2 8176 39368 8176 39368 0 _0346_
rlabel metal2 7560 39144 7560 39144 0 _0347_
rlabel metal2 8008 35952 8008 35952 0 _0348_
rlabel metal2 11592 36064 11592 36064 0 _0349_
rlabel metal3 11928 36680 11928 36680 0 _0350_
rlabel metal3 12320 35672 12320 35672 0 _0351_
rlabel metal2 12152 33432 12152 33432 0 _0352_
rlabel metal2 17640 30576 17640 30576 0 _0353_
rlabel metal3 18816 26824 18816 26824 0 _0354_
rlabel metal2 18088 31192 18088 31192 0 _0355_
rlabel metal2 16408 28448 16408 28448 0 _0356_
rlabel metal2 17416 28896 17416 28896 0 _0357_
rlabel metal2 19096 28224 19096 28224 0 _0358_
rlabel metal3 19432 28672 19432 28672 0 _0359_
rlabel metal2 18200 30800 18200 30800 0 _0360_
rlabel metal3 18592 29624 18592 29624 0 _0361_
rlabel metal2 15400 29008 15400 29008 0 _0362_
rlabel metal2 15064 31416 15064 31416 0 _0363_
rlabel metal2 13832 30184 13832 30184 0 _0364_
rlabel metal2 15624 27944 15624 27944 0 _0365_
rlabel metal2 13944 30912 13944 30912 0 _0366_
rlabel metal3 15260 31528 15260 31528 0 _0367_
rlabel metal2 12600 33936 12600 33936 0 _0368_
rlabel metal2 12936 33320 12936 33320 0 _0369_
rlabel metal2 17976 25816 17976 25816 0 _0370_
rlabel metal2 16072 25648 16072 25648 0 _0371_
rlabel metal2 15624 31248 15624 31248 0 _0372_
rlabel metal2 15288 31752 15288 31752 0 _0373_
rlabel metal2 14616 32256 14616 32256 0 _0374_
rlabel metal2 15176 10304 15176 10304 0 _0375_
rlabel metal2 16688 16184 16688 16184 0 _0376_
rlabel metal2 14952 9968 14952 9968 0 _0377_
rlabel metal2 17976 9744 17976 9744 0 _0378_
rlabel metal3 16856 9016 16856 9016 0 _0379_
rlabel metal2 16968 16296 16968 16296 0 _0380_
rlabel metal2 14392 10248 14392 10248 0 _0381_
rlabel metal3 13440 13832 13440 13832 0 _0382_
rlabel metal2 6776 17192 6776 17192 0 _0383_
rlabel metal3 9408 15288 9408 15288 0 _0384_
rlabel metal3 6944 15400 6944 15400 0 _0385_
rlabel metal2 7448 17192 7448 17192 0 _0386_
rlabel metal2 7168 15400 7168 15400 0 _0387_
rlabel metal2 8064 16632 8064 16632 0 _0388_
rlabel metal2 7784 14056 7784 14056 0 _0389_
rlabel metal3 7056 13720 7056 13720 0 _0390_
rlabel metal2 7448 14000 7448 14000 0 _0391_
rlabel metal2 7112 14896 7112 14896 0 _0392_
rlabel metal2 11032 21952 11032 21952 0 _0393_
rlabel metal2 12712 14336 12712 14336 0 _0394_
rlabel metal2 6328 15792 6328 15792 0 _0395_
rlabel metal2 2968 15568 2968 15568 0 _0396_
rlabel metal2 11480 18704 11480 18704 0 _0397_
rlabel metal2 11368 14168 11368 14168 0 _0398_
rlabel metal2 15624 16576 15624 16576 0 _0399_
rlabel metal2 14056 13104 14056 13104 0 _0400_
rlabel metal2 10136 15596 10136 15596 0 _0401_
rlabel metal2 12936 15204 12936 15204 0 _0402_
rlabel metal3 12208 15512 12208 15512 0 _0403_
rlabel metal2 12376 14000 12376 14000 0 _0404_
rlabel metal3 12880 13160 12880 13160 0 _0405_
rlabel metal2 11816 10976 11816 10976 0 _0406_
rlabel metal2 12264 15204 12264 15204 0 _0407_
rlabel metal2 12376 14896 12376 14896 0 _0408_
rlabel metal2 14336 16744 14336 16744 0 _0409_
rlabel metal2 13664 18536 13664 18536 0 _0410_
rlabel metal3 11480 18424 11480 18424 0 _0411_
rlabel metal2 9912 19544 9912 19544 0 _0412_
rlabel metal3 15484 12824 15484 12824 0 _0413_
rlabel metal2 10136 12992 10136 12992 0 _0414_
rlabel metal2 10472 13328 10472 13328 0 _0415_
rlabel metal2 9912 13104 9912 13104 0 _0416_
rlabel metal2 13944 16660 13944 16660 0 _0417_
rlabel metal2 15176 8008 15176 8008 0 _0418_
rlabel metal2 14392 9352 14392 9352 0 _0419_
rlabel metal2 44296 17248 44296 17248 0 _0420_
rlabel metal2 44968 17248 44968 17248 0 _0421_
rlabel metal2 42840 17136 42840 17136 0 _0422_
rlabel metal2 44352 18536 44352 18536 0 _0423_
rlabel metal2 43232 19992 43232 19992 0 _0424_
rlabel metal2 41832 20384 41832 20384 0 _0425_
rlabel metal2 43400 16632 43400 16632 0 _0426_
rlabel metal2 32312 12992 32312 12992 0 _0427_
rlabel metal2 35336 9856 35336 9856 0 _0428_
rlabel metal2 33488 11256 33488 11256 0 _0429_
rlabel metal2 34104 17136 34104 17136 0 _0430_
rlabel metal3 34552 12264 34552 12264 0 _0431_
rlabel metal3 33040 14504 33040 14504 0 _0432_
rlabel metal3 36792 11144 36792 11144 0 _0433_
rlabel metal2 37576 6776 37576 6776 0 _0434_
rlabel metal3 38808 12040 38808 12040 0 _0435_
rlabel metal2 37016 12320 37016 12320 0 _0436_
rlabel metal2 37184 11368 37184 11368 0 _0437_
rlabel metal3 35056 11256 35056 11256 0 _0438_
rlabel metal2 32088 13104 32088 13104 0 _0439_
rlabel metal2 27832 10976 27832 10976 0 _0440_
rlabel metal2 28616 10584 28616 10584 0 _0441_
rlabel metal2 27608 9576 27608 9576 0 _0442_
rlabel metal3 23632 9800 23632 9800 0 _0443_
rlabel metal2 29512 11312 29512 11312 0 _0444_
rlabel metal2 27776 16968 27776 16968 0 _0445_
rlabel metal3 25032 14504 25032 14504 0 _0446_
rlabel metal3 29120 12152 29120 12152 0 _0447_
rlabel metal2 33768 11480 33768 11480 0 _0448_
rlabel metal2 33992 12936 33992 12936 0 _0449_
rlabel metal2 31080 12544 31080 12544 0 _0450_
rlabel metal2 31416 12768 31416 12768 0 _0451_
rlabel metal3 25368 15288 25368 15288 0 _0452_
rlabel metal2 24136 12824 24136 12824 0 _0453_
rlabel metal2 27720 16688 27720 16688 0 _0454_
rlabel metal2 24248 12656 24248 12656 0 _0455_
rlabel metal2 26488 12264 26488 12264 0 _0456_
rlabel metal3 28336 9800 28336 9800 0 _0457_
rlabel metal3 25144 12936 25144 12936 0 _0458_
rlabel metal2 25256 13608 25256 13608 0 _0459_
rlabel metal2 23128 16576 23128 16576 0 _0460_
rlabel metal2 26600 13272 26600 13272 0 _0461_
rlabel metal2 29512 13384 29512 13384 0 _0462_
rlabel metal2 29960 13440 29960 13440 0 _0463_
rlabel metal2 13440 18424 13440 18424 0 _0464_
rlabel metal2 37128 18536 37128 18536 0 _0465_
rlabel metal2 39144 11424 39144 11424 0 _0466_
rlabel metal2 36120 13048 36120 13048 0 _0467_
rlabel metal3 33600 10696 33600 10696 0 _0468_
rlabel metal2 29176 10864 29176 10864 0 _0469_
rlabel metal3 30408 11368 30408 11368 0 _0470_
rlabel metal3 26236 12040 26236 12040 0 _0471_
rlabel metal2 30520 11648 30520 11648 0 _0472_
rlabel metal3 31416 11368 31416 11368 0 _0473_
rlabel metal2 36008 13048 36008 13048 0 _0474_
rlabel metal3 36624 15848 36624 15848 0 _0475_
rlabel metal3 36792 19880 36792 19880 0 _0476_
rlabel metal2 10024 32984 10024 32984 0 _0477_
rlabel metal2 13720 32480 13720 32480 0 _0478_
rlabel metal3 9744 38808 9744 38808 0 _0479_
rlabel metal3 9408 38136 9408 38136 0 _0480_
rlabel metal2 5768 33376 5768 33376 0 _0481_
rlabel metal2 9912 33600 9912 33600 0 _0482_
rlabel metal2 11480 33768 11480 33768 0 _0483_
rlabel metal2 11816 32872 11816 32872 0 _0484_
rlabel metal2 13440 30968 13440 30968 0 _0485_
rlabel metal3 21000 30968 21000 30968 0 _0486_
rlabel metal2 37240 30464 37240 30464 0 _0487_
rlabel metal2 37688 38724 37688 38724 0 _0488_
rlabel metal2 36232 40320 36232 40320 0 _0489_
rlabel metal2 48160 44744 48160 44744 0 _0490_
rlabel metal3 31696 38696 31696 38696 0 _0491_
rlabel metal2 10920 6776 10920 6776 0 _0492_
rlabel metal2 12712 21896 12712 21896 0 _0493_
rlabel metal2 12432 21784 12432 21784 0 _0494_
rlabel metal3 13384 21448 13384 21448 0 _0495_
rlabel metal3 16688 25480 16688 25480 0 _0496_
rlabel metal2 26824 32032 26824 32032 0 _0497_
rlabel metal2 18536 35560 18536 35560 0 _0498_
rlabel metal3 20328 29288 20328 29288 0 _0499_
rlabel metal3 13440 22232 13440 22232 0 _0500_
rlabel metal2 12040 21784 12040 21784 0 _0501_
rlabel metal2 11592 21840 11592 21840 0 _0502_
rlabel metal2 7000 6664 7000 6664 0 _0503_
rlabel metal2 23016 9240 23016 9240 0 _0504_
rlabel metal2 11480 7392 11480 7392 0 _0505_
rlabel metal3 8008 6552 8008 6552 0 _0506_
rlabel metal3 8960 8232 8960 8232 0 _0507_
rlabel metal2 7112 8232 7112 8232 0 _0508_
rlabel metal3 9744 8008 9744 8008 0 _0509_
rlabel metal2 8120 8232 8120 8232 0 _0510_
rlabel metal2 7896 4592 7896 4592 0 _0511_
rlabel metal2 8624 4424 8624 4424 0 _0512_
rlabel metal2 9688 8232 9688 8232 0 _0513_
rlabel metal2 10920 7896 10920 7896 0 _0514_
rlabel metal3 10136 4312 10136 4312 0 _0515_
rlabel metal2 17080 7000 17080 7000 0 _0516_
rlabel metal2 11256 4760 11256 4760 0 _0517_
rlabel metal2 13048 7616 13048 7616 0 _0518_
rlabel metal3 13440 7448 13440 7448 0 _0519_
rlabel metal2 26600 5936 26600 5936 0 _0520_
rlabel metal2 20328 5936 20328 5936 0 _0521_
rlabel metal2 19544 4648 19544 4648 0 _0522_
rlabel metal2 26376 6328 26376 6328 0 _0523_
rlabel metal2 20104 4480 20104 4480 0 _0524_
rlabel metal2 21112 4592 21112 4592 0 _0525_
rlabel metal2 23688 17024 23688 17024 0 _0526_
rlabel metal2 20552 4760 20552 4760 0 _0527_
rlabel metal2 23576 5880 23576 5880 0 _0528_
rlabel metal2 26152 6944 26152 6944 0 _0529_
rlabel metal2 29624 6608 29624 6608 0 _0530_
rlabel metal2 24360 6384 24360 6384 0 _0531_
rlabel metal2 26824 5544 26824 5544 0 _0532_
rlabel metal2 27272 5376 27272 5376 0 _0533_
rlabel metal3 32648 6440 32648 6440 0 _0534_
rlabel metal2 27944 5768 27944 5768 0 _0535_
rlabel metal2 29064 5376 29064 5376 0 _0536_
rlabel metal2 29624 5264 29624 5264 0 _0537_
rlabel metal2 30296 5376 30296 5376 0 _0538_
rlabel metal2 31416 5992 31416 5992 0 _0539_
rlabel metal2 33432 5208 33432 5208 0 _0540_
rlabel metal2 43176 7224 43176 7224 0 _0541_
rlabel metal2 34216 6216 34216 6216 0 _0542_
rlabel metal2 35000 6216 35000 6216 0 _0543_
rlabel metal2 35224 6384 35224 6384 0 _0544_
rlabel metal2 47824 17640 47824 17640 0 _0545_
rlabel metal2 43848 10808 43848 10808 0 _0546_
rlabel metal2 41720 6664 41720 6664 0 _0547_
rlabel metal2 46424 14112 46424 14112 0 _0548_
rlabel metal2 42672 6664 42672 6664 0 _0549_
rlabel metal2 42280 8232 42280 8232 0 _0550_
rlabel metal3 43456 8120 43456 8120 0 _0551_
rlabel metal2 44632 10024 44632 10024 0 _0552_
rlabel metal2 44072 34216 44072 34216 0 _0553_
rlabel metal2 47936 23912 47936 23912 0 _0554_
rlabel metal2 43624 11872 43624 11872 0 _0555_
rlabel metal2 46536 24304 46536 24304 0 _0556_
rlabel metal3 45472 17640 45472 17640 0 _0557_
rlabel metal2 47096 17024 47096 17024 0 _0558_
rlabel metal2 39256 20272 39256 20272 0 _0559_
rlabel metal2 47208 17976 47208 17976 0 _0560_
rlabel metal3 45808 19992 45808 19992 0 _0561_
rlabel metal2 46760 19656 46760 19656 0 _0562_
rlabel metal2 44968 23576 44968 23576 0 _0563_
rlabel metal2 46984 23912 46984 23912 0 _0564_
rlabel metal2 46088 24696 46088 24696 0 _0565_
rlabel metal2 45864 25536 45864 25536 0 _0566_
rlabel metal2 47656 24192 47656 24192 0 _0567_
rlabel metal3 47096 24696 47096 24696 0 _0568_
rlabel metal3 44744 12264 44744 12264 0 _0569_
rlabel metal2 45304 12936 45304 12936 0 _0570_
rlabel metal3 26824 37352 26824 37352 0 _0571_
rlabel metal2 15344 27832 15344 27832 0 _0572_
rlabel metal2 3080 28728 3080 28728 0 _0573_
rlabel metal3 9184 36456 9184 36456 0 _0574_
rlabel metal3 6216 38920 6216 38920 0 _0575_
rlabel metal2 7560 37632 7560 37632 0 _0576_
rlabel metal3 7224 38808 7224 38808 0 _0577_
rlabel metal3 7672 38696 7672 38696 0 _0578_
rlabel metal3 7672 38024 7672 38024 0 _0579_
rlabel metal2 8904 28896 8904 28896 0 _0580_
rlabel metal2 4872 30296 4872 30296 0 _0581_
rlabel metal2 7168 31192 7168 31192 0 _0582_
rlabel metal2 7784 35784 7784 35784 0 _0583_
rlabel metal2 10808 28056 10808 28056 0 _0584_
rlabel metal2 9688 27608 9688 27608 0 _0585_
rlabel metal3 10192 27832 10192 27832 0 _0586_
rlabel metal3 10304 25480 10304 25480 0 _0587_
rlabel metal3 10080 27160 10080 27160 0 _0588_
rlabel metal2 10584 19488 10584 19488 0 _0589_
rlabel metal2 3304 20832 3304 20832 0 _0590_
rlabel metal2 5992 21112 5992 21112 0 _0591_
rlabel metal3 7896 18648 7896 18648 0 _0592_
rlabel metal2 6888 17976 6888 17976 0 _0593_
rlabel metal3 10136 19432 10136 19432 0 _0594_
rlabel metal3 7560 22904 7560 22904 0 _0595_
rlabel metal2 8232 23408 8232 23408 0 _0596_
rlabel metal2 8568 19208 8568 19208 0 _0597_
rlabel metal2 11368 25704 11368 25704 0 _0598_
rlabel metal2 10808 21728 10808 21728 0 _0599_
rlabel metal3 13048 19208 13048 19208 0 _0600_
rlabel metal3 7168 20104 7168 20104 0 _0601_
rlabel metal2 10584 18704 10584 18704 0 _0602_
rlabel metal3 11424 19320 11424 19320 0 _0603_
rlabel metal2 8568 20160 8568 20160 0 _0604_
rlabel metal3 9632 19992 9632 19992 0 _0605_
rlabel metal2 11200 19432 11200 19432 0 _0606_
rlabel metal2 10304 18424 10304 18424 0 _0607_
rlabel metal2 8288 18312 8288 18312 0 _0608_
rlabel metal3 9240 18424 9240 18424 0 _0609_
rlabel metal2 10472 18872 10472 18872 0 _0610_
rlabel metal2 17640 18760 17640 18760 0 _0611_
rlabel metal2 17416 17696 17416 17696 0 _0612_
rlabel metal2 16856 20272 16856 20272 0 _0613_
rlabel metal2 17472 16856 17472 16856 0 _0614_
rlabel metal3 15680 20776 15680 20776 0 _0615_
rlabel metal2 16128 17080 16128 17080 0 _0616_
rlabel metal3 16800 16744 16800 16744 0 _0617_
rlabel metal2 18032 17080 18032 17080 0 _0618_
rlabel metal2 16744 17248 16744 17248 0 _0619_
rlabel metal2 29624 17976 29624 17976 0 _0620_
rlabel metal2 29344 20440 29344 20440 0 _0621_
rlabel metal2 27384 18200 27384 18200 0 _0622_
rlabel metal3 25704 18200 25704 18200 0 _0623_
rlabel metal2 24360 18256 24360 18256 0 _0624_
rlabel metal2 25592 16520 25592 16520 0 _0625_
rlabel metal2 22904 22232 22904 22232 0 _0626_
rlabel metal2 22680 19208 22680 19208 0 _0627_
rlabel metal2 25368 16744 25368 16744 0 _0628_
rlabel metal3 24640 17640 24640 17640 0 _0629_
rlabel metal2 26600 17752 26600 17752 0 _0630_
rlabel metal2 29456 20888 29456 20888 0 _0631_
rlabel metal2 30296 16408 30296 16408 0 _0632_
rlabel metal2 29568 15960 29568 15960 0 _0633_
rlabel metal2 27832 22064 27832 22064 0 _0634_
rlabel metal3 28896 15848 28896 15848 0 _0635_
rlabel metal2 30520 17416 30520 17416 0 _0636_
rlabel metal2 31752 23240 31752 23240 0 _0637_
rlabel metal2 30352 19208 30352 19208 0 _0638_
rlabel metal2 29736 16408 29736 16408 0 _0639_
rlabel metal2 29960 17024 29960 17024 0 _0640_
rlabel metal2 25144 16912 25144 16912 0 _0641_
rlabel metal2 27048 16520 27048 16520 0 _0642_
rlabel metal2 27608 16464 27608 16464 0 _0643_
rlabel metal2 27944 17024 27944 17024 0 _0644_
rlabel metal2 30184 18312 30184 18312 0 _0645_
rlabel metal2 30968 17696 30968 17696 0 _0646_
rlabel metal2 38472 24528 38472 24528 0 _0647_
rlabel metal2 37016 25032 37016 25032 0 _0648_
rlabel metal2 39368 25536 39368 25536 0 _0649_
rlabel metal3 38136 22232 38136 22232 0 _0650_
rlabel metal2 39424 23352 39424 23352 0 _0651_
rlabel metal2 41160 24472 41160 24472 0 _0652_
rlabel metal2 40936 25872 40936 25872 0 _0653_
rlabel metal2 41048 24752 41048 24752 0 _0654_
rlabel metal2 38808 25032 38808 25032 0 _0655_
rlabel metal2 38360 23912 38360 23912 0 _0656_
rlabel metal2 38248 25088 38248 25088 0 _0657_
rlabel metal2 39200 27832 39200 27832 0 _0658_
rlabel metal2 39032 20048 39032 20048 0 _0659_
rlabel metal2 37912 20888 37912 20888 0 _0660_
rlabel metal2 38248 20888 38248 20888 0 _0661_
rlabel metal2 39088 20216 39088 20216 0 _0662_
rlabel metal3 38976 20664 38976 20664 0 _0663_
rlabel metal2 38472 21168 38472 21168 0 _0664_
rlabel metal2 42896 26264 42896 26264 0 _0665_
rlabel metal2 38920 28952 38920 28952 0 _0666_
rlabel metal2 37912 28840 37912 28840 0 _0667_
rlabel metal2 38696 28280 38696 28280 0 _0668_
rlabel metal2 39984 27608 39984 27608 0 _0669_
rlabel metal2 39592 27384 39592 27384 0 _0670_
rlabel metal2 36904 26936 36904 26936 0 _0671_
rlabel metal2 39424 21560 39424 21560 0 _0672_
rlabel metal2 38976 21784 38976 21784 0 _0673_
rlabel metal2 38920 25144 38920 25144 0 _0674_
rlabel metal3 39816 26264 39816 26264 0 _0675_
rlabel metal3 37184 29400 37184 29400 0 _0676_
rlabel metal3 37688 27832 37688 27832 0 _0677_
rlabel metal3 31024 26488 31024 26488 0 _0678_
rlabel metal3 24192 40600 24192 40600 0 _0679_
rlabel metal3 23688 40936 23688 40936 0 _0680_
rlabel metal2 24248 32312 24248 32312 0 _0681_
rlabel metal3 25032 32312 25032 32312 0 _0682_
rlabel metal2 25256 40824 25256 40824 0 _0683_
rlabel metal2 24416 36232 24416 36232 0 _0684_
rlabel metal2 25536 33208 25536 33208 0 _0685_
rlabel metal3 22512 38808 22512 38808 0 _0686_
rlabel metal3 26208 23912 26208 23912 0 _0687_
rlabel metal2 26600 42000 26600 42000 0 _0688_
rlabel metal2 26488 38696 26488 38696 0 _0689_
rlabel metal3 21728 39592 21728 39592 0 _0690_
rlabel metal2 23576 42672 23576 42672 0 _0691_
rlabel metal2 27384 40488 27384 40488 0 _0692_
rlabel metal2 26880 41384 26880 41384 0 _0693_
rlabel metal2 26712 39816 26712 39816 0 _0694_
rlabel metal2 25032 41104 25032 41104 0 _0695_
rlabel metal2 26152 41216 26152 41216 0 _0696_
rlabel metal2 27608 41216 27608 41216 0 _0697_
rlabel metal2 23464 43232 23464 43232 0 _0698_
rlabel metal3 28448 43512 28448 43512 0 _0699_
rlabel metal2 27328 42728 27328 42728 0 _0700_
rlabel metal2 27160 43232 27160 43232 0 _0701_
rlabel metal2 27608 43736 27608 43736 0 _0702_
rlabel metal2 25032 42952 25032 42952 0 _0703_
rlabel metal2 19376 42728 19376 42728 0 _0704_
rlabel metal2 25816 43008 25816 43008 0 _0705_
rlabel metal2 25592 43176 25592 43176 0 _0706_
rlabel metal2 25200 43624 25200 43624 0 _0707_
rlabel metal2 23240 42504 23240 42504 0 _0708_
rlabel metal2 19880 43008 19880 43008 0 _0709_
rlabel metal2 22680 42896 22680 42896 0 _0710_
rlabel metal2 20328 43064 20328 43064 0 _0711_
rlabel metal2 22512 42840 22512 42840 0 _0712_
rlabel metal2 22624 43736 22624 43736 0 _0713_
rlabel metal3 17584 43400 17584 43400 0 _0714_
rlabel metal2 18424 43904 18424 43904 0 _0715_
rlabel metal2 21056 44296 21056 44296 0 _0716_
rlabel metal3 20328 44296 20328 44296 0 _0717_
rlabel metal2 18592 44296 18592 44296 0 _0718_
rlabel metal2 19712 39368 19712 39368 0 _0719_
rlabel metal3 17192 43512 17192 43512 0 _0720_
rlabel metal2 20048 42168 20048 42168 0 _0721_
rlabel metal2 20216 41776 20216 41776 0 _0722_
rlabel metal2 17416 43176 17416 43176 0 _0723_
rlabel metal2 17640 41104 17640 41104 0 _0724_
rlabel metal2 20944 41944 20944 41944 0 _0725_
rlabel metal2 21336 41496 21336 41496 0 _0726_
rlabel metal2 17416 41888 17416 41888 0 _0727_
rlabel metal2 19992 39648 19992 39648 0 _0728_
rlabel metal2 20272 39592 20272 39592 0 _0729_
rlabel metal2 18648 38724 18648 38724 0 _0730_
rlabel metal2 19768 36624 19768 36624 0 _0731_
rlabel metal2 23800 35896 23800 35896 0 _0732_
rlabel metal2 25032 34328 25032 34328 0 _0733_
rlabel metal2 24696 35784 24696 35784 0 _0734_
rlabel metal2 23128 34104 23128 34104 0 _0735_
rlabel metal2 24360 36624 24360 36624 0 _0736_
rlabel metal2 20272 36680 20272 36680 0 _0737_
rlabel metal2 26656 35560 26656 35560 0 _0738_
rlabel metal2 23240 35896 23240 35896 0 _0739_
rlabel metal3 22680 35448 22680 35448 0 _0740_
rlabel metal2 19880 35168 19880 35168 0 _0741_
rlabel metal2 19712 35000 19712 35000 0 _0742_
rlabel metal2 22904 31304 22904 31304 0 _0743_
rlabel metal2 23128 24248 23128 24248 0 _0744_
rlabel metal2 22680 31080 22680 31080 0 _0745_
rlabel metal3 18424 37352 18424 37352 0 _0746_
rlabel metal2 19152 26488 19152 26488 0 _0747_
rlabel metal2 19432 32536 19432 32536 0 _0748_
rlabel metal2 35672 31080 35672 31080 0 _0749_
rlabel metal2 34216 30464 34216 30464 0 _0750_
rlabel metal2 42280 30016 42280 30016 0 _0751_
rlabel metal3 36736 29960 36736 29960 0 _0752_
rlabel metal2 42616 25928 42616 25928 0 _0753_
rlabel metal3 43568 27160 43568 27160 0 _0754_
rlabel metal2 42616 27496 42616 27496 0 _0755_
rlabel metal2 41496 27608 41496 27608 0 _0756_
rlabel metal3 15680 25256 15680 25256 0 _0757_
rlabel metal2 15960 26320 15960 26320 0 _0758_
rlabel metal2 16968 26600 16968 26600 0 _0759_
rlabel metal2 16408 24920 16408 24920 0 _0760_
rlabel metal3 17248 26264 17248 26264 0 _0761_
rlabel metal2 15512 27832 15512 27832 0 _0762_
rlabel metal3 15428 15176 15428 15176 0 _0763_
rlabel metal2 15232 26824 15232 26824 0 _0764_
rlabel metal2 15512 25368 15512 25368 0 _0765_
rlabel metal2 13496 34608 13496 34608 0 _0766_
rlabel metal2 9240 36064 9240 36064 0 _0767_
rlabel metal2 10696 35000 10696 35000 0 _0768_
rlabel metal2 15064 26544 15064 26544 0 _0769_
rlabel metal2 15512 16240 15512 16240 0 _0770_
rlabel metal2 16072 11536 16072 11536 0 _0771_
rlabel metal2 15624 10976 15624 10976 0 _0772_
rlabel metal3 13160 11256 13160 11256 0 _0773_
rlabel metal2 13720 11592 13720 11592 0 _0774_
rlabel metal2 13664 15848 13664 15848 0 _0775_
rlabel metal2 10024 16016 10024 16016 0 _0776_
rlabel metal2 7896 16408 7896 16408 0 _0777_
rlabel metal2 8904 17584 8904 17584 0 _0778_
rlabel metal2 10920 16744 10920 16744 0 _0779_
rlabel metal2 10584 16520 10584 16520 0 _0780_
rlabel metal2 11592 15736 11592 15736 0 _0781_
rlabel metal2 12824 15960 12824 15960 0 _0782_
rlabel metal2 13496 16520 13496 16520 0 _0783_
rlabel metal3 15008 16184 15008 16184 0 _0784_
rlabel metal3 17248 11480 17248 11480 0 _0785_
rlabel metal2 18200 12880 18200 12880 0 _0786_
rlabel metal2 15512 11536 15512 11536 0 _0787_
rlabel metal2 15848 11760 15848 11760 0 _0788_
rlabel metal2 16408 15596 16408 15596 0 _0789_
rlabel metal2 16184 15736 16184 15736 0 _0790_
rlabel metal2 35896 14000 35896 14000 0 _0791_
rlabel metal2 35784 10192 35784 10192 0 _0792_
rlabel metal2 35112 12880 35112 12880 0 _0793_
rlabel metal2 36120 14280 36120 14280 0 _0794_
rlabel metal2 34440 13440 34440 13440 0 _0795_
rlabel metal2 34888 14168 34888 14168 0 _0796_
rlabel metal3 33712 14392 33712 14392 0 _0797_
rlabel metal2 27384 15344 27384 15344 0 _0798_
rlabel metal2 27496 15204 27496 15204 0 _0799_
rlabel metal2 25592 15120 25592 15120 0 _0800_
rlabel metal2 24808 14728 24808 14728 0 _0801_
rlabel metal2 26824 14672 26824 14672 0 _0802_
rlabel metal2 26376 15064 26376 15064 0 _0803_
rlabel metal2 28168 14000 28168 14000 0 _0804_
rlabel metal2 33208 14896 33208 14896 0 _0805_
rlabel metal2 27384 14784 27384 14784 0 _0806_
rlabel metal2 25816 9408 25816 9408 0 _0807_
rlabel metal2 26376 12712 26376 12712 0 _0808_
rlabel metal3 30856 14280 30856 14280 0 _0809_
rlabel metal2 35336 14224 35336 14224 0 _0810_
rlabel metal3 35168 14616 35168 14616 0 _0811_
rlabel metal2 34104 15512 34104 15512 0 _0812_
rlabel metal2 33320 15736 33320 15736 0 _0813_
rlabel metal3 44184 16072 44184 16072 0 _0814_
rlabel metal2 42504 15624 42504 15624 0 _0815_
rlabel metal2 43344 12376 43344 12376 0 _0816_
rlabel metal3 42784 15288 42784 15288 0 _0817_
rlabel metal2 38024 16800 38024 16800 0 _0818_
rlabel metal2 36008 16184 36008 16184 0 _0819_
rlabel metal2 42168 16800 42168 16800 0 _0820_
rlabel metal2 39368 16072 39368 16072 0 _0821_
rlabel metal2 41048 16016 41048 16016 0 _0822_
rlabel metal2 40824 15792 40824 15792 0 _0823_
rlabel metal3 42168 16184 42168 16184 0 _0824_
rlabel metal2 42056 15904 42056 15904 0 _0825_
rlabel metal2 41496 16408 41496 16408 0 _0826_
rlabel metal2 40936 16408 40936 16408 0 _0827_
rlabel metal2 42168 27384 42168 27384 0 _0828_
rlabel metal2 32424 29400 32424 29400 0 _0829_
rlabel metal3 32200 30072 32200 30072 0 _0830_
rlabel metal2 34664 34104 34664 34104 0 _0831_
rlabel metal2 33320 30912 33320 30912 0 _0832_
rlabel metal2 31360 31752 31360 31752 0 _0833_
rlabel metal2 30464 30408 30464 30408 0 _0834_
rlabel metal2 29512 30744 29512 30744 0 _0835_
rlabel metal3 28560 30856 28560 30856 0 _0836_
rlabel metal2 27720 31136 27720 31136 0 _0837_
rlabel metal3 32592 33208 32592 33208 0 _0838_
rlabel metal3 29848 31528 29848 31528 0 _0839_
rlabel metal3 29848 31864 29848 31864 0 _0840_
rlabel metal2 29736 32984 29736 32984 0 _0841_
rlabel metal2 30968 33936 30968 33936 0 _0842_
rlabel metal2 30912 35560 30912 35560 0 _0843_
rlabel metal3 33712 31976 33712 31976 0 _0844_
rlabel metal2 34104 32648 34104 32648 0 _0845_
rlabel metal2 34720 31528 34720 31528 0 _0846_
rlabel metal2 35056 31864 35056 31864 0 _0847_
rlabel metal2 2632 39144 2632 39144 0 _0848_
rlabel metal2 24080 28056 24080 28056 0 _0849_
rlabel metal3 20160 23912 20160 23912 0 _0850_
rlabel metal2 2856 29344 2856 29344 0 _0851_
rlabel metal3 4704 39816 4704 39816 0 _0852_
rlabel metal2 2408 38528 2408 38528 0 _0853_
rlabel metal2 3192 37856 3192 37856 0 _0854_
rlabel metal3 3584 38808 3584 38808 0 _0855_
rlabel metal2 25032 25536 25032 25536 0 _0856_
rlabel metal2 2856 30576 2856 30576 0 _0857_
rlabel metal2 5264 35560 5264 35560 0 _0858_
rlabel metal2 4984 36120 4984 36120 0 _0859_
rlabel metal2 3024 30408 3024 30408 0 _0860_
rlabel metal2 3304 31024 3304 31024 0 _0861_
rlabel metal2 2520 29008 2520 29008 0 _0862_
rlabel metal2 5992 25984 5992 25984 0 _0863_
rlabel metal2 4648 28672 4648 28672 0 _0864_
rlabel metal3 6440 23912 6440 23912 0 _0865_
rlabel metal2 5600 25704 5600 25704 0 _0866_
rlabel metal2 7896 25032 7896 25032 0 _0867_
rlabel metal2 2968 23184 2968 23184 0 _0868_
rlabel metal2 5544 23408 5544 23408 0 _0869_
rlabel metal3 3920 23016 3920 23016 0 _0870_
rlabel metal2 18872 21280 18872 21280 0 _0871_
rlabel metal2 5712 21560 5712 21560 0 _0872_
rlabel metal2 4872 20440 4872 20440 0 _0873_
rlabel metal2 4984 21168 4984 21168 0 _0874_
rlabel metal2 2856 20412 2856 20412 0 _0875_
rlabel metal2 6328 21392 6328 21392 0 _0876_
rlabel metal2 15400 20720 15400 20720 0 _0877_
rlabel metal2 6440 20776 6440 20776 0 _0878_
rlabel metal2 14616 21056 14616 21056 0 _0879_
rlabel metal2 18312 21112 18312 21112 0 _0880_
rlabel metal2 17416 22568 17416 22568 0 _0881_
rlabel metal2 19880 20832 19880 20832 0 _0882_
rlabel metal3 20496 20664 20496 20664 0 _0883_
rlabel metal3 21672 21000 21672 21000 0 _0884_
rlabel metal2 22232 22960 22232 22960 0 _0885_
rlabel metal2 22344 23520 22344 23520 0 _0886_
rlabel metal2 22120 25144 22120 25144 0 _0887_
rlabel metal2 23576 20776 23576 20776 0 _0888_
rlabel metal2 23352 20440 23352 20440 0 _0889_
rlabel metal2 20384 19432 20384 19432 0 _0890_
rlabel metal2 30744 20496 30744 20496 0 _0891_
rlabel metal3 25312 19432 25312 19432 0 _0892_
rlabel metal2 27160 19544 27160 19544 0 _0893_
rlabel metal2 29512 20412 29512 20412 0 _0894_
rlabel metal3 24976 24696 24976 24696 0 clk
rlabel metal2 29848 22484 29848 22484 0 clknet_0_clk
rlabel metal2 1848 12544 1848 12544 0 clknet_4_0_0_clk
rlabel metal2 40264 16436 40264 16436 0 clknet_4_10_0_clk
rlabel metal2 39704 22736 39704 22736 0 clknet_4_11_0_clk
rlabel metal2 33544 26040 33544 26040 0 clknet_4_12_0_clk
rlabel metal2 31976 43904 31976 43904 0 clknet_4_13_0_clk
rlabel metal2 45248 26264 45248 26264 0 clknet_4_14_0_clk
rlabel metal2 46536 38752 46536 38752 0 clknet_4_15_0_clk
rlabel metal2 1960 23912 1960 23912 0 clknet_4_1_0_clk
rlabel metal2 20048 16744 20048 16744 0 clknet_4_2_0_clk
rlabel metal2 20552 23184 20552 23184 0 clknet_4_3_0_clk
rlabel metal2 1848 29400 1848 29400 0 clknet_4_4_0_clk
rlabel metal2 1848 35616 1848 35616 0 clknet_4_5_0_clk
rlabel metal3 22288 27832 22288 27832 0 clknet_4_6_0_clk
rlabel metal2 21000 45080 21000 45080 0 clknet_4_7_0_clk
rlabel metal2 31864 16072 31864 16072 0 clknet_4_8_0_clk
rlabel metal2 31192 17696 31192 17696 0 clknet_4_9_0_clk
rlabel metal2 27272 40712 27272 40712 0 net1
rlabel metal2 24528 39816 24528 39816 0 net10
rlabel metal2 47096 15148 47096 15148 0 net100
rlabel metal2 45640 16744 45640 16744 0 net101
rlabel metal2 46088 21224 46088 21224 0 net102
rlabel via2 45864 23016 45864 23016 0 net103
rlabel metal2 10920 40488 10920 40488 0 net104
rlabel metal3 47096 27048 47096 27048 0 net105
rlabel metal2 43064 23660 43064 23660 0 net106
rlabel metal2 9016 40432 9016 40432 0 net107
rlabel metal2 15848 36344 15848 36344 0 net108
rlabel metal2 17640 39872 17640 39872 0 net109
rlabel metal3 13048 45640 13048 45640 0 net11
rlabel metal2 18088 35000 18088 35000 0 net110
rlabel metal3 17920 32424 17920 32424 0 net111
rlabel metal2 12600 24192 12600 24192 0 net112
rlabel metal3 10696 22456 10696 22456 0 net113
rlabel metal2 29176 42280 29176 42280 0 net114
rlabel metal3 46648 40376 46648 40376 0 net115
rlabel metal2 48272 45080 48272 45080 0 net116
rlabel metal2 38248 45024 38248 45024 0 net117
rlabel metal2 38920 44688 38920 44688 0 net118
rlabel metal2 34328 42616 34328 42616 0 net119
rlabel metal2 7112 3976 7112 3976 0 net12
rlabel metal2 32536 45080 32536 45080 0 net120
rlabel metal3 31360 45192 31360 45192 0 net121
rlabel metal2 46872 44632 46872 44632 0 net122
rlabel metal3 43568 34888 43568 34888 0 net123
rlabel metal3 31304 43512 31304 43512 0 net124
rlabel metal2 44240 33096 44240 33096 0 net125
rlabel metal2 47096 32816 47096 32816 0 net126
rlabel metal2 31528 43960 31528 43960 0 net127
rlabel metal2 45304 34944 45304 34944 0 net128
rlabel metal2 21224 30968 21224 30968 0 net129
rlabel metal3 4480 8120 4480 8120 0 net13
rlabel metal2 17976 39088 17976 39088 0 net130
rlabel metal3 17976 29904 17976 29904 0 net131
rlabel metal2 10696 40488 10696 40488 0 net132
rlabel metal2 10136 39088 10136 39088 0 net133
rlabel metal2 43848 23128 43848 23128 0 net134
rlabel metal3 42896 16968 42896 16968 0 net135
rlabel metal2 43624 7504 43624 7504 0 net136
rlabel metal2 26656 10584 26656 10584 0 net137
rlabel metal2 15960 7000 15960 7000 0 net138
rlabel metal3 12544 9800 12544 9800 0 net139
rlabel metal2 7728 3416 7728 3416 0 net14
rlabel metal2 7168 16072 7168 16072 0 net140
rlabel metal3 6384 21560 6384 21560 0 net141
rlabel metal2 41048 2058 41048 2058 0 net142
rlabel metal2 47208 45864 47208 45864 0 net143
rlabel metal3 47306 47096 47306 47096 0 net144
rlabel metal2 8792 5768 8792 5768 0 net15
rlabel metal2 9632 3416 9632 3416 0 net16
rlabel metal2 13160 4144 13160 4144 0 net17
rlabel metal2 19264 4536 19264 4536 0 net18
rlabel metal2 20216 3388 20216 3388 0 net19
rlabel metal2 28840 44464 28840 44464 0 net2
rlabel metal2 23688 3976 23688 3976 0 net20
rlabel metal2 24920 4592 24920 4592 0 net21
rlabel metal2 14504 44240 14504 44240 0 net22
rlabel metal2 31304 3976 31304 3976 0 net23
rlabel metal2 32200 4760 32200 4760 0 net24
rlabel metal2 35112 3808 35112 3808 0 net25
rlabel metal3 36400 4536 36400 4536 0 net26
rlabel metal2 42728 4200 42728 4200 0 net27
rlabel metal2 42056 8456 42056 8456 0 net28
rlabel metal2 44968 10304 44968 10304 0 net29
rlabel metal2 24808 43008 24808 43008 0 net3
rlabel metal3 45976 15960 45976 15960 0 net30
rlabel metal2 47880 19992 47880 19992 0 net31
rlabel metal2 44856 23688 44856 23688 0 net32
rlabel metal2 10024 42840 10024 42840 0 net33
rlabel metal2 45808 24696 45808 24696 0 net34
rlabel metal2 44296 12376 44296 12376 0 net35
rlabel metal2 9800 43064 9800 43064 0 net36
rlabel metal2 12096 40488 12096 40488 0 net37
rlabel metal2 15176 43064 15176 43064 0 net38
rlabel metal2 15008 37352 15008 37352 0 net39
rlabel metal2 23240 43344 23240 43344 0 net4
rlabel metal2 2072 34384 2072 34384 0 net40
rlabel metal2 2072 22456 2072 22456 0 net41
rlabel metal2 2072 20832 2072 20832 0 net42
rlabel metal2 21392 42168 21392 42168 0 net43
rlabel metal2 10304 4536 10304 4536 0 net44
rlabel metal2 27832 5376 27832 5376 0 net45
rlabel metal2 47544 18088 47544 18088 0 net46
rlabel metal2 28112 43680 28112 43680 0 net47
rlabel metal2 33824 40152 33824 40152 0 net48
rlabel metal2 48160 38920 48160 38920 0 net49
rlabel metal2 18536 43848 18536 43848 0 net5
rlabel metal2 35112 42840 35112 42840 0 net50
rlabel metal3 45080 34776 45080 34776 0 net51
rlabel metal2 32536 43792 32536 43792 0 net52
rlabel metal2 32200 44352 32200 44352 0 net53
rlabel metal2 40152 45808 40152 45808 0 net54
rlabel metal2 31584 41944 31584 41944 0 net55
rlabel metal3 35672 42616 35672 42616 0 net56
rlabel metal2 36456 41104 36456 41104 0 net57
rlabel metal2 38472 44632 38472 44632 0 net58
rlabel metal2 32872 45024 32872 45024 0 net59
rlabel metal2 16520 44352 16520 44352 0 net6
rlabel metal3 45528 36344 45528 36344 0 net60
rlabel metal2 38808 44184 38808 44184 0 net61
rlabel metal2 41496 42392 41496 42392 0 net62
rlabel metal2 42392 35280 42392 35280 0 net63
rlabel metal2 46536 44660 46536 44660 0 net64
rlabel metal2 30632 45192 30632 45192 0 net65
rlabel metal2 41720 40208 41720 40208 0 net66
rlabel metal2 41272 44632 41272 44632 0 net67
rlabel metal2 39256 45808 39256 45808 0 net68
rlabel metal2 44856 43904 44856 43904 0 net69
rlabel metal2 17416 40488 17416 40488 0 net7
rlabel metal2 32872 42672 32872 42672 0 net70
rlabel metal2 45696 42168 45696 42168 0 net71
rlabel metal2 37072 40600 37072 40600 0 net72
rlabel metal2 44800 39368 44800 39368 0 net73
rlabel metal3 42056 37912 42056 37912 0 net74
rlabel metal2 45360 40376 45360 40376 0 net75
rlabel metal2 40376 41944 40376 41944 0 net76
rlabel metal2 48104 41832 48104 41832 0 net77
rlabel metal3 35392 42168 35392 42168 0 net78
rlabel metal2 38024 43456 38024 43456 0 net79
rlabel metal2 18928 40600 18928 40600 0 net8
rlabel metal3 41440 39816 41440 39816 0 net80
rlabel metal2 23856 39592 23856 39592 0 net81
rlabel metal2 9688 37184 9688 37184 0 net82
rlabel metal2 4312 5768 4312 5768 0 net83
rlabel metal2 6440 17360 6440 17360 0 net84
rlabel metal3 10192 11256 10192 11256 0 net85
rlabel metal2 12320 9800 12320 9800 0 net86
rlabel metal2 15680 5096 15680 5096 0 net87
rlabel metal2 16408 8736 16408 8736 0 net88
rlabel metal2 19432 5600 19432 5600 0 net89
rlabel metal2 33768 39424 33768 39424 0 net9
rlabel metal3 25200 12264 25200 12264 0 net90
rlabel metal2 25704 9464 25704 9464 0 net91
rlabel metal2 25480 3864 25480 3864 0 net92
rlabel metal2 15288 42224 15288 42224 0 net93
rlabel metal3 31920 4200 31920 4200 0 net94
rlabel metal2 33544 5152 33544 5152 0 net95
rlabel metal2 34440 11704 34440 11704 0 net96
rlabel metal2 38472 4648 38472 4648 0 net97
rlabel metal2 43960 7056 43960 7056 0 net98
rlabel metal2 43568 16856 43568 16856 0 net99
rlabel metal2 48216 35784 48216 35784 0 recv_buf_data\[0\]
rlabel metal2 42840 36232 42840 36232 0 recv_buf_data\[1\]
rlabel metal2 47768 42336 47768 42336 0 recv_buf_data\[2\]
rlabel metal2 42392 39536 42392 39536 0 recv_buf_data\[3\]
rlabel metal3 42000 38920 42000 38920 0 recv_buf_data\[4\]
rlabel metal2 42056 42504 42056 42504 0 recv_buf_data\[5\]
rlabel metal2 39256 42392 39256 42392 0 recv_buf_data\[6\]
rlabel metal2 34664 41216 34664 41216 0 recv_buf_data\[7\]
rlabel metal2 31976 38752 31976 38752 0 recv_buf_valid
rlabel metal2 8792 35224 8792 35224 0 recv_divcnt\[0\]
rlabel metal2 5320 12600 5320 12600 0 recv_divcnt\[10\]
rlabel metal2 7168 11368 7168 11368 0 recv_divcnt\[11\]
rlabel metal2 10080 11144 10080 11144 0 recv_divcnt\[12\]
rlabel metal2 16408 11256 16408 11256 0 recv_divcnt\[13\]
rlabel metal2 15736 10640 15736 10640 0 recv_divcnt\[14\]
rlabel metal2 17864 9800 17864 9800 0 recv_divcnt\[15\]
rlabel metal3 23800 14280 23800 14280 0 recv_divcnt\[16\]
rlabel metal2 22792 12488 22792 12488 0 recv_divcnt\[17\]
rlabel metal2 23632 10696 23632 10696 0 recv_divcnt\[18\]
rlabel metal2 28504 12432 28504 12432 0 recv_divcnt\[19\]
rlabel metal2 11088 34888 11088 34888 0 recv_divcnt\[1\]
rlabel metal2 31864 9576 31864 9576 0 recv_divcnt\[20\]
rlabel metal3 33488 12152 33488 12152 0 recv_divcnt\[21\]
rlabel metal3 37576 8904 37576 8904 0 recv_divcnt\[22\]
rlabel metal2 39256 9968 39256 9968 0 recv_divcnt\[23\]
rlabel metal2 37688 18088 37688 18088 0 recv_divcnt\[24\]
rlabel metal2 43064 18424 43064 18424 0 recv_divcnt\[25\]
rlabel metal2 44968 16856 44968 16856 0 recv_divcnt\[26\]
rlabel metal3 45360 15176 45360 15176 0 recv_divcnt\[27\]
rlabel metal2 44240 27272 44240 27272 0 recv_divcnt\[28\]
rlabel metal3 46760 28616 46760 28616 0 recv_divcnt\[29\]
rlabel metal2 8232 32760 8232 32760 0 recv_divcnt\[2\]
rlabel metal3 41944 24920 41944 24920 0 recv_divcnt\[30\]
rlabel metal2 43736 23352 43736 23352 0 recv_divcnt\[31\]
rlabel metal2 12712 30352 12712 30352 0 recv_divcnt\[3\]
rlabel metal3 16856 26936 16856 26936 0 recv_divcnt\[4\]
rlabel via2 18536 28056 18536 28056 0 recv_divcnt\[5\]
rlabel metal2 18592 24920 18592 24920 0 recv_divcnt\[6\]
rlabel metal3 16352 23016 16352 23016 0 recv_divcnt\[7\]
rlabel metal2 6216 15568 6216 15568 0 recv_divcnt\[8\]
rlabel metal3 5320 14392 5320 14392 0 recv_divcnt\[9\]
rlabel metal2 46200 32816 46200 32816 0 recv_pattern\[0\]
rlabel metal2 45752 33768 45752 33768 0 recv_pattern\[1\]
rlabel metal3 44184 33320 44184 33320 0 recv_pattern\[2\]
rlabel metal2 42056 32368 42056 32368 0 recv_pattern\[3\]
rlabel metal2 40600 34552 40600 34552 0 recv_pattern\[4\]
rlabel metal2 40040 36848 40040 36848 0 recv_pattern\[5\]
rlabel metal3 36568 38136 36568 38136 0 recv_pattern\[6\]
rlabel metal2 36344 35728 36344 35728 0 recv_pattern\[7\]
rlabel metal2 31080 30128 31080 30128 0 recv_state\[0\]
rlabel metal3 32872 34104 32872 34104 0 recv_state\[1\]
rlabel metal2 32816 34888 32816 34888 0 recv_state\[2\]
rlabel metal3 34104 33320 34104 33320 0 recv_state\[3\]
rlabel metal2 28616 46312 28616 46312 0 reg_dat_di[0]
rlabel metal2 28504 45696 28504 45696 0 reg_dat_di[1]
rlabel metal2 23800 46144 23800 46144 0 reg_dat_di[2]
rlabel metal2 22960 45864 22960 45864 0 reg_dat_di[3]
rlabel metal2 21000 45584 21000 45584 0 reg_dat_di[4]
rlabel metal2 16856 47250 16856 47250 0 reg_dat_di[5]
rlabel metal2 16072 46312 16072 46312 0 reg_dat_di[6]
rlabel metal2 20104 46200 20104 46200 0 reg_dat_di[7]
rlabel metal3 48146 34328 48146 34328 0 reg_dat_do[0]
rlabel metal3 47026 49784 47026 49784 0 reg_dat_do[10]
rlabel metal2 47768 36400 47768 36400 0 reg_dat_do[11]
rlabel metal2 45192 46928 45192 46928 0 reg_dat_do[12]
rlabel metal2 45080 47082 45080 47082 0 reg_dat_do[13]
rlabel metal2 40376 47698 40376 47698 0 reg_dat_do[14]
rlabel metal3 46914 48440 46914 48440 0 reg_dat_do[15]
rlabel metal2 40152 43176 40152 43176 0 reg_dat_do[16]
rlabel metal3 46634 44408 46634 44408 0 reg_dat_do[17]
rlabel metal2 42392 47138 42392 47138 0 reg_dat_do[18]
rlabel metal3 45640 45192 45640 45192 0 reg_dat_do[19]
rlabel metal3 48482 38360 48482 38360 0 reg_dat_do[1]
rlabel metal2 44408 47250 44408 47250 0 reg_dat_do[20]
rlabel metal2 44072 41888 44072 41888 0 reg_dat_do[21]
rlabel metal2 47992 35784 47992 35784 0 reg_dat_do[22]
rlabel metal2 47432 37128 47432 37128 0 reg_dat_do[23]
rlabel metal3 46522 45752 46522 45752 0 reg_dat_do[24]
rlabel metal3 46578 43736 46578 43736 0 reg_dat_do[25]
rlabel metal2 41048 47306 41048 47306 0 reg_dat_do[26]
rlabel metal2 41720 47698 41720 47698 0 reg_dat_do[27]
rlabel metal2 43064 46914 43064 46914 0 reg_dat_do[28]
rlabel metal3 46690 47768 46690 47768 0 reg_dat_do[29]
rlabel metal2 47880 41888 47880 41888 0 reg_dat_do[2]
rlabel metal2 45752 46970 45752 46970 0 reg_dat_do[30]
rlabel metal3 48538 37688 48538 37688 0 reg_dat_do[31]
rlabel metal2 45080 39592 45080 39592 0 reg_dat_do[3]
rlabel metal2 47992 41272 47992 41272 0 reg_dat_do[4]
rlabel metal2 44968 42560 44968 42560 0 reg_dat_do[5]
rlabel metal3 47978 37016 47978 37016 0 reg_dat_do[6]
rlabel metal2 35000 47698 35000 47698 0 reg_dat_do[7]
rlabel metal2 43848 45640 43848 45640 0 reg_dat_do[8]
rlabel metal2 45080 41440 45080 41440 0 reg_dat_do[9]
rlabel metal2 33096 45192 33096 45192 0 reg_dat_re
rlabel metal2 23576 47698 23576 47698 0 reg_dat_wait
rlabel metal2 24584 45360 24584 45360 0 reg_dat_we
rlabel metal2 12376 45920 12376 45920 0 reg_div_di[0]
rlabel metal2 7392 3416 7392 3416 0 reg_div_di[10]
rlabel metal3 1246 8120 1246 8120 0 reg_div_di[11]
rlabel metal2 7840 3192 7840 3192 0 reg_div_di[12]
rlabel metal3 7672 3528 7672 3528 0 reg_div_di[13]
rlabel metal2 9352 3864 9352 3864 0 reg_div_di[14]
rlabel metal2 13608 4872 13608 4872 0 reg_div_di[15]
rlabel metal2 18872 4144 18872 4144 0 reg_div_di[16]
rlabel metal3 19264 3528 19264 3528 0 reg_div_di[17]
rlabel metal2 23744 2744 23744 2744 0 reg_div_di[18]
rlabel metal2 26264 2058 26264 2058 0 reg_div_di[19]
rlabel metal2 13496 47642 13496 47642 0 reg_div_di[1]
rlabel metal2 31696 3528 31696 3528 0 reg_div_di[20]
rlabel metal3 31696 4312 31696 4312 0 reg_div_di[21]
rlabel metal3 36736 3528 36736 3528 0 reg_div_di[22]
rlabel metal3 36568 4312 36568 4312 0 reg_div_di[23]
rlabel metal2 42952 3472 42952 3472 0 reg_div_di[24]
rlabel metal2 48216 8904 48216 8904 0 reg_div_di[25]
rlabel metal2 48216 10752 48216 10752 0 reg_div_di[26]
rlabel metal3 48762 17528 48762 17528 0 reg_div_di[27]
rlabel metal2 48104 19824 48104 19824 0 reg_div_di[28]
rlabel metal2 47544 24528 47544 24528 0 reg_div_di[29]
rlabel metal2 10584 46312 10584 46312 0 reg_div_di[2]
rlabel metal2 48216 25144 48216 25144 0 reg_div_di[30]
rlabel metal2 48216 12936 48216 12936 0 reg_div_di[31]
rlabel metal2 9576 45864 9576 45864 0 reg_div_di[3]
rlabel metal2 11704 46312 11704 46312 0 reg_div_di[4]
rlabel metal2 15568 45864 15568 45864 0 reg_div_di[5]
rlabel metal2 14840 47586 14840 47586 0 reg_div_di[6]
rlabel metal2 1736 34272 1736 34272 0 reg_div_di[7]
rlabel metal2 1736 23016 1736 23016 0 reg_div_di[8]
rlabel metal2 1736 21504 1736 21504 0 reg_div_di[9]
rlabel metal3 1358 37016 1358 37016 0 reg_div_do[0]
rlabel metal2 1960 18032 1960 18032 0 reg_div_do[10]
rlabel metal2 1960 16912 1960 16912 0 reg_div_do[11]
rlabel metal2 10808 1806 10808 1806 0 reg_div_do[12]
rlabel metal2 12152 854 12152 854 0 reg_div_do[13]
rlabel metal2 14840 2086 14840 2086 0 reg_div_do[14]
rlabel metal3 17024 3416 17024 3416 0 reg_div_do[15]
rlabel metal3 20384 3640 20384 3640 0 reg_div_do[16]
rlabel metal2 24248 1582 24248 1582 0 reg_div_do[17]
rlabel metal2 25592 2198 25592 2198 0 reg_div_do[18]
rlabel metal3 28504 3640 28504 3640 0 reg_div_do[19]
rlabel metal3 1358 42392 1358 42392 0 reg_div_do[1]
rlabel metal3 31696 3416 31696 3416 0 reg_div_do[20]
rlabel metal3 33936 5208 33936 5208 0 reg_div_do[21]
rlabel metal3 35672 3640 35672 3640 0 reg_div_do[22]
rlabel metal2 37688 2058 37688 2058 0 reg_div_do[23]
rlabel metal2 47320 6328 47320 6328 0 reg_div_do[24]
rlabel metal2 47992 9688 47992 9688 0 reg_div_do[25]
rlabel metal3 48650 11480 48650 11480 0 reg_div_do[26]
rlabel metal2 47992 16408 47992 16408 0 reg_div_do[27]
rlabel metal2 47992 20776 47992 20776 0 reg_div_do[28]
rlabel metal2 47992 22736 47992 22736 0 reg_div_do[29]
rlabel metal3 1414 41720 1414 41720 0 reg_div_do[2]
rlabel metal3 48594 26264 48594 26264 0 reg_div_do[30]
rlabel metal2 47992 12432 47992 12432 0 reg_div_do[31]
rlabel metal3 1358 40376 1358 40376 0 reg_div_do[3]
rlabel metal3 1358 39704 1358 39704 0 reg_div_do[4]
rlabel metal2 16184 47698 16184 47698 0 reg_div_do[5]
rlabel metal3 1358 36344 1358 36344 0 reg_div_do[6]
rlabel metal3 1358 33656 1358 33656 0 reg_div_do[7]
rlabel metal3 1358 24248 1358 24248 0 reg_div_do[8]
rlabel metal3 1358 21560 1358 21560 0 reg_div_do[9]
rlabel metal2 21672 46144 21672 46144 0 reg_div_we[0]
rlabel metal2 10136 2058 10136 2058 0 reg_div_we[1]
rlabel metal2 28504 5040 28504 5040 0 reg_div_we[2]
rlabel metal2 45640 18312 45640 18312 0 reg_div_we[3]
rlabel metal2 27496 46144 27496 46144 0 resetn
rlabel metal2 22904 35196 22904 35196 0 send_bitcnt\[0\]
rlabel metal2 22680 35672 22680 35672 0 send_bitcnt\[1\]
rlabel metal3 21896 35784 21896 35784 0 send_bitcnt\[2\]
rlabel metal2 24472 30968 24472 30968 0 send_bitcnt\[3\]
rlabel metal2 6440 37688 6440 37688 0 send_divcnt\[0\]
rlabel metal2 6216 18032 6216 18032 0 send_divcnt\[10\]
rlabel metal3 6104 19208 6104 19208 0 send_divcnt\[11\]
rlabel metal3 6720 22232 6720 22232 0 send_divcnt\[12\]
rlabel metal2 14728 19600 14728 19600 0 send_divcnt\[13\]
rlabel metal2 16688 19880 16688 19880 0 send_divcnt\[14\]
rlabel metal2 17752 19992 17752 19992 0 send_divcnt\[15\]
rlabel metal2 28056 17248 28056 17248 0 send_divcnt\[16\]
rlabel metal2 23352 22680 23352 22680 0 send_divcnt\[17\]
rlabel metal2 22904 18256 22904 18256 0 send_divcnt\[18\]
rlabel metal2 28168 19264 28168 19264 0 send_divcnt\[19\]
rlabel metal3 7168 40600 7168 40600 0 send_divcnt\[1\]
rlabel metal2 28112 22344 28112 22344 0 send_divcnt\[20\]
rlabel metal2 28952 15232 28952 15232 0 send_divcnt\[21\]
rlabel metal2 31472 20552 31472 20552 0 send_divcnt\[22\]
rlabel metal2 33880 17640 33880 17640 0 send_divcnt\[23\]
rlabel metal2 28616 25368 28616 25368 0 send_divcnt\[24\]
rlabel metal2 37800 22960 37800 22960 0 send_divcnt\[25\]
rlabel metal2 35336 22400 35336 22400 0 send_divcnt\[26\]
rlabel metal2 31752 22680 31752 22680 0 send_divcnt\[27\]
rlabel metal3 37744 25480 37744 25480 0 send_divcnt\[28\]
rlabel metal3 36232 26824 36232 26824 0 send_divcnt\[29\]
rlabel metal2 5208 37688 5208 37688 0 send_divcnt\[2\]
rlabel metal3 32760 27720 32760 27720 0 send_divcnt\[30\]
rlabel metal2 28952 27776 28952 27776 0 send_divcnt\[31\]
rlabel metal2 5712 36456 5712 36456 0 send_divcnt\[3\]
rlabel metal2 5656 29400 5656 29400 0 send_divcnt\[4\]
rlabel metal3 4984 28616 4984 28616 0 send_divcnt\[5\]
rlabel metal2 5376 28616 5376 28616 0 send_divcnt\[6\]
rlabel metal2 6328 24976 6328 24976 0 send_divcnt\[7\]
rlabel metal2 6888 24248 6888 24248 0 send_divcnt\[8\]
rlabel metal2 6440 24024 6440 24024 0 send_divcnt\[9\]
rlabel metal2 21448 32368 21448 32368 0 send_dummy
rlabel metal2 26376 40096 26376 40096 0 send_pattern\[1\]
rlabel metal2 27608 42392 27608 42392 0 send_pattern\[2\]
rlabel metal2 26824 44296 26824 44296 0 send_pattern\[3\]
rlabel metal3 23800 44184 23800 44184 0 send_pattern\[4\]
rlabel metal2 21448 44464 21448 44464 0 send_pattern\[5\]
rlabel metal2 19544 44352 19544 44352 0 send_pattern\[6\]
rlabel via2 19656 41944 19656 41944 0 send_pattern\[7\]
rlabel metal2 22288 40264 22288 40264 0 send_pattern\[8\]
rlabel metal2 34104 45640 34104 45640 0 uart_in[1]
rlabel metal2 28952 47698 28952 47698 0 uart_out[0]
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ctrl
  CLASS BLOCK ;
  FOREIGN ctrl ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN ctrl_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END ctrl_in[0]
  PIN ctrl_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 117.600 250.000 118.160 ;
    END
  END ctrl_in[1]
  PIN ctrl_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END ctrl_oeb[0]
  PIN ctrl_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 127.680 250.000 128.240 ;
    END
  END ctrl_oeb[1]
  PIN ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 4.000 ;
    END
  END ctrl_out[0]
  PIN ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 0.000 121.520 4.000 ;
    END
  END ctrl_out[1]
  PIN reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 120.960 250.000 121.520 ;
    END
  END reset
  PIN resetn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 124.320 250.000 124.880 ;
    END
  END resetn
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 231.580 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 231.580 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 243.040 231.580 ;
      LAYER Metal2 ;
        RECT 22.380 4.300 241.220 231.470 ;
        RECT 22.380 4.000 120.660 4.300 ;
        RECT 121.820 4.000 124.020 4.300 ;
        RECT 125.180 4.000 127.380 4.300 ;
        RECT 128.540 4.000 241.220 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 128.540 246.000 231.420 ;
        RECT 4.000 127.380 245.700 128.540 ;
        RECT 4.000 125.180 246.000 127.380 ;
        RECT 4.300 124.020 245.700 125.180 ;
        RECT 4.000 121.820 246.000 124.020 ;
        RECT 4.000 120.660 245.700 121.820 ;
        RECT 4.000 118.460 246.000 120.660 ;
        RECT 4.000 117.300 245.700 118.460 ;
        RECT 4.000 15.540 246.000 117.300 ;
  END
END ctrl
END LIBRARY


magic
tech gf180mcuD
magscale 1 10
timestamp 1702206060
<< metal1 >>
rect 19170 56590 19182 56642
rect 19234 56639 19246 56642
rect 20066 56639 20078 56642
rect 19234 56593 20078 56639
rect 19234 56590 19246 56593
rect 20066 56590 20078 56593
rect 20130 56590 20142 56642
rect 23986 56590 23998 56642
rect 24050 56639 24062 56642
rect 24994 56639 25006 56642
rect 24050 56593 25006 56639
rect 24050 56590 24062 56593
rect 24994 56590 25006 56593
rect 25058 56590 25070 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 19182 56306 19234 56318
rect 19182 56242 19234 56254
rect 33182 56306 33234 56318
rect 33182 56242 33234 56254
rect 46622 56082 46674 56094
rect 50430 56082 50482 56094
rect 20178 56030 20190 56082
rect 20242 56030 20254 56082
rect 23986 56030 23998 56082
rect 24050 56030 24062 56082
rect 27346 56030 27358 56082
rect 27410 56030 27422 56082
rect 29474 56030 29486 56082
rect 29538 56030 29550 56082
rect 32386 56030 32398 56082
rect 32450 56030 32462 56082
rect 35970 56030 35982 56082
rect 36034 56030 36046 56082
rect 42802 56030 42814 56082
rect 42866 56030 42878 56082
rect 46162 56030 46174 56082
rect 46226 56030 46238 56082
rect 49522 56030 49534 56082
rect 49586 56030 49598 56082
rect 46622 56018 46674 56030
rect 50430 56018 50482 56030
rect 24670 55970 24722 55982
rect 35310 55970 35362 55982
rect 40014 55970 40066 55982
rect 47630 55970 47682 55982
rect 30930 55918 30942 55970
rect 30994 55918 31006 55970
rect 36754 55918 36766 55970
rect 36818 55918 36830 55970
rect 38994 55918 39006 55970
rect 39058 55918 39070 55970
rect 42130 55918 42142 55970
rect 42194 55918 42206 55970
rect 24670 55906 24722 55918
rect 35310 55906 35362 55918
rect 40014 55906 40066 55918
rect 47630 55906 47682 55918
rect 22990 55858 23042 55870
rect 22990 55794 23042 55806
rect 24558 55858 24610 55870
rect 24558 55794 24610 55806
rect 26798 55858 26850 55870
rect 26798 55794 26850 55806
rect 43822 55858 43874 55870
rect 43822 55794 43874 55806
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 35758 55522 35810 55534
rect 35758 55458 35810 55470
rect 37102 55410 37154 55422
rect 14578 55358 14590 55410
rect 14642 55358 14654 55410
rect 20738 55358 20750 55410
rect 20802 55358 20814 55410
rect 24210 55358 24222 55410
rect 24274 55358 24286 55410
rect 26338 55358 26350 55410
rect 26402 55358 26414 55410
rect 33730 55358 33742 55410
rect 33794 55358 33806 55410
rect 40562 55358 40574 55410
rect 40626 55358 40638 55410
rect 42130 55358 42142 55410
rect 42194 55358 42206 55410
rect 45490 55358 45502 55410
rect 45554 55358 45566 55410
rect 51650 55358 51662 55410
rect 51714 55358 51726 55410
rect 37102 55346 37154 55358
rect 17490 55246 17502 55298
rect 17554 55246 17566 55298
rect 17938 55246 17950 55298
rect 18002 55246 18014 55298
rect 23538 55246 23550 55298
rect 23602 55246 23614 55298
rect 30930 55246 30942 55298
rect 30994 55246 31006 55298
rect 37650 55246 37662 55298
rect 37714 55246 37726 55298
rect 40898 55246 40910 55298
rect 40962 55246 40974 55298
rect 48402 55246 48414 55298
rect 48466 55246 48478 55298
rect 48738 55246 48750 55298
rect 48802 55246 48814 55298
rect 28478 55186 28530 55198
rect 35646 55186 35698 55198
rect 16706 55134 16718 55186
rect 16770 55134 16782 55186
rect 18610 55134 18622 55186
rect 18674 55134 18686 55186
rect 31602 55134 31614 55186
rect 31666 55134 31678 55186
rect 28478 55122 28530 55134
rect 35646 55122 35698 55134
rect 36318 55186 36370 55198
rect 43934 55186 43986 55198
rect 38434 55134 38446 55186
rect 38498 55134 38510 55186
rect 47618 55134 47630 55186
rect 47682 55134 47694 55186
rect 49522 55134 49534 55186
rect 49586 55134 49598 55186
rect 36318 55122 36370 55134
rect 43934 55122 43986 55134
rect 28366 55074 28418 55086
rect 28366 55010 28418 55022
rect 34190 55074 34242 55086
rect 34190 55010 34242 55022
rect 34638 55074 34690 55086
rect 34638 55010 34690 55022
rect 35086 55074 35138 55086
rect 35086 55010 35138 55022
rect 36206 55074 36258 55086
rect 36206 55010 36258 55022
rect 43822 55074 43874 55086
rect 43822 55010 43874 55022
rect 44942 55074 44994 55086
rect 44942 55010 44994 55022
rect 52110 55074 52162 55086
rect 52110 55010 52162 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 16718 54738 16770 54750
rect 16718 54674 16770 54686
rect 17726 54738 17778 54750
rect 17726 54674 17778 54686
rect 18510 54738 18562 54750
rect 18510 54674 18562 54686
rect 23662 54738 23714 54750
rect 31390 54738 31442 54750
rect 25666 54686 25678 54738
rect 25730 54686 25742 54738
rect 23662 54674 23714 54686
rect 31390 54674 31442 54686
rect 34190 54738 34242 54750
rect 34190 54674 34242 54686
rect 38334 54738 38386 54750
rect 38334 54674 38386 54686
rect 39006 54738 39058 54750
rect 39006 54674 39058 54686
rect 39790 54738 39842 54750
rect 39790 54674 39842 54686
rect 41246 54738 41298 54750
rect 41246 54674 41298 54686
rect 42030 54738 42082 54750
rect 42030 54674 42082 54686
rect 46286 54738 46338 54750
rect 46286 54674 46338 54686
rect 46398 54738 46450 54750
rect 46398 54674 46450 54686
rect 48078 54738 48130 54750
rect 48078 54674 48130 54686
rect 48862 54738 48914 54750
rect 48862 54674 48914 54686
rect 49422 54738 49474 54750
rect 49422 54674 49474 54686
rect 16830 54626 16882 54638
rect 33630 54626 33682 54638
rect 38222 54626 38274 54638
rect 25554 54574 25566 54626
rect 25618 54574 25630 54626
rect 27010 54574 27022 54626
rect 27074 54574 27086 54626
rect 28354 54574 28366 54626
rect 28418 54574 28430 54626
rect 32162 54574 32174 54626
rect 32226 54574 32238 54626
rect 35522 54574 35534 54626
rect 35586 54574 35598 54626
rect 16830 54562 16882 54574
rect 33630 54562 33682 54574
rect 38222 54562 38274 54574
rect 39118 54626 39170 54638
rect 39118 54562 39170 54574
rect 40126 54626 40178 54638
rect 40126 54562 40178 54574
rect 41918 54626 41970 54638
rect 43362 54574 43374 54626
rect 43426 54574 43438 54626
rect 41918 54562 41970 54574
rect 17502 54514 17554 54526
rect 17502 54450 17554 54462
rect 17614 54514 17666 54526
rect 17614 54450 17666 54462
rect 17838 54514 17890 54526
rect 26574 54514 26626 54526
rect 32510 54514 32562 54526
rect 18050 54462 18062 54514
rect 18114 54462 18126 54514
rect 18946 54462 18958 54514
rect 19010 54462 19022 54514
rect 24658 54462 24670 54514
rect 24722 54462 24734 54514
rect 25442 54462 25454 54514
rect 25506 54462 25518 54514
rect 27682 54462 27694 54514
rect 27746 54462 27758 54514
rect 17838 54450 17890 54462
rect 26574 54450 26626 54462
rect 32510 54450 32562 54462
rect 33182 54514 33234 54526
rect 33182 54450 33234 54462
rect 33294 54514 33346 54526
rect 38446 54514 38498 54526
rect 34738 54462 34750 54514
rect 34802 54462 34814 54514
rect 37986 54462 37998 54514
rect 38050 54462 38062 54514
rect 33294 54450 33346 54462
rect 38446 54450 38498 54462
rect 38558 54514 38610 54526
rect 38558 54450 38610 54462
rect 39566 54514 39618 54526
rect 39566 54450 39618 54462
rect 39678 54514 39730 54526
rect 39678 54450 39730 54462
rect 39902 54514 39954 54526
rect 41134 54514 41186 54526
rect 40898 54462 40910 54514
rect 40962 54462 40974 54514
rect 39902 54450 39954 54462
rect 41134 54450 41186 54462
rect 41358 54514 41410 54526
rect 46510 54514 46562 54526
rect 41570 54462 41582 54514
rect 41634 54462 41646 54514
rect 42578 54462 42590 54514
rect 42642 54462 42654 54514
rect 46050 54462 46062 54514
rect 46114 54462 46126 54514
rect 41358 54450 41410 54462
rect 46510 54450 46562 54462
rect 46622 54514 46674 54526
rect 47294 54514 47346 54526
rect 47058 54462 47070 54514
rect 47122 54462 47134 54514
rect 46622 54450 46674 54462
rect 47294 54450 47346 54462
rect 47518 54514 47570 54526
rect 53566 54514 53618 54526
rect 47730 54462 47742 54514
rect 47794 54462 47806 54514
rect 52994 54462 53006 54514
rect 53058 54462 53070 54514
rect 47518 54450 47570 54462
rect 53566 54450 53618 54462
rect 18398 54402 18450 54414
rect 30942 54402 30994 54414
rect 33518 54402 33570 54414
rect 19618 54350 19630 54402
rect 19682 54350 19694 54402
rect 21746 54350 21758 54402
rect 21810 54350 21822 54402
rect 30482 54350 30494 54402
rect 30546 54350 30558 54402
rect 31378 54350 31390 54402
rect 31442 54350 31454 54402
rect 18398 54338 18450 54350
rect 30942 54338 30994 54350
rect 33518 54338 33570 54350
rect 33966 54402 34018 54414
rect 45502 54402 45554 54414
rect 34178 54350 34190 54402
rect 34242 54350 34254 54402
rect 37650 54350 37662 54402
rect 37714 54350 37726 54402
rect 33966 54338 34018 54350
rect 45502 54338 45554 54350
rect 47406 54402 47458 54414
rect 47406 54338 47458 54350
rect 48190 54402 48242 54414
rect 48190 54338 48242 54350
rect 49310 54402 49362 54414
rect 49310 54338 49362 54350
rect 49870 54402 49922 54414
rect 50194 54350 50206 54402
rect 50258 54350 50270 54402
rect 52322 54350 52334 54402
rect 52386 54350 52398 54402
rect 49870 54338 49922 54350
rect 31614 54290 31666 54302
rect 31614 54226 31666 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 17390 53842 17442 53854
rect 27246 53842 27298 53854
rect 44942 53842 44994 53854
rect 48974 53842 49026 53854
rect 50766 53842 50818 53854
rect 16706 53790 16718 53842
rect 16770 53790 16782 53842
rect 19842 53790 19854 53842
rect 19906 53790 19918 53842
rect 26562 53790 26574 53842
rect 26626 53790 26638 53842
rect 27794 53790 27806 53842
rect 27858 53790 27870 53842
rect 29250 53790 29262 53842
rect 29314 53790 29326 53842
rect 31378 53790 31390 53842
rect 31442 53790 31454 53842
rect 33506 53790 33518 53842
rect 33570 53790 33582 53842
rect 37650 53790 37662 53842
rect 37714 53790 37726 53842
rect 41906 53790 41918 53842
rect 41970 53790 41982 53842
rect 44146 53790 44158 53842
rect 44210 53790 44222 53842
rect 45602 53790 45614 53842
rect 45666 53790 45678 53842
rect 49522 53790 49534 53842
rect 49586 53790 49598 53842
rect 17390 53778 17442 53790
rect 27246 53778 27298 53790
rect 44942 53778 44994 53790
rect 48974 53778 49026 53790
rect 50766 53778 50818 53790
rect 51438 53842 51490 53854
rect 51438 53778 51490 53790
rect 17614 53730 17666 53742
rect 13794 53678 13806 53730
rect 13858 53678 13870 53730
rect 17614 53666 17666 53678
rect 18846 53730 18898 53742
rect 18846 53666 18898 53678
rect 19294 53730 19346 53742
rect 29374 53730 29426 53742
rect 37774 53730 37826 53742
rect 43822 53730 43874 53742
rect 49646 53730 49698 53742
rect 51550 53730 51602 53742
rect 19730 53678 19742 53730
rect 19794 53678 19806 53730
rect 23202 53678 23214 53730
rect 23266 53678 23278 53730
rect 23762 53678 23774 53730
rect 23826 53678 23838 53730
rect 28354 53678 28366 53730
rect 28418 53678 28430 53730
rect 29138 53678 29150 53730
rect 29202 53678 29214 53730
rect 29810 53678 29822 53730
rect 29874 53678 29886 53730
rect 30706 53678 30718 53730
rect 30770 53678 30782 53730
rect 33842 53678 33854 53730
rect 33906 53678 33918 53730
rect 39106 53678 39118 53730
rect 39170 53678 39182 53730
rect 43138 53678 43150 53730
rect 43202 53678 43214 53730
rect 43586 53678 43598 53730
rect 43650 53678 43662 53730
rect 48402 53678 48414 53730
rect 48466 53678 48478 53730
rect 50418 53678 50430 53730
rect 50482 53678 50494 53730
rect 19294 53666 19346 53678
rect 29374 53666 29426 53678
rect 37774 53666 37826 53678
rect 43822 53666 43874 53678
rect 49646 53666 49698 53678
rect 51550 53666 51602 53678
rect 17054 53618 17106 53630
rect 18958 53618 19010 53630
rect 14578 53566 14590 53618
rect 14642 53566 14654 53618
rect 18386 53566 18398 53618
rect 18450 53566 18462 53618
rect 17054 53554 17106 53566
rect 18958 53554 19010 53566
rect 19182 53618 19234 53630
rect 19182 53554 19234 53566
rect 20190 53618 20242 53630
rect 20190 53554 20242 53566
rect 20414 53618 20466 53630
rect 27806 53618 27858 53630
rect 38222 53618 38274 53630
rect 44158 53618 44210 53630
rect 50094 53618 50146 53630
rect 22642 53566 22654 53618
rect 22706 53566 22718 53618
rect 24434 53566 24446 53618
rect 24498 53566 24510 53618
rect 35410 53566 35422 53618
rect 35474 53566 35486 53618
rect 39778 53566 39790 53618
rect 39842 53566 39854 53618
rect 42242 53566 42254 53618
rect 42306 53566 42318 53618
rect 42914 53566 42926 53618
rect 42978 53566 42990 53618
rect 47730 53566 47742 53618
rect 47794 53566 47806 53618
rect 20414 53554 20466 53566
rect 27806 53554 27858 53566
rect 38222 53554 38274 53566
rect 44158 53554 44210 53566
rect 50094 53554 50146 53566
rect 50878 53618 50930 53630
rect 50878 53554 50930 53566
rect 51102 53618 51154 53630
rect 51102 53554 51154 53566
rect 17278 53506 17330 53518
rect 17278 53442 17330 53454
rect 17502 53506 17554 53518
rect 17502 53442 17554 53454
rect 18062 53506 18114 53518
rect 18062 53442 18114 53454
rect 19070 53506 19122 53518
rect 19070 53442 19122 53454
rect 19966 53506 20018 53518
rect 19966 53442 20018 53454
rect 21646 53506 21698 53518
rect 21646 53442 21698 53454
rect 22094 53506 22146 53518
rect 22094 53442 22146 53454
rect 22318 53506 22370 53518
rect 27358 53506 27410 53518
rect 22978 53454 22990 53506
rect 23042 53454 23054 53506
rect 22318 53442 22370 53454
rect 27358 53442 27410 53454
rect 27918 53506 27970 53518
rect 27918 53442 27970 53454
rect 28142 53506 28194 53518
rect 28142 53442 28194 53454
rect 29598 53506 29650 53518
rect 29598 53442 29650 53454
rect 37214 53506 37266 53518
rect 37214 53442 37266 53454
rect 37662 53506 37714 53518
rect 37662 53442 37714 53454
rect 37998 53506 38050 53518
rect 37998 53442 38050 53454
rect 38670 53506 38722 53518
rect 38670 53442 38722 53454
rect 42590 53506 42642 53518
rect 42590 53442 42642 53454
rect 44046 53506 44098 53518
rect 44046 53442 44098 53454
rect 44830 53506 44882 53518
rect 44830 53442 44882 53454
rect 49534 53506 49586 53518
rect 49534 53442 49586 53454
rect 49870 53506 49922 53518
rect 49870 53442 49922 53454
rect 50654 53506 50706 53518
rect 50654 53442 50706 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 15486 53170 15538 53182
rect 15486 53106 15538 53118
rect 19630 53170 19682 53182
rect 19630 53106 19682 53118
rect 24110 53170 24162 53182
rect 24110 53106 24162 53118
rect 24334 53170 24386 53182
rect 24334 53106 24386 53118
rect 25342 53170 25394 53182
rect 25342 53106 25394 53118
rect 30158 53170 30210 53182
rect 30158 53106 30210 53118
rect 30718 53170 30770 53182
rect 30718 53106 30770 53118
rect 31614 53170 31666 53182
rect 31614 53106 31666 53118
rect 32510 53170 32562 53182
rect 32510 53106 32562 53118
rect 34078 53170 34130 53182
rect 34078 53106 34130 53118
rect 36990 53170 37042 53182
rect 36990 53106 37042 53118
rect 41022 53170 41074 53182
rect 41022 53106 41074 53118
rect 41470 53170 41522 53182
rect 46174 53170 46226 53182
rect 41906 53118 41918 53170
rect 41970 53118 41982 53170
rect 45602 53118 45614 53170
rect 45666 53118 45678 53170
rect 41470 53106 41522 53118
rect 46174 53106 46226 53118
rect 46286 53170 46338 53182
rect 46286 53106 46338 53118
rect 46510 53170 46562 53182
rect 47742 53170 47794 53182
rect 46946 53118 46958 53170
rect 47010 53118 47022 53170
rect 49074 53118 49086 53170
rect 49138 53118 49150 53170
rect 46510 53106 46562 53118
rect 47742 53106 47794 53118
rect 15598 53058 15650 53070
rect 17726 53058 17778 53070
rect 17378 53006 17390 53058
rect 17442 53006 17454 53058
rect 15598 52994 15650 53006
rect 17726 52994 17778 53006
rect 18174 53058 18226 53070
rect 18174 52994 18226 53006
rect 24446 53058 24498 53070
rect 24446 52994 24498 53006
rect 25678 53058 25730 53070
rect 25678 52994 25730 53006
rect 25902 53058 25954 53070
rect 31838 53058 31890 53070
rect 27570 53006 27582 53058
rect 27634 53006 27646 53058
rect 25902 52994 25954 53006
rect 31838 52994 31890 53006
rect 40238 53058 40290 53070
rect 47630 53058 47682 53070
rect 44146 53006 44158 53058
rect 44210 53006 44222 53058
rect 40238 52994 40290 53006
rect 47630 52994 47682 53006
rect 19742 52946 19794 52958
rect 24222 52946 24274 52958
rect 25454 52946 25506 52958
rect 31502 52946 31554 52958
rect 20738 52894 20750 52946
rect 20802 52894 20814 52946
rect 24658 52894 24670 52946
rect 24722 52894 24734 52946
rect 26898 52894 26910 52946
rect 26962 52894 26974 52946
rect 19742 52882 19794 52894
rect 24222 52882 24274 52894
rect 25454 52882 25506 52894
rect 31502 52882 31554 52894
rect 31950 52946 32002 52958
rect 39230 52946 39282 52958
rect 33506 52894 33518 52946
rect 33570 52894 33582 52946
rect 35970 52894 35982 52946
rect 36034 52894 36046 52946
rect 31950 52882 32002 52894
rect 39230 52882 39282 52894
rect 39566 52946 39618 52958
rect 39566 52882 39618 52894
rect 39790 52946 39842 52958
rect 46062 52946 46114 52958
rect 44930 52894 44942 52946
rect 44994 52894 45006 52946
rect 45378 52894 45390 52946
rect 45442 52894 45454 52946
rect 39790 52882 39842 52894
rect 46062 52882 46114 52894
rect 46398 52946 46450 52958
rect 48750 52946 48802 52958
rect 47170 52894 47182 52946
rect 47234 52894 47246 52946
rect 46398 52882 46450 52894
rect 48750 52882 48802 52894
rect 50878 52946 50930 52958
rect 50878 52882 50930 52894
rect 51326 52946 51378 52958
rect 51650 52894 51662 52946
rect 51714 52894 51726 52946
rect 52434 52894 52446 52946
rect 52498 52894 52510 52946
rect 51326 52882 51378 52894
rect 18622 52834 18674 52846
rect 30606 52834 30658 52846
rect 21410 52782 21422 52834
rect 21474 52782 21486 52834
rect 23538 52782 23550 52834
rect 23602 52782 23614 52834
rect 25330 52782 25342 52834
rect 25394 52782 25406 52834
rect 29698 52782 29710 52834
rect 29762 52782 29774 52834
rect 18622 52770 18674 52782
rect 30606 52770 30658 52782
rect 39342 52834 39394 52846
rect 48190 52834 48242 52846
rect 39890 52782 39902 52834
rect 39954 52831 39966 52834
rect 40114 52831 40126 52834
rect 39954 52785 40126 52831
rect 39954 52782 39966 52785
rect 40114 52782 40126 52785
rect 40178 52782 40190 52834
rect 39342 52770 39394 52782
rect 48190 52770 48242 52782
rect 49534 52834 49586 52846
rect 49534 52770 49586 52782
rect 50430 52834 50482 52846
rect 50430 52770 50482 52782
rect 51214 52834 51266 52846
rect 54562 52782 54574 52834
rect 54626 52782 54638 52834
rect 51214 52770 51266 52782
rect 30494 52722 30546 52734
rect 30494 52658 30546 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 18174 52386 18226 52398
rect 18174 52322 18226 52334
rect 18398 52386 18450 52398
rect 18398 52322 18450 52334
rect 24558 52386 24610 52398
rect 24558 52322 24610 52334
rect 26798 52386 26850 52398
rect 26798 52322 26850 52334
rect 31390 52386 31442 52398
rect 48738 52334 48750 52386
rect 48802 52383 48814 52386
rect 49522 52383 49534 52386
rect 48802 52337 49534 52383
rect 48802 52334 48814 52337
rect 49522 52334 49534 52337
rect 49586 52334 49598 52386
rect 31390 52322 31442 52334
rect 18958 52274 19010 52286
rect 16370 52222 16382 52274
rect 16434 52222 16446 52274
rect 18958 52210 19010 52222
rect 20638 52274 20690 52286
rect 20638 52210 20690 52222
rect 24222 52274 24274 52286
rect 24222 52210 24274 52222
rect 24670 52274 24722 52286
rect 24670 52210 24722 52222
rect 46622 52274 46674 52286
rect 46622 52210 46674 52222
rect 48750 52274 48802 52286
rect 51202 52222 51214 52274
rect 51266 52222 51278 52274
rect 48750 52210 48802 52222
rect 16830 52162 16882 52174
rect 13570 52110 13582 52162
rect 13634 52110 13646 52162
rect 16830 52098 16882 52110
rect 17838 52162 17890 52174
rect 17838 52098 17890 52110
rect 17950 52162 18002 52174
rect 20750 52162 20802 52174
rect 19170 52110 19182 52162
rect 19234 52110 19246 52162
rect 20402 52110 20414 52162
rect 20466 52110 20478 52162
rect 17950 52098 18002 52110
rect 20750 52098 20802 52110
rect 21982 52162 22034 52174
rect 21982 52098 22034 52110
rect 22094 52162 22146 52174
rect 22094 52098 22146 52110
rect 22430 52162 22482 52174
rect 29374 52162 29426 52174
rect 25218 52110 25230 52162
rect 25282 52110 25294 52162
rect 26226 52110 26238 52162
rect 26290 52110 26302 52162
rect 22430 52098 22482 52110
rect 29374 52098 29426 52110
rect 29598 52162 29650 52174
rect 29598 52098 29650 52110
rect 29822 52162 29874 52174
rect 37326 52162 37378 52174
rect 45166 52162 45218 52174
rect 30370 52110 30382 52162
rect 30434 52110 30446 52162
rect 33282 52110 33294 52162
rect 33346 52110 33358 52162
rect 39554 52110 39566 52162
rect 39618 52110 39630 52162
rect 40002 52110 40014 52162
rect 40066 52110 40078 52162
rect 29822 52098 29874 52110
rect 37326 52098 37378 52110
rect 45166 52098 45218 52110
rect 49310 52162 49362 52174
rect 50318 52162 50370 52174
rect 51326 52162 51378 52174
rect 49746 52110 49758 52162
rect 49810 52110 49822 52162
rect 50754 52110 50766 52162
rect 50818 52110 50830 52162
rect 49310 52098 49362 52110
rect 50318 52098 50370 52110
rect 51326 52098 51378 52110
rect 18846 52050 18898 52062
rect 14242 51998 14254 52050
rect 14306 51998 14318 52050
rect 18846 51986 18898 51998
rect 21870 52050 21922 52062
rect 21870 51986 21922 51998
rect 30046 52050 30098 52062
rect 38558 52050 38610 52062
rect 51214 52050 51266 52062
rect 34066 51998 34078 52050
rect 34130 51998 34142 52050
rect 37650 51998 37662 52050
rect 37714 51998 37726 52050
rect 41794 51998 41806 52050
rect 41858 51998 41870 52050
rect 30046 51986 30098 51998
rect 38558 51986 38610 51998
rect 51214 51986 51266 51998
rect 17838 51938 17890 51950
rect 40238 51938 40290 51950
rect 25442 51886 25454 51938
rect 25506 51886 25518 51938
rect 36306 51886 36318 51938
rect 36370 51886 36382 51938
rect 17838 51874 17890 51886
rect 40238 51874 40290 51886
rect 49982 51938 50034 51950
rect 49982 51874 50034 51886
rect 50094 51938 50146 51950
rect 50094 51874 50146 51886
rect 50206 51938 50258 51950
rect 50206 51874 50258 51886
rect 50990 51938 51042 51950
rect 50990 51874 51042 51886
rect 52782 51938 52834 51950
rect 52782 51874 52834 51886
rect 53230 51938 53282 51950
rect 53230 51874 53282 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 14478 51602 14530 51614
rect 14478 51538 14530 51550
rect 16046 51602 16098 51614
rect 16046 51538 16098 51550
rect 29150 51602 29202 51614
rect 34638 51602 34690 51614
rect 33058 51550 33070 51602
rect 33122 51550 33134 51602
rect 29150 51538 29202 51550
rect 34638 51538 34690 51550
rect 39006 51602 39058 51614
rect 44146 51550 44158 51602
rect 44210 51550 44222 51602
rect 39006 51538 39058 51550
rect 16494 51490 16546 51502
rect 33854 51490 33906 51502
rect 18386 51438 18398 51490
rect 18450 51438 18462 51490
rect 23650 51438 23662 51490
rect 23714 51438 23726 51490
rect 30370 51438 30382 51490
rect 30434 51438 30446 51490
rect 16494 51426 16546 51438
rect 33854 51426 33906 51438
rect 34974 51490 35026 51502
rect 34974 51426 35026 51438
rect 39118 51490 39170 51502
rect 39118 51426 39170 51438
rect 39454 51490 39506 51502
rect 39454 51426 39506 51438
rect 39790 51490 39842 51502
rect 46062 51490 46114 51502
rect 42466 51438 42478 51490
rect 42530 51438 42542 51490
rect 45378 51438 45390 51490
rect 45442 51438 45454 51490
rect 39790 51426 39842 51438
rect 46062 51426 46114 51438
rect 47182 51490 47234 51502
rect 47182 51426 47234 51438
rect 47854 51490 47906 51502
rect 47854 51426 47906 51438
rect 52446 51490 52498 51502
rect 52446 51426 52498 51438
rect 16270 51378 16322 51390
rect 21870 51378 21922 51390
rect 15810 51326 15822 51378
rect 15874 51326 15886 51378
rect 17602 51326 17614 51378
rect 17666 51326 17678 51378
rect 16270 51314 16322 51326
rect 21870 51314 21922 51326
rect 22206 51378 22258 51390
rect 22206 51314 22258 51326
rect 22542 51378 22594 51390
rect 33966 51378 34018 51390
rect 34526 51378 34578 51390
rect 23426 51326 23438 51378
rect 23490 51326 23502 51378
rect 25666 51326 25678 51378
rect 25730 51326 25742 51378
rect 29698 51326 29710 51378
rect 29762 51326 29774 51378
rect 33282 51326 33294 51378
rect 33346 51326 33358 51378
rect 34290 51326 34302 51378
rect 34354 51326 34366 51378
rect 22542 51314 22594 51326
rect 33966 51314 34018 51326
rect 34526 51314 34578 51326
rect 34750 51378 34802 51390
rect 40014 51378 40066 51390
rect 43822 51378 43874 51390
rect 35410 51326 35422 51378
rect 35474 51326 35486 51378
rect 38770 51326 38782 51378
rect 38834 51326 38846 51378
rect 40898 51326 40910 51378
rect 40962 51326 40974 51378
rect 34750 51314 34802 51326
rect 40014 51314 40066 51326
rect 43822 51314 43874 51326
rect 45054 51378 45106 51390
rect 45054 51314 45106 51326
rect 46622 51378 46674 51390
rect 46622 51314 46674 51326
rect 46958 51378 47010 51390
rect 52670 51378 52722 51390
rect 51986 51326 51998 51378
rect 52050 51326 52062 51378
rect 46958 51314 47010 51326
rect 52670 51314 52722 51326
rect 53118 51378 53170 51390
rect 53118 51314 53170 51326
rect 53342 51378 53394 51390
rect 53342 51314 53394 51326
rect 53566 51378 53618 51390
rect 53566 51314 53618 51326
rect 53902 51378 53954 51390
rect 53902 51314 53954 51326
rect 14590 51266 14642 51278
rect 14590 51202 14642 51214
rect 16158 51266 16210 51278
rect 22094 51266 22146 51278
rect 20514 51214 20526 51266
rect 20578 51214 20590 51266
rect 16158 51202 16210 51214
rect 22094 51202 22146 51214
rect 22990 51266 23042 51278
rect 39566 51266 39618 51278
rect 46734 51266 46786 51278
rect 26338 51214 26350 51266
rect 26402 51214 26414 51266
rect 28578 51214 28590 51266
rect 28642 51214 28654 51266
rect 32498 51214 32510 51266
rect 32562 51214 32574 51266
rect 36082 51214 36094 51266
rect 36146 51214 36158 51266
rect 38322 51214 38334 51266
rect 38386 51214 38398 51266
rect 46050 51214 46062 51266
rect 46114 51214 46126 51266
rect 22990 51202 23042 51214
rect 39566 51202 39618 51214
rect 46734 51202 46786 51214
rect 47966 51266 48018 51278
rect 47966 51202 48018 51214
rect 49198 51266 49250 51278
rect 52894 51266 52946 51278
rect 51314 51214 51326 51266
rect 51378 51214 51390 51266
rect 49198 51202 49250 51214
rect 52894 51202 52946 51214
rect 53790 51266 53842 51278
rect 53790 51202 53842 51214
rect 46286 51154 46338 51166
rect 46286 51090 46338 51102
rect 48078 51154 48130 51166
rect 48078 51090 48130 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 41134 50818 41186 50830
rect 41134 50754 41186 50766
rect 51886 50818 51938 50830
rect 51886 50754 51938 50766
rect 1934 50706 1986 50718
rect 1934 50642 1986 50654
rect 13694 50706 13746 50718
rect 18622 50706 18674 50718
rect 51998 50706 52050 50718
rect 15810 50654 15822 50706
rect 15874 50654 15886 50706
rect 17042 50654 17054 50706
rect 17106 50654 17118 50706
rect 24210 50654 24222 50706
rect 24274 50654 24286 50706
rect 27570 50654 27582 50706
rect 27634 50654 27646 50706
rect 32050 50654 32062 50706
rect 32114 50654 32126 50706
rect 50418 50654 50430 50706
rect 50482 50654 50494 50706
rect 55570 50654 55582 50706
rect 55634 50654 55646 50706
rect 13694 50642 13746 50654
rect 18622 50642 18674 50654
rect 51998 50642 52050 50654
rect 15374 50594 15426 50606
rect 3826 50542 3838 50594
rect 3890 50542 3902 50594
rect 15374 50530 15426 50542
rect 15710 50594 15762 50606
rect 15710 50530 15762 50542
rect 16158 50594 16210 50606
rect 17502 50594 17554 50606
rect 18734 50594 18786 50606
rect 17154 50542 17166 50594
rect 17218 50542 17230 50594
rect 17826 50542 17838 50594
rect 17890 50542 17902 50594
rect 16158 50530 16210 50542
rect 17502 50530 17554 50542
rect 18734 50530 18786 50542
rect 19070 50594 19122 50606
rect 39118 50594 39170 50606
rect 21410 50542 21422 50594
rect 21474 50542 21486 50594
rect 24546 50542 24558 50594
rect 24610 50542 24622 50594
rect 29138 50542 29150 50594
rect 29202 50542 29214 50594
rect 32610 50542 32622 50594
rect 32674 50542 32686 50594
rect 36418 50542 36430 50594
rect 36482 50542 36494 50594
rect 36978 50542 36990 50594
rect 37042 50542 37054 50594
rect 19070 50530 19122 50542
rect 39118 50530 39170 50542
rect 41918 50594 41970 50606
rect 46386 50542 46398 50594
rect 46450 50542 46462 50594
rect 46834 50542 46846 50594
rect 46898 50542 46910 50594
rect 49522 50542 49534 50594
rect 49586 50542 49598 50594
rect 52658 50542 52670 50594
rect 52722 50542 52734 50594
rect 41918 50530 41970 50542
rect 13582 50482 13634 50494
rect 13582 50418 13634 50430
rect 14926 50482 14978 50494
rect 14926 50418 14978 50430
rect 15822 50482 15874 50494
rect 18510 50482 18562 50494
rect 28366 50482 28418 50494
rect 18050 50430 18062 50482
rect 18114 50430 18126 50482
rect 19730 50430 19742 50482
rect 19794 50430 19806 50482
rect 22082 50430 22094 50482
rect 22146 50430 22158 50482
rect 25330 50430 25342 50482
rect 25394 50430 25406 50482
rect 15822 50418 15874 50430
rect 18510 50418 18562 50430
rect 28366 50418 28418 50430
rect 28478 50482 28530 50494
rect 28478 50418 28530 50430
rect 28590 50482 28642 50494
rect 35310 50482 35362 50494
rect 41246 50482 41298 50494
rect 29922 50430 29934 50482
rect 29986 50430 29998 50482
rect 32722 50430 32734 50482
rect 32786 50430 32798 50482
rect 37090 50430 37102 50482
rect 37154 50430 37166 50482
rect 40786 50430 40798 50482
rect 40850 50430 40862 50482
rect 28590 50418 28642 50430
rect 35310 50418 35362 50430
rect 41246 50418 41298 50430
rect 41358 50482 41410 50494
rect 41358 50418 41410 50430
rect 42254 50482 42306 50494
rect 42254 50418 42306 50430
rect 42590 50482 42642 50494
rect 42590 50418 42642 50430
rect 43038 50482 43090 50494
rect 47406 50482 47458 50494
rect 44930 50430 44942 50482
rect 44994 50430 45006 50482
rect 53442 50430 53454 50482
rect 53506 50430 53518 50482
rect 43038 50418 43090 50430
rect 47406 50418 47458 50430
rect 16046 50370 16098 50382
rect 16046 50306 16098 50318
rect 16942 50370 16994 50382
rect 16942 50306 16994 50318
rect 19406 50370 19458 50382
rect 34850 50318 34862 50370
rect 34914 50318 34926 50370
rect 39778 50318 39790 50370
rect 39842 50318 39854 50370
rect 45042 50318 45054 50370
rect 45106 50318 45118 50370
rect 19406 50306 19458 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 18398 50034 18450 50046
rect 18398 49970 18450 49982
rect 20638 50034 20690 50046
rect 20638 49970 20690 49982
rect 21758 50034 21810 50046
rect 25342 50034 25394 50046
rect 23202 49982 23214 50034
rect 23266 49982 23278 50034
rect 21758 49970 21810 49982
rect 25342 49970 25394 49982
rect 26462 50034 26514 50046
rect 26462 49970 26514 49982
rect 27246 50034 27298 50046
rect 27246 49970 27298 49982
rect 27358 50034 27410 50046
rect 27358 49970 27410 49982
rect 30494 50034 30546 50046
rect 34750 50034 34802 50046
rect 34402 49982 34414 50034
rect 34466 49982 34478 50034
rect 30494 49970 30546 49982
rect 34750 49970 34802 49982
rect 35982 50034 36034 50046
rect 35982 49970 36034 49982
rect 36318 50034 36370 50046
rect 36318 49970 36370 49982
rect 36878 50034 36930 50046
rect 36878 49970 36930 49982
rect 48862 50034 48914 50046
rect 54014 50034 54066 50046
rect 50754 49982 50766 50034
rect 50818 49982 50830 50034
rect 48862 49970 48914 49982
rect 54014 49970 54066 49982
rect 54126 50034 54178 50046
rect 54126 49970 54178 49982
rect 54798 50034 54850 50046
rect 54798 49970 54850 49982
rect 2046 49922 2098 49934
rect 17390 49922 17442 49934
rect 12898 49870 12910 49922
rect 12962 49870 12974 49922
rect 15698 49870 15710 49922
rect 15762 49870 15774 49922
rect 16818 49870 16830 49922
rect 16882 49870 16894 49922
rect 2046 49858 2098 49870
rect 17390 49858 17442 49870
rect 21982 49922 22034 49934
rect 21982 49858 22034 49870
rect 24670 49922 24722 49934
rect 24670 49858 24722 49870
rect 26574 49922 26626 49934
rect 26574 49858 26626 49870
rect 27582 49922 27634 49934
rect 27582 49858 27634 49870
rect 29486 49922 29538 49934
rect 48750 49922 48802 49934
rect 30146 49870 30158 49922
rect 30210 49870 30222 49922
rect 32498 49870 32510 49922
rect 32562 49870 32574 49922
rect 38210 49870 38222 49922
rect 38274 49870 38286 49922
rect 46050 49870 46062 49922
rect 46114 49870 46126 49922
rect 29486 49858 29538 49870
rect 48750 49858 48802 49870
rect 49086 49922 49138 49934
rect 52334 49922 52386 49934
rect 49746 49870 49758 49922
rect 49810 49870 49822 49922
rect 49086 49858 49138 49870
rect 52334 49858 52386 49870
rect 53902 49922 53954 49934
rect 53902 49858 53954 49870
rect 54574 49922 54626 49934
rect 54574 49858 54626 49870
rect 1710 49810 1762 49822
rect 15374 49810 15426 49822
rect 12226 49758 12238 49810
rect 12290 49758 12302 49810
rect 1710 49746 1762 49758
rect 15374 49746 15426 49758
rect 16494 49810 16546 49822
rect 16494 49746 16546 49758
rect 17502 49810 17554 49822
rect 19518 49810 19570 49822
rect 17938 49758 17950 49810
rect 18002 49758 18014 49810
rect 17502 49746 17554 49758
rect 19518 49746 19570 49758
rect 19742 49810 19794 49822
rect 19742 49746 19794 49758
rect 20078 49810 20130 49822
rect 25790 49810 25842 49822
rect 26350 49810 26402 49822
rect 27694 49810 27746 49822
rect 23426 49758 23438 49810
rect 23490 49758 23502 49810
rect 26114 49758 26126 49810
rect 26178 49758 26190 49810
rect 26786 49758 26798 49810
rect 26850 49758 26862 49810
rect 20078 49746 20130 49758
rect 25790 49746 25842 49758
rect 26350 49746 26402 49758
rect 27694 49746 27746 49758
rect 28814 49810 28866 49822
rect 28814 49746 28866 49758
rect 29262 49810 29314 49822
rect 29262 49746 29314 49758
rect 32174 49810 32226 49822
rect 36094 49810 36146 49822
rect 44942 49810 44994 49822
rect 49198 49810 49250 49822
rect 33618 49758 33630 49810
rect 33682 49758 33694 49810
rect 36530 49758 36542 49810
rect 36594 49758 36606 49810
rect 37426 49758 37438 49810
rect 37490 49758 37502 49810
rect 41682 49758 41694 49810
rect 41746 49758 41758 49810
rect 45378 49758 45390 49810
rect 45442 49758 45454 49810
rect 32174 49746 32226 49758
rect 36094 49746 36146 49758
rect 44942 49746 44994 49758
rect 49198 49746 49250 49758
rect 51438 49810 51490 49822
rect 51438 49746 51490 49758
rect 51886 49810 51938 49822
rect 51886 49746 51938 49758
rect 2494 49698 2546 49710
rect 2494 49634 2546 49646
rect 11566 49698 11618 49710
rect 16158 49698 16210 49710
rect 15026 49646 15038 49698
rect 15090 49646 15102 49698
rect 11566 49634 11618 49646
rect 16158 49634 16210 49646
rect 19070 49698 19122 49710
rect 19070 49634 19122 49646
rect 19630 49698 19682 49710
rect 19630 49634 19682 49646
rect 20414 49698 20466 49710
rect 20414 49634 20466 49646
rect 20526 49698 20578 49710
rect 25230 49698 25282 49710
rect 21634 49646 21646 49698
rect 21698 49646 21710 49698
rect 20526 49634 20578 49646
rect 25230 49634 25282 49646
rect 25678 49698 25730 49710
rect 25678 49634 25730 49646
rect 27470 49698 27522 49710
rect 27470 49634 27522 49646
rect 28254 49698 28306 49710
rect 28254 49634 28306 49646
rect 29038 49698 29090 49710
rect 29038 49634 29090 49646
rect 31838 49698 31890 49710
rect 34078 49698 34130 49710
rect 33282 49646 33294 49698
rect 33346 49646 33358 49698
rect 31838 49634 31890 49646
rect 34078 49634 34130 49646
rect 35198 49698 35250 49710
rect 35198 49634 35250 49646
rect 36206 49698 36258 49710
rect 36206 49634 36258 49646
rect 36990 49698 37042 49710
rect 40338 49646 40350 49698
rect 40402 49646 40414 49698
rect 42354 49646 42366 49698
rect 42418 49646 42430 49698
rect 44482 49646 44494 49698
rect 44546 49646 44558 49698
rect 48178 49646 48190 49698
rect 48242 49646 48254 49698
rect 54786 49646 54798 49698
rect 54850 49646 54862 49698
rect 36990 49634 37042 49646
rect 11454 49586 11506 49598
rect 11454 49522 11506 49534
rect 17726 49586 17778 49598
rect 17726 49522 17778 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 42366 49250 42418 49262
rect 42366 49186 42418 49198
rect 27582 49138 27634 49150
rect 37214 49138 37266 49150
rect 10770 49086 10782 49138
rect 10834 49086 10846 49138
rect 12898 49086 12910 49138
rect 12962 49086 12974 49138
rect 27010 49086 27022 49138
rect 27074 49086 27086 49138
rect 33730 49086 33742 49138
rect 33794 49086 33806 49138
rect 27582 49074 27634 49086
rect 37214 49074 37266 49086
rect 37550 49138 37602 49150
rect 37550 49074 37602 49086
rect 42702 49138 42754 49150
rect 42702 49074 42754 49086
rect 43150 49138 43202 49150
rect 43150 49074 43202 49086
rect 47070 49138 47122 49150
rect 48066 49086 48078 49138
rect 48130 49086 48142 49138
rect 50194 49086 50206 49138
rect 50258 49086 50270 49138
rect 52658 49086 52670 49138
rect 52722 49086 52734 49138
rect 54786 49086 54798 49138
rect 54850 49086 54862 49138
rect 47070 49074 47122 49086
rect 14814 49026 14866 49038
rect 15822 49026 15874 49038
rect 10098 48974 10110 49026
rect 10162 48974 10174 49026
rect 14690 48974 14702 49026
rect 14754 48974 14766 49026
rect 15138 48974 15150 49026
rect 15202 48974 15214 49026
rect 14814 48962 14866 48974
rect 15822 48962 15874 48974
rect 17054 49026 17106 49038
rect 17054 48962 17106 48974
rect 17390 49026 17442 49038
rect 38110 49026 38162 49038
rect 43374 49026 43426 49038
rect 22754 48974 22766 49026
rect 22818 48974 22830 49026
rect 24098 48974 24110 49026
rect 24162 48974 24174 49026
rect 30706 48974 30718 49026
rect 30770 48974 30782 49026
rect 32946 48974 32958 49026
rect 33010 48974 33022 49026
rect 39778 48974 39790 49026
rect 39842 48974 39854 49026
rect 41458 48974 41470 49026
rect 41522 48974 41534 49026
rect 17390 48962 17442 48974
rect 38110 48962 38162 48974
rect 43374 48962 43426 48974
rect 44830 49026 44882 49038
rect 47282 48974 47294 49026
rect 47346 48974 47358 49026
rect 55458 48974 55470 49026
rect 55522 48974 55534 49026
rect 44830 48962 44882 48974
rect 1710 48914 1762 48926
rect 1710 48850 1762 48862
rect 16830 48914 16882 48926
rect 30942 48914 30994 48926
rect 43038 48914 43090 48926
rect 22530 48862 22542 48914
rect 22594 48862 22606 48914
rect 24882 48862 24894 48914
rect 24946 48862 24958 48914
rect 39890 48862 39902 48914
rect 39954 48862 39966 48914
rect 40562 48862 40574 48914
rect 40626 48862 40638 48914
rect 16830 48850 16882 48862
rect 30942 48850 30994 48862
rect 43038 48850 43090 48862
rect 43598 48914 43650 48926
rect 50866 48862 50878 48914
rect 50930 48862 50942 48914
rect 43598 48850 43650 48862
rect 2046 48802 2098 48814
rect 2046 48738 2098 48750
rect 2494 48802 2546 48814
rect 2494 48738 2546 48750
rect 13918 48802 13970 48814
rect 13918 48738 13970 48750
rect 17166 48802 17218 48814
rect 17166 48738 17218 48750
rect 29374 48802 29426 48814
rect 29374 48738 29426 48750
rect 30382 48802 30434 48814
rect 30382 48738 30434 48750
rect 31390 48802 31442 48814
rect 31390 48738 31442 48750
rect 35534 48802 35586 48814
rect 35534 48738 35586 48750
rect 36318 48802 36370 48814
rect 36318 48738 36370 48750
rect 42478 48802 42530 48814
rect 50542 48802 50594 48814
rect 45154 48750 45166 48802
rect 45218 48750 45230 48802
rect 42478 48738 42530 48750
rect 50542 48738 50594 48750
rect 51326 48802 51378 48814
rect 51326 48738 51378 48750
rect 51774 48802 51826 48814
rect 51774 48738 51826 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 12126 48466 12178 48478
rect 12126 48402 12178 48414
rect 12238 48466 12290 48478
rect 12238 48402 12290 48414
rect 13358 48466 13410 48478
rect 13358 48402 13410 48414
rect 25454 48466 25506 48478
rect 25454 48402 25506 48414
rect 30718 48466 30770 48478
rect 30718 48402 30770 48414
rect 36542 48466 36594 48478
rect 36542 48402 36594 48414
rect 38782 48466 38834 48478
rect 42814 48466 42866 48478
rect 41122 48414 41134 48466
rect 41186 48414 41198 48466
rect 38782 48402 38834 48414
rect 42814 48402 42866 48414
rect 45726 48466 45778 48478
rect 45726 48402 45778 48414
rect 51886 48466 51938 48478
rect 51886 48402 51938 48414
rect 2046 48354 2098 48366
rect 2046 48290 2098 48302
rect 17838 48354 17890 48366
rect 25790 48354 25842 48366
rect 20290 48302 20302 48354
rect 20354 48302 20366 48354
rect 17838 48290 17890 48302
rect 25790 48290 25842 48302
rect 31502 48354 31554 48366
rect 31502 48290 31554 48302
rect 42142 48354 42194 48366
rect 42142 48290 42194 48302
rect 43038 48354 43090 48366
rect 45838 48354 45890 48366
rect 43586 48302 43598 48354
rect 43650 48302 43662 48354
rect 43038 48290 43090 48302
rect 45838 48290 45890 48302
rect 46846 48354 46898 48366
rect 47730 48302 47742 48354
rect 47794 48302 47806 48354
rect 46846 48290 46898 48302
rect 1710 48242 1762 48254
rect 12014 48242 12066 48254
rect 25230 48242 25282 48254
rect 11778 48190 11790 48242
rect 11842 48190 11854 48242
rect 12450 48190 12462 48242
rect 12514 48190 12526 48242
rect 14018 48190 14030 48242
rect 14082 48190 14094 48242
rect 19506 48190 19518 48242
rect 19570 48190 19582 48242
rect 1710 48178 1762 48190
rect 12014 48178 12066 48190
rect 25230 48178 25282 48190
rect 25566 48242 25618 48254
rect 30382 48242 30434 48254
rect 30034 48190 30046 48242
rect 30098 48190 30110 48242
rect 25566 48178 25618 48190
rect 30382 48178 30434 48190
rect 30830 48242 30882 48254
rect 30830 48178 30882 48190
rect 30942 48242 30994 48254
rect 30942 48178 30994 48190
rect 31726 48242 31778 48254
rect 31726 48178 31778 48190
rect 31950 48242 32002 48254
rect 36878 48242 36930 48254
rect 33170 48190 33182 48242
rect 33234 48190 33246 48242
rect 31950 48178 32002 48190
rect 36878 48178 36930 48190
rect 37102 48242 37154 48254
rect 37102 48178 37154 48190
rect 37438 48242 37490 48254
rect 37438 48178 37490 48190
rect 37662 48242 37714 48254
rect 37662 48178 37714 48190
rect 37998 48242 38050 48254
rect 37998 48178 38050 48190
rect 38334 48242 38386 48254
rect 42590 48242 42642 48254
rect 41346 48190 41358 48242
rect 41410 48190 41422 48242
rect 41794 48190 41806 48242
rect 41858 48190 41870 48242
rect 38334 48178 38386 48190
rect 42590 48178 42642 48190
rect 42814 48242 42866 48254
rect 42814 48178 42866 48190
rect 43934 48242 43986 48254
rect 43934 48178 43986 48190
rect 45390 48242 45442 48254
rect 45390 48178 45442 48190
rect 46062 48242 46114 48254
rect 46062 48178 46114 48190
rect 46398 48242 46450 48254
rect 46398 48178 46450 48190
rect 47070 48242 47122 48254
rect 47070 48178 47122 48190
rect 47406 48242 47458 48254
rect 48738 48190 48750 48242
rect 48802 48190 48814 48242
rect 52658 48190 52670 48242
rect 52722 48190 52734 48242
rect 47406 48178 47458 48190
rect 2494 48130 2546 48142
rect 2494 48066 2546 48078
rect 12910 48130 12962 48142
rect 24670 48130 24722 48142
rect 36990 48130 37042 48142
rect 14690 48078 14702 48130
rect 14754 48078 14766 48130
rect 16818 48078 16830 48130
rect 16882 48078 16894 48130
rect 17826 48078 17838 48130
rect 17890 48078 17902 48130
rect 22418 48078 22430 48130
rect 22482 48078 22494 48130
rect 27234 48078 27246 48130
rect 27298 48078 27310 48130
rect 29362 48078 29374 48130
rect 29426 48078 29438 48130
rect 33954 48078 33966 48130
rect 34018 48078 34030 48130
rect 36082 48078 36094 48130
rect 36146 48078 36158 48130
rect 12910 48066 12962 48078
rect 24670 48066 24722 48078
rect 36990 48066 37042 48078
rect 37886 48130 37938 48142
rect 37886 48066 37938 48078
rect 40014 48130 40066 48142
rect 40014 48066 40066 48078
rect 40350 48130 40402 48142
rect 40350 48066 40402 48078
rect 42030 48130 42082 48142
rect 42030 48066 42082 48078
rect 46622 48130 46674 48142
rect 46622 48066 46674 48078
rect 48190 48130 48242 48142
rect 53118 48130 53170 48142
rect 49858 48078 49870 48130
rect 49922 48078 49934 48130
rect 48190 48066 48242 48078
rect 53118 48066 53170 48078
rect 17614 48018 17666 48030
rect 17614 47954 17666 47966
rect 32174 48018 32226 48030
rect 32174 47954 32226 47966
rect 32622 48018 32674 48030
rect 32622 47954 32674 47966
rect 51662 48018 51714 48030
rect 51662 47954 51714 47966
rect 51998 48018 52050 48030
rect 51998 47954 52050 47966
rect 52334 48018 52386 48030
rect 52334 47954 52386 47966
rect 52670 48018 52722 48030
rect 52670 47954 52722 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 16382 47682 16434 47694
rect 16382 47618 16434 47630
rect 16718 47682 16770 47694
rect 16718 47618 16770 47630
rect 26798 47682 26850 47694
rect 26798 47618 26850 47630
rect 29262 47682 29314 47694
rect 29262 47618 29314 47630
rect 33294 47682 33346 47694
rect 33294 47618 33346 47630
rect 36430 47682 36482 47694
rect 36430 47618 36482 47630
rect 45838 47682 45890 47694
rect 45838 47618 45890 47630
rect 12910 47570 12962 47582
rect 26910 47570 26962 47582
rect 12450 47518 12462 47570
rect 12514 47518 12526 47570
rect 17826 47518 17838 47570
rect 17890 47518 17902 47570
rect 19954 47518 19966 47570
rect 20018 47518 20030 47570
rect 12910 47506 12962 47518
rect 26910 47506 26962 47518
rect 27806 47570 27858 47582
rect 40350 47570 40402 47582
rect 50206 47570 50258 47582
rect 30706 47518 30718 47570
rect 30770 47518 30782 47570
rect 32834 47518 32846 47570
rect 32898 47518 32910 47570
rect 39890 47518 39902 47570
rect 39954 47518 39966 47570
rect 42130 47518 42142 47570
rect 42194 47518 42206 47570
rect 44258 47518 44270 47570
rect 44322 47518 44334 47570
rect 46834 47518 46846 47570
rect 46898 47518 46910 47570
rect 27806 47506 27858 47518
rect 40350 47506 40402 47518
rect 50206 47506 50258 47518
rect 51102 47570 51154 47582
rect 51102 47506 51154 47518
rect 57934 47570 57986 47582
rect 57934 47506 57986 47518
rect 20302 47458 20354 47470
rect 9650 47406 9662 47458
rect 9714 47406 9726 47458
rect 17154 47406 17166 47458
rect 17218 47406 17230 47458
rect 20302 47394 20354 47406
rect 24334 47458 24386 47470
rect 28366 47458 28418 47470
rect 33182 47458 33234 47470
rect 24882 47406 24894 47458
rect 24946 47406 24958 47458
rect 30034 47406 30046 47458
rect 30098 47406 30110 47458
rect 24334 47394 24386 47406
rect 28366 47394 28418 47406
rect 33182 47394 33234 47406
rect 34078 47458 34130 47470
rect 40126 47458 40178 47470
rect 50990 47458 51042 47470
rect 35186 47406 35198 47458
rect 35250 47406 35262 47458
rect 36082 47406 36094 47458
rect 36146 47406 36158 47458
rect 36978 47406 36990 47458
rect 37042 47406 37054 47458
rect 41458 47406 41470 47458
rect 41522 47406 41534 47458
rect 48962 47406 48974 47458
rect 49026 47406 49038 47458
rect 49634 47406 49646 47458
rect 49698 47406 49710 47458
rect 34078 47394 34130 47406
rect 40126 47394 40178 47406
rect 50990 47394 51042 47406
rect 51214 47458 51266 47470
rect 51214 47394 51266 47406
rect 51438 47458 51490 47470
rect 51438 47394 51490 47406
rect 51886 47458 51938 47470
rect 55570 47406 55582 47458
rect 55634 47406 55646 47458
rect 51886 47394 51938 47406
rect 1710 47346 1762 47358
rect 16494 47346 16546 47358
rect 25342 47346 25394 47358
rect 10322 47294 10334 47346
rect 10386 47294 10398 47346
rect 21298 47294 21310 47346
rect 21362 47294 21374 47346
rect 22754 47294 22766 47346
rect 22818 47294 22830 47346
rect 1710 47282 1762 47294
rect 16494 47282 16546 47294
rect 25342 47282 25394 47294
rect 27022 47346 27074 47358
rect 27022 47282 27074 47294
rect 29150 47346 29202 47358
rect 29150 47282 29202 47294
rect 29262 47346 29314 47358
rect 36318 47346 36370 47358
rect 50654 47346 50706 47358
rect 34962 47294 34974 47346
rect 35026 47294 35038 47346
rect 37762 47294 37774 47346
rect 37826 47294 37838 47346
rect 29262 47282 29314 47294
rect 36318 47282 36370 47294
rect 50654 47282 50706 47294
rect 52110 47346 52162 47358
rect 52110 47282 52162 47294
rect 2046 47234 2098 47246
rect 2046 47170 2098 47182
rect 2494 47234 2546 47246
rect 21646 47234 21698 47246
rect 27694 47234 27746 47246
rect 20626 47182 20638 47234
rect 20690 47182 20702 47234
rect 26338 47182 26350 47234
rect 26402 47182 26414 47234
rect 2494 47170 2546 47182
rect 21646 47170 21698 47182
rect 27694 47170 27746 47182
rect 27918 47234 27970 47246
rect 27918 47170 27970 47182
rect 33294 47234 33346 47246
rect 33294 47170 33346 47182
rect 34190 47234 34242 47246
rect 34190 47170 34242 47182
rect 34302 47234 34354 47246
rect 34302 47170 34354 47182
rect 34526 47234 34578 47246
rect 34526 47170 34578 47182
rect 35758 47234 35810 47246
rect 35758 47170 35810 47182
rect 40462 47234 40514 47246
rect 40462 47170 40514 47182
rect 40686 47234 40738 47246
rect 40686 47170 40738 47182
rect 44942 47234 44994 47246
rect 44942 47170 44994 47182
rect 45950 47234 46002 47246
rect 45950 47170 46002 47182
rect 46062 47234 46114 47246
rect 46062 47170 46114 47182
rect 51774 47234 51826 47246
rect 51774 47170 51826 47182
rect 55246 47234 55298 47246
rect 55246 47170 55298 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 10894 46898 10946 46910
rect 10894 46834 10946 46846
rect 11902 46898 11954 46910
rect 11902 46834 11954 46846
rect 17614 46898 17666 46910
rect 17614 46834 17666 46846
rect 31838 46898 31890 46910
rect 31838 46834 31890 46846
rect 33742 46898 33794 46910
rect 36542 46898 36594 46910
rect 35522 46846 35534 46898
rect 35586 46846 35598 46898
rect 33742 46834 33794 46846
rect 36542 46834 36594 46846
rect 44270 46898 44322 46910
rect 49534 46898 49586 46910
rect 48738 46846 48750 46898
rect 48802 46846 48814 46898
rect 44270 46834 44322 46846
rect 49534 46834 49586 46846
rect 50206 46898 50258 46910
rect 50206 46834 50258 46846
rect 53902 46898 53954 46910
rect 53902 46834 53954 46846
rect 2046 46786 2098 46798
rect 2046 46722 2098 46734
rect 11006 46786 11058 46798
rect 11006 46722 11058 46734
rect 11790 46786 11842 46798
rect 17390 46786 17442 46798
rect 26238 46786 26290 46798
rect 16706 46734 16718 46786
rect 16770 46734 16782 46786
rect 21074 46734 21086 46786
rect 21138 46734 21150 46786
rect 11790 46722 11842 46734
rect 17390 46722 17442 46734
rect 26238 46722 26290 46734
rect 32174 46786 32226 46798
rect 32174 46722 32226 46734
rect 32286 46786 32338 46798
rect 32286 46722 32338 46734
rect 34078 46786 34130 46798
rect 34078 46722 34130 46734
rect 36766 46786 36818 46798
rect 36766 46722 36818 46734
rect 41246 46786 41298 46798
rect 41246 46722 41298 46734
rect 42366 46786 42418 46798
rect 49422 46786 49474 46798
rect 45826 46734 45838 46786
rect 45890 46734 45902 46786
rect 52658 46734 52670 46786
rect 52722 46734 52734 46786
rect 42366 46722 42418 46734
rect 49422 46722 49474 46734
rect 1710 46674 1762 46686
rect 1710 46610 1762 46622
rect 11566 46674 11618 46686
rect 11566 46610 11618 46622
rect 11678 46674 11730 46686
rect 11678 46610 11730 46622
rect 12014 46674 12066 46686
rect 16382 46674 16434 46686
rect 13234 46622 13246 46674
rect 13298 46622 13310 46674
rect 12014 46610 12066 46622
rect 16382 46610 16434 46622
rect 17614 46674 17666 46686
rect 17614 46610 17666 46622
rect 17950 46674 18002 46686
rect 17950 46610 18002 46622
rect 19854 46674 19906 46686
rect 19854 46610 19906 46622
rect 20078 46674 20130 46686
rect 20078 46610 20130 46622
rect 20526 46674 20578 46686
rect 26574 46674 26626 46686
rect 23650 46622 23662 46674
rect 23714 46622 23726 46674
rect 25666 46622 25678 46674
rect 25730 46622 25742 46674
rect 20526 46610 20578 46622
rect 26574 46610 26626 46622
rect 26798 46674 26850 46686
rect 26798 46610 26850 46622
rect 27022 46674 27074 46686
rect 30942 46674 30994 46686
rect 27570 46622 27582 46674
rect 27634 46622 27646 46674
rect 27022 46610 27074 46622
rect 30942 46610 30994 46622
rect 33966 46674 34018 46686
rect 33966 46610 34018 46622
rect 35198 46674 35250 46686
rect 35198 46610 35250 46622
rect 36654 46674 36706 46686
rect 40910 46674 40962 46686
rect 37090 46622 37102 46674
rect 37154 46622 37166 46674
rect 37874 46622 37886 46674
rect 37938 46622 37950 46674
rect 36654 46610 36706 46622
rect 40910 46610 40962 46622
rect 41134 46674 41186 46686
rect 41134 46610 41186 46622
rect 41694 46674 41746 46686
rect 41694 46610 41746 46622
rect 42254 46674 42306 46686
rect 45042 46622 45054 46674
rect 45106 46622 45118 46674
rect 48962 46622 48974 46674
rect 49026 46622 49038 46674
rect 49746 46622 49758 46674
rect 49810 46622 49822 46674
rect 53330 46622 53342 46674
rect 53394 46622 53406 46674
rect 42254 46610 42306 46622
rect 2494 46562 2546 46574
rect 2494 46498 2546 46510
rect 2942 46562 2994 46574
rect 2942 46498 2994 46510
rect 9886 46562 9938 46574
rect 9886 46498 9938 46510
rect 12686 46562 12738 46574
rect 24446 46562 24498 46574
rect 26686 46562 26738 46574
rect 33182 46562 33234 46574
rect 13906 46510 13918 46562
rect 13970 46510 13982 46562
rect 16034 46510 16046 46562
rect 16098 46510 16110 46562
rect 21858 46510 21870 46562
rect 21922 46510 21934 46562
rect 25330 46510 25342 46562
rect 25394 46510 25406 46562
rect 28242 46510 28254 46562
rect 28306 46510 28318 46562
rect 30370 46510 30382 46562
rect 30434 46510 30446 46562
rect 12686 46498 12738 46510
rect 24446 46498 24498 46510
rect 26686 46498 26738 46510
rect 33182 46498 33234 46510
rect 34862 46562 34914 46574
rect 34862 46498 34914 46510
rect 36206 46562 36258 46574
rect 44382 46562 44434 46574
rect 40002 46510 40014 46562
rect 40066 46510 40078 46562
rect 47954 46510 47966 46562
rect 48018 46510 48030 46562
rect 50530 46510 50542 46562
rect 50594 46510 50606 46562
rect 36206 46498 36258 46510
rect 44382 46498 44434 46510
rect 9774 46450 9826 46462
rect 2258 46398 2270 46450
rect 2322 46447 2334 46450
rect 3042 46447 3054 46450
rect 2322 46401 3054 46447
rect 2322 46398 2334 46401
rect 3042 46398 3054 46401
rect 3106 46398 3118 46450
rect 9774 46386 9826 46398
rect 20302 46450 20354 46462
rect 20302 46386 20354 46398
rect 32286 46450 32338 46462
rect 32286 46386 32338 46398
rect 41918 46450 41970 46462
rect 41918 46386 41970 46398
rect 42142 46450 42194 46462
rect 42142 46386 42194 46398
rect 44494 46450 44546 46462
rect 44494 46386 44546 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 13582 46114 13634 46126
rect 13582 46050 13634 46062
rect 14590 46114 14642 46126
rect 14590 46050 14642 46062
rect 20190 46114 20242 46126
rect 20190 46050 20242 46062
rect 26686 46114 26738 46126
rect 26686 46050 26738 46062
rect 48302 46114 48354 46126
rect 48302 46050 48354 46062
rect 48526 46114 48578 46126
rect 48526 46050 48578 46062
rect 13022 46002 13074 46014
rect 9090 45950 9102 46002
rect 9154 45950 9166 46002
rect 11218 45950 11230 46002
rect 11282 45950 11294 46002
rect 11778 45950 11790 46002
rect 11842 45950 11854 46002
rect 13022 45938 13074 45950
rect 14142 46002 14194 46014
rect 14142 45938 14194 45950
rect 14702 46002 14754 46014
rect 19630 46002 19682 46014
rect 15138 45950 15150 46002
rect 15202 45950 15214 46002
rect 14702 45938 14754 45950
rect 19630 45938 19682 45950
rect 20750 46002 20802 46014
rect 31726 46002 31778 46014
rect 37998 46002 38050 46014
rect 23874 45950 23886 46002
rect 23938 45950 23950 46002
rect 26002 45950 26014 46002
rect 26066 45950 26078 46002
rect 26450 45950 26462 46002
rect 26514 45950 26526 46002
rect 33954 45950 33966 46002
rect 34018 45950 34030 46002
rect 20750 45938 20802 45950
rect 31726 45938 31778 45950
rect 37998 45938 38050 45950
rect 40238 46002 40290 46014
rect 42142 46002 42194 46014
rect 40786 45950 40798 46002
rect 40850 45950 40862 46002
rect 40238 45938 40290 45950
rect 42142 45938 42194 45950
rect 48078 46002 48130 46014
rect 48078 45938 48130 45950
rect 49198 46002 49250 46014
rect 49198 45938 49250 45950
rect 50430 46002 50482 46014
rect 54898 45950 54910 46002
rect 54962 45950 54974 46002
rect 57698 45950 57710 46002
rect 57762 45950 57774 46002
rect 50430 45938 50482 45950
rect 13694 45890 13746 45902
rect 1810 45838 1822 45890
rect 1874 45838 1886 45890
rect 8418 45838 8430 45890
rect 8482 45838 8494 45890
rect 11554 45838 11566 45890
rect 11618 45838 11630 45890
rect 13694 45826 13746 45838
rect 13918 45890 13970 45902
rect 13918 45826 13970 45838
rect 15262 45890 15314 45902
rect 19966 45890 20018 45902
rect 15698 45838 15710 45890
rect 15762 45838 15774 45890
rect 15262 45826 15314 45838
rect 19966 45826 20018 45838
rect 20414 45890 20466 45902
rect 20414 45826 20466 45838
rect 20526 45890 20578 45902
rect 20526 45826 20578 45838
rect 21870 45890 21922 45902
rect 28142 45890 28194 45902
rect 22082 45838 22094 45890
rect 22146 45838 22158 45890
rect 23202 45838 23214 45890
rect 23266 45838 23278 45890
rect 26338 45838 26350 45890
rect 26402 45838 26414 45890
rect 21870 45826 21922 45838
rect 28142 45826 28194 45838
rect 28702 45890 28754 45902
rect 28702 45826 28754 45838
rect 32286 45890 32338 45902
rect 40126 45890 40178 45902
rect 45166 45890 45218 45902
rect 33394 45838 33406 45890
rect 33458 45838 33470 45890
rect 41010 45838 41022 45890
rect 41074 45838 41086 45890
rect 43698 45838 43710 45890
rect 43762 45838 43774 45890
rect 32286 45826 32338 45838
rect 40126 45826 40178 45838
rect 45166 45826 45218 45838
rect 45278 45890 45330 45902
rect 48638 45890 48690 45902
rect 47506 45838 47518 45890
rect 47570 45838 47582 45890
rect 52658 45838 52670 45890
rect 52722 45838 52734 45890
rect 55794 45838 55806 45890
rect 55858 45838 55870 45890
rect 45278 45826 45330 45838
rect 48638 45826 48690 45838
rect 2382 45778 2434 45790
rect 2382 45714 2434 45726
rect 3166 45778 3218 45790
rect 3166 45714 3218 45726
rect 11790 45778 11842 45790
rect 11790 45714 11842 45726
rect 12238 45778 12290 45790
rect 12238 45714 12290 45726
rect 14254 45778 14306 45790
rect 14254 45714 14306 45726
rect 18062 45778 18114 45790
rect 18062 45714 18114 45726
rect 18286 45778 18338 45790
rect 18286 45714 18338 45726
rect 22766 45778 22818 45790
rect 22766 45714 22818 45726
rect 32062 45778 32114 45790
rect 32062 45714 32114 45726
rect 41694 45778 41746 45790
rect 41694 45714 41746 45726
rect 45390 45778 45442 45790
rect 47966 45778 48018 45790
rect 47282 45726 47294 45778
rect 47346 45726 47358 45778
rect 45390 45714 45442 45726
rect 47966 45714 48018 45726
rect 51886 45778 51938 45790
rect 51886 45714 51938 45726
rect 2046 45666 2098 45678
rect 2046 45602 2098 45614
rect 2718 45666 2770 45678
rect 2718 45602 2770 45614
rect 12014 45666 12066 45678
rect 12014 45602 12066 45614
rect 15150 45666 15202 45678
rect 15150 45602 15202 45614
rect 15486 45666 15538 45678
rect 15486 45602 15538 45614
rect 18174 45666 18226 45678
rect 18174 45602 18226 45614
rect 21422 45666 21474 45678
rect 21422 45602 21474 45614
rect 27134 45666 27186 45678
rect 27134 45602 27186 45614
rect 28030 45666 28082 45678
rect 28030 45602 28082 45614
rect 28254 45666 28306 45678
rect 28254 45602 28306 45614
rect 29262 45666 29314 45678
rect 29262 45602 29314 45614
rect 32398 45666 32450 45678
rect 32398 45602 32450 45614
rect 32510 45666 32562 45678
rect 32510 45602 32562 45614
rect 35870 45666 35922 45678
rect 35870 45602 35922 45614
rect 39566 45666 39618 45678
rect 39566 45602 39618 45614
rect 39902 45666 39954 45678
rect 39902 45602 39954 45614
rect 40350 45666 40402 45678
rect 51998 45666 52050 45678
rect 43474 45614 43486 45666
rect 43538 45614 43550 45666
rect 45826 45614 45838 45666
rect 45890 45614 45902 45666
rect 40350 45602 40402 45614
rect 51998 45602 52050 45614
rect 52222 45666 52274 45678
rect 52222 45602 52274 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 10670 45330 10722 45342
rect 20638 45330 20690 45342
rect 16594 45278 16606 45330
rect 16658 45278 16670 45330
rect 10670 45266 10722 45278
rect 20638 45266 20690 45278
rect 21422 45330 21474 45342
rect 21422 45266 21474 45278
rect 25342 45330 25394 45342
rect 25342 45266 25394 45278
rect 27022 45330 27074 45342
rect 50878 45330 50930 45342
rect 38322 45278 38334 45330
rect 38386 45278 38398 45330
rect 27022 45266 27074 45278
rect 50878 45266 50930 45278
rect 54686 45330 54738 45342
rect 54686 45266 54738 45278
rect 2046 45218 2098 45230
rect 2046 45154 2098 45166
rect 11230 45218 11282 45230
rect 11230 45154 11282 45166
rect 14926 45218 14978 45230
rect 26238 45218 26290 45230
rect 31390 45218 31442 45230
rect 18162 45166 18174 45218
rect 18226 45166 18238 45218
rect 20962 45166 20974 45218
rect 21026 45166 21038 45218
rect 21746 45166 21758 45218
rect 21810 45166 21822 45218
rect 30594 45166 30606 45218
rect 30658 45166 30670 45218
rect 14926 45154 14978 45166
rect 26238 45154 26290 45166
rect 31390 45154 31442 45166
rect 34414 45218 34466 45230
rect 34414 45154 34466 45166
rect 34526 45218 34578 45230
rect 34526 45154 34578 45166
rect 45054 45218 45106 45230
rect 45054 45154 45106 45166
rect 45166 45218 45218 45230
rect 45166 45154 45218 45166
rect 47182 45218 47234 45230
rect 53330 45166 53342 45218
rect 53394 45166 53406 45218
rect 47182 45154 47234 45166
rect 1710 45106 1762 45118
rect 1710 45042 1762 45054
rect 10782 45106 10834 45118
rect 10782 45042 10834 45054
rect 11006 45106 11058 45118
rect 14366 45106 14418 45118
rect 15262 45106 15314 45118
rect 12114 45054 12126 45106
rect 12178 45054 12190 45106
rect 14690 45054 14702 45106
rect 14754 45054 14766 45106
rect 11006 45042 11058 45054
rect 14366 45042 14418 45054
rect 15262 45042 15314 45054
rect 16270 45106 16322 45118
rect 26798 45106 26850 45118
rect 17490 45054 17502 45106
rect 17554 45054 17566 45106
rect 22082 45054 22094 45106
rect 22146 45054 22158 45106
rect 26002 45054 26014 45106
rect 26066 45054 26078 45106
rect 16270 45042 16322 45054
rect 26798 45042 26850 45054
rect 27470 45106 27522 45118
rect 31166 45106 31218 45118
rect 29474 45054 29486 45106
rect 29538 45054 29550 45106
rect 30370 45054 30382 45106
rect 30434 45054 30446 45106
rect 27470 45042 27522 45054
rect 31166 45042 31218 45054
rect 31726 45106 31778 45118
rect 31726 45042 31778 45054
rect 31950 45106 32002 45118
rect 34750 45106 34802 45118
rect 33394 45054 33406 45106
rect 33458 45054 33470 45106
rect 33842 45054 33854 45106
rect 33906 45054 33918 45106
rect 31950 45042 32002 45054
rect 34750 45042 34802 45054
rect 35086 45106 35138 45118
rect 35086 45042 35138 45054
rect 35758 45106 35810 45118
rect 35758 45042 35810 45054
rect 36318 45106 36370 45118
rect 37886 45106 37938 45118
rect 37314 45054 37326 45106
rect 37378 45054 37390 45106
rect 36318 45042 36370 45054
rect 37886 45042 37938 45054
rect 38670 45106 38722 45118
rect 42814 45106 42866 45118
rect 41570 45054 41582 45106
rect 41634 45054 41646 45106
rect 38670 45042 38722 45054
rect 42814 45042 42866 45054
rect 43150 45106 43202 45118
rect 43150 45042 43202 45054
rect 43486 45106 43538 45118
rect 47630 45106 47682 45118
rect 54462 45106 54514 45118
rect 44258 45054 44270 45106
rect 44322 45054 44334 45106
rect 54002 45054 54014 45106
rect 54066 45054 54078 45106
rect 43486 45042 43538 45054
rect 47630 45042 47682 45054
rect 54462 45042 54514 45054
rect 55134 45106 55186 45118
rect 55134 45042 55186 45054
rect 55470 45106 55522 45118
rect 55470 45042 55522 45054
rect 2494 44994 2546 45006
rect 2494 44930 2546 44942
rect 9774 44994 9826 45006
rect 9774 44930 9826 44942
rect 10894 44994 10946 45006
rect 15374 44994 15426 45006
rect 13234 44942 13246 44994
rect 13298 44942 13310 44994
rect 14802 44942 14814 44994
rect 14866 44942 14878 44994
rect 10894 44930 10946 44942
rect 15374 44930 15426 44942
rect 15822 44994 15874 45006
rect 26910 44994 26962 45006
rect 20290 44942 20302 44994
rect 20354 44942 20366 44994
rect 23202 44942 23214 44994
rect 23266 44942 23278 44994
rect 15822 44930 15874 44942
rect 26910 44930 26962 44942
rect 29934 44994 29986 45006
rect 34078 44994 34130 45006
rect 31490 44942 31502 44994
rect 31554 44942 31566 44994
rect 29934 44930 29986 44942
rect 34078 44930 34130 44942
rect 37998 44994 38050 45006
rect 37998 44930 38050 44942
rect 38894 44994 38946 45006
rect 42254 44994 42306 45006
rect 41794 44942 41806 44994
rect 41858 44942 41870 44994
rect 38894 44930 38946 44942
rect 42254 44930 42306 44942
rect 43262 44994 43314 45006
rect 44718 44994 44770 45006
rect 43810 44942 43822 44994
rect 43874 44942 43886 44994
rect 43262 44930 43314 44942
rect 44718 44930 44770 44942
rect 47406 44994 47458 45006
rect 54574 44994 54626 45006
rect 51202 44942 51214 44994
rect 51266 44942 51278 44994
rect 47406 44930 47458 44942
rect 54574 44930 54626 44942
rect 9662 44882 9714 44894
rect 9662 44818 9714 44830
rect 45166 44882 45218 44894
rect 45166 44818 45218 44830
rect 47854 44882 47906 44894
rect 47854 44818 47906 44830
rect 48302 44882 48354 44894
rect 48302 44818 48354 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 25902 44546 25954 44558
rect 24322 44494 24334 44546
rect 24386 44543 24398 44546
rect 24546 44543 24558 44546
rect 24386 44497 24558 44543
rect 24386 44494 24398 44497
rect 24546 44494 24558 44497
rect 24610 44494 24622 44546
rect 25902 44482 25954 44494
rect 38110 44546 38162 44558
rect 38110 44482 38162 44494
rect 38782 44546 38834 44558
rect 38782 44482 38834 44494
rect 43710 44546 43762 44558
rect 43710 44482 43762 44494
rect 46286 44546 46338 44558
rect 46286 44482 46338 44494
rect 46510 44546 46562 44558
rect 51662 44546 51714 44558
rect 49410 44494 49422 44546
rect 49474 44494 49486 44546
rect 46510 44482 46562 44494
rect 51662 44482 51714 44494
rect 1934 44434 1986 44446
rect 18510 44434 18562 44446
rect 8866 44382 8878 44434
rect 8930 44382 8942 44434
rect 10994 44382 11006 44434
rect 11058 44382 11070 44434
rect 15586 44382 15598 44434
rect 15650 44382 15662 44434
rect 1934 44370 1986 44382
rect 18510 44370 18562 44382
rect 20750 44434 20802 44446
rect 20750 44370 20802 44382
rect 23662 44434 23714 44446
rect 23662 44370 23714 44382
rect 24558 44434 24610 44446
rect 24558 44370 24610 44382
rect 25006 44434 25058 44446
rect 25006 44370 25058 44382
rect 25678 44434 25730 44446
rect 27918 44434 27970 44446
rect 39006 44434 39058 44446
rect 27234 44382 27246 44434
rect 27298 44382 27310 44434
rect 32050 44382 32062 44434
rect 32114 44382 32126 44434
rect 32946 44382 32958 44434
rect 33010 44382 33022 44434
rect 25678 44370 25730 44382
rect 27918 44370 27970 44382
rect 39006 44370 39058 44382
rect 43822 44434 43874 44446
rect 43822 44370 43874 44382
rect 45390 44434 45442 44446
rect 45390 44370 45442 44382
rect 45726 44434 45778 44446
rect 50878 44434 50930 44446
rect 49074 44382 49086 44434
rect 49138 44382 49150 44434
rect 45726 44370 45778 44382
rect 50878 44370 50930 44382
rect 51886 44434 51938 44446
rect 51886 44370 51938 44382
rect 52110 44434 52162 44446
rect 52110 44370 52162 44382
rect 55022 44434 55074 44446
rect 57810 44382 57822 44434
rect 57874 44382 57886 44434
rect 55022 44370 55074 44382
rect 12462 44322 12514 44334
rect 4274 44270 4286 44322
rect 4338 44270 4350 44322
rect 8194 44270 8206 44322
rect 8258 44270 8270 44322
rect 12462 44258 12514 44270
rect 12574 44322 12626 44334
rect 12574 44258 12626 44270
rect 13022 44322 13074 44334
rect 13022 44258 13074 44270
rect 13918 44322 13970 44334
rect 13918 44258 13970 44270
rect 14254 44322 14306 44334
rect 14254 44258 14306 44270
rect 17614 44322 17666 44334
rect 17614 44258 17666 44270
rect 18622 44322 18674 44334
rect 18622 44258 18674 44270
rect 21422 44322 21474 44334
rect 24222 44322 24274 44334
rect 21858 44270 21870 44322
rect 21922 44270 21934 44322
rect 23090 44270 23102 44322
rect 23154 44270 23166 44322
rect 21422 44258 21474 44270
rect 24222 44258 24274 44270
rect 26126 44322 26178 44334
rect 32510 44322 32562 44334
rect 35310 44322 35362 44334
rect 38558 44322 38610 44334
rect 27122 44270 27134 44322
rect 27186 44270 27198 44322
rect 29138 44270 29150 44322
rect 29202 44270 29214 44322
rect 33170 44270 33182 44322
rect 33234 44270 33246 44322
rect 35634 44270 35646 44322
rect 35698 44270 35710 44322
rect 26126 44258 26178 44270
rect 32510 44258 32562 44270
rect 35310 44258 35362 44270
rect 38558 44258 38610 44270
rect 39566 44322 39618 44334
rect 39566 44258 39618 44270
rect 40014 44322 40066 44334
rect 40014 44258 40066 44270
rect 41470 44322 41522 44334
rect 41470 44258 41522 44270
rect 41806 44322 41858 44334
rect 41806 44258 41858 44270
rect 42926 44322 42978 44334
rect 42926 44258 42978 44270
rect 43038 44322 43090 44334
rect 43038 44258 43090 44270
rect 45950 44322 46002 44334
rect 45950 44258 46002 44270
rect 47070 44322 47122 44334
rect 47506 44270 47518 44322
rect 47570 44270 47582 44322
rect 48962 44270 48974 44322
rect 49026 44270 49038 44322
rect 52658 44270 52670 44322
rect 52722 44270 52734 44322
rect 55682 44270 55694 44322
rect 55746 44270 55758 44322
rect 47070 44258 47122 44270
rect 13582 44210 13634 44222
rect 13582 44146 13634 44158
rect 14478 44210 14530 44222
rect 14478 44146 14530 44158
rect 14926 44210 14978 44222
rect 14926 44146 14978 44158
rect 15262 44210 15314 44222
rect 15262 44146 15314 44158
rect 15486 44210 15538 44222
rect 15486 44146 15538 44158
rect 16270 44210 16322 44222
rect 16270 44146 16322 44158
rect 18398 44210 18450 44222
rect 18398 44146 18450 44158
rect 18958 44210 19010 44222
rect 18958 44146 19010 44158
rect 19406 44210 19458 44222
rect 19406 44146 19458 44158
rect 22318 44210 22370 44222
rect 22318 44146 22370 44158
rect 22654 44210 22706 44222
rect 22654 44146 22706 44158
rect 23550 44210 23602 44222
rect 23550 44146 23602 44158
rect 23774 44210 23826 44222
rect 33854 44210 33906 44222
rect 29922 44158 29934 44210
rect 29986 44158 29998 44210
rect 23774 44146 23826 44158
rect 33854 44146 33906 44158
rect 34190 44210 34242 44222
rect 34190 44146 34242 44158
rect 34414 44210 34466 44222
rect 34414 44146 34466 44158
rect 34750 44210 34802 44222
rect 34750 44146 34802 44158
rect 35086 44210 35138 44222
rect 35086 44146 35138 44158
rect 39342 44210 39394 44222
rect 39342 44146 39394 44158
rect 43262 44210 43314 44222
rect 43262 44146 43314 44158
rect 47966 44210 48018 44222
rect 47966 44146 48018 44158
rect 50766 44210 50818 44222
rect 50766 44146 50818 44158
rect 50990 44210 51042 44222
rect 50990 44146 51042 44158
rect 51214 44210 51266 44222
rect 51214 44146 51266 44158
rect 11454 44098 11506 44110
rect 11454 44034 11506 44046
rect 12798 44098 12850 44110
rect 12798 44034 12850 44046
rect 14030 44098 14082 44110
rect 18062 44098 18114 44110
rect 15922 44046 15934 44098
rect 15986 44046 15998 44098
rect 17266 44046 17278 44098
rect 17330 44046 17342 44098
rect 14030 44034 14082 44046
rect 18062 44034 18114 44046
rect 20414 44098 20466 44110
rect 20414 44034 20466 44046
rect 26574 44098 26626 44110
rect 26574 44034 26626 44046
rect 34638 44098 34690 44110
rect 34638 44034 34690 44046
rect 35198 44098 35250 44110
rect 35198 44034 35250 44046
rect 39454 44098 39506 44110
rect 39454 44034 39506 44046
rect 41582 44098 41634 44110
rect 41582 44034 41634 44046
rect 42814 44098 42866 44110
rect 42814 44034 42866 44046
rect 46622 44098 46674 44110
rect 46622 44034 46674 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 27470 43762 27522 43774
rect 10210 43710 10222 43762
rect 10274 43710 10286 43762
rect 27470 43698 27522 43710
rect 29710 43762 29762 43774
rect 29710 43698 29762 43710
rect 33630 43762 33682 43774
rect 33630 43698 33682 43710
rect 42926 43762 42978 43774
rect 42926 43698 42978 43710
rect 49086 43762 49138 43774
rect 49086 43698 49138 43710
rect 2046 43650 2098 43662
rect 2046 43586 2098 43598
rect 4846 43650 4898 43662
rect 4846 43586 4898 43598
rect 5294 43650 5346 43662
rect 19630 43650 19682 43662
rect 17490 43598 17502 43650
rect 17554 43598 17566 43650
rect 5294 43586 5346 43598
rect 19630 43586 19682 43598
rect 19854 43650 19906 43662
rect 19854 43586 19906 43598
rect 19966 43650 20018 43662
rect 19966 43586 20018 43598
rect 20078 43650 20130 43662
rect 20078 43586 20130 43598
rect 22318 43650 22370 43662
rect 22318 43586 22370 43598
rect 23214 43650 23266 43662
rect 23214 43586 23266 43598
rect 23438 43650 23490 43662
rect 23438 43586 23490 43598
rect 23662 43650 23714 43662
rect 23662 43586 23714 43598
rect 24334 43650 24386 43662
rect 24334 43586 24386 43598
rect 27022 43650 27074 43662
rect 27022 43586 27074 43598
rect 29038 43650 29090 43662
rect 29038 43586 29090 43598
rect 29150 43650 29202 43662
rect 29150 43586 29202 43598
rect 33406 43650 33458 43662
rect 33406 43586 33458 43598
rect 33518 43650 33570 43662
rect 37774 43650 37826 43662
rect 35186 43598 35198 43650
rect 35250 43598 35262 43650
rect 33518 43586 33570 43598
rect 37774 43586 37826 43598
rect 40126 43650 40178 43662
rect 40126 43586 40178 43598
rect 40238 43650 40290 43662
rect 40238 43586 40290 43598
rect 43374 43650 43426 43662
rect 43374 43586 43426 43598
rect 48750 43650 48802 43662
rect 48750 43586 48802 43598
rect 48862 43650 48914 43662
rect 48862 43586 48914 43598
rect 49870 43650 49922 43662
rect 49870 43586 49922 43598
rect 49982 43650 50034 43662
rect 49982 43586 50034 43598
rect 53006 43650 53058 43662
rect 53006 43586 53058 43598
rect 53118 43650 53170 43662
rect 53118 43586 53170 43598
rect 1710 43538 1762 43550
rect 17838 43538 17890 43550
rect 23998 43538 24050 43550
rect 27246 43538 27298 43550
rect 8642 43486 8654 43538
rect 8706 43486 8718 43538
rect 9986 43486 9998 43538
rect 10050 43486 10062 43538
rect 10546 43486 10558 43538
rect 10610 43486 10622 43538
rect 13906 43486 13918 43538
rect 13970 43486 13982 43538
rect 20738 43486 20750 43538
rect 20802 43486 20814 43538
rect 25778 43486 25790 43538
rect 25842 43486 25854 43538
rect 1710 43474 1762 43486
rect 17838 43474 17890 43486
rect 23998 43474 24050 43486
rect 27246 43474 27298 43486
rect 29598 43538 29650 43550
rect 29598 43474 29650 43486
rect 29822 43538 29874 43550
rect 32958 43538 33010 43550
rect 37662 43538 37714 43550
rect 42142 43538 42194 43550
rect 30146 43486 30158 43538
rect 30210 43486 30222 43538
rect 34514 43486 34526 43538
rect 34578 43486 34590 43538
rect 38994 43486 39006 43538
rect 39058 43486 39070 43538
rect 29822 43474 29874 43486
rect 32958 43474 33010 43486
rect 37662 43474 37714 43486
rect 42142 43474 42194 43486
rect 42590 43538 42642 43550
rect 42590 43474 42642 43486
rect 42814 43538 42866 43550
rect 51214 43538 51266 43550
rect 46050 43486 46062 43538
rect 46114 43486 46126 43538
rect 47394 43486 47406 43538
rect 47458 43486 47470 43538
rect 50866 43486 50878 43538
rect 50930 43486 50942 43538
rect 42814 43474 42866 43486
rect 51214 43474 51266 43486
rect 51774 43538 51826 43550
rect 52098 43486 52110 43538
rect 52162 43486 52174 43538
rect 53442 43486 53454 43538
rect 53506 43486 53518 43538
rect 51774 43474 51826 43486
rect 2494 43426 2546 43438
rect 21422 43426 21474 43438
rect 5730 43374 5742 43426
rect 5794 43374 5806 43426
rect 7858 43374 7870 43426
rect 7922 43374 7934 43426
rect 11330 43374 11342 43426
rect 11394 43374 11406 43426
rect 13458 43374 13470 43426
rect 13522 43374 13534 43426
rect 14690 43374 14702 43426
rect 14754 43374 14766 43426
rect 16818 43374 16830 43426
rect 16882 43374 16894 43426
rect 20514 43374 20526 43426
rect 20578 43374 20590 43426
rect 2494 43362 2546 43374
rect 21422 43362 21474 43374
rect 22878 43426 22930 43438
rect 27134 43426 27186 43438
rect 23538 43374 23550 43426
rect 23602 43374 23614 43426
rect 26450 43374 26462 43426
rect 26514 43374 26526 43426
rect 22878 43362 22930 43374
rect 27134 43362 27186 43374
rect 28702 43426 28754 43438
rect 38222 43426 38274 43438
rect 41022 43426 41074 43438
rect 37314 43374 37326 43426
rect 37378 43374 37390 43426
rect 39330 43374 39342 43426
rect 39394 43374 39406 43426
rect 28702 43362 28754 43374
rect 38222 43362 38274 43374
rect 41022 43362 41074 43374
rect 43822 43426 43874 43438
rect 46734 43426 46786 43438
rect 51326 43426 51378 43438
rect 46274 43374 46286 43426
rect 46338 43374 46350 43426
rect 47506 43374 47518 43426
rect 47570 43374 47582 43426
rect 43822 43362 43874 43374
rect 46734 43362 46786 43374
rect 51326 43362 51378 43374
rect 51662 43426 51714 43438
rect 51662 43362 51714 43374
rect 4622 43314 4674 43326
rect 4622 43250 4674 43262
rect 4958 43314 5010 43326
rect 4958 43250 5010 43262
rect 5406 43314 5458 43326
rect 5406 43250 5458 43262
rect 22542 43314 22594 43326
rect 29150 43314 29202 43326
rect 40126 43314 40178 43326
rect 26562 43262 26574 43314
rect 26626 43262 26638 43314
rect 38994 43262 39006 43314
rect 39058 43262 39070 43314
rect 22542 43250 22594 43262
rect 29150 43250 29202 43262
rect 40126 43250 40178 43262
rect 42030 43314 42082 43326
rect 42030 43250 42082 43262
rect 43262 43314 43314 43326
rect 49870 43314 49922 43326
rect 48066 43262 48078 43314
rect 48130 43262 48142 43314
rect 55346 43262 55358 43314
rect 55410 43262 55422 43314
rect 43262 43250 43314 43262
rect 49870 43250 49922 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 4062 42978 4114 42990
rect 4062 42914 4114 42926
rect 11230 42978 11282 42990
rect 11230 42914 11282 42926
rect 12014 42978 12066 42990
rect 12014 42914 12066 42926
rect 13470 42978 13522 42990
rect 13470 42914 13522 42926
rect 14366 42978 14418 42990
rect 14366 42914 14418 42926
rect 14702 42978 14754 42990
rect 14702 42914 14754 42926
rect 17950 42978 18002 42990
rect 17950 42914 18002 42926
rect 18174 42978 18226 42990
rect 18174 42914 18226 42926
rect 20526 42978 20578 42990
rect 20526 42914 20578 42926
rect 46286 42978 46338 42990
rect 46286 42914 46338 42926
rect 6078 42866 6130 42878
rect 6078 42802 6130 42814
rect 8878 42866 8930 42878
rect 8878 42802 8930 42814
rect 10446 42866 10498 42878
rect 10446 42802 10498 42814
rect 13582 42866 13634 42878
rect 13582 42802 13634 42814
rect 18286 42866 18338 42878
rect 18286 42802 18338 42814
rect 20078 42866 20130 42878
rect 20078 42802 20130 42814
rect 47518 42866 47570 42878
rect 51202 42814 51214 42866
rect 51266 42814 51278 42866
rect 47518 42802 47570 42814
rect 3390 42754 3442 42766
rect 5854 42754 5906 42766
rect 15486 42754 15538 42766
rect 23326 42754 23378 42766
rect 3714 42702 3726 42754
rect 3778 42702 3790 42754
rect 5618 42702 5630 42754
rect 5682 42702 5694 42754
rect 6738 42702 6750 42754
rect 6802 42702 6814 42754
rect 8306 42702 8318 42754
rect 8370 42702 8382 42754
rect 14690 42702 14702 42754
rect 14754 42702 14766 42754
rect 22530 42702 22542 42754
rect 22594 42702 22606 42754
rect 22754 42702 22766 42754
rect 22818 42702 22830 42754
rect 3390 42690 3442 42702
rect 5854 42690 5906 42702
rect 15486 42690 15538 42702
rect 23326 42690 23378 42702
rect 23886 42754 23938 42766
rect 25118 42754 25170 42766
rect 24322 42702 24334 42754
rect 24386 42702 24398 42754
rect 24546 42702 24558 42754
rect 24610 42702 24622 42754
rect 23886 42690 23938 42702
rect 25118 42690 25170 42702
rect 25678 42754 25730 42766
rect 25678 42690 25730 42702
rect 26910 42754 26962 42766
rect 26910 42690 26962 42702
rect 28142 42754 28194 42766
rect 35422 42754 35474 42766
rect 32498 42702 32510 42754
rect 32562 42702 32574 42754
rect 28142 42690 28194 42702
rect 35422 42690 35474 42702
rect 35534 42754 35586 42766
rect 35534 42690 35586 42702
rect 39006 42754 39058 42766
rect 42590 42754 42642 42766
rect 46398 42754 46450 42766
rect 39666 42702 39678 42754
rect 39730 42702 39742 42754
rect 40114 42702 40126 42754
rect 40178 42702 40190 42754
rect 42130 42702 42142 42754
rect 42194 42702 42206 42754
rect 42802 42702 42814 42754
rect 42866 42702 42878 42754
rect 39006 42690 39058 42702
rect 42590 42690 42642 42702
rect 46398 42690 46450 42702
rect 47406 42754 47458 42766
rect 47406 42690 47458 42702
rect 47630 42754 47682 42766
rect 47630 42690 47682 42702
rect 49422 42754 49474 42766
rect 49422 42690 49474 42702
rect 50430 42754 50482 42766
rect 50430 42690 50482 42702
rect 50766 42754 50818 42766
rect 51426 42702 51438 42754
rect 51490 42702 51502 42754
rect 54786 42702 54798 42754
rect 54850 42702 54862 42754
rect 55570 42702 55582 42754
rect 55634 42702 55646 42754
rect 50766 42690 50818 42702
rect 1710 42642 1762 42654
rect 1710 42578 1762 42590
rect 2046 42642 2098 42654
rect 2046 42578 2098 42590
rect 6190 42642 6242 42654
rect 8094 42642 8146 42654
rect 6850 42590 6862 42642
rect 6914 42590 6926 42642
rect 7522 42590 7534 42642
rect 7586 42590 7598 42642
rect 6190 42578 6242 42590
rect 8094 42578 8146 42590
rect 8766 42642 8818 42654
rect 8766 42578 8818 42590
rect 11342 42642 11394 42654
rect 11342 42578 11394 42590
rect 11566 42642 11618 42654
rect 11566 42578 11618 42590
rect 11902 42642 11954 42654
rect 11902 42578 11954 42590
rect 17838 42642 17890 42654
rect 17838 42578 17890 42590
rect 19070 42642 19122 42654
rect 19070 42578 19122 42590
rect 19406 42642 19458 42654
rect 20526 42642 20578 42654
rect 19406 42578 19458 42590
rect 20414 42586 20466 42598
rect 2494 42530 2546 42542
rect 2494 42466 2546 42478
rect 3950 42530 4002 42542
rect 13694 42530 13746 42542
rect 18734 42530 18786 42542
rect 7634 42478 7646 42530
rect 7698 42478 7710 42530
rect 15138 42478 15150 42530
rect 15202 42478 15214 42530
rect 3950 42466 4002 42478
rect 13694 42466 13746 42478
rect 18734 42466 18786 42478
rect 19518 42530 19570 42542
rect 20526 42578 20578 42590
rect 23774 42642 23826 42654
rect 23774 42578 23826 42590
rect 25342 42642 25394 42654
rect 25342 42578 25394 42590
rect 26350 42642 26402 42654
rect 26350 42578 26402 42590
rect 26574 42642 26626 42654
rect 26574 42578 26626 42590
rect 28254 42642 28306 42654
rect 28254 42578 28306 42590
rect 29262 42642 29314 42654
rect 29262 42578 29314 42590
rect 30382 42642 30434 42654
rect 30382 42578 30434 42590
rect 30718 42642 30770 42654
rect 30718 42578 30770 42590
rect 31278 42642 31330 42654
rect 34078 42642 34130 42654
rect 35870 42642 35922 42654
rect 32722 42590 32734 42642
rect 32786 42590 32798 42642
rect 33730 42590 33742 42642
rect 33794 42590 33806 42642
rect 34402 42590 34414 42642
rect 34466 42590 34478 42642
rect 31278 42578 31330 42590
rect 34078 42578 34130 42590
rect 35870 42578 35922 42590
rect 40350 42642 40402 42654
rect 40350 42578 40402 42590
rect 42366 42642 42418 42654
rect 42366 42578 42418 42590
rect 46286 42642 46338 42654
rect 46286 42578 46338 42590
rect 47854 42642 47906 42654
rect 47854 42578 47906 42590
rect 50654 42642 50706 42654
rect 50654 42578 50706 42590
rect 52110 42642 52162 42654
rect 53666 42590 53678 42642
rect 53730 42590 53742 42642
rect 57362 42590 57374 42642
rect 57426 42590 57438 42642
rect 52110 42578 52162 42590
rect 20414 42522 20466 42534
rect 21870 42530 21922 42542
rect 19518 42466 19570 42478
rect 21870 42466 21922 42478
rect 22318 42530 22370 42542
rect 22318 42466 22370 42478
rect 22990 42530 23042 42542
rect 22990 42466 23042 42478
rect 23102 42530 23154 42542
rect 23102 42466 23154 42478
rect 23662 42530 23714 42542
rect 23662 42466 23714 42478
rect 24782 42530 24834 42542
rect 24782 42466 24834 42478
rect 24894 42530 24946 42542
rect 24894 42466 24946 42478
rect 25566 42530 25618 42542
rect 25566 42466 25618 42478
rect 26686 42530 26738 42542
rect 26686 42466 26738 42478
rect 28478 42530 28530 42542
rect 28478 42466 28530 42478
rect 34750 42530 34802 42542
rect 34750 42466 34802 42478
rect 35758 42530 35810 42542
rect 35758 42466 35810 42478
rect 38446 42530 38498 42542
rect 38446 42466 38498 42478
rect 38670 42530 38722 42542
rect 38670 42466 38722 42478
rect 38894 42530 38946 42542
rect 38894 42466 38946 42478
rect 42478 42530 42530 42542
rect 42478 42466 42530 42478
rect 43486 42530 43538 42542
rect 43486 42466 43538 42478
rect 45054 42530 45106 42542
rect 45054 42466 45106 42478
rect 48862 42530 48914 42542
rect 48862 42466 48914 42478
rect 49086 42530 49138 42542
rect 49086 42466 49138 42478
rect 49310 42530 49362 42542
rect 49310 42466 49362 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 2046 42194 2098 42206
rect 2046 42130 2098 42142
rect 3950 42194 4002 42206
rect 12126 42194 12178 42206
rect 5842 42142 5854 42194
rect 5906 42142 5918 42194
rect 3950 42130 4002 42142
rect 12126 42130 12178 42142
rect 25902 42194 25954 42206
rect 25902 42130 25954 42142
rect 26126 42194 26178 42206
rect 31950 42194 32002 42206
rect 29362 42142 29374 42194
rect 29426 42142 29438 42194
rect 26126 42130 26178 42142
rect 31950 42130 32002 42142
rect 33742 42194 33794 42206
rect 33742 42130 33794 42142
rect 34750 42194 34802 42206
rect 49534 42194 49586 42206
rect 41570 42142 41582 42194
rect 41634 42142 41646 42194
rect 45714 42142 45726 42194
rect 45778 42142 45790 42194
rect 34750 42130 34802 42142
rect 49534 42130 49586 42142
rect 51214 42194 51266 42206
rect 51214 42130 51266 42142
rect 51326 42194 51378 42206
rect 51326 42130 51378 42142
rect 51438 42194 51490 42206
rect 51438 42130 51490 42142
rect 6190 42082 6242 42094
rect 8206 42082 8258 42094
rect 4386 42030 4398 42082
rect 4450 42030 4462 42082
rect 5954 42030 5966 42082
rect 6018 42030 6030 42082
rect 6514 42030 6526 42082
rect 6578 42030 6590 42082
rect 7074 42030 7086 42082
rect 7138 42030 7150 42082
rect 6190 42018 6242 42030
rect 8206 42018 8258 42030
rect 10334 42082 10386 42094
rect 12574 42082 12626 42094
rect 11442 42030 11454 42082
rect 11506 42030 11518 42082
rect 10334 42018 10386 42030
rect 12574 42018 12626 42030
rect 12686 42082 12738 42094
rect 23214 42082 23266 42094
rect 13794 42030 13806 42082
rect 13858 42030 13870 42082
rect 21298 42030 21310 42082
rect 21362 42030 21374 42082
rect 21634 42030 21646 42082
rect 21698 42030 21710 42082
rect 12686 42018 12738 42030
rect 23214 42018 23266 42030
rect 23550 42082 23602 42094
rect 23550 42018 23602 42030
rect 23662 42082 23714 42094
rect 23662 42018 23714 42030
rect 26350 42082 26402 42094
rect 26350 42018 26402 42030
rect 26798 42082 26850 42094
rect 26798 42018 26850 42030
rect 30718 42082 30770 42094
rect 39678 42082 39730 42094
rect 47966 42082 48018 42094
rect 35858 42030 35870 42082
rect 35922 42030 35934 42082
rect 43138 42030 43150 42082
rect 43202 42030 43214 42082
rect 30718 42018 30770 42030
rect 39678 42018 39730 42030
rect 47966 42018 48018 42030
rect 48078 42082 48130 42094
rect 48078 42018 48130 42030
rect 49310 42082 49362 42094
rect 49310 42018 49362 42030
rect 1710 41970 1762 41982
rect 1710 41906 1762 41918
rect 3838 41970 3890 41982
rect 5406 41970 5458 41982
rect 4274 41918 4286 41970
rect 4338 41918 4350 41970
rect 3838 41906 3890 41918
rect 5406 41906 5458 41918
rect 6302 41970 6354 41982
rect 6302 41906 6354 41918
rect 8094 41970 8146 41982
rect 11118 41970 11170 41982
rect 10546 41918 10558 41970
rect 10610 41918 10622 41970
rect 8094 41906 8146 41918
rect 11118 41906 11170 41918
rect 12014 41970 12066 41982
rect 12014 41906 12066 41918
rect 12350 41970 12402 41982
rect 12350 41906 12402 41918
rect 12910 41970 12962 41982
rect 12910 41906 12962 41918
rect 13470 41970 13522 41982
rect 20750 41970 20802 41982
rect 17378 41918 17390 41970
rect 17442 41918 17454 41970
rect 18162 41918 18174 41970
rect 18226 41918 18238 41970
rect 13470 41906 13522 41918
rect 20750 41906 20802 41918
rect 21086 41970 21138 41982
rect 21086 41906 21138 41918
rect 22542 41970 22594 41982
rect 22542 41906 22594 41918
rect 22990 41970 23042 41982
rect 22990 41906 23042 41918
rect 26686 41970 26738 41982
rect 26686 41906 26738 41918
rect 29038 41970 29090 41982
rect 29038 41906 29090 41918
rect 30270 41970 30322 41982
rect 30270 41906 30322 41918
rect 30494 41970 30546 41982
rect 30494 41906 30546 41918
rect 30942 41970 30994 41982
rect 39230 41970 39282 41982
rect 35074 41918 35086 41970
rect 35138 41918 35150 41970
rect 30942 41906 30994 41918
rect 39230 41906 39282 41918
rect 39902 41970 39954 41982
rect 39902 41906 39954 41918
rect 41246 41970 41298 41982
rect 46062 41970 46114 41982
rect 42354 41918 42366 41970
rect 42418 41918 42430 41970
rect 41246 41906 41298 41918
rect 46062 41906 46114 41918
rect 47518 41970 47570 41982
rect 47518 41906 47570 41918
rect 49086 41970 49138 41982
rect 49086 41906 49138 41918
rect 51886 41970 51938 41982
rect 53006 41970 53058 41982
rect 52546 41918 52558 41970
rect 52610 41918 52622 41970
rect 53442 41918 53454 41970
rect 53506 41918 53518 41970
rect 51886 41906 51938 41918
rect 53006 41906 53058 41918
rect 2494 41858 2546 41870
rect 2494 41794 2546 41806
rect 2942 41858 2994 41870
rect 2942 41794 2994 41806
rect 8654 41858 8706 41870
rect 8654 41794 8706 41806
rect 14254 41858 14306 41870
rect 14254 41794 14306 41806
rect 14926 41858 14978 41870
rect 14926 41794 14978 41806
rect 16942 41858 16994 41870
rect 22766 41858 22818 41870
rect 20290 41806 20302 41858
rect 20354 41806 20366 41858
rect 16942 41794 16994 41806
rect 22766 41794 22818 41806
rect 24222 41858 24274 41870
rect 24222 41794 24274 41806
rect 24670 41858 24722 41870
rect 24670 41794 24722 41806
rect 27358 41858 27410 41870
rect 27358 41794 27410 41806
rect 30830 41858 30882 41870
rect 30830 41794 30882 41806
rect 31390 41858 31442 41870
rect 38446 41858 38498 41870
rect 37986 41806 37998 41858
rect 38050 41806 38062 41858
rect 31390 41794 31442 41806
rect 38446 41794 38498 41806
rect 38894 41858 38946 41870
rect 38894 41794 38946 41806
rect 39790 41858 39842 41870
rect 39790 41794 39842 41806
rect 40350 41858 40402 41870
rect 46510 41858 46562 41870
rect 45266 41806 45278 41858
rect 45330 41806 45342 41858
rect 40350 41794 40402 41806
rect 46510 41794 46562 41806
rect 49198 41858 49250 41870
rect 49198 41794 49250 41806
rect 50878 41858 50930 41870
rect 50878 41794 50930 41806
rect 53118 41858 53170 41870
rect 55234 41806 55246 41858
rect 55298 41806 55310 41858
rect 53118 41794 53170 41806
rect 8206 41746 8258 41758
rect 8206 41682 8258 41694
rect 8766 41746 8818 41758
rect 8766 41682 8818 41694
rect 23662 41746 23714 41758
rect 23662 41682 23714 41694
rect 26238 41746 26290 41758
rect 26238 41682 26290 41694
rect 26798 41746 26850 41758
rect 26798 41682 26850 41694
rect 47966 41746 48018 41758
rect 47966 41682 48018 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 13582 41410 13634 41422
rect 13582 41346 13634 41358
rect 20190 41298 20242 41310
rect 12674 41246 12686 41298
rect 12738 41246 12750 41298
rect 20190 41234 20242 41246
rect 22094 41298 22146 41310
rect 36430 41298 36482 41310
rect 42142 41298 42194 41310
rect 55022 41298 55074 41310
rect 28578 41246 28590 41298
rect 28642 41246 28654 41298
rect 31378 41246 31390 41298
rect 31442 41246 31454 41298
rect 33506 41246 33518 41298
rect 33570 41246 33582 41298
rect 37426 41246 37438 41298
rect 37490 41246 37502 41298
rect 39554 41246 39566 41298
rect 39618 41246 39630 41298
rect 41682 41246 41694 41298
rect 41746 41246 41758 41298
rect 43586 41246 43598 41298
rect 43650 41246 43662 41298
rect 51202 41246 51214 41298
rect 51266 41246 51278 41298
rect 22094 41234 22146 41246
rect 36430 41234 36482 41246
rect 42142 41234 42194 41246
rect 55022 41234 55074 41246
rect 57934 41298 57986 41310
rect 57934 41234 57986 41246
rect 8206 41186 8258 41198
rect 13694 41186 13746 41198
rect 1810 41134 1822 41186
rect 1874 41134 1886 41186
rect 7634 41134 7646 41186
rect 7698 41134 7710 41186
rect 10882 41134 10894 41186
rect 10946 41134 10958 41186
rect 8206 41122 8258 41134
rect 13694 41122 13746 41134
rect 14030 41186 14082 41198
rect 14030 41122 14082 41134
rect 14366 41186 14418 41198
rect 14366 41122 14418 41134
rect 15038 41186 15090 41198
rect 15038 41122 15090 41134
rect 15150 41186 15202 41198
rect 15150 41122 15202 41134
rect 15822 41186 15874 41198
rect 15822 41122 15874 41134
rect 19182 41186 19234 41198
rect 19182 41122 19234 41134
rect 19518 41186 19570 41198
rect 22542 41186 22594 41198
rect 22418 41134 22430 41186
rect 22482 41134 22494 41186
rect 19518 41122 19570 41134
rect 22542 41122 22594 41134
rect 23326 41186 23378 41198
rect 23326 41122 23378 41134
rect 23550 41186 23602 41198
rect 23550 41122 23602 41134
rect 23774 41186 23826 41198
rect 23774 41122 23826 41134
rect 23998 41186 24050 41198
rect 23998 41122 24050 41134
rect 24334 41186 24386 41198
rect 30046 41186 30098 41198
rect 34190 41186 34242 41198
rect 42254 41186 42306 41198
rect 45166 41186 45218 41198
rect 25778 41134 25790 41186
rect 25842 41134 25854 41186
rect 30706 41134 30718 41186
rect 30770 41134 30782 41186
rect 38210 41134 38222 41186
rect 38274 41134 38286 41186
rect 38770 41134 38782 41186
rect 38834 41134 38846 41186
rect 42802 41134 42814 41186
rect 42866 41134 42878 41186
rect 43922 41134 43934 41186
rect 43986 41134 43998 41186
rect 24334 41122 24386 41134
rect 30046 41122 30098 41134
rect 34190 41122 34242 41134
rect 42254 41122 42306 41134
rect 45166 41122 45218 41134
rect 47630 41186 47682 41198
rect 47954 41134 47966 41186
rect 48018 41134 48030 41186
rect 48402 41134 48414 41186
rect 48466 41134 48478 41186
rect 52658 41134 52670 41186
rect 52722 41134 52734 41186
rect 55906 41134 55918 41186
rect 55970 41134 55982 41186
rect 47630 41122 47682 41134
rect 2046 41074 2098 41086
rect 2046 41010 2098 41022
rect 2382 41074 2434 41086
rect 2382 41010 2434 41022
rect 2718 41074 2770 41086
rect 2718 41010 2770 41022
rect 3166 41074 3218 41086
rect 8654 41074 8706 41086
rect 6178 41022 6190 41074
rect 6242 41022 6254 41074
rect 3166 41010 3218 41022
rect 8654 41010 8706 41022
rect 13582 41074 13634 41086
rect 13582 41010 13634 41022
rect 14590 41074 14642 41086
rect 14590 41010 14642 41022
rect 14926 41074 14978 41086
rect 14926 41010 14978 41022
rect 15486 41074 15538 41086
rect 15486 41010 15538 41022
rect 16046 41074 16098 41086
rect 16046 41010 16098 41022
rect 19630 41074 19682 41086
rect 19630 41010 19682 41022
rect 19854 41074 19906 41086
rect 19854 41010 19906 41022
rect 24670 41074 24722 41086
rect 24670 41010 24722 41022
rect 25006 41074 25058 41086
rect 45278 41074 45330 41086
rect 47518 41074 47570 41086
rect 26450 41022 26462 41074
rect 26514 41022 26526 41074
rect 38434 41022 38446 41074
rect 38498 41022 38510 41074
rect 46722 41022 46734 41074
rect 46786 41022 46798 41074
rect 49074 41022 49086 41074
rect 49138 41022 49150 41074
rect 25006 41010 25058 41022
rect 45278 41010 45330 41022
rect 47518 41010 47570 41022
rect 14142 40962 14194 40974
rect 6290 40910 6302 40962
rect 6354 40910 6366 40962
rect 14142 40898 14194 40910
rect 15934 40962 15986 40974
rect 15934 40898 15986 40910
rect 16606 40962 16658 40974
rect 16606 40898 16658 40910
rect 18398 40962 18450 40974
rect 18398 40898 18450 40910
rect 18734 40962 18786 40974
rect 18734 40898 18786 40910
rect 18958 40962 19010 40974
rect 18958 40898 19010 40910
rect 19070 40962 19122 40974
rect 19070 40898 19122 40910
rect 21646 40962 21698 40974
rect 21646 40898 21698 40910
rect 22654 40962 22706 40974
rect 22654 40898 22706 40910
rect 22766 40962 22818 40974
rect 22766 40898 22818 40910
rect 23438 40962 23490 40974
rect 23438 40898 23490 40910
rect 24446 40962 24498 40974
rect 24446 40898 24498 40910
rect 29486 40962 29538 40974
rect 29486 40898 29538 40910
rect 34750 40962 34802 40974
rect 34750 40898 34802 40910
rect 35646 40962 35698 40974
rect 35646 40898 35698 40910
rect 36990 40962 37042 40974
rect 36990 40898 37042 40910
rect 45502 40962 45554 40974
rect 45502 40898 45554 40910
rect 45950 40962 46002 40974
rect 45950 40898 46002 40910
rect 46398 40962 46450 40974
rect 46398 40898 46450 40910
rect 47406 40962 47458 40974
rect 47406 40898 47458 40910
rect 51662 40962 51714 40974
rect 51662 40898 51714 40910
rect 52110 40962 52162 40974
rect 52110 40898 52162 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 8654 40626 8706 40638
rect 8654 40562 8706 40574
rect 13358 40626 13410 40638
rect 25342 40626 25394 40638
rect 21410 40574 21422 40626
rect 21474 40574 21486 40626
rect 13358 40562 13410 40574
rect 25342 40562 25394 40574
rect 26686 40626 26738 40638
rect 26686 40562 26738 40574
rect 26798 40626 26850 40638
rect 26798 40562 26850 40574
rect 26910 40626 26962 40638
rect 26910 40562 26962 40574
rect 27918 40626 27970 40638
rect 27918 40562 27970 40574
rect 28814 40626 28866 40638
rect 28814 40562 28866 40574
rect 29934 40626 29986 40638
rect 29934 40562 29986 40574
rect 30942 40626 30994 40638
rect 30942 40562 30994 40574
rect 31614 40626 31666 40638
rect 31614 40562 31666 40574
rect 31950 40626 32002 40638
rect 31950 40562 32002 40574
rect 38110 40626 38162 40638
rect 38110 40562 38162 40574
rect 38670 40626 38722 40638
rect 38670 40562 38722 40574
rect 41470 40626 41522 40638
rect 41470 40562 41522 40574
rect 41694 40626 41746 40638
rect 41694 40562 41746 40574
rect 42030 40626 42082 40638
rect 42030 40562 42082 40574
rect 56590 40626 56642 40638
rect 56590 40562 56642 40574
rect 2046 40514 2098 40526
rect 12798 40514 12850 40526
rect 10322 40462 10334 40514
rect 10386 40462 10398 40514
rect 2046 40450 2098 40462
rect 12798 40450 12850 40462
rect 13582 40514 13634 40526
rect 25678 40514 25730 40526
rect 14690 40462 14702 40514
rect 14754 40462 14766 40514
rect 22530 40462 22542 40514
rect 22594 40462 22606 40514
rect 13582 40450 13634 40462
rect 25678 40450 25730 40462
rect 25790 40514 25842 40526
rect 25790 40450 25842 40462
rect 29822 40514 29874 40526
rect 29822 40450 29874 40462
rect 30718 40514 30770 40526
rect 41022 40514 41074 40526
rect 39554 40462 39566 40514
rect 39618 40462 39630 40514
rect 30718 40450 30770 40462
rect 41022 40450 41074 40462
rect 41358 40514 41410 40526
rect 41358 40450 41410 40462
rect 42590 40514 42642 40526
rect 50082 40462 50094 40514
rect 50146 40462 50158 40514
rect 42590 40450 42642 40462
rect 1710 40402 1762 40414
rect 1710 40338 1762 40350
rect 2494 40402 2546 40414
rect 7870 40402 7922 40414
rect 19406 40402 19458 40414
rect 30046 40402 30098 40414
rect 4610 40350 4622 40402
rect 4674 40350 4686 40402
rect 9538 40350 9550 40402
rect 9602 40350 9614 40402
rect 14018 40350 14030 40402
rect 14082 40350 14094 40402
rect 18834 40350 18846 40402
rect 18898 40350 18910 40402
rect 21186 40350 21198 40402
rect 21250 40350 21262 40402
rect 21858 40350 21870 40402
rect 21922 40350 21934 40402
rect 2494 40338 2546 40350
rect 7870 40338 7922 40350
rect 19406 40338 19458 40350
rect 30046 40338 30098 40350
rect 30382 40402 30434 40414
rect 30382 40338 30434 40350
rect 31278 40402 31330 40414
rect 31278 40338 31330 40350
rect 32510 40402 32562 40414
rect 37774 40402 37826 40414
rect 33842 40350 33854 40402
rect 33906 40350 33918 40402
rect 32510 40338 32562 40350
rect 37774 40338 37826 40350
rect 39902 40402 39954 40414
rect 39902 40338 39954 40350
rect 42814 40402 42866 40414
rect 42814 40338 42866 40350
rect 43262 40402 43314 40414
rect 43262 40338 43314 40350
rect 43486 40402 43538 40414
rect 48862 40402 48914 40414
rect 56814 40402 56866 40414
rect 44370 40350 44382 40402
rect 44434 40350 44446 40402
rect 45266 40350 45278 40402
rect 45330 40350 45342 40402
rect 49298 40350 49310 40402
rect 49362 40350 49374 40402
rect 52770 40350 52782 40402
rect 52834 40350 52846 40402
rect 53442 40350 53454 40402
rect 53506 40350 53518 40402
rect 57138 40350 57150 40402
rect 57202 40350 57214 40402
rect 43486 40338 43538 40350
rect 48862 40338 48914 40350
rect 56814 40338 56866 40350
rect 12910 40290 12962 40302
rect 5282 40238 5294 40290
rect 5346 40238 5358 40290
rect 7410 40238 7422 40290
rect 7474 40238 7486 40290
rect 12450 40238 12462 40290
rect 12514 40238 12526 40290
rect 12910 40226 12962 40238
rect 13470 40290 13522 40302
rect 19518 40290 19570 40302
rect 26238 40290 26290 40302
rect 16818 40238 16830 40290
rect 16882 40238 16894 40290
rect 24658 40238 24670 40290
rect 24722 40238 24734 40290
rect 13470 40226 13522 40238
rect 19518 40226 19570 40238
rect 26238 40226 26290 40238
rect 26462 40290 26514 40302
rect 37438 40290 37490 40302
rect 43374 40290 43426 40302
rect 44830 40290 44882 40302
rect 56030 40290 56082 40302
rect 34514 40238 34526 40290
rect 34578 40238 34590 40290
rect 36642 40238 36654 40290
rect 36706 40238 36718 40290
rect 39106 40238 39118 40290
rect 39170 40238 39182 40290
rect 43922 40238 43934 40290
rect 43986 40238 43998 40290
rect 45938 40238 45950 40290
rect 46002 40238 46014 40290
rect 48066 40238 48078 40290
rect 48130 40238 48142 40290
rect 52210 40238 52222 40290
rect 52274 40238 52286 40290
rect 55570 40238 55582 40290
rect 55634 40238 55646 40290
rect 26462 40226 26514 40238
rect 37438 40226 37490 40238
rect 43374 40226 43426 40238
rect 44830 40226 44882 40238
rect 56030 40226 56082 40238
rect 56702 40290 56754 40302
rect 56702 40226 56754 40238
rect 7758 40178 7810 40190
rect 7758 40114 7810 40126
rect 8318 40178 8370 40190
rect 8318 40114 8370 40126
rect 8542 40178 8594 40190
rect 8542 40114 8594 40126
rect 25790 40178 25842 40190
rect 25790 40114 25842 40126
rect 31054 40178 31106 40190
rect 31054 40114 31106 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 10670 39842 10722 39854
rect 10322 39790 10334 39842
rect 10386 39790 10398 39842
rect 10670 39778 10722 39790
rect 12126 39842 12178 39854
rect 12126 39778 12178 39790
rect 32398 39842 32450 39854
rect 32398 39778 32450 39790
rect 1934 39730 1986 39742
rect 1934 39666 1986 39678
rect 6526 39730 6578 39742
rect 10894 39730 10946 39742
rect 7074 39678 7086 39730
rect 7138 39678 7150 39730
rect 9202 39678 9214 39730
rect 9266 39678 9278 39730
rect 6526 39666 6578 39678
rect 10894 39666 10946 39678
rect 11566 39730 11618 39742
rect 29262 39730 29314 39742
rect 14242 39678 14254 39730
rect 14306 39678 14318 39730
rect 16370 39678 16382 39730
rect 16434 39678 16446 39730
rect 22082 39678 22094 39730
rect 22146 39678 22158 39730
rect 24210 39678 24222 39730
rect 24274 39678 24286 39730
rect 24770 39678 24782 39730
rect 24834 39678 24846 39730
rect 11566 39666 11618 39678
rect 29262 39666 29314 39678
rect 30606 39730 30658 39742
rect 30606 39666 30658 39678
rect 34078 39730 34130 39742
rect 44942 39730 44994 39742
rect 44258 39678 44270 39730
rect 44322 39678 44334 39730
rect 34078 39666 34130 39678
rect 44942 39666 44994 39678
rect 45726 39730 45778 39742
rect 45726 39666 45778 39678
rect 48974 39730 49026 39742
rect 48974 39666 49026 39678
rect 51214 39730 51266 39742
rect 51214 39666 51266 39678
rect 51662 39730 51714 39742
rect 51662 39666 51714 39678
rect 52782 39730 52834 39742
rect 53218 39678 53230 39730
rect 53282 39678 53294 39730
rect 55346 39678 55358 39730
rect 55410 39678 55422 39730
rect 52782 39666 52834 39678
rect 6078 39618 6130 39630
rect 11902 39618 11954 39630
rect 4274 39566 4286 39618
rect 4338 39566 4350 39618
rect 9986 39566 9998 39618
rect 10050 39566 10062 39618
rect 6078 39554 6130 39566
rect 11902 39554 11954 39566
rect 12910 39618 12962 39630
rect 18958 39618 19010 39630
rect 28254 39618 28306 39630
rect 32286 39618 32338 39630
rect 35870 39618 35922 39630
rect 13570 39566 13582 39618
rect 13634 39566 13646 39618
rect 18386 39566 18398 39618
rect 18450 39566 18462 39618
rect 21298 39566 21310 39618
rect 21362 39566 21374 39618
rect 27682 39566 27694 39618
rect 27746 39566 27758 39618
rect 28578 39566 28590 39618
rect 28642 39566 28654 39618
rect 34514 39566 34526 39618
rect 34578 39566 34590 39618
rect 35074 39566 35086 39618
rect 35138 39566 35150 39618
rect 12910 39554 12962 39566
rect 18958 39554 19010 39566
rect 28254 39554 28306 39566
rect 32286 39554 32338 39566
rect 35870 39554 35922 39566
rect 37214 39618 37266 39630
rect 37214 39554 37266 39566
rect 38446 39618 38498 39630
rect 45838 39618 45890 39630
rect 41458 39566 41470 39618
rect 41522 39566 41534 39618
rect 45266 39566 45278 39618
rect 45330 39566 45342 39618
rect 38446 39554 38498 39566
rect 45838 39554 45890 39566
rect 51550 39618 51602 39630
rect 51550 39554 51602 39566
rect 52222 39618 52274 39630
rect 56018 39566 56030 39618
rect 56082 39566 56094 39618
rect 52222 39554 52274 39566
rect 5966 39506 6018 39518
rect 5966 39442 6018 39454
rect 19070 39506 19122 39518
rect 31614 39506 31666 39518
rect 26898 39454 26910 39506
rect 26962 39454 26974 39506
rect 19070 39442 19122 39454
rect 31614 39442 31666 39454
rect 31950 39506 32002 39518
rect 31950 39442 32002 39454
rect 33966 39506 34018 39518
rect 37538 39454 37550 39506
rect 37602 39454 37614 39506
rect 42130 39454 42142 39506
rect 42194 39454 42206 39506
rect 33966 39442 34018 39454
rect 5742 39394 5794 39406
rect 5742 39330 5794 39342
rect 6414 39394 6466 39406
rect 28030 39394 28082 39406
rect 12450 39342 12462 39394
rect 12514 39342 12526 39394
rect 6414 39330 6466 39342
rect 28030 39330 28082 39342
rect 28142 39394 28194 39406
rect 28142 39330 28194 39342
rect 31390 39394 31442 39406
rect 31390 39330 31442 39342
rect 32398 39394 32450 39406
rect 32398 39330 32450 39342
rect 33742 39394 33794 39406
rect 33742 39330 33794 39342
rect 34190 39394 34242 39406
rect 34190 39330 34242 39342
rect 34862 39394 34914 39406
rect 34862 39330 34914 39342
rect 36206 39394 36258 39406
rect 36206 39330 36258 39342
rect 37998 39394 38050 39406
rect 37998 39330 38050 39342
rect 38894 39394 38946 39406
rect 38894 39330 38946 39342
rect 45614 39394 45666 39406
rect 45614 39330 45666 39342
rect 50318 39394 50370 39406
rect 50318 39330 50370 39342
rect 50766 39394 50818 39406
rect 50766 39330 50818 39342
rect 51774 39394 51826 39406
rect 51774 39330 51826 39342
rect 56590 39394 56642 39406
rect 56590 39330 56642 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 7646 39058 7698 39070
rect 7646 38994 7698 39006
rect 8990 39058 9042 39070
rect 8990 38994 9042 39006
rect 10222 39058 10274 39070
rect 10222 38994 10274 39006
rect 11118 39058 11170 39070
rect 11118 38994 11170 39006
rect 13022 39058 13074 39070
rect 13022 38994 13074 39006
rect 13582 39058 13634 39070
rect 13582 38994 13634 39006
rect 14142 39058 14194 39070
rect 14142 38994 14194 39006
rect 15598 39058 15650 39070
rect 15598 38994 15650 39006
rect 24446 39058 24498 39070
rect 24446 38994 24498 39006
rect 25678 39058 25730 39070
rect 25678 38994 25730 39006
rect 25902 39058 25954 39070
rect 25902 38994 25954 39006
rect 33182 39058 33234 39070
rect 33182 38994 33234 39006
rect 33966 39058 34018 39070
rect 33966 38994 34018 39006
rect 34302 39058 34354 39070
rect 34302 38994 34354 39006
rect 34526 39058 34578 39070
rect 34526 38994 34578 39006
rect 35758 39058 35810 39070
rect 35758 38994 35810 39006
rect 41806 39058 41858 39070
rect 41806 38994 41858 39006
rect 41918 39058 41970 39070
rect 41918 38994 41970 39006
rect 43822 39058 43874 39070
rect 43822 38994 43874 39006
rect 52222 39058 52274 39070
rect 52222 38994 52274 39006
rect 53230 39058 53282 39070
rect 53230 38994 53282 39006
rect 2046 38946 2098 38958
rect 2046 38882 2098 38894
rect 4622 38946 4674 38958
rect 4622 38882 4674 38894
rect 6414 38946 6466 38958
rect 13358 38946 13410 38958
rect 35422 38946 35474 38958
rect 12674 38894 12686 38946
rect 12738 38894 12750 38946
rect 15922 38894 15934 38946
rect 15986 38894 15998 38946
rect 21410 38894 21422 38946
rect 21474 38894 21486 38946
rect 27122 38894 27134 38946
rect 27186 38894 27198 38946
rect 6414 38882 6466 38894
rect 13358 38882 13410 38894
rect 35422 38882 35474 38894
rect 35982 38946 36034 38958
rect 35982 38882 36034 38894
rect 36654 38946 36706 38958
rect 36654 38882 36706 38894
rect 36990 38946 37042 38958
rect 36990 38882 37042 38894
rect 42590 38946 42642 38958
rect 42590 38882 42642 38894
rect 42814 38946 42866 38958
rect 52446 38946 52498 38958
rect 45490 38894 45502 38946
rect 45554 38894 45566 38946
rect 42814 38882 42866 38894
rect 52446 38882 52498 38894
rect 53006 38946 53058 38958
rect 53006 38882 53058 38894
rect 56702 38946 56754 38958
rect 56702 38882 56754 38894
rect 1710 38834 1762 38846
rect 1710 38770 1762 38782
rect 4734 38834 4786 38846
rect 4734 38770 4786 38782
rect 5966 38834 6018 38846
rect 5966 38770 6018 38782
rect 6862 38834 6914 38846
rect 6862 38770 6914 38782
rect 20862 38834 20914 38846
rect 21870 38834 21922 38846
rect 21186 38782 21198 38834
rect 21250 38782 21262 38834
rect 20862 38770 20914 38782
rect 21870 38770 21922 38782
rect 22430 38834 22482 38846
rect 22430 38770 22482 38782
rect 25230 38834 25282 38846
rect 25230 38770 25282 38782
rect 25790 38834 25842 38846
rect 34190 38834 34242 38846
rect 26450 38782 26462 38834
rect 26514 38782 26526 38834
rect 25790 38770 25842 38782
rect 29586 38770 29598 38822
rect 29650 38770 29662 38822
rect 34190 38770 34242 38782
rect 35534 38834 35586 38846
rect 35534 38770 35586 38782
rect 36094 38834 36146 38846
rect 36094 38770 36146 38782
rect 36878 38834 36930 38846
rect 41582 38834 41634 38846
rect 37426 38782 37438 38834
rect 37490 38782 37502 38834
rect 36878 38770 36930 38782
rect 41582 38770 41634 38782
rect 42030 38834 42082 38846
rect 42030 38770 42082 38782
rect 42478 38834 42530 38846
rect 42478 38770 42530 38782
rect 42926 38834 42978 38846
rect 42926 38770 42978 38782
rect 45838 38834 45890 38846
rect 52558 38834 52610 38846
rect 48850 38782 48862 38834
rect 48914 38782 48926 38834
rect 45838 38770 45890 38782
rect 52558 38770 52610 38782
rect 52894 38834 52946 38846
rect 53442 38782 53454 38834
rect 53506 38782 53518 38834
rect 52894 38770 52946 38782
rect 2494 38722 2546 38734
rect 2494 38658 2546 38670
rect 5070 38722 5122 38734
rect 5070 38658 5122 38670
rect 6750 38722 6802 38734
rect 6750 38658 6802 38670
rect 25454 38722 25506 38734
rect 35086 38722 35138 38734
rect 44158 38722 44210 38734
rect 29250 38670 29262 38722
rect 29314 38670 29326 38722
rect 30370 38670 30382 38722
rect 30434 38670 30446 38722
rect 32498 38670 32510 38722
rect 32562 38670 32574 38722
rect 38210 38670 38222 38722
rect 38274 38670 38286 38722
rect 40338 38670 40350 38722
rect 40402 38670 40414 38722
rect 25454 38658 25506 38670
rect 35086 38658 35138 38670
rect 44158 38658 44210 38670
rect 46510 38722 46562 38734
rect 49522 38670 49534 38722
rect 49586 38670 49598 38722
rect 51650 38670 51662 38722
rect 51714 38670 51726 38722
rect 46510 38658 46562 38670
rect 5182 38610 5234 38622
rect 5182 38546 5234 38558
rect 5518 38610 5570 38622
rect 5518 38546 5570 38558
rect 5630 38610 5682 38622
rect 5630 38546 5682 38558
rect 5854 38610 5906 38622
rect 5854 38546 5906 38558
rect 6526 38610 6578 38622
rect 6526 38546 6578 38558
rect 13694 38610 13746 38622
rect 35422 38610 35474 38622
rect 13906 38558 13918 38610
rect 13970 38607 13982 38610
rect 14242 38607 14254 38610
rect 13970 38561 14254 38607
rect 13970 38558 13982 38561
rect 14242 38558 14254 38561
rect 14306 38558 14318 38610
rect 13694 38546 13746 38558
rect 35422 38546 35474 38558
rect 36990 38610 37042 38622
rect 36990 38546 37042 38558
rect 46622 38610 46674 38622
rect 55346 38558 55358 38610
rect 55410 38558 55422 38610
rect 46622 38546 46674 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 5854 38274 5906 38286
rect 5854 38210 5906 38222
rect 6190 38274 6242 38286
rect 6190 38210 6242 38222
rect 12574 38274 12626 38286
rect 12574 38210 12626 38222
rect 36542 38274 36594 38286
rect 36542 38210 36594 38222
rect 37326 38274 37378 38286
rect 39666 38222 39678 38274
rect 39730 38271 39742 38274
rect 40002 38271 40014 38274
rect 39730 38225 40014 38271
rect 39730 38222 39742 38225
rect 40002 38222 40014 38225
rect 40066 38222 40078 38274
rect 37326 38210 37378 38222
rect 14814 38162 14866 38174
rect 23774 38162 23826 38174
rect 10882 38110 10894 38162
rect 10946 38110 10958 38162
rect 18722 38110 18734 38162
rect 18786 38110 18798 38162
rect 14814 38098 14866 38110
rect 23774 38098 23826 38110
rect 29486 38162 29538 38174
rect 29486 38098 29538 38110
rect 30270 38162 30322 38174
rect 30270 38098 30322 38110
rect 30830 38162 30882 38174
rect 30830 38098 30882 38110
rect 31838 38162 31890 38174
rect 31838 38098 31890 38110
rect 37886 38162 37938 38174
rect 45054 38162 45106 38174
rect 44146 38110 44158 38162
rect 44210 38110 44222 38162
rect 37886 38098 37938 38110
rect 45054 38098 45106 38110
rect 47182 38162 47234 38174
rect 51650 38110 51662 38162
rect 51714 38110 51726 38162
rect 55906 38110 55918 38162
rect 55970 38110 55982 38162
rect 47182 38098 47234 38110
rect 5966 38050 6018 38062
rect 5966 37986 6018 37998
rect 6414 38050 6466 38062
rect 12014 38050 12066 38062
rect 8082 37998 8094 38050
rect 8146 37998 8158 38050
rect 6414 37986 6466 37998
rect 12014 37986 12066 37998
rect 12238 38050 12290 38062
rect 12238 37986 12290 37998
rect 13806 38050 13858 38062
rect 13806 37986 13858 37998
rect 14366 38050 14418 38062
rect 19966 38050 20018 38062
rect 15250 37998 15262 38050
rect 15314 37998 15326 38050
rect 15810 37998 15822 38050
rect 15874 37998 15886 38050
rect 14366 37986 14418 37998
rect 19966 37986 20018 37998
rect 21870 38050 21922 38062
rect 29710 38050 29762 38062
rect 22306 37998 22318 38050
rect 22370 37998 22382 38050
rect 21870 37986 21922 37998
rect 29710 37986 29762 37998
rect 30158 38050 30210 38062
rect 30158 37986 30210 37998
rect 32174 38050 32226 38062
rect 32174 37986 32226 37998
rect 35646 38050 35698 38062
rect 35646 37986 35698 37998
rect 37550 38050 37602 38062
rect 37550 37986 37602 37998
rect 37774 38050 37826 38062
rect 37774 37986 37826 37998
rect 37998 38050 38050 38062
rect 40686 38050 40738 38062
rect 46622 38050 46674 38062
rect 40226 37998 40238 38050
rect 40290 37998 40302 38050
rect 40898 37998 40910 38050
rect 40962 37998 40974 38050
rect 41346 37998 41358 38050
rect 41410 37998 41422 38050
rect 37998 37986 38050 37998
rect 40686 37986 40738 37998
rect 46622 37986 46674 37998
rect 46958 38050 47010 38062
rect 46958 37986 47010 37998
rect 47070 38050 47122 38062
rect 47070 37986 47122 37998
rect 47294 38050 47346 38062
rect 48738 37998 48750 38050
rect 48802 37998 48814 38050
rect 52994 37998 53006 38050
rect 53058 37998 53070 38050
rect 47294 37986 47346 37998
rect 1710 37938 1762 37950
rect 1710 37874 1762 37886
rect 2046 37938 2098 37950
rect 2046 37874 2098 37886
rect 6526 37938 6578 37950
rect 6526 37874 6578 37886
rect 7310 37938 7362 37950
rect 7310 37874 7362 37886
rect 7646 37938 7698 37950
rect 11342 37938 11394 37950
rect 8754 37886 8766 37938
rect 8818 37886 8830 37938
rect 7646 37874 7698 37886
rect 11342 37874 11394 37886
rect 11566 37938 11618 37950
rect 11566 37874 11618 37886
rect 14030 37938 14082 37950
rect 14030 37874 14082 37886
rect 15486 37938 15538 37950
rect 20190 37938 20242 37950
rect 16594 37886 16606 37938
rect 16658 37886 16670 37938
rect 15486 37874 15538 37886
rect 20190 37874 20242 37886
rect 20862 37938 20914 37950
rect 35982 37938 36034 37950
rect 34290 37886 34302 37938
rect 34354 37886 34366 37938
rect 34962 37886 34974 37938
rect 35026 37886 35038 37938
rect 20862 37874 20914 37886
rect 35982 37874 36034 37886
rect 36430 37938 36482 37950
rect 36430 37874 36482 37886
rect 40574 37938 40626 37950
rect 46286 37938 46338 37950
rect 42018 37886 42030 37938
rect 42082 37886 42094 37938
rect 40574 37874 40626 37886
rect 46286 37874 46338 37886
rect 47518 37938 47570 37950
rect 49522 37886 49534 37938
rect 49586 37886 49598 37938
rect 53778 37886 53790 37938
rect 53842 37886 53854 37938
rect 47518 37874 47570 37886
rect 2494 37826 2546 37838
rect 2494 37762 2546 37774
rect 11454 37826 11506 37838
rect 11454 37762 11506 37774
rect 14254 37826 14306 37838
rect 21310 37826 21362 37838
rect 23214 37826 23266 37838
rect 19618 37774 19630 37826
rect 19682 37774 19694 37826
rect 22530 37774 22542 37826
rect 22594 37774 22606 37826
rect 14254 37762 14306 37774
rect 21310 37762 21362 37774
rect 23214 37762 23266 37774
rect 27806 37826 27858 37838
rect 27806 37762 27858 37774
rect 28590 37826 28642 37838
rect 28590 37762 28642 37774
rect 30382 37826 30434 37838
rect 30382 37762 30434 37774
rect 32510 37826 32562 37838
rect 32510 37762 32562 37774
rect 33182 37826 33234 37838
rect 33182 37762 33234 37774
rect 33630 37826 33682 37838
rect 33630 37762 33682 37774
rect 33966 37826 34018 37838
rect 33966 37762 34018 37774
rect 34638 37826 34690 37838
rect 36206 37826 36258 37838
rect 35298 37774 35310 37826
rect 35362 37774 35374 37826
rect 34638 37762 34690 37774
rect 36206 37762 36258 37774
rect 40014 37826 40066 37838
rect 40014 37762 40066 37774
rect 40462 37826 40514 37838
rect 40462 37762 40514 37774
rect 46398 37826 46450 37838
rect 46398 37762 46450 37774
rect 52222 37826 52274 37838
rect 52222 37762 52274 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 2046 37490 2098 37502
rect 2046 37426 2098 37438
rect 6302 37490 6354 37502
rect 6302 37426 6354 37438
rect 15374 37490 15426 37502
rect 15374 37426 15426 37438
rect 28366 37490 28418 37502
rect 28366 37426 28418 37438
rect 28926 37490 28978 37502
rect 28926 37426 28978 37438
rect 29038 37490 29090 37502
rect 29038 37426 29090 37438
rect 30382 37490 30434 37502
rect 30382 37426 30434 37438
rect 30718 37490 30770 37502
rect 30718 37426 30770 37438
rect 31390 37490 31442 37502
rect 31390 37426 31442 37438
rect 33406 37490 33458 37502
rect 33406 37426 33458 37438
rect 34414 37490 34466 37502
rect 34414 37426 34466 37438
rect 37326 37490 37378 37502
rect 37326 37426 37378 37438
rect 39454 37490 39506 37502
rect 39454 37426 39506 37438
rect 40126 37490 40178 37502
rect 40126 37426 40178 37438
rect 41358 37490 41410 37502
rect 41358 37426 41410 37438
rect 45838 37490 45890 37502
rect 45838 37426 45890 37438
rect 46174 37490 46226 37502
rect 46174 37426 46226 37438
rect 50430 37490 50482 37502
rect 50430 37426 50482 37438
rect 50878 37490 50930 37502
rect 50878 37426 50930 37438
rect 51438 37490 51490 37502
rect 51438 37426 51490 37438
rect 52446 37490 52498 37502
rect 52446 37426 52498 37438
rect 6974 37378 7026 37390
rect 6974 37314 7026 37326
rect 7310 37378 7362 37390
rect 12462 37378 12514 37390
rect 11218 37326 11230 37378
rect 11282 37326 11294 37378
rect 7310 37314 7362 37326
rect 12462 37314 12514 37326
rect 14814 37378 14866 37390
rect 24334 37378 24386 37390
rect 15922 37326 15934 37378
rect 15986 37326 15998 37378
rect 16482 37326 16494 37378
rect 16546 37326 16558 37378
rect 14814 37314 14866 37326
rect 24334 37314 24386 37326
rect 25230 37378 25282 37390
rect 25230 37314 25282 37326
rect 26910 37378 26962 37390
rect 26910 37314 26962 37326
rect 29262 37378 29314 37390
rect 37102 37378 37154 37390
rect 34738 37326 34750 37378
rect 34802 37326 34814 37378
rect 29262 37314 29314 37326
rect 37102 37314 37154 37326
rect 37438 37378 37490 37390
rect 37438 37314 37490 37326
rect 39902 37378 39954 37390
rect 39902 37314 39954 37326
rect 41134 37378 41186 37390
rect 46286 37378 46338 37390
rect 42130 37326 42142 37378
rect 42194 37326 42206 37378
rect 41134 37314 41186 37326
rect 46286 37314 46338 37326
rect 47630 37378 47682 37390
rect 47630 37314 47682 37326
rect 51214 37378 51266 37390
rect 51214 37314 51266 37326
rect 52222 37378 52274 37390
rect 52222 37314 52274 37326
rect 1710 37266 1762 37278
rect 1710 37202 1762 37214
rect 5854 37266 5906 37278
rect 5854 37202 5906 37214
rect 5966 37266 6018 37278
rect 5966 37202 6018 37214
rect 6190 37266 6242 37278
rect 6190 37202 6242 37214
rect 11566 37266 11618 37278
rect 13806 37266 13858 37278
rect 13346 37214 13358 37266
rect 13410 37214 13422 37266
rect 11566 37202 11618 37214
rect 13806 37202 13858 37214
rect 14366 37266 14418 37278
rect 21310 37266 21362 37278
rect 20962 37214 20974 37266
rect 21026 37214 21038 37266
rect 14366 37202 14418 37214
rect 21310 37202 21362 37214
rect 21422 37266 21474 37278
rect 21422 37202 21474 37214
rect 21646 37266 21698 37278
rect 21646 37202 21698 37214
rect 21870 37266 21922 37278
rect 21870 37202 21922 37214
rect 22318 37266 22370 37278
rect 26686 37266 26738 37278
rect 23650 37214 23662 37266
rect 23714 37214 23726 37266
rect 25666 37214 25678 37266
rect 25730 37214 25742 37266
rect 22318 37202 22370 37214
rect 26686 37202 26738 37214
rect 27022 37266 27074 37278
rect 27022 37202 27074 37214
rect 27582 37266 27634 37278
rect 27582 37202 27634 37214
rect 27918 37266 27970 37278
rect 27918 37202 27970 37214
rect 28030 37266 28082 37278
rect 28030 37202 28082 37214
rect 28142 37266 28194 37278
rect 28142 37202 28194 37214
rect 28814 37266 28866 37278
rect 28814 37202 28866 37214
rect 36878 37266 36930 37278
rect 36878 37202 36930 37214
rect 37774 37266 37826 37278
rect 39790 37266 39842 37278
rect 38210 37214 38222 37266
rect 38274 37214 38286 37266
rect 37774 37202 37826 37214
rect 39790 37202 39842 37214
rect 40910 37266 40962 37278
rect 40910 37202 40962 37214
rect 41806 37266 41858 37278
rect 41806 37202 41858 37214
rect 46062 37266 46114 37278
rect 48078 37266 48130 37278
rect 47058 37214 47070 37266
rect 47122 37214 47134 37266
rect 46062 37202 46114 37214
rect 48078 37202 48130 37214
rect 48862 37266 48914 37278
rect 48862 37202 48914 37214
rect 51550 37266 51602 37278
rect 51550 37202 51602 37214
rect 51662 37266 51714 37278
rect 51662 37202 51714 37214
rect 51774 37266 51826 37278
rect 51774 37202 51826 37214
rect 52670 37266 52722 37278
rect 52670 37202 52722 37214
rect 52782 37266 52834 37278
rect 56018 37214 56030 37266
rect 56082 37214 56094 37266
rect 52782 37202 52834 37214
rect 2494 37154 2546 37166
rect 2494 37090 2546 37102
rect 2942 37154 2994 37166
rect 12910 37154 12962 37166
rect 12562 37102 12574 37154
rect 12626 37102 12638 37154
rect 2942 37090 2994 37102
rect 12910 37090 12962 37102
rect 17502 37154 17554 37166
rect 35310 37154 35362 37166
rect 18050 37102 18062 37154
rect 18114 37102 18126 37154
rect 20178 37102 20190 37154
rect 20242 37102 20254 37154
rect 23986 37102 23998 37154
rect 24050 37102 24062 37154
rect 25554 37102 25566 37154
rect 25618 37102 25630 37154
rect 31826 37102 31838 37154
rect 31890 37102 31902 37154
rect 33842 37102 33854 37154
rect 33906 37102 33918 37154
rect 17502 37090 17554 37102
rect 35310 37090 35362 37102
rect 35758 37154 35810 37166
rect 35758 37090 35810 37102
rect 36094 37154 36146 37166
rect 36094 37090 36146 37102
rect 36542 37154 36594 37166
rect 36542 37090 36594 37102
rect 39342 37154 39394 37166
rect 39342 37090 39394 37102
rect 41022 37154 41074 37166
rect 41022 37090 41074 37102
rect 45390 37154 45442 37166
rect 52558 37154 52610 37166
rect 46834 37102 46846 37154
rect 46898 37102 46910 37154
rect 45390 37090 45442 37102
rect 52558 37090 52610 37102
rect 6414 37042 6466 37054
rect 6414 36978 6466 36990
rect 12238 37042 12290 37054
rect 12238 36978 12290 36990
rect 15710 37042 15762 37054
rect 55022 37042 55074 37054
rect 36082 36990 36094 37042
rect 36146 37039 36158 37042
rect 36418 37039 36430 37042
rect 36146 36993 36430 37039
rect 36146 36990 36158 36993
rect 36418 36990 36430 36993
rect 36482 37039 36494 37042
rect 36754 37039 36766 37042
rect 36482 36993 36766 37039
rect 36482 36990 36494 36993
rect 36754 36990 36766 36993
rect 36818 36990 36830 37042
rect 15710 36978 15762 36990
rect 55022 36978 55074 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 23102 36706 23154 36718
rect 23102 36642 23154 36654
rect 23550 36706 23602 36718
rect 23550 36642 23602 36654
rect 25566 36706 25618 36718
rect 25566 36642 25618 36654
rect 51326 36706 51378 36718
rect 51326 36642 51378 36654
rect 17838 36594 17890 36606
rect 20638 36594 20690 36606
rect 8418 36542 8430 36594
rect 8482 36542 8494 36594
rect 10546 36542 10558 36594
rect 10610 36542 10622 36594
rect 20066 36542 20078 36594
rect 20130 36542 20142 36594
rect 17838 36530 17890 36542
rect 20638 36530 20690 36542
rect 21422 36594 21474 36606
rect 21422 36530 21474 36542
rect 24782 36594 24834 36606
rect 24782 36530 24834 36542
rect 26238 36594 26290 36606
rect 26238 36530 26290 36542
rect 28478 36594 28530 36606
rect 28478 36530 28530 36542
rect 30942 36594 30994 36606
rect 30942 36530 30994 36542
rect 32734 36594 32786 36606
rect 37102 36594 37154 36606
rect 35074 36542 35086 36594
rect 35138 36542 35150 36594
rect 32734 36530 32786 36542
rect 37102 36530 37154 36542
rect 39790 36594 39842 36606
rect 39790 36530 39842 36542
rect 42590 36594 42642 36606
rect 42590 36530 42642 36542
rect 47070 36594 47122 36606
rect 47070 36530 47122 36542
rect 47854 36594 47906 36606
rect 47854 36530 47906 36542
rect 49534 36594 49586 36606
rect 49534 36530 49586 36542
rect 49982 36594 50034 36606
rect 49982 36530 50034 36542
rect 50430 36594 50482 36606
rect 50430 36530 50482 36542
rect 52782 36594 52834 36606
rect 54450 36542 54462 36594
rect 54514 36542 54526 36594
rect 56578 36542 56590 36594
rect 56642 36542 56654 36594
rect 52782 36530 52834 36542
rect 11790 36482 11842 36494
rect 13806 36482 13858 36494
rect 7746 36430 7758 36482
rect 7810 36430 7822 36482
rect 12674 36430 12686 36482
rect 12738 36430 12750 36482
rect 11790 36418 11842 36430
rect 13806 36418 13858 36430
rect 16718 36482 16770 36494
rect 19966 36482 20018 36494
rect 23102 36482 23154 36494
rect 17154 36430 17166 36482
rect 17218 36430 17230 36482
rect 19506 36430 19518 36482
rect 19570 36430 19582 36482
rect 20178 36430 20190 36482
rect 20242 36430 20254 36482
rect 22194 36430 22206 36482
rect 22258 36430 22270 36482
rect 16718 36418 16770 36430
rect 19966 36418 20018 36430
rect 23102 36418 23154 36430
rect 23774 36482 23826 36494
rect 28702 36482 28754 36494
rect 24322 36430 24334 36482
rect 24386 36430 24398 36482
rect 26450 36430 26462 36482
rect 26514 36430 26526 36482
rect 26786 36430 26798 36482
rect 26850 36430 26862 36482
rect 23774 36418 23826 36430
rect 28702 36418 28754 36430
rect 30382 36482 30434 36494
rect 30382 36418 30434 36430
rect 30830 36482 30882 36494
rect 34638 36482 34690 36494
rect 33282 36430 33294 36482
rect 33346 36430 33358 36482
rect 30830 36418 30882 36430
rect 34638 36418 34690 36430
rect 34750 36482 34802 36494
rect 34750 36418 34802 36430
rect 36094 36482 36146 36494
rect 40238 36482 40290 36494
rect 42702 36482 42754 36494
rect 39106 36430 39118 36482
rect 39170 36430 39182 36482
rect 39554 36430 39566 36482
rect 39618 36430 39630 36482
rect 41682 36430 41694 36482
rect 41746 36430 41758 36482
rect 42242 36430 42254 36482
rect 42306 36430 42318 36482
rect 36094 36418 36146 36430
rect 40238 36418 40290 36430
rect 42702 36418 42754 36430
rect 42814 36482 42866 36494
rect 42814 36418 42866 36430
rect 45278 36482 45330 36494
rect 45278 36418 45330 36430
rect 45502 36482 45554 36494
rect 45502 36418 45554 36430
rect 45726 36482 45778 36494
rect 47742 36482 47794 36494
rect 47506 36430 47518 36482
rect 47570 36430 47582 36482
rect 45726 36418 45778 36430
rect 47742 36418 47794 36430
rect 50654 36482 50706 36494
rect 51438 36482 51490 36494
rect 50978 36430 50990 36482
rect 51042 36430 51054 36482
rect 50654 36418 50706 36430
rect 51438 36418 51490 36430
rect 53118 36482 53170 36494
rect 53778 36430 53790 36482
rect 53842 36430 53854 36482
rect 53118 36418 53170 36430
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 2382 36370 2434 36382
rect 2382 36306 2434 36318
rect 2718 36370 2770 36382
rect 2718 36306 2770 36318
rect 3166 36370 3218 36382
rect 22654 36370 22706 36382
rect 12898 36318 12910 36370
rect 12962 36318 12974 36370
rect 16370 36318 16382 36370
rect 16434 36318 16446 36370
rect 17378 36318 17390 36370
rect 17442 36318 17454 36370
rect 3166 36306 3218 36318
rect 22654 36306 22706 36318
rect 22990 36370 23042 36382
rect 22990 36306 23042 36318
rect 25454 36370 25506 36382
rect 25454 36306 25506 36318
rect 27806 36370 27858 36382
rect 27806 36306 27858 36318
rect 28030 36370 28082 36382
rect 28030 36306 28082 36318
rect 28254 36370 28306 36382
rect 28254 36306 28306 36318
rect 30046 36370 30098 36382
rect 33966 36370 34018 36382
rect 33058 36318 33070 36370
rect 33122 36318 33134 36370
rect 30046 36306 30098 36318
rect 33966 36306 34018 36318
rect 34078 36370 34130 36382
rect 34078 36306 34130 36318
rect 34302 36370 34354 36382
rect 34302 36306 34354 36318
rect 35534 36370 35586 36382
rect 35534 36306 35586 36318
rect 35870 36370 35922 36382
rect 46734 36370 46786 36382
rect 41906 36318 41918 36370
rect 41970 36318 41982 36370
rect 35870 36306 35922 36318
rect 46734 36306 46786 36318
rect 48526 36370 48578 36382
rect 48526 36306 48578 36318
rect 48862 36370 48914 36382
rect 48862 36306 48914 36318
rect 49086 36370 49138 36382
rect 49086 36306 49138 36318
rect 51886 36370 51938 36382
rect 51886 36306 51938 36318
rect 52110 36370 52162 36382
rect 52110 36306 52162 36318
rect 52670 36370 52722 36382
rect 52670 36306 52722 36318
rect 53006 36370 53058 36382
rect 53006 36306 53058 36318
rect 2046 36258 2098 36270
rect 2046 36194 2098 36206
rect 11006 36258 11058 36270
rect 11006 36194 11058 36206
rect 12238 36258 12290 36270
rect 16046 36258 16098 36270
rect 13458 36206 13470 36258
rect 13522 36206 13534 36258
rect 12238 36194 12290 36206
rect 16046 36194 16098 36206
rect 19742 36258 19794 36270
rect 19742 36194 19794 36206
rect 25566 36258 25618 36270
rect 25566 36194 25618 36206
rect 29710 36258 29762 36270
rect 29710 36194 29762 36206
rect 30270 36258 30322 36270
rect 30270 36194 30322 36206
rect 30494 36258 30546 36270
rect 30494 36194 30546 36206
rect 31054 36258 31106 36270
rect 31054 36194 31106 36206
rect 31278 36258 31330 36270
rect 31278 36194 31330 36206
rect 31838 36258 31890 36270
rect 31838 36194 31890 36206
rect 34974 36258 35026 36270
rect 34974 36194 35026 36206
rect 35086 36258 35138 36270
rect 35086 36194 35138 36206
rect 35646 36258 35698 36270
rect 35646 36194 35698 36206
rect 40126 36258 40178 36270
rect 40126 36194 40178 36206
rect 40350 36258 40402 36270
rect 40350 36194 40402 36206
rect 40574 36258 40626 36270
rect 40574 36194 40626 36206
rect 41134 36258 41186 36270
rect 41134 36194 41186 36206
rect 42478 36258 42530 36270
rect 42478 36194 42530 36206
rect 43486 36258 43538 36270
rect 43486 36194 43538 36206
rect 44942 36258 44994 36270
rect 44942 36194 44994 36206
rect 46174 36258 46226 36270
rect 46174 36194 46226 36206
rect 46958 36258 47010 36270
rect 46958 36194 47010 36206
rect 47182 36258 47234 36270
rect 47182 36194 47234 36206
rect 47966 36258 48018 36270
rect 47966 36194 48018 36206
rect 48078 36258 48130 36270
rect 48078 36194 48130 36206
rect 48638 36258 48690 36270
rect 48638 36194 48690 36206
rect 51214 36258 51266 36270
rect 51214 36194 51266 36206
rect 51774 36258 51826 36270
rect 51774 36194 51826 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 13470 35922 13522 35934
rect 13470 35858 13522 35870
rect 15598 35922 15650 35934
rect 15598 35858 15650 35870
rect 18510 35922 18562 35934
rect 18510 35858 18562 35870
rect 18734 35922 18786 35934
rect 18734 35858 18786 35870
rect 23326 35922 23378 35934
rect 23326 35858 23378 35870
rect 23774 35922 23826 35934
rect 23774 35858 23826 35870
rect 24110 35922 24162 35934
rect 24110 35858 24162 35870
rect 24670 35922 24722 35934
rect 24670 35858 24722 35870
rect 26686 35922 26738 35934
rect 26686 35858 26738 35870
rect 28702 35922 28754 35934
rect 28702 35858 28754 35870
rect 30830 35922 30882 35934
rect 34526 35922 34578 35934
rect 32162 35870 32174 35922
rect 32226 35870 32238 35922
rect 30830 35858 30882 35870
rect 34526 35858 34578 35870
rect 39678 35922 39730 35934
rect 39678 35858 39730 35870
rect 39902 35922 39954 35934
rect 39902 35858 39954 35870
rect 40238 35922 40290 35934
rect 40238 35858 40290 35870
rect 41246 35922 41298 35934
rect 41246 35858 41298 35870
rect 41918 35922 41970 35934
rect 41918 35858 41970 35870
rect 51326 35922 51378 35934
rect 51326 35858 51378 35870
rect 51662 35922 51714 35934
rect 51662 35858 51714 35870
rect 52222 35922 52274 35934
rect 52222 35858 52274 35870
rect 52670 35922 52722 35934
rect 52670 35858 52722 35870
rect 25230 35810 25282 35822
rect 5842 35758 5854 35810
rect 5906 35758 5918 35810
rect 19058 35758 19070 35810
rect 19122 35758 19134 35810
rect 25230 35746 25282 35758
rect 27246 35810 27298 35822
rect 27246 35746 27298 35758
rect 30270 35810 30322 35822
rect 30270 35746 30322 35758
rect 30606 35810 30658 35822
rect 30606 35746 30658 35758
rect 31166 35810 31218 35822
rect 31166 35746 31218 35758
rect 31614 35810 31666 35822
rect 31614 35746 31666 35758
rect 33070 35810 33122 35822
rect 33070 35746 33122 35758
rect 33406 35810 33458 35822
rect 33406 35746 33458 35758
rect 34414 35810 34466 35822
rect 41470 35810 41522 35822
rect 35522 35758 35534 35810
rect 35586 35758 35598 35810
rect 34414 35746 34466 35758
rect 41470 35746 41522 35758
rect 42254 35810 42306 35822
rect 47854 35810 47906 35822
rect 43362 35758 43374 35810
rect 43426 35758 43438 35810
rect 42254 35746 42306 35758
rect 47854 35746 47906 35758
rect 47966 35810 48018 35822
rect 47966 35746 48018 35758
rect 48750 35810 48802 35822
rect 51550 35810 51602 35822
rect 50082 35758 50094 35810
rect 50146 35758 50158 35810
rect 48750 35746 48802 35758
rect 51550 35746 51602 35758
rect 52894 35810 52946 35822
rect 52894 35746 52946 35758
rect 14142 35698 14194 35710
rect 4274 35646 4286 35698
rect 4338 35646 4350 35698
rect 5170 35646 5182 35698
rect 5234 35646 5246 35698
rect 9538 35646 9550 35698
rect 9602 35646 9614 35698
rect 14142 35634 14194 35646
rect 14366 35698 14418 35710
rect 14366 35634 14418 35646
rect 14590 35698 14642 35710
rect 14590 35634 14642 35646
rect 23662 35698 23714 35710
rect 23662 35634 23714 35646
rect 23886 35698 23938 35710
rect 26126 35698 26178 35710
rect 25890 35646 25902 35698
rect 25954 35646 25966 35698
rect 23886 35634 23938 35646
rect 26126 35634 26178 35646
rect 26462 35698 26514 35710
rect 26462 35634 26514 35646
rect 26798 35698 26850 35710
rect 28142 35698 28194 35710
rect 27906 35646 27918 35698
rect 27970 35646 27982 35698
rect 26798 35634 26850 35646
rect 28142 35634 28194 35646
rect 28478 35698 28530 35710
rect 28478 35634 28530 35646
rect 28814 35698 28866 35710
rect 30830 35698 30882 35710
rect 29810 35646 29822 35698
rect 29874 35646 29886 35698
rect 30034 35646 30046 35698
rect 30098 35646 30110 35698
rect 28814 35634 28866 35646
rect 30830 35634 30882 35646
rect 32510 35698 32562 35710
rect 39566 35698 39618 35710
rect 33954 35646 33966 35698
rect 34018 35646 34030 35698
rect 34178 35646 34190 35698
rect 34242 35646 34254 35698
rect 34850 35646 34862 35698
rect 34914 35646 34926 35698
rect 32510 35634 32562 35646
rect 39566 35634 39618 35646
rect 41134 35698 41186 35710
rect 41134 35634 41186 35646
rect 41582 35698 41634 35710
rect 41582 35634 41634 35646
rect 42030 35698 42082 35710
rect 47182 35698 47234 35710
rect 42690 35646 42702 35698
rect 42754 35646 42766 35698
rect 42030 35634 42082 35646
rect 47182 35634 47234 35646
rect 48862 35698 48914 35710
rect 50990 35698 51042 35710
rect 49186 35646 49198 35698
rect 49250 35646 49262 35698
rect 50306 35646 50318 35698
rect 50370 35646 50382 35698
rect 48862 35634 48914 35646
rect 50990 35634 51042 35646
rect 51774 35698 51826 35710
rect 51774 35634 51826 35646
rect 52446 35698 52498 35710
rect 52446 35634 52498 35646
rect 53006 35698 53058 35710
rect 53442 35646 53454 35698
rect 53506 35646 53518 35698
rect 53006 35634 53058 35646
rect 8430 35586 8482 35598
rect 12910 35586 12962 35598
rect 7970 35534 7982 35586
rect 8034 35534 8046 35586
rect 10322 35534 10334 35586
rect 10386 35534 10398 35586
rect 12450 35534 12462 35586
rect 12514 35534 12526 35586
rect 8430 35522 8482 35534
rect 12910 35522 12962 35534
rect 14254 35586 14306 35598
rect 14254 35522 14306 35534
rect 15150 35586 15202 35598
rect 15150 35522 15202 35534
rect 16158 35586 16210 35598
rect 38110 35586 38162 35598
rect 45950 35586 46002 35598
rect 37650 35534 37662 35586
rect 37714 35534 37726 35586
rect 45490 35534 45502 35586
rect 45554 35534 45566 35586
rect 16158 35522 16210 35534
rect 38110 35522 38162 35534
rect 45950 35522 46002 35534
rect 46398 35586 46450 35598
rect 46398 35522 46450 35534
rect 46734 35586 46786 35598
rect 46734 35522 46786 35534
rect 52334 35586 52386 35598
rect 52334 35522 52386 35534
rect 1934 35474 1986 35486
rect 1934 35410 1986 35422
rect 16046 35474 16098 35486
rect 46958 35474 47010 35486
rect 45714 35422 45726 35474
rect 45778 35471 45790 35474
rect 46386 35471 46398 35474
rect 45778 35425 46398 35471
rect 45778 35422 45790 35425
rect 46386 35422 46398 35425
rect 46450 35422 46462 35474
rect 16046 35410 16098 35422
rect 46958 35410 47010 35422
rect 47630 35474 47682 35486
rect 47630 35410 47682 35422
rect 47966 35474 48018 35486
rect 55346 35422 55358 35474
rect 55410 35422 55422 35474
rect 47966 35410 48018 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 10894 35138 10946 35150
rect 10894 35074 10946 35086
rect 22990 35138 23042 35150
rect 22990 35074 23042 35086
rect 23438 35138 23490 35150
rect 23438 35074 23490 35086
rect 26798 35138 26850 35150
rect 26798 35074 26850 35086
rect 29038 35138 29090 35150
rect 29038 35074 29090 35086
rect 41806 35138 41858 35150
rect 41806 35074 41858 35086
rect 11006 35026 11058 35038
rect 25118 35026 25170 35038
rect 15810 34974 15822 35026
rect 15874 34974 15886 35026
rect 17938 34974 17950 35026
rect 18002 34974 18014 35026
rect 11006 34962 11058 34974
rect 25118 34962 25170 34974
rect 29934 35026 29986 35038
rect 29934 34962 29986 34974
rect 30382 35026 30434 35038
rect 32958 35026 33010 35038
rect 30930 34974 30942 35026
rect 30994 35023 31006 35026
rect 30994 34977 31215 35023
rect 30994 34974 31006 34977
rect 30382 34962 30434 34974
rect 23214 34914 23266 34926
rect 15138 34862 15150 34914
rect 15202 34862 15214 34914
rect 22194 34862 22206 34914
rect 22258 34862 22270 34914
rect 23214 34850 23266 34862
rect 24110 34914 24162 34926
rect 24110 34850 24162 34862
rect 26462 34914 26514 34926
rect 26462 34850 26514 34862
rect 28142 34914 28194 34926
rect 28142 34850 28194 34862
rect 29486 34914 29538 34926
rect 29486 34850 29538 34862
rect 29710 34914 29762 34926
rect 29710 34850 29762 34862
rect 30942 34914 30994 34926
rect 31169 34914 31215 34977
rect 32958 34962 33010 34974
rect 33630 35026 33682 35038
rect 33630 34962 33682 34974
rect 36094 35026 36146 35038
rect 36094 34962 36146 34974
rect 37102 35026 37154 35038
rect 37102 34962 37154 34974
rect 39678 35026 39730 35038
rect 39678 34962 39730 34974
rect 40910 35026 40962 35038
rect 40910 34962 40962 34974
rect 44942 35026 44994 35038
rect 52670 35026 52722 35038
rect 48178 34974 48190 35026
rect 48242 34974 48254 35026
rect 44942 34962 44994 34974
rect 52670 34962 52722 34974
rect 54126 35026 54178 35038
rect 54126 34962 54178 34974
rect 57934 35026 57986 35038
rect 57934 34962 57986 34974
rect 31726 34914 31778 34926
rect 31154 34862 31166 34914
rect 31218 34862 31230 34914
rect 30942 34850 30994 34862
rect 31726 34850 31778 34862
rect 32062 34914 32114 34926
rect 34638 34914 34690 34926
rect 32274 34862 32286 34914
rect 32338 34862 32350 34914
rect 32062 34850 32114 34862
rect 34638 34850 34690 34862
rect 35198 34914 35250 34926
rect 39230 34914 39282 34926
rect 35634 34862 35646 34914
rect 35698 34862 35710 34914
rect 35198 34850 35250 34862
rect 39230 34850 39282 34862
rect 39454 34914 39506 34926
rect 41134 34914 41186 34926
rect 42254 34914 42306 34926
rect 40114 34862 40126 34914
rect 40178 34862 40190 34914
rect 41458 34862 41470 34914
rect 41522 34862 41534 34914
rect 39454 34850 39506 34862
rect 41134 34850 41186 34862
rect 42254 34850 42306 34862
rect 42702 34914 42754 34926
rect 42702 34850 42754 34862
rect 42926 34914 42978 34926
rect 42926 34850 42978 34862
rect 43486 34914 43538 34926
rect 50654 34914 50706 34926
rect 46946 34862 46958 34914
rect 47010 34862 47022 34914
rect 43486 34850 43538 34862
rect 50654 34850 50706 34862
rect 50990 34914 51042 34926
rect 50990 34850 51042 34862
rect 51326 34914 51378 34926
rect 51326 34850 51378 34862
rect 51662 34914 51714 34926
rect 51662 34850 51714 34862
rect 51774 34914 51826 34926
rect 52782 34914 52834 34926
rect 52098 34862 52110 34914
rect 52162 34862 52174 34914
rect 53330 34862 53342 34914
rect 53394 34862 53406 34914
rect 55570 34862 55582 34914
rect 55634 34862 55646 34914
rect 51774 34850 51826 34862
rect 52782 34850 52834 34862
rect 5854 34802 5906 34814
rect 5854 34738 5906 34750
rect 14254 34802 14306 34814
rect 14254 34738 14306 34750
rect 21646 34802 21698 34814
rect 21646 34738 21698 34750
rect 22766 34802 22818 34814
rect 22766 34738 22818 34750
rect 23886 34802 23938 34814
rect 23886 34738 23938 34750
rect 26238 34802 26290 34814
rect 26238 34738 26290 34750
rect 31390 34802 31442 34814
rect 31390 34738 31442 34750
rect 31502 34802 31554 34814
rect 31502 34738 31554 34750
rect 38558 34802 38610 34814
rect 38558 34738 38610 34750
rect 49982 34802 50034 34814
rect 49982 34738 50034 34750
rect 5518 34690 5570 34702
rect 5518 34626 5570 34638
rect 5742 34690 5794 34702
rect 5742 34626 5794 34638
rect 14142 34690 14194 34702
rect 14142 34626 14194 34638
rect 14702 34690 14754 34702
rect 14702 34626 14754 34638
rect 21310 34690 21362 34702
rect 21310 34626 21362 34638
rect 22430 34690 22482 34702
rect 25902 34690 25954 34702
rect 24434 34638 24446 34690
rect 24498 34638 24510 34690
rect 22430 34626 22482 34638
rect 25902 34626 25954 34638
rect 27246 34690 27298 34702
rect 27246 34626 27298 34638
rect 27694 34690 27746 34702
rect 27694 34626 27746 34638
rect 30270 34690 30322 34702
rect 30270 34626 30322 34638
rect 30494 34690 30546 34702
rect 30494 34626 30546 34638
rect 34302 34690 34354 34702
rect 34302 34626 34354 34638
rect 34526 34690 34578 34702
rect 34526 34626 34578 34638
rect 34750 34690 34802 34702
rect 34750 34626 34802 34638
rect 37662 34690 37714 34702
rect 37662 34626 37714 34638
rect 38222 34690 38274 34702
rect 38222 34626 38274 34638
rect 38782 34690 38834 34702
rect 41694 34690 41746 34702
rect 40338 34638 40350 34690
rect 40402 34638 40414 34690
rect 38782 34626 38834 34638
rect 41694 34626 41746 34638
rect 42030 34690 42082 34702
rect 42030 34626 42082 34638
rect 42142 34690 42194 34702
rect 42142 34626 42194 34638
rect 44046 34690 44098 34702
rect 44046 34626 44098 34638
rect 45950 34690 46002 34702
rect 46622 34690 46674 34702
rect 46274 34638 46286 34690
rect 46338 34638 46350 34690
rect 45950 34626 46002 34638
rect 46622 34626 46674 34638
rect 49870 34690 49922 34702
rect 49870 34626 49922 34638
rect 50542 34690 50594 34702
rect 50542 34626 50594 34638
rect 51102 34690 51154 34702
rect 51102 34626 51154 34638
rect 51550 34690 51602 34702
rect 51550 34626 51602 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 7982 34354 8034 34366
rect 7982 34290 8034 34302
rect 12238 34354 12290 34366
rect 12238 34290 12290 34302
rect 16270 34354 16322 34366
rect 16270 34290 16322 34302
rect 16494 34354 16546 34366
rect 16494 34290 16546 34302
rect 18398 34354 18450 34366
rect 18398 34290 18450 34302
rect 22878 34354 22930 34366
rect 22878 34290 22930 34302
rect 24782 34354 24834 34366
rect 24782 34290 24834 34302
rect 25230 34354 25282 34366
rect 25230 34290 25282 34302
rect 31166 34354 31218 34366
rect 46958 34354 47010 34366
rect 37090 34302 37102 34354
rect 37154 34302 37166 34354
rect 43250 34302 43262 34354
rect 43314 34302 43326 34354
rect 31166 34290 31218 34302
rect 46958 34290 47010 34302
rect 48078 34354 48130 34366
rect 48078 34290 48130 34302
rect 48302 34354 48354 34366
rect 48302 34290 48354 34302
rect 48862 34354 48914 34366
rect 48862 34290 48914 34302
rect 50206 34354 50258 34366
rect 50206 34290 50258 34302
rect 51326 34354 51378 34366
rect 51326 34290 51378 34302
rect 8542 34242 8594 34254
rect 16158 34242 16210 34254
rect 42590 34242 42642 34254
rect 47182 34242 47234 34254
rect 10546 34190 10558 34242
rect 10610 34190 10622 34242
rect 13346 34190 13358 34242
rect 13410 34190 13422 34242
rect 20178 34190 20190 34242
rect 20242 34190 20254 34242
rect 23538 34190 23550 34242
rect 23602 34190 23614 34242
rect 23762 34190 23774 34242
rect 23826 34190 23838 34242
rect 25554 34190 25566 34242
rect 25618 34190 25630 34242
rect 29922 34190 29934 34242
rect 29986 34190 29998 34242
rect 38210 34190 38222 34242
rect 38274 34190 38286 34242
rect 45378 34190 45390 34242
rect 45442 34190 45454 34242
rect 45826 34190 45838 34242
rect 45890 34190 45902 34242
rect 8542 34178 8594 34190
rect 16158 34178 16210 34190
rect 42590 34178 42642 34190
rect 47182 34178 47234 34190
rect 47630 34242 47682 34254
rect 47630 34178 47682 34190
rect 47966 34242 48018 34254
rect 47966 34178 48018 34190
rect 48750 34242 48802 34254
rect 48750 34178 48802 34190
rect 52782 34242 52834 34254
rect 52782 34178 52834 34190
rect 4286 34130 4338 34142
rect 8318 34130 8370 34142
rect 4722 34078 4734 34130
rect 4786 34078 4798 34130
rect 4286 34066 4338 34078
rect 8318 34066 8370 34078
rect 8654 34130 8706 34142
rect 8654 34066 8706 34078
rect 10222 34130 10274 34142
rect 16382 34130 16434 34142
rect 12674 34078 12686 34130
rect 12738 34078 12750 34130
rect 15922 34078 15934 34130
rect 15986 34078 15998 34130
rect 10222 34066 10274 34078
rect 16382 34066 16434 34078
rect 18286 34130 18338 34142
rect 18286 34066 18338 34078
rect 18622 34130 18674 34142
rect 29598 34130 29650 34142
rect 18834 34078 18846 34130
rect 18898 34078 18910 34130
rect 19506 34078 19518 34130
rect 19570 34078 19582 34130
rect 18622 34066 18674 34078
rect 29598 34066 29650 34078
rect 35534 34130 35586 34142
rect 35534 34066 35586 34078
rect 35982 34130 36034 34142
rect 35982 34066 36034 34078
rect 36206 34130 36258 34142
rect 48974 34130 49026 34142
rect 37538 34078 37550 34130
rect 37602 34078 37614 34130
rect 42018 34078 42030 34130
rect 42082 34078 42094 34130
rect 43026 34078 43038 34130
rect 43090 34078 43102 34130
rect 47394 34078 47406 34130
rect 47458 34078 47470 34130
rect 36206 34066 36258 34078
rect 48974 34066 49026 34078
rect 49422 34130 49474 34142
rect 49422 34066 49474 34078
rect 50654 34130 50706 34142
rect 50654 34066 50706 34078
rect 50878 34130 50930 34142
rect 50878 34066 50930 34078
rect 51998 34130 52050 34142
rect 51998 34066 52050 34078
rect 52894 34130 52946 34142
rect 53218 34078 53230 34130
rect 53282 34078 53294 34130
rect 52894 34066 52946 34078
rect 1822 34018 1874 34030
rect 11006 34018 11058 34030
rect 17726 34018 17778 34030
rect 5394 33966 5406 34018
rect 5458 33966 5470 34018
rect 7522 33966 7534 34018
rect 7586 33966 7598 34018
rect 15474 33966 15486 34018
rect 15538 33966 15550 34018
rect 1822 33954 1874 33966
rect 11006 33954 11058 33966
rect 17726 33954 17778 33966
rect 18510 34018 18562 34030
rect 26462 34018 26514 34030
rect 22306 33966 22318 34018
rect 22370 33966 22382 34018
rect 18510 33954 18562 33966
rect 26462 33954 26514 33966
rect 31614 34018 31666 34030
rect 31614 33954 31666 33966
rect 33742 34018 33794 34030
rect 33742 33954 33794 33966
rect 34190 34018 34242 34030
rect 34190 33954 34242 33966
rect 34750 34018 34802 34030
rect 34750 33954 34802 33966
rect 36094 34018 36146 34030
rect 36094 33954 36146 33966
rect 36542 34018 36594 34030
rect 43710 34018 43762 34030
rect 40338 33966 40350 34018
rect 40402 33966 40414 34018
rect 42130 33966 42142 34018
rect 42194 33966 42206 34018
rect 36542 33954 36594 33966
rect 43710 33954 43762 33966
rect 47518 34018 47570 34030
rect 47518 33954 47570 33966
rect 49870 34018 49922 34030
rect 49870 33954 49922 33966
rect 51102 34018 51154 34030
rect 51102 33954 51154 33966
rect 52222 34018 52274 34030
rect 52222 33954 52274 33966
rect 17838 33906 17890 33918
rect 17838 33842 17890 33854
rect 23214 33906 23266 33918
rect 23214 33842 23266 33854
rect 34974 33906 35026 33918
rect 34974 33842 35026 33854
rect 35310 33906 35362 33918
rect 35310 33842 35362 33854
rect 36766 33906 36818 33918
rect 36766 33842 36818 33854
rect 44830 33906 44882 33918
rect 44830 33842 44882 33854
rect 45166 33906 45218 33918
rect 45166 33842 45218 33854
rect 51774 33906 51826 33918
rect 51774 33842 51826 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 34302 33570 34354 33582
rect 5506 33518 5518 33570
rect 5570 33567 5582 33570
rect 5842 33567 5854 33570
rect 5570 33521 5854 33567
rect 5570 33518 5582 33521
rect 5842 33518 5854 33521
rect 5906 33518 5918 33570
rect 34302 33506 34354 33518
rect 38558 33570 38610 33582
rect 52782 33570 52834 33582
rect 42690 33518 42702 33570
rect 42754 33567 42766 33570
rect 43026 33567 43038 33570
rect 42754 33521 43038 33567
rect 42754 33518 42766 33521
rect 43026 33518 43038 33521
rect 43090 33518 43102 33570
rect 38558 33506 38610 33518
rect 52782 33506 52834 33518
rect 57934 33570 57986 33582
rect 57934 33506 57986 33518
rect 6190 33458 6242 33470
rect 10894 33458 10946 33470
rect 15934 33458 15986 33470
rect 4722 33406 4734 33458
rect 4786 33406 4798 33458
rect 10434 33406 10446 33458
rect 10498 33406 10510 33458
rect 15474 33406 15486 33458
rect 15538 33406 15550 33458
rect 6190 33394 6242 33406
rect 10894 33394 10946 33406
rect 15934 33394 15986 33406
rect 16606 33458 16658 33470
rect 24110 33458 24162 33470
rect 35758 33458 35810 33470
rect 18162 33406 18174 33458
rect 18226 33406 18238 33458
rect 20290 33406 20302 33458
rect 20354 33406 20366 33458
rect 27794 33406 27806 33458
rect 27858 33406 27870 33458
rect 29138 33406 29150 33458
rect 29202 33406 29214 33458
rect 34850 33406 34862 33458
rect 34914 33406 34926 33458
rect 16606 33394 16658 33406
rect 24110 33394 24162 33406
rect 35758 33394 35810 33406
rect 37662 33458 37714 33470
rect 37662 33394 37714 33406
rect 42702 33458 42754 33470
rect 51438 33458 51490 33470
rect 47730 33406 47742 33458
rect 47794 33406 47806 33458
rect 50978 33406 50990 33458
rect 51042 33406 51054 33458
rect 42702 33394 42754 33406
rect 51438 33394 51490 33406
rect 6862 33346 6914 33358
rect 1922 33294 1934 33346
rect 1986 33294 1998 33346
rect 6626 33294 6638 33346
rect 6690 33294 6702 33346
rect 6862 33282 6914 33294
rect 7198 33346 7250 33358
rect 11566 33346 11618 33358
rect 7634 33294 7646 33346
rect 7698 33294 7710 33346
rect 7198 33282 7250 33294
rect 11566 33282 11618 33294
rect 12350 33346 12402 33358
rect 12350 33282 12402 33294
rect 12910 33346 12962 33358
rect 12910 33282 12962 33294
rect 15374 33346 15426 33358
rect 15374 33282 15426 33294
rect 17054 33346 17106 33358
rect 22990 33346 23042 33358
rect 38894 33346 38946 33358
rect 43038 33346 43090 33358
rect 52670 33346 52722 33358
rect 17378 33294 17390 33346
rect 17442 33294 17454 33346
rect 21858 33294 21870 33346
rect 21922 33294 21934 33346
rect 22306 33294 22318 33346
rect 22370 33294 22382 33346
rect 24882 33294 24894 33346
rect 24946 33294 24958 33346
rect 32050 33294 32062 33346
rect 32114 33294 32126 33346
rect 35298 33294 35310 33346
rect 35362 33294 35374 33346
rect 39442 33294 39454 33346
rect 39506 33294 39518 33346
rect 44034 33294 44046 33346
rect 44098 33294 44110 33346
rect 44930 33294 44942 33346
rect 44994 33294 45006 33346
rect 48178 33294 48190 33346
rect 48242 33294 48254 33346
rect 55570 33294 55582 33346
rect 55634 33294 55646 33346
rect 17054 33282 17106 33294
rect 22990 33282 23042 33294
rect 38894 33282 38946 33294
rect 43038 33282 43090 33294
rect 52670 33282 52722 33294
rect 14254 33234 14306 33246
rect 2594 33182 2606 33234
rect 2658 33182 2670 33234
rect 8306 33182 8318 33234
rect 8370 33182 8382 33234
rect 14254 33170 14306 33182
rect 14926 33234 14978 33246
rect 14926 33170 14978 33182
rect 15486 33234 15538 33246
rect 15486 33170 15538 33182
rect 22542 33234 22594 33246
rect 22542 33170 22594 33182
rect 24446 33234 24498 33246
rect 24446 33170 24498 33182
rect 24558 33234 24610 33246
rect 28478 33234 28530 33246
rect 25666 33182 25678 33234
rect 25730 33182 25742 33234
rect 24558 33170 24610 33182
rect 28478 33170 28530 33182
rect 28590 33234 28642 33246
rect 32510 33234 32562 33246
rect 31266 33182 31278 33234
rect 31330 33182 31342 33234
rect 28590 33170 28642 33182
rect 32510 33170 32562 33182
rect 34414 33234 34466 33246
rect 34414 33170 34466 33182
rect 36094 33234 36146 33246
rect 36094 33170 36146 33182
rect 36430 33234 36482 33246
rect 44270 33234 44322 33246
rect 51326 33234 51378 33246
rect 39666 33182 39678 33234
rect 39730 33182 39742 33234
rect 45602 33182 45614 33234
rect 45666 33182 45678 33234
rect 48850 33182 48862 33234
rect 48914 33182 48926 33234
rect 36430 33170 36482 33182
rect 44270 33170 44322 33182
rect 51326 33170 51378 33182
rect 54462 33234 54514 33246
rect 54462 33170 54514 33182
rect 5854 33122 5906 33134
rect 5854 33058 5906 33070
rect 6078 33122 6130 33134
rect 6078 33058 6130 33070
rect 6302 33122 6354 33134
rect 6302 33058 6354 33070
rect 7086 33122 7138 33134
rect 7086 33058 7138 33070
rect 11678 33122 11730 33134
rect 11678 33058 11730 33070
rect 11902 33122 11954 33134
rect 13806 33122 13858 33134
rect 13458 33070 13470 33122
rect 13522 33070 13534 33122
rect 11902 33058 11954 33070
rect 13806 33058 13858 33070
rect 15150 33122 15202 33134
rect 15150 33058 15202 33070
rect 16046 33122 16098 33134
rect 16046 33058 16098 33070
rect 32398 33122 32450 33134
rect 32398 33058 32450 33070
rect 32958 33122 33010 33134
rect 32958 33058 33010 33070
rect 33854 33122 33906 33134
rect 33854 33058 33906 33070
rect 34302 33122 34354 33134
rect 34302 33058 34354 33070
rect 37102 33122 37154 33134
rect 37102 33058 37154 33070
rect 37998 33122 38050 33134
rect 37998 33058 38050 33070
rect 51886 33122 51938 33134
rect 51886 33058 51938 33070
rect 53230 33122 53282 33134
rect 53230 33058 53282 33070
rect 54574 33122 54626 33134
rect 54574 33058 54626 33070
rect 55358 33122 55410 33134
rect 55358 33058 55410 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 8094 32786 8146 32798
rect 8094 32722 8146 32734
rect 8430 32786 8482 32798
rect 8430 32722 8482 32734
rect 14366 32786 14418 32798
rect 14366 32722 14418 32734
rect 15822 32786 15874 32798
rect 15822 32722 15874 32734
rect 16494 32786 16546 32798
rect 16494 32722 16546 32734
rect 16830 32786 16882 32798
rect 25566 32786 25618 32798
rect 20850 32734 20862 32786
rect 20914 32734 20926 32786
rect 16830 32722 16882 32734
rect 25566 32722 25618 32734
rect 25678 32786 25730 32798
rect 25678 32722 25730 32734
rect 29822 32786 29874 32798
rect 29822 32722 29874 32734
rect 31726 32786 31778 32798
rect 31726 32722 31778 32734
rect 38894 32786 38946 32798
rect 38894 32722 38946 32734
rect 39342 32786 39394 32798
rect 39342 32722 39394 32734
rect 50542 32786 50594 32798
rect 52546 32734 52558 32786
rect 52610 32734 52622 32786
rect 50542 32722 50594 32734
rect 9774 32674 9826 32686
rect 5394 32622 5406 32674
rect 5458 32622 5470 32674
rect 6850 32622 6862 32674
rect 6914 32622 6926 32674
rect 9774 32610 9826 32622
rect 15710 32674 15762 32686
rect 15710 32610 15762 32622
rect 25230 32674 25282 32686
rect 25230 32610 25282 32622
rect 26462 32674 26514 32686
rect 26462 32610 26514 32622
rect 29486 32674 29538 32686
rect 29486 32610 29538 32622
rect 30046 32674 30098 32686
rect 30046 32610 30098 32622
rect 51774 32674 51826 32686
rect 55234 32622 55246 32674
rect 55298 32622 55310 32674
rect 51774 32610 51826 32622
rect 8318 32562 8370 32574
rect 1810 32510 1822 32562
rect 1874 32510 1886 32562
rect 5282 32510 5294 32562
rect 5346 32510 5358 32562
rect 6962 32510 6974 32562
rect 7026 32510 7038 32562
rect 8318 32498 8370 32510
rect 8542 32562 8594 32574
rect 8542 32498 8594 32510
rect 9550 32562 9602 32574
rect 9550 32498 9602 32510
rect 9998 32562 10050 32574
rect 9998 32498 10050 32510
rect 10222 32562 10274 32574
rect 14702 32562 14754 32574
rect 10546 32510 10558 32562
rect 10610 32510 10622 32562
rect 10222 32498 10274 32510
rect 14702 32498 14754 32510
rect 15038 32562 15090 32574
rect 15038 32498 15090 32510
rect 15374 32562 15426 32574
rect 25454 32562 25506 32574
rect 26798 32562 26850 32574
rect 19730 32510 19742 32562
rect 19794 32510 19806 32562
rect 21074 32510 21086 32562
rect 21138 32510 21150 32562
rect 25890 32510 25902 32562
rect 25954 32510 25966 32562
rect 15374 32498 15426 32510
rect 25454 32498 25506 32510
rect 26798 32498 26850 32510
rect 29710 32562 29762 32574
rect 29710 32498 29762 32510
rect 29934 32562 29986 32574
rect 31614 32562 31666 32574
rect 31378 32510 31390 32562
rect 31442 32510 31454 32562
rect 29934 32498 29986 32510
rect 31614 32498 31666 32510
rect 31838 32562 31890 32574
rect 31838 32498 31890 32510
rect 31950 32562 32002 32574
rect 31950 32498 32002 32510
rect 34750 32562 34802 32574
rect 34750 32498 34802 32510
rect 35310 32562 35362 32574
rect 36206 32562 36258 32574
rect 35970 32510 35982 32562
rect 36034 32510 36046 32562
rect 35310 32498 35362 32510
rect 36206 32498 36258 32510
rect 38782 32562 38834 32574
rect 45054 32562 45106 32574
rect 41682 32510 41694 32562
rect 41746 32510 41758 32562
rect 38782 32498 38834 32510
rect 45054 32498 45106 32510
rect 47966 32562 48018 32574
rect 47966 32498 48018 32510
rect 51886 32562 51938 32574
rect 51886 32498 51938 32510
rect 52222 32562 52274 32574
rect 55906 32510 55918 32562
rect 55970 32510 55982 32562
rect 52222 32498 52274 32510
rect 7646 32450 7698 32462
rect 2482 32398 2494 32450
rect 2546 32398 2558 32450
rect 4610 32398 4622 32450
rect 4674 32398 4686 32450
rect 5842 32398 5854 32450
rect 5906 32398 5918 32450
rect 7646 32386 7698 32398
rect 9102 32450 9154 32462
rect 13918 32450 13970 32462
rect 11218 32398 11230 32450
rect 11282 32398 11294 32450
rect 13346 32398 13358 32450
rect 13410 32398 13422 32450
rect 9102 32386 9154 32398
rect 13918 32386 13970 32398
rect 14926 32450 14978 32462
rect 14926 32386 14978 32398
rect 27246 32450 27298 32462
rect 27246 32386 27298 32398
rect 29150 32450 29202 32462
rect 29150 32386 29202 32398
rect 31054 32450 31106 32462
rect 31054 32386 31106 32398
rect 33966 32450 34018 32462
rect 33966 32386 34018 32398
rect 36766 32450 36818 32462
rect 36766 32386 36818 32398
rect 37214 32450 37266 32462
rect 37214 32386 37266 32398
rect 39454 32450 39506 32462
rect 42466 32398 42478 32450
rect 42530 32398 42542 32450
rect 44594 32398 44606 32450
rect 44658 32398 44670 32450
rect 53106 32398 53118 32450
rect 53170 32398 53182 32450
rect 39454 32386 39506 32398
rect 14142 32338 14194 32350
rect 14142 32274 14194 32286
rect 14478 32338 14530 32350
rect 14478 32274 14530 32286
rect 15822 32338 15874 32350
rect 15822 32274 15874 32286
rect 19742 32338 19794 32350
rect 19742 32274 19794 32286
rect 20078 32338 20130 32350
rect 38894 32338 38946 32350
rect 34626 32286 34638 32338
rect 34690 32335 34702 32338
rect 35074 32335 35086 32338
rect 34690 32289 35086 32335
rect 34690 32286 34702 32289
rect 35074 32286 35086 32289
rect 35138 32286 35150 32338
rect 20078 32274 20130 32286
rect 38894 32274 38946 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 15150 32002 15202 32014
rect 15150 31938 15202 31950
rect 42142 32002 42194 32014
rect 42142 31938 42194 31950
rect 51886 32002 51938 32014
rect 51886 31938 51938 31950
rect 2830 31890 2882 31902
rect 2830 31826 2882 31838
rect 6078 31890 6130 31902
rect 6078 31826 6130 31838
rect 7646 31890 7698 31902
rect 11230 31890 11282 31902
rect 8866 31838 8878 31890
rect 8930 31838 8942 31890
rect 9426 31838 9438 31890
rect 9490 31838 9502 31890
rect 7646 31826 7698 31838
rect 11230 31826 11282 31838
rect 12910 31890 12962 31902
rect 12910 31826 12962 31838
rect 15822 31890 15874 31902
rect 15822 31826 15874 31838
rect 22542 31890 22594 31902
rect 22542 31826 22594 31838
rect 23998 31890 24050 31902
rect 23998 31826 24050 31838
rect 25454 31890 25506 31902
rect 29710 31890 29762 31902
rect 40686 31890 40738 31902
rect 42030 31890 42082 31902
rect 51550 31890 51602 31902
rect 26450 31838 26462 31890
rect 26514 31838 26526 31890
rect 28578 31838 28590 31890
rect 28642 31838 28654 31890
rect 38994 31838 39006 31890
rect 39058 31838 39070 31890
rect 41570 31838 41582 31890
rect 41634 31838 41646 31890
rect 43586 31838 43598 31890
rect 43650 31838 43662 31890
rect 50306 31838 50318 31890
rect 50370 31838 50382 31890
rect 54338 31838 54350 31890
rect 54402 31838 54414 31890
rect 25454 31826 25506 31838
rect 29710 31826 29762 31838
rect 40686 31826 40738 31838
rect 42030 31826 42082 31838
rect 51550 31826 51602 31838
rect 1710 31778 1762 31790
rect 1710 31714 1762 31726
rect 4622 31778 4674 31790
rect 4622 31714 4674 31726
rect 4846 31778 4898 31790
rect 4846 31714 4898 31726
rect 6190 31778 6242 31790
rect 6190 31714 6242 31726
rect 6526 31778 6578 31790
rect 14590 31778 14642 31790
rect 8530 31726 8542 31778
rect 8594 31726 8606 31778
rect 11666 31726 11678 31778
rect 11730 31726 11742 31778
rect 14130 31726 14142 31778
rect 14194 31726 14206 31778
rect 6526 31714 6578 31726
rect 14590 31714 14642 31726
rect 15598 31778 15650 31790
rect 15598 31714 15650 31726
rect 16270 31778 16322 31790
rect 16270 31714 16322 31726
rect 19182 31778 19234 31790
rect 19182 31714 19234 31726
rect 19630 31778 19682 31790
rect 22654 31778 22706 31790
rect 19842 31726 19854 31778
rect 19906 31726 19918 31778
rect 19630 31714 19682 31726
rect 22654 31714 22706 31726
rect 23214 31778 23266 31790
rect 29486 31778 29538 31790
rect 41246 31778 41298 31790
rect 24210 31726 24222 31778
rect 24274 31726 24286 31778
rect 25666 31726 25678 31778
rect 25730 31726 25742 31778
rect 30146 31726 30158 31778
rect 30210 31726 30222 31778
rect 38546 31726 38558 31778
rect 38610 31726 38622 31778
rect 39890 31726 39902 31778
rect 39954 31726 39966 31778
rect 23214 31714 23266 31726
rect 29486 31714 29538 31726
rect 41246 31714 41298 31726
rect 41470 31778 41522 31790
rect 50878 31778 50930 31790
rect 47506 31726 47518 31778
rect 47570 31726 47582 31778
rect 41470 31714 41522 31726
rect 50878 31714 50930 31726
rect 52558 31778 52610 31790
rect 52558 31714 52610 31726
rect 53230 31778 53282 31790
rect 53778 31726 53790 31778
rect 53842 31726 53854 31778
rect 55010 31726 55022 31778
rect 55074 31726 55086 31778
rect 53230 31714 53282 31726
rect 2942 31666 2994 31678
rect 2942 31602 2994 31614
rect 3614 31666 3666 31678
rect 3614 31602 3666 31614
rect 3838 31666 3890 31678
rect 3838 31602 3890 31614
rect 4062 31666 4114 31678
rect 4062 31602 4114 31614
rect 4510 31666 4562 31678
rect 4510 31602 4562 31614
rect 5070 31666 5122 31678
rect 5070 31602 5122 31614
rect 5966 31666 6018 31678
rect 5966 31602 6018 31614
rect 7758 31666 7810 31678
rect 7758 31602 7810 31614
rect 8094 31666 8146 31678
rect 8094 31602 8146 31614
rect 9774 31666 9826 31678
rect 9774 31602 9826 31614
rect 10110 31666 10162 31678
rect 10110 31602 10162 31614
rect 10334 31666 10386 31678
rect 10334 31602 10386 31614
rect 11342 31666 11394 31678
rect 11342 31602 11394 31614
rect 14702 31666 14754 31678
rect 14702 31602 14754 31614
rect 15038 31666 15090 31678
rect 15038 31602 15090 31614
rect 15262 31666 15314 31678
rect 15262 31602 15314 31614
rect 16606 31666 16658 31678
rect 16606 31602 16658 31614
rect 16830 31666 16882 31678
rect 16830 31602 16882 31614
rect 17054 31666 17106 31678
rect 17054 31602 17106 31614
rect 17390 31666 17442 31678
rect 17390 31602 17442 31614
rect 18622 31666 18674 31678
rect 18622 31602 18674 31614
rect 18734 31666 18786 31678
rect 18734 31602 18786 31614
rect 18958 31666 19010 31678
rect 18958 31602 19010 31614
rect 20526 31666 20578 31678
rect 20526 31602 20578 31614
rect 22990 31666 23042 31678
rect 22990 31602 23042 31614
rect 23550 31666 23602 31678
rect 23550 31602 23602 31614
rect 23886 31666 23938 31678
rect 23886 31602 23938 31614
rect 24782 31666 24834 31678
rect 38110 31666 38162 31678
rect 41022 31666 41074 31678
rect 52110 31666 52162 31678
rect 32162 31614 32174 31666
rect 32226 31614 32238 31666
rect 39666 31614 39678 31666
rect 39730 31614 39742 31666
rect 48178 31614 48190 31666
rect 48242 31614 48254 31666
rect 24782 31602 24834 31614
rect 38110 31602 38162 31614
rect 41022 31602 41074 31614
rect 52110 31602 52162 31614
rect 2718 31554 2770 31566
rect 2034 31502 2046 31554
rect 2098 31502 2110 31554
rect 2718 31490 2770 31502
rect 3166 31554 3218 31566
rect 3166 31490 3218 31502
rect 3726 31554 3778 31566
rect 3726 31490 3778 31502
rect 7198 31554 7250 31566
rect 7198 31490 7250 31502
rect 7534 31554 7586 31566
rect 7534 31490 7586 31502
rect 9550 31554 9602 31566
rect 9550 31490 9602 31502
rect 10222 31554 10274 31566
rect 10222 31490 10274 31502
rect 11118 31554 11170 31566
rect 11118 31490 11170 31502
rect 12126 31554 12178 31566
rect 12126 31490 12178 31502
rect 16382 31554 16434 31566
rect 16382 31490 16434 31502
rect 17166 31554 17218 31566
rect 17166 31490 17218 31502
rect 17726 31554 17778 31566
rect 23214 31554 23266 31566
rect 18050 31502 18062 31554
rect 18114 31502 18126 31554
rect 17726 31490 17778 31502
rect 23214 31490 23266 31502
rect 24446 31554 24498 31566
rect 24446 31490 24498 31502
rect 24670 31554 24722 31566
rect 24670 31490 24722 31502
rect 29822 31554 29874 31566
rect 29822 31490 29874 31502
rect 36206 31554 36258 31566
rect 36206 31490 36258 31502
rect 41582 31554 41634 31566
rect 41582 31490 41634 31502
rect 42702 31554 42754 31566
rect 42702 31490 42754 31502
rect 43150 31554 43202 31566
rect 43150 31490 43202 31502
rect 44158 31554 44210 31566
rect 44158 31490 44210 31502
rect 50990 31554 51042 31566
rect 50990 31490 51042 31502
rect 53006 31554 53058 31566
rect 53006 31490 53058 31502
rect 53118 31554 53170 31566
rect 53118 31490 53170 31502
rect 54014 31554 54066 31566
rect 54014 31490 54066 31502
rect 54238 31554 54290 31566
rect 54238 31490 54290 31502
rect 54350 31554 54402 31566
rect 55694 31554 55746 31566
rect 54786 31502 54798 31554
rect 54850 31502 54862 31554
rect 54350 31490 54402 31502
rect 55694 31490 55746 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 4734 31218 4786 31230
rect 4734 31154 4786 31166
rect 4958 31218 5010 31230
rect 4958 31154 5010 31166
rect 5630 31218 5682 31230
rect 5630 31154 5682 31166
rect 5966 31218 6018 31230
rect 5966 31154 6018 31166
rect 12574 31218 12626 31230
rect 12574 31154 12626 31166
rect 14926 31218 14978 31230
rect 14926 31154 14978 31166
rect 18846 31218 18898 31230
rect 18846 31154 18898 31166
rect 19406 31218 19458 31230
rect 19406 31154 19458 31166
rect 19966 31218 20018 31230
rect 19966 31154 20018 31166
rect 20302 31218 20354 31230
rect 20302 31154 20354 31166
rect 21534 31218 21586 31230
rect 21534 31154 21586 31166
rect 25454 31218 25506 31230
rect 25454 31154 25506 31166
rect 26798 31218 26850 31230
rect 26798 31154 26850 31166
rect 34302 31218 34354 31230
rect 34302 31154 34354 31166
rect 34974 31218 35026 31230
rect 34974 31154 35026 31166
rect 49422 31218 49474 31230
rect 49422 31154 49474 31166
rect 54910 31218 54962 31230
rect 54910 31154 54962 31166
rect 56702 31218 56754 31230
rect 56702 31154 56754 31166
rect 2046 31106 2098 31118
rect 2046 31042 2098 31054
rect 2718 31106 2770 31118
rect 2718 31042 2770 31054
rect 3390 31106 3442 31118
rect 8990 31106 9042 31118
rect 4498 31054 4510 31106
rect 4562 31054 4574 31106
rect 3390 31042 3442 31054
rect 8990 31042 9042 31054
rect 9550 31106 9602 31118
rect 9550 31042 9602 31054
rect 16494 31106 16546 31118
rect 16494 31042 16546 31054
rect 18734 31106 18786 31118
rect 18734 31042 18786 31054
rect 19518 31106 19570 31118
rect 25230 31106 25282 31118
rect 29710 31106 29762 31118
rect 22194 31054 22206 31106
rect 22258 31054 22270 31106
rect 27794 31054 27806 31106
rect 27858 31054 27870 31106
rect 19518 31042 19570 31054
rect 25230 31042 25282 31054
rect 29710 31042 29762 31054
rect 31726 31106 31778 31118
rect 31726 31042 31778 31054
rect 33182 31106 33234 31118
rect 33182 31042 33234 31054
rect 36654 31106 36706 31118
rect 44606 31106 44658 31118
rect 54350 31106 54402 31118
rect 39330 31054 39342 31106
rect 39394 31054 39406 31106
rect 39666 31054 39678 31106
rect 39730 31054 39742 31106
rect 45714 31054 45726 31106
rect 45778 31054 45790 31106
rect 36654 31042 36706 31054
rect 44606 31042 44658 31054
rect 54350 31042 54402 31054
rect 2382 30994 2434 31006
rect 1810 30942 1822 30994
rect 1874 30942 1886 30994
rect 2382 30930 2434 30942
rect 3054 30994 3106 31006
rect 3054 30930 3106 30942
rect 4174 30994 4226 31006
rect 4174 30930 4226 30942
rect 5070 30994 5122 31006
rect 11342 30994 11394 31006
rect 12238 30994 12290 31006
rect 8418 30942 8430 30994
rect 8482 30942 8494 30994
rect 9986 30942 9998 30994
rect 10050 30942 10062 30994
rect 11890 30942 11902 30994
rect 11954 30942 11966 30994
rect 5070 30930 5122 30942
rect 11342 30930 11394 30942
rect 12238 30930 12290 30942
rect 12462 30994 12514 31006
rect 12462 30930 12514 30942
rect 12798 30994 12850 31006
rect 19854 30994 19906 31006
rect 16034 30942 16046 30994
rect 16098 30942 16110 30994
rect 17714 30942 17726 30994
rect 17778 30942 17790 30994
rect 12798 30930 12850 30942
rect 19854 30930 19906 30942
rect 20078 30994 20130 31006
rect 20078 30930 20130 30942
rect 21870 30994 21922 31006
rect 23774 30994 23826 31006
rect 22978 30942 22990 30994
rect 23042 30942 23054 30994
rect 21870 30930 21922 30942
rect 23774 30930 23826 30942
rect 24222 30994 24274 31006
rect 24222 30930 24274 30942
rect 24446 30994 24498 31006
rect 29486 30994 29538 31006
rect 27906 30942 27918 30994
rect 27970 30942 27982 30994
rect 24446 30930 24498 30942
rect 29486 30930 29538 30942
rect 29822 30994 29874 31006
rect 31838 30994 31890 31006
rect 30706 30942 30718 30994
rect 30770 30942 30782 30994
rect 31490 30942 31502 30994
rect 31554 30942 31566 30994
rect 29822 30930 29874 30942
rect 31838 30930 31890 30942
rect 31950 30994 32002 31006
rect 34190 30994 34242 31006
rect 32162 30942 32174 30994
rect 32226 30942 32238 30994
rect 33506 30942 33518 30994
rect 33570 30942 33582 30994
rect 31950 30930 32002 30942
rect 34190 30930 34242 30942
rect 35422 30994 35474 31006
rect 54574 30994 54626 31006
rect 38098 30942 38110 30994
rect 38162 30942 38174 30994
rect 43810 30942 43822 30994
rect 43874 30942 43886 30994
rect 44370 30942 44382 30994
rect 44434 30942 44446 30994
rect 45042 30942 45054 30994
rect 45106 30942 45118 30994
rect 49746 30942 49758 30994
rect 49810 30942 49822 30994
rect 52994 30942 53006 30994
rect 53058 30942 53070 30994
rect 53666 30942 53678 30994
rect 53730 30942 53742 30994
rect 35422 30930 35474 30942
rect 54574 30930 54626 30942
rect 54686 30994 54738 31006
rect 54686 30930 54738 30942
rect 54798 30994 54850 31006
rect 54798 30930 54850 30942
rect 55582 30994 55634 31006
rect 55582 30930 55634 30942
rect 3838 30882 3890 30894
rect 3838 30818 3890 30830
rect 6414 30882 6466 30894
rect 11118 30882 11170 30894
rect 8194 30830 8206 30882
rect 8258 30830 8270 30882
rect 9874 30830 9886 30882
rect 9938 30830 9950 30882
rect 6414 30818 6466 30830
rect 11118 30818 11170 30830
rect 13246 30882 13298 30894
rect 18398 30882 18450 30894
rect 15586 30830 15598 30882
rect 15650 30830 15662 30882
rect 17490 30830 17502 30882
rect 17554 30830 17566 30882
rect 13246 30818 13298 30830
rect 18398 30818 18450 30830
rect 22542 30882 22594 30894
rect 24334 30882 24386 30894
rect 23314 30830 23326 30882
rect 23378 30830 23390 30882
rect 22542 30818 22594 30830
rect 24334 30818 24386 30830
rect 25342 30882 25394 30894
rect 31166 30882 31218 30894
rect 30370 30830 30382 30882
rect 30434 30830 30446 30882
rect 25342 30818 25394 30830
rect 31166 30818 31218 30830
rect 33854 30882 33906 30894
rect 33854 30818 33906 30830
rect 35870 30882 35922 30894
rect 35870 30818 35922 30830
rect 37214 30882 37266 30894
rect 37214 30818 37266 30830
rect 37662 30882 37714 30894
rect 48862 30882 48914 30894
rect 38546 30830 38558 30882
rect 38610 30830 38622 30882
rect 37662 30818 37714 30830
rect 40898 30803 40910 30855
rect 40962 30803 40974 30855
rect 43026 30830 43038 30882
rect 43090 30830 43102 30882
rect 47842 30830 47854 30882
rect 47906 30830 47918 30882
rect 51986 30830 51998 30882
rect 52050 30830 52062 30882
rect 53106 30830 53118 30882
rect 53170 30830 53182 30882
rect 48862 30818 48914 30830
rect 11566 30770 11618 30782
rect 11566 30706 11618 30718
rect 18846 30770 18898 30782
rect 18846 30706 18898 30718
rect 27134 30770 27186 30782
rect 27134 30706 27186 30718
rect 33070 30770 33122 30782
rect 33070 30706 33122 30718
rect 33518 30770 33570 30782
rect 33518 30706 33570 30718
rect 34302 30770 34354 30782
rect 34302 30706 34354 30718
rect 35646 30770 35698 30782
rect 35646 30706 35698 30718
rect 36542 30770 36594 30782
rect 36542 30706 36594 30718
rect 39902 30770 39954 30782
rect 39902 30706 39954 30718
rect 40238 30770 40290 30782
rect 55694 30770 55746 30782
rect 52994 30718 53006 30770
rect 53058 30718 53070 30770
rect 40238 30706 40290 30718
rect 55694 30706 55746 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 8878 30434 8930 30446
rect 8878 30370 8930 30382
rect 9102 30434 9154 30446
rect 9102 30370 9154 30382
rect 9326 30434 9378 30446
rect 9326 30370 9378 30382
rect 10782 30434 10834 30446
rect 10782 30370 10834 30382
rect 11006 30434 11058 30446
rect 11006 30370 11058 30382
rect 18734 30434 18786 30446
rect 18734 30370 18786 30382
rect 22430 30434 22482 30446
rect 22430 30370 22482 30382
rect 22878 30434 22930 30446
rect 22878 30370 22930 30382
rect 37102 30434 37154 30446
rect 37102 30370 37154 30382
rect 39678 30434 39730 30446
rect 39678 30370 39730 30382
rect 44942 30434 44994 30446
rect 44942 30370 44994 30382
rect 10222 30322 10274 30334
rect 4610 30270 4622 30322
rect 4674 30270 4686 30322
rect 10222 30258 10274 30270
rect 16158 30322 16210 30334
rect 16158 30258 16210 30270
rect 17054 30322 17106 30334
rect 17054 30258 17106 30270
rect 18958 30322 19010 30334
rect 23550 30322 23602 30334
rect 23090 30270 23102 30322
rect 23154 30270 23166 30322
rect 18958 30258 19010 30270
rect 23550 30258 23602 30270
rect 23774 30322 23826 30334
rect 23774 30258 23826 30270
rect 24110 30322 24162 30334
rect 24110 30258 24162 30270
rect 30158 30322 30210 30334
rect 37214 30322 37266 30334
rect 44046 30322 44098 30334
rect 34402 30270 34414 30322
rect 34466 30270 34478 30322
rect 39330 30270 39342 30322
rect 39394 30270 39406 30322
rect 49074 30270 49086 30322
rect 49138 30270 49150 30322
rect 49634 30270 49646 30322
rect 49698 30270 49710 30322
rect 56018 30270 56030 30322
rect 56082 30270 56094 30322
rect 58146 30270 58158 30322
rect 58210 30270 58222 30322
rect 30158 30258 30210 30270
rect 37214 30258 37266 30270
rect 44046 30258 44098 30270
rect 5518 30210 5570 30222
rect 1810 30158 1822 30210
rect 1874 30158 1886 30210
rect 5518 30146 5570 30158
rect 5742 30210 5794 30222
rect 5742 30146 5794 30158
rect 6078 30210 6130 30222
rect 6078 30146 6130 30158
rect 7982 30210 8034 30222
rect 7982 30146 8034 30158
rect 8654 30210 8706 30222
rect 8654 30146 8706 30158
rect 10558 30210 10610 30222
rect 10558 30146 10610 30158
rect 16942 30210 16994 30222
rect 16942 30146 16994 30158
rect 17166 30210 17218 30222
rect 17166 30146 17218 30158
rect 17838 30210 17890 30222
rect 17838 30146 17890 30158
rect 18062 30210 18114 30222
rect 18062 30146 18114 30158
rect 22542 30210 22594 30222
rect 30046 30210 30098 30222
rect 37886 30210 37938 30222
rect 27122 30158 27134 30210
rect 27186 30158 27198 30210
rect 30818 30158 30830 30210
rect 30882 30158 30894 30210
rect 31602 30158 31614 30210
rect 31666 30158 31678 30210
rect 32274 30158 32286 30210
rect 32338 30158 32350 30210
rect 34850 30158 34862 30210
rect 34914 30158 34926 30210
rect 35858 30158 35870 30210
rect 35922 30158 35934 30210
rect 37426 30158 37438 30210
rect 37490 30158 37502 30210
rect 22542 30146 22594 30158
rect 30046 30146 30098 30158
rect 37886 30146 37938 30158
rect 38222 30210 38274 30222
rect 38222 30146 38274 30158
rect 38670 30210 38722 30222
rect 38670 30146 38722 30158
rect 39006 30210 39058 30222
rect 39006 30146 39058 30158
rect 40126 30210 40178 30222
rect 40126 30146 40178 30158
rect 40686 30210 40738 30222
rect 40686 30146 40738 30158
rect 45278 30210 45330 30222
rect 52670 30210 52722 30222
rect 48738 30158 48750 30210
rect 48802 30158 48814 30210
rect 50082 30158 50094 30210
rect 50146 30158 50158 30210
rect 51538 30158 51550 30210
rect 51602 30158 51614 30210
rect 45278 30146 45330 30158
rect 52670 30146 52722 30158
rect 53230 30210 53282 30222
rect 53230 30146 53282 30158
rect 53566 30210 53618 30222
rect 53566 30146 53618 30158
rect 54462 30210 54514 30222
rect 54462 30146 54514 30158
rect 54910 30210 54962 30222
rect 55234 30158 55246 30210
rect 55298 30158 55310 30210
rect 54910 30146 54962 30158
rect 5966 30098 6018 30110
rect 2482 30046 2494 30098
rect 2546 30046 2558 30098
rect 5966 30034 6018 30046
rect 10446 30098 10498 30110
rect 13806 30098 13858 30110
rect 11666 30046 11678 30098
rect 11730 30046 11742 30098
rect 10446 30034 10498 30046
rect 13806 30034 13858 30046
rect 16270 30098 16322 30110
rect 16270 30034 16322 30046
rect 16606 30098 16658 30110
rect 16606 30034 16658 30046
rect 21646 30098 21698 30110
rect 21646 30034 21698 30046
rect 22430 30098 22482 30110
rect 22430 30034 22482 30046
rect 23102 30098 23154 30110
rect 23102 30034 23154 30046
rect 30270 30098 30322 30110
rect 30270 30034 30322 30046
rect 30382 30098 30434 30110
rect 36318 30098 36370 30110
rect 35410 30046 35422 30098
rect 35474 30046 35486 30098
rect 30382 30034 30434 30046
rect 36318 30034 36370 30046
rect 36430 30098 36482 30110
rect 36430 30034 36482 30046
rect 38446 30098 38498 30110
rect 38446 30034 38498 30046
rect 41022 30098 41074 30110
rect 48190 30098 48242 30110
rect 45490 30046 45502 30098
rect 45554 30046 45566 30098
rect 46050 30046 46062 30098
rect 46114 30046 46126 30098
rect 41022 30034 41074 30046
rect 48190 30034 48242 30046
rect 50542 30098 50594 30110
rect 53006 30098 53058 30110
rect 51986 30046 51998 30098
rect 52050 30046 52062 30098
rect 50542 30034 50594 30046
rect 53006 30034 53058 30046
rect 53342 30098 53394 30110
rect 54114 30046 54126 30098
rect 54178 30046 54190 30098
rect 53342 30034 53394 30046
rect 5070 29986 5122 29998
rect 9774 29986 9826 29998
rect 8306 29934 8318 29986
rect 8370 29934 8382 29986
rect 5070 29922 5122 29934
rect 9774 29922 9826 29934
rect 12014 29986 12066 29998
rect 12014 29922 12066 29934
rect 12574 29986 12626 29998
rect 12574 29922 12626 29934
rect 13470 29986 13522 29998
rect 13470 29922 13522 29934
rect 17614 29986 17666 29998
rect 17614 29922 17666 29934
rect 17950 29986 18002 29998
rect 19518 29986 19570 29998
rect 18386 29934 18398 29986
rect 18450 29934 18462 29986
rect 17950 29922 18002 29934
rect 19518 29922 19570 29934
rect 21310 29986 21362 29998
rect 21310 29922 21362 29934
rect 23998 29986 24050 29998
rect 23998 29922 24050 29934
rect 24222 29986 24274 29998
rect 24222 29922 24274 29934
rect 24894 29986 24946 29998
rect 24894 29922 24946 29934
rect 27358 29986 27410 29998
rect 36094 29986 36146 29998
rect 34850 29934 34862 29986
rect 34914 29934 34926 29986
rect 27358 29922 27410 29934
rect 36094 29922 36146 29934
rect 37998 29986 38050 29998
rect 37998 29922 38050 29934
rect 38558 29986 38610 29998
rect 38558 29922 38610 29934
rect 39454 29986 39506 29998
rect 39454 29922 39506 29934
rect 40014 29986 40066 29998
rect 52782 29986 52834 29998
rect 51426 29934 51438 29986
rect 51490 29934 51502 29986
rect 40014 29922 40066 29934
rect 52782 29922 52834 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 2046 29650 2098 29662
rect 2046 29586 2098 29598
rect 3166 29650 3218 29662
rect 3166 29586 3218 29598
rect 3614 29650 3666 29662
rect 3614 29586 3666 29598
rect 3726 29650 3778 29662
rect 3726 29586 3778 29598
rect 6078 29650 6130 29662
rect 6078 29586 6130 29598
rect 7982 29650 8034 29662
rect 7982 29586 8034 29598
rect 8654 29650 8706 29662
rect 8654 29586 8706 29598
rect 8878 29650 8930 29662
rect 8878 29586 8930 29598
rect 9998 29650 10050 29662
rect 9998 29586 10050 29598
rect 10110 29650 10162 29662
rect 10110 29586 10162 29598
rect 17502 29650 17554 29662
rect 17502 29586 17554 29598
rect 22430 29650 22482 29662
rect 22430 29586 22482 29598
rect 25342 29650 25394 29662
rect 25342 29586 25394 29598
rect 34078 29650 34130 29662
rect 34078 29586 34130 29598
rect 34302 29650 34354 29662
rect 34302 29586 34354 29598
rect 37438 29650 37490 29662
rect 37438 29586 37490 29598
rect 39006 29650 39058 29662
rect 39006 29586 39058 29598
rect 39230 29650 39282 29662
rect 39230 29586 39282 29598
rect 45278 29650 45330 29662
rect 45278 29586 45330 29598
rect 45950 29650 46002 29662
rect 45950 29586 46002 29598
rect 47966 29650 48018 29662
rect 47966 29586 48018 29598
rect 50990 29650 51042 29662
rect 50990 29586 51042 29598
rect 52446 29650 52498 29662
rect 52446 29586 52498 29598
rect 52558 29650 52610 29662
rect 52558 29586 52610 29598
rect 53118 29650 53170 29662
rect 53118 29586 53170 29598
rect 54014 29650 54066 29662
rect 54014 29586 54066 29598
rect 54238 29650 54290 29662
rect 54238 29586 54290 29598
rect 55806 29650 55858 29662
rect 55806 29586 55858 29598
rect 57150 29650 57202 29662
rect 57150 29586 57202 29598
rect 58158 29650 58210 29662
rect 58158 29586 58210 29598
rect 2718 29538 2770 29550
rect 2718 29474 2770 29486
rect 4286 29538 4338 29550
rect 4286 29474 4338 29486
rect 4510 29538 4562 29550
rect 4510 29474 4562 29486
rect 5966 29538 6018 29550
rect 5966 29474 6018 29486
rect 9662 29538 9714 29550
rect 33294 29538 33346 29550
rect 13010 29486 13022 29538
rect 13074 29486 13086 29538
rect 18050 29486 18062 29538
rect 18114 29486 18126 29538
rect 18610 29486 18622 29538
rect 18674 29486 18686 29538
rect 21186 29486 21198 29538
rect 21250 29486 21262 29538
rect 23314 29486 23326 29538
rect 23378 29486 23390 29538
rect 27346 29486 27358 29538
rect 27410 29486 27422 29538
rect 9662 29474 9714 29486
rect 33294 29474 33346 29486
rect 35086 29538 35138 29550
rect 35086 29474 35138 29486
rect 35422 29538 35474 29550
rect 35422 29474 35474 29486
rect 35646 29538 35698 29550
rect 35646 29474 35698 29486
rect 36542 29538 36594 29550
rect 36542 29474 36594 29486
rect 38110 29538 38162 29550
rect 38110 29474 38162 29486
rect 43262 29538 43314 29550
rect 43262 29474 43314 29486
rect 43710 29538 43762 29550
rect 47182 29538 47234 29550
rect 44370 29486 44382 29538
rect 44434 29486 44446 29538
rect 43710 29474 43762 29486
rect 47182 29474 47234 29486
rect 47854 29538 47906 29550
rect 47854 29474 47906 29486
rect 51214 29538 51266 29550
rect 51214 29474 51266 29486
rect 53790 29538 53842 29550
rect 53790 29474 53842 29486
rect 54686 29538 54738 29550
rect 54686 29474 54738 29486
rect 55134 29538 55186 29550
rect 55134 29474 55186 29486
rect 55246 29538 55298 29550
rect 55246 29474 55298 29486
rect 55582 29538 55634 29550
rect 55582 29474 55634 29486
rect 55918 29538 55970 29550
rect 57810 29486 57822 29538
rect 57874 29486 57886 29538
rect 55918 29474 55970 29486
rect 1710 29426 1762 29438
rect 1710 29362 1762 29374
rect 2382 29426 2434 29438
rect 2382 29362 2434 29374
rect 3502 29426 3554 29438
rect 3502 29362 3554 29374
rect 4174 29426 4226 29438
rect 4174 29362 4226 29374
rect 4622 29426 4674 29438
rect 7422 29426 7474 29438
rect 6962 29374 6974 29426
rect 7026 29374 7038 29426
rect 4622 29362 4674 29374
rect 7422 29362 7474 29374
rect 7758 29426 7810 29438
rect 7758 29362 7810 29374
rect 8094 29426 8146 29438
rect 8094 29362 8146 29374
rect 8990 29426 9042 29438
rect 8990 29362 9042 29374
rect 9886 29426 9938 29438
rect 30942 29426 30994 29438
rect 33182 29426 33234 29438
rect 12226 29374 12238 29426
rect 12290 29374 12302 29426
rect 21970 29374 21982 29426
rect 22034 29374 22046 29426
rect 23426 29374 23438 29426
rect 23490 29374 23502 29426
rect 26562 29374 26574 29426
rect 26626 29374 26638 29426
rect 30370 29374 30382 29426
rect 30434 29374 30446 29426
rect 31826 29374 31838 29426
rect 31890 29374 31902 29426
rect 9886 29362 9938 29374
rect 30942 29362 30994 29374
rect 33182 29362 33234 29374
rect 33406 29426 33458 29438
rect 33854 29426 33906 29438
rect 33506 29374 33518 29426
rect 33570 29374 33582 29426
rect 33406 29362 33458 29374
rect 33854 29362 33906 29374
rect 34414 29426 34466 29438
rect 34414 29362 34466 29374
rect 35198 29426 35250 29438
rect 35198 29362 35250 29374
rect 36318 29426 36370 29438
rect 36990 29426 37042 29438
rect 36642 29374 36654 29426
rect 36706 29374 36718 29426
rect 36318 29362 36370 29374
rect 36990 29362 37042 29374
rect 37214 29426 37266 29438
rect 37214 29362 37266 29374
rect 37550 29426 37602 29438
rect 37550 29362 37602 29374
rect 38446 29426 38498 29438
rect 38446 29362 38498 29374
rect 38782 29426 38834 29438
rect 42702 29426 42754 29438
rect 43374 29426 43426 29438
rect 47406 29426 47458 29438
rect 39442 29374 39454 29426
rect 39506 29374 39518 29426
rect 43026 29374 43038 29426
rect 43090 29374 43102 29426
rect 44146 29374 44158 29426
rect 44210 29374 44222 29426
rect 38782 29362 38834 29374
rect 42702 29362 42754 29374
rect 43374 29362 43426 29374
rect 47406 29362 47458 29374
rect 48078 29426 48130 29438
rect 49982 29426 50034 29438
rect 49746 29374 49758 29426
rect 49810 29374 49822 29426
rect 48078 29362 48130 29374
rect 49982 29362 50034 29374
rect 50878 29426 50930 29438
rect 50878 29362 50930 29374
rect 51326 29426 51378 29438
rect 52222 29426 52274 29438
rect 51986 29374 51998 29426
rect 52050 29374 52062 29426
rect 51326 29362 51378 29374
rect 52222 29362 52274 29374
rect 53230 29426 53282 29438
rect 53230 29362 53282 29374
rect 54126 29426 54178 29438
rect 54126 29362 54178 29374
rect 54798 29426 54850 29438
rect 54798 29362 54850 29374
rect 57486 29426 57538 29438
rect 57486 29362 57538 29374
rect 5070 29314 5122 29326
rect 5070 29250 5122 29262
rect 5518 29314 5570 29326
rect 5518 29250 5570 29262
rect 6190 29314 6242 29326
rect 6190 29250 6242 29262
rect 6526 29314 6578 29326
rect 6526 29250 6578 29262
rect 10670 29314 10722 29326
rect 10670 29250 10722 29262
rect 11902 29314 11954 29326
rect 26350 29314 26402 29326
rect 31054 29314 31106 29326
rect 32398 29314 32450 29326
rect 15138 29262 15150 29314
rect 15202 29262 15214 29314
rect 19058 29262 19070 29314
rect 19122 29262 19134 29314
rect 29474 29262 29486 29314
rect 29538 29262 29550 29314
rect 31602 29262 31614 29314
rect 31666 29262 31678 29314
rect 11902 29250 11954 29262
rect 26350 29250 26402 29262
rect 31054 29250 31106 29262
rect 32398 29250 32450 29262
rect 36430 29314 36482 29326
rect 36430 29250 36482 29262
rect 38558 29314 38610 29326
rect 38558 29250 38610 29262
rect 41470 29314 41522 29326
rect 41470 29250 41522 29262
rect 42478 29314 42530 29326
rect 42478 29250 42530 29262
rect 49086 29314 49138 29326
rect 56926 29314 56978 29326
rect 52546 29262 52558 29314
rect 52610 29262 52622 29314
rect 49086 29250 49138 29262
rect 56926 29250 56978 29262
rect 17838 29202 17890 29214
rect 17838 29138 17890 29150
rect 22766 29202 22818 29214
rect 22766 29138 22818 29150
rect 38894 29202 38946 29214
rect 38894 29138 38946 29150
rect 44942 29202 44994 29214
rect 44942 29138 44994 29150
rect 53118 29202 53170 29214
rect 53118 29138 53170 29150
rect 54686 29202 54738 29214
rect 54686 29138 54738 29150
rect 55246 29202 55298 29214
rect 55246 29138 55298 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 18062 28866 18114 28878
rect 18062 28802 18114 28814
rect 25678 28866 25730 28878
rect 25678 28802 25730 28814
rect 27246 28866 27298 28878
rect 27246 28802 27298 28814
rect 32510 28866 32562 28878
rect 37202 28814 37214 28866
rect 37266 28863 37278 28866
rect 37762 28863 37774 28866
rect 37266 28817 37774 28863
rect 37266 28814 37278 28817
rect 37762 28814 37774 28817
rect 37826 28814 37838 28866
rect 32510 28802 32562 28814
rect 8094 28754 8146 28766
rect 4610 28702 4622 28754
rect 4674 28702 4686 28754
rect 5954 28702 5966 28754
rect 6018 28702 6030 28754
rect 7522 28702 7534 28754
rect 7586 28702 7598 28754
rect 8094 28690 8146 28702
rect 13918 28754 13970 28766
rect 13918 28690 13970 28702
rect 18286 28754 18338 28766
rect 18286 28690 18338 28702
rect 18622 28754 18674 28766
rect 18622 28690 18674 28702
rect 19294 28754 19346 28766
rect 19294 28690 19346 28702
rect 22206 28754 22258 28766
rect 30830 28754 30882 28766
rect 25106 28702 25118 28754
rect 25170 28702 25182 28754
rect 22206 28690 22258 28702
rect 30830 28690 30882 28702
rect 31614 28754 31666 28766
rect 31614 28690 31666 28702
rect 32398 28754 32450 28766
rect 32398 28690 32450 28702
rect 33294 28754 33346 28766
rect 33294 28690 33346 28702
rect 33406 28754 33458 28766
rect 33406 28690 33458 28702
rect 33854 28754 33906 28766
rect 33854 28690 33906 28702
rect 34750 28754 34802 28766
rect 37214 28754 37266 28766
rect 35634 28702 35646 28754
rect 35698 28702 35710 28754
rect 34750 28690 34802 28702
rect 37214 28690 37266 28702
rect 37998 28754 38050 28766
rect 37998 28690 38050 28702
rect 40686 28754 40738 28766
rect 44270 28754 44322 28766
rect 42242 28702 42254 28754
rect 42306 28702 42318 28754
rect 40686 28690 40738 28702
rect 44270 28690 44322 28702
rect 47966 28754 48018 28766
rect 47966 28690 48018 28702
rect 48526 28754 48578 28766
rect 48526 28690 48578 28702
rect 49870 28754 49922 28766
rect 49870 28690 49922 28702
rect 51326 28754 51378 28766
rect 55806 28754 55858 28766
rect 55234 28702 55246 28754
rect 55298 28702 55310 28754
rect 51326 28690 51378 28702
rect 55806 28690 55858 28702
rect 56366 28754 56418 28766
rect 56366 28690 56418 28702
rect 57598 28754 57650 28766
rect 57598 28690 57650 28702
rect 6302 28642 6354 28654
rect 1810 28590 1822 28642
rect 1874 28590 1886 28642
rect 6302 28578 6354 28590
rect 6638 28642 6690 28654
rect 7982 28642 8034 28654
rect 7298 28590 7310 28642
rect 7362 28590 7374 28642
rect 6638 28578 6690 28590
rect 7982 28578 8034 28590
rect 8206 28642 8258 28654
rect 8206 28578 8258 28590
rect 8654 28642 8706 28654
rect 8654 28578 8706 28590
rect 9438 28642 9490 28654
rect 9438 28578 9490 28590
rect 12462 28642 12514 28654
rect 12462 28578 12514 28590
rect 13358 28642 13410 28654
rect 13358 28578 13410 28590
rect 18510 28642 18562 28654
rect 18510 28578 18562 28590
rect 26462 28642 26514 28654
rect 26462 28578 26514 28590
rect 27582 28642 27634 28654
rect 29934 28642 29986 28654
rect 31502 28642 31554 28654
rect 28018 28590 28030 28642
rect 28082 28590 28094 28642
rect 30370 28590 30382 28642
rect 30434 28590 30446 28642
rect 27582 28578 27634 28590
rect 29934 28578 29986 28590
rect 31502 28578 31554 28590
rect 31726 28642 31778 28654
rect 31726 28578 31778 28590
rect 32062 28642 32114 28654
rect 32062 28578 32114 28590
rect 35198 28642 35250 28654
rect 35870 28642 35922 28654
rect 35522 28590 35534 28642
rect 35586 28590 35598 28642
rect 35198 28578 35250 28590
rect 35870 28578 35922 28590
rect 36542 28642 36594 28654
rect 36542 28578 36594 28590
rect 40798 28642 40850 28654
rect 42590 28642 42642 28654
rect 41122 28590 41134 28642
rect 41186 28590 41198 28642
rect 41906 28590 41918 28642
rect 41970 28590 41982 28642
rect 40798 28578 40850 28590
rect 42590 28578 42642 28590
rect 43262 28642 43314 28654
rect 43262 28578 43314 28590
rect 43486 28642 43538 28654
rect 43486 28578 43538 28590
rect 45950 28642 46002 28654
rect 45950 28578 46002 28590
rect 46174 28642 46226 28654
rect 46174 28578 46226 28590
rect 47406 28642 47458 28654
rect 50766 28642 50818 28654
rect 50418 28590 50430 28642
rect 50482 28590 50494 28642
rect 47406 28578 47458 28590
rect 50766 28578 50818 28590
rect 51886 28642 51938 28654
rect 51886 28578 51938 28590
rect 53342 28642 53394 28654
rect 53342 28578 53394 28590
rect 53902 28642 53954 28654
rect 53902 28578 53954 28590
rect 54126 28642 54178 28654
rect 55134 28642 55186 28654
rect 54674 28590 54686 28642
rect 54738 28590 54750 28642
rect 54126 28578 54178 28590
rect 55134 28578 55186 28590
rect 57150 28642 57202 28654
rect 57150 28578 57202 28590
rect 58158 28642 58210 28654
rect 58158 28578 58210 28590
rect 6078 28530 6130 28542
rect 12798 28530 12850 28542
rect 2482 28478 2494 28530
rect 2546 28478 2558 28530
rect 9090 28478 9102 28530
rect 9154 28478 9166 28530
rect 6078 28466 6130 28478
rect 12798 28466 12850 28478
rect 18734 28530 18786 28542
rect 18734 28466 18786 28478
rect 25902 28530 25954 28542
rect 33182 28530 33234 28542
rect 28354 28478 28366 28530
rect 28418 28478 28430 28530
rect 29586 28478 29598 28530
rect 29650 28478 29662 28530
rect 25902 28466 25954 28478
rect 33182 28466 33234 28478
rect 34862 28530 34914 28542
rect 34862 28466 34914 28478
rect 35086 28530 35138 28542
rect 35086 28466 35138 28478
rect 36206 28530 36258 28542
rect 36206 28466 36258 28478
rect 36318 28530 36370 28542
rect 36318 28466 36370 28478
rect 43710 28530 43762 28542
rect 43710 28466 43762 28478
rect 43822 28530 43874 28542
rect 43822 28466 43874 28478
rect 46622 28530 46674 28542
rect 46622 28466 46674 28478
rect 51438 28530 51490 28542
rect 51438 28466 51490 28478
rect 52894 28530 52946 28542
rect 52894 28466 52946 28478
rect 5070 28418 5122 28430
rect 5070 28354 5122 28366
rect 12686 28418 12738 28430
rect 12686 28354 12738 28366
rect 13806 28418 13858 28430
rect 13806 28354 13858 28366
rect 14030 28418 14082 28430
rect 14030 28354 14082 28366
rect 17838 28418 17890 28430
rect 17838 28354 17890 28366
rect 19854 28418 19906 28430
rect 19854 28354 19906 28366
rect 20302 28418 20354 28430
rect 20302 28354 20354 28366
rect 23662 28418 23714 28430
rect 23662 28354 23714 28366
rect 23998 28418 24050 28430
rect 23998 28354 24050 28366
rect 24670 28418 24722 28430
rect 24670 28354 24722 28366
rect 25790 28418 25842 28430
rect 25790 28354 25842 28366
rect 37550 28418 37602 28430
rect 37550 28354 37602 28366
rect 38558 28418 38610 28430
rect 38558 28354 38610 28366
rect 39006 28418 39058 28430
rect 39006 28354 39058 28366
rect 40574 28418 40626 28430
rect 40574 28354 40626 28366
rect 45278 28418 45330 28430
rect 45278 28354 45330 28366
rect 45390 28418 45442 28430
rect 45390 28354 45442 28366
rect 45502 28418 45554 28430
rect 45502 28354 45554 28366
rect 46734 28418 46786 28430
rect 46734 28354 46786 28366
rect 46846 28418 46898 28430
rect 46846 28354 46898 28366
rect 47854 28418 47906 28430
rect 47854 28354 47906 28366
rect 48078 28418 48130 28430
rect 48078 28354 48130 28366
rect 51214 28418 51266 28430
rect 51214 28354 51266 28366
rect 52670 28418 52722 28430
rect 52670 28354 52722 28366
rect 52782 28418 52834 28430
rect 54910 28418 54962 28430
rect 53554 28366 53566 28418
rect 53618 28366 53630 28418
rect 52782 28354 52834 28366
rect 54910 28354 54962 28366
rect 55246 28418 55298 28430
rect 55246 28354 55298 28366
rect 55918 28418 55970 28430
rect 55918 28354 55970 28366
rect 57822 28418 57874 28430
rect 57822 28354 57874 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 2718 28082 2770 28094
rect 2718 28018 2770 28030
rect 3166 28082 3218 28094
rect 3166 28018 3218 28030
rect 3614 28082 3666 28094
rect 3614 28018 3666 28030
rect 3726 28082 3778 28094
rect 3726 28018 3778 28030
rect 4622 28082 4674 28094
rect 4622 28018 4674 28030
rect 13022 28082 13074 28094
rect 13022 28018 13074 28030
rect 13582 28082 13634 28094
rect 13582 28018 13634 28030
rect 14254 28082 14306 28094
rect 14254 28018 14306 28030
rect 18062 28082 18114 28094
rect 18062 28018 18114 28030
rect 22094 28082 22146 28094
rect 22094 28018 22146 28030
rect 26686 28082 26738 28094
rect 26686 28018 26738 28030
rect 28366 28082 28418 28094
rect 28366 28018 28418 28030
rect 29262 28082 29314 28094
rect 29262 28018 29314 28030
rect 30270 28082 30322 28094
rect 30270 28018 30322 28030
rect 31838 28082 31890 28094
rect 31838 28018 31890 28030
rect 39006 28082 39058 28094
rect 39006 28018 39058 28030
rect 42254 28082 42306 28094
rect 42254 28018 42306 28030
rect 42366 28082 42418 28094
rect 42366 28018 42418 28030
rect 43150 28082 43202 28094
rect 43150 28018 43202 28030
rect 44158 28082 44210 28094
rect 44158 28018 44210 28030
rect 44270 28082 44322 28094
rect 44270 28018 44322 28030
rect 48862 28082 48914 28094
rect 49970 28030 49982 28082
rect 50034 28030 50046 28082
rect 55346 28030 55358 28082
rect 55410 28030 55422 28082
rect 48862 28018 48914 28030
rect 1710 27970 1762 27982
rect 1710 27906 1762 27918
rect 2046 27970 2098 27982
rect 2046 27906 2098 27918
rect 5070 27970 5122 27982
rect 5070 27906 5122 27918
rect 5518 27970 5570 27982
rect 5518 27906 5570 27918
rect 5630 27970 5682 27982
rect 5630 27906 5682 27918
rect 8430 27970 8482 27982
rect 8430 27906 8482 27918
rect 11566 27970 11618 27982
rect 11566 27906 11618 27918
rect 12798 27970 12850 27982
rect 12798 27906 12850 27918
rect 13246 27970 13298 27982
rect 13246 27906 13298 27918
rect 13806 27970 13858 27982
rect 13806 27906 13858 27918
rect 13918 27970 13970 27982
rect 19182 27970 19234 27982
rect 23662 27970 23714 27982
rect 14578 27918 14590 27970
rect 14642 27918 14654 27970
rect 17378 27918 17390 27970
rect 17442 27918 17454 27970
rect 22978 27918 22990 27970
rect 23042 27918 23054 27970
rect 13918 27906 13970 27918
rect 19182 27906 19234 27918
rect 23662 27906 23714 27918
rect 28590 27970 28642 27982
rect 28590 27906 28642 27918
rect 29710 27970 29762 27982
rect 29710 27906 29762 27918
rect 33294 27970 33346 27982
rect 33294 27906 33346 27918
rect 35870 27970 35922 27982
rect 35870 27906 35922 27918
rect 40238 27970 40290 27982
rect 40238 27906 40290 27918
rect 42590 27970 42642 27982
rect 42590 27906 42642 27918
rect 44046 27970 44098 27982
rect 50430 27970 50482 27982
rect 46050 27918 46062 27970
rect 46114 27918 46126 27970
rect 44046 27906 44098 27918
rect 50430 27906 50482 27918
rect 53006 27970 53058 27982
rect 57810 27918 57822 27970
rect 57874 27918 57886 27970
rect 53006 27906 53058 27918
rect 3502 27858 3554 27870
rect 2482 27806 2494 27858
rect 2546 27806 2558 27858
rect 3502 27794 3554 27806
rect 4174 27858 4226 27870
rect 4174 27794 4226 27806
rect 4398 27858 4450 27870
rect 4398 27794 4450 27806
rect 4846 27858 4898 27870
rect 4846 27794 4898 27806
rect 5294 27858 5346 27870
rect 5294 27794 5346 27806
rect 7646 27858 7698 27870
rect 7646 27794 7698 27806
rect 9550 27858 9602 27870
rect 9550 27794 9602 27806
rect 9774 27858 9826 27870
rect 9774 27794 9826 27806
rect 10222 27858 10274 27870
rect 10222 27794 10274 27806
rect 11790 27858 11842 27870
rect 11790 27794 11842 27806
rect 12462 27858 12514 27870
rect 12462 27794 12514 27806
rect 13358 27858 13410 27870
rect 13358 27794 13410 27806
rect 18286 27858 18338 27870
rect 21646 27858 21698 27870
rect 18610 27806 18622 27858
rect 18674 27806 18686 27858
rect 19618 27806 19630 27858
rect 19682 27806 19694 27858
rect 21074 27806 21086 27858
rect 21138 27806 21150 27858
rect 18286 27794 18338 27806
rect 21646 27794 21698 27806
rect 22430 27858 22482 27870
rect 25566 27858 25618 27870
rect 23202 27806 23214 27858
rect 23266 27806 23278 27858
rect 24098 27806 24110 27858
rect 24162 27806 24174 27858
rect 22430 27794 22482 27806
rect 25566 27794 25618 27806
rect 25902 27858 25954 27870
rect 25902 27794 25954 27806
rect 26014 27858 26066 27870
rect 26014 27794 26066 27806
rect 28702 27858 28754 27870
rect 28702 27794 28754 27806
rect 28814 27858 28866 27870
rect 28814 27794 28866 27806
rect 29038 27858 29090 27870
rect 29038 27794 29090 27806
rect 29374 27858 29426 27870
rect 29374 27794 29426 27806
rect 31950 27858 32002 27870
rect 31950 27794 32002 27806
rect 32062 27858 32114 27870
rect 38558 27858 38610 27870
rect 33954 27806 33966 27858
rect 34018 27806 34030 27858
rect 36082 27806 36094 27858
rect 36146 27806 36158 27858
rect 36306 27806 36318 27858
rect 36370 27806 36382 27858
rect 37650 27806 37662 27858
rect 37714 27806 37726 27858
rect 32062 27794 32114 27806
rect 38558 27794 38610 27806
rect 39230 27858 39282 27870
rect 39230 27794 39282 27806
rect 40126 27858 40178 27870
rect 40126 27794 40178 27806
rect 40462 27858 40514 27870
rect 40462 27794 40514 27806
rect 41358 27858 41410 27870
rect 41358 27794 41410 27806
rect 41582 27858 41634 27870
rect 41582 27794 41634 27806
rect 41806 27858 41858 27870
rect 41806 27794 41858 27806
rect 42142 27858 42194 27870
rect 51550 27858 51602 27870
rect 43474 27806 43486 27858
rect 43538 27806 43550 27858
rect 43810 27806 43822 27858
rect 43874 27806 43886 27858
rect 45378 27806 45390 27858
rect 45442 27806 45454 27858
rect 42142 27794 42194 27806
rect 51550 27794 51602 27806
rect 51998 27858 52050 27870
rect 55694 27858 55746 27870
rect 54226 27806 54238 27858
rect 54290 27806 54302 27858
rect 54674 27806 54686 27858
rect 54738 27806 54750 27858
rect 51998 27794 52050 27806
rect 55694 27794 55746 27806
rect 58158 27858 58210 27870
rect 58158 27794 58210 27806
rect 7422 27746 7474 27758
rect 7422 27682 7474 27694
rect 9662 27746 9714 27758
rect 9662 27682 9714 27694
rect 17726 27746 17778 27758
rect 17726 27682 17778 27694
rect 18174 27746 18226 27758
rect 25678 27746 25730 27758
rect 20066 27694 20078 27746
rect 20130 27694 20142 27746
rect 21186 27694 21198 27746
rect 21250 27694 21262 27746
rect 24546 27694 24558 27746
rect 24610 27694 24622 27746
rect 18174 27682 18226 27694
rect 25678 27682 25730 27694
rect 31054 27746 31106 27758
rect 31054 27682 31106 27694
rect 32286 27746 32338 27758
rect 34750 27746 34802 27758
rect 34178 27694 34190 27746
rect 34242 27694 34254 27746
rect 32286 27682 32338 27694
rect 34750 27682 34802 27694
rect 35198 27746 35250 27758
rect 38222 27746 38274 27758
rect 37314 27694 37326 27746
rect 37378 27694 37390 27746
rect 35198 27682 35250 27694
rect 38222 27682 38274 27694
rect 38782 27746 38834 27758
rect 38782 27682 38834 27694
rect 39118 27746 39170 27758
rect 39118 27682 39170 27694
rect 44718 27746 44770 27758
rect 54014 27746 54066 27758
rect 48178 27694 48190 27746
rect 48242 27694 48254 27746
rect 44718 27682 44770 27694
rect 54014 27682 54066 27694
rect 57150 27746 57202 27758
rect 57150 27682 57202 27694
rect 57598 27746 57650 27758
rect 57598 27682 57650 27694
rect 7982 27634 8034 27646
rect 7982 27570 8034 27582
rect 8654 27634 8706 27646
rect 8654 27570 8706 27582
rect 8990 27634 9042 27646
rect 8990 27570 9042 27582
rect 12126 27634 12178 27646
rect 12126 27570 12178 27582
rect 32510 27634 32562 27646
rect 32510 27570 32562 27582
rect 40910 27634 40962 27646
rect 40910 27570 40962 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 18622 27298 18674 27310
rect 18622 27234 18674 27246
rect 19742 27298 19794 27310
rect 19742 27234 19794 27246
rect 20190 27298 20242 27310
rect 20190 27234 20242 27246
rect 24110 27298 24162 27310
rect 24110 27234 24162 27246
rect 33070 27298 33122 27310
rect 33070 27234 33122 27246
rect 38670 27298 38722 27310
rect 54350 27298 54402 27310
rect 51202 27246 51214 27298
rect 51266 27246 51278 27298
rect 54562 27246 54574 27298
rect 54626 27295 54638 27298
rect 55010 27295 55022 27298
rect 54626 27249 55022 27295
rect 54626 27246 54638 27249
rect 55010 27246 55022 27249
rect 55074 27246 55086 27298
rect 38670 27234 38722 27246
rect 54350 27234 54402 27246
rect 14142 27186 14194 27198
rect 21422 27186 21474 27198
rect 6402 27134 6414 27186
rect 6466 27134 6478 27186
rect 18162 27134 18174 27186
rect 18226 27134 18238 27186
rect 14142 27122 14194 27134
rect 21422 27122 21474 27134
rect 22430 27186 22482 27198
rect 22430 27122 22482 27134
rect 23214 27186 23266 27198
rect 32510 27186 32562 27198
rect 25442 27134 25454 27186
rect 25506 27134 25518 27186
rect 27570 27134 27582 27186
rect 27634 27134 27646 27186
rect 23214 27122 23266 27134
rect 32510 27122 32562 27134
rect 33630 27186 33682 27198
rect 33630 27122 33682 27134
rect 34190 27186 34242 27198
rect 34190 27122 34242 27134
rect 35310 27186 35362 27198
rect 35310 27122 35362 27134
rect 36318 27186 36370 27198
rect 36318 27122 36370 27134
rect 37550 27186 37602 27198
rect 37550 27122 37602 27134
rect 40238 27186 40290 27198
rect 40238 27122 40290 27134
rect 41134 27186 41186 27198
rect 44942 27186 44994 27198
rect 43026 27134 43038 27186
rect 43090 27134 43102 27186
rect 43922 27134 43934 27186
rect 43986 27134 43998 27186
rect 41134 27122 41186 27134
rect 44942 27122 44994 27134
rect 46174 27186 46226 27198
rect 52782 27186 52834 27198
rect 47730 27134 47742 27186
rect 47794 27134 47806 27186
rect 51090 27134 51102 27186
rect 51154 27134 51166 27186
rect 46174 27122 46226 27134
rect 52782 27122 52834 27134
rect 54910 27186 54962 27198
rect 56018 27134 56030 27186
rect 56082 27134 56094 27186
rect 58146 27134 58158 27186
rect 58210 27134 58222 27186
rect 54910 27122 54962 27134
rect 1710 27074 1762 27086
rect 3950 27074 4002 27086
rect 2482 27022 2494 27074
rect 2546 27022 2558 27074
rect 3490 27022 3502 27074
rect 3554 27022 3566 27074
rect 1710 27010 1762 27022
rect 3950 27010 4002 27022
rect 4398 27074 4450 27086
rect 4398 27010 4450 27022
rect 4622 27074 4674 27086
rect 4622 27010 4674 27022
rect 4734 27074 4786 27086
rect 4734 27010 4786 27022
rect 5070 27074 5122 27086
rect 12574 27074 12626 27086
rect 8418 27022 8430 27074
rect 8482 27022 8494 27074
rect 10434 27022 10446 27074
rect 10498 27022 10510 27074
rect 5070 27010 5122 27022
rect 12574 27010 12626 27022
rect 13806 27074 13858 27086
rect 13806 27010 13858 27022
rect 14030 27074 14082 27086
rect 14030 27010 14082 27022
rect 14366 27074 14418 27086
rect 19294 27074 19346 27086
rect 15250 27022 15262 27074
rect 15314 27022 15326 27074
rect 18946 27022 18958 27074
rect 19010 27022 19022 27074
rect 14366 27010 14418 27022
rect 19294 27010 19346 27022
rect 19854 27074 19906 27086
rect 19854 27010 19906 27022
rect 20414 27074 20466 27086
rect 20414 27010 20466 27022
rect 21310 27074 21362 27086
rect 23438 27074 23490 27086
rect 22754 27022 22766 27074
rect 22818 27022 22830 27074
rect 21310 27010 21362 27022
rect 23438 27010 23490 27022
rect 23886 27074 23938 27086
rect 23886 27010 23938 27022
rect 24334 27074 24386 27086
rect 30494 27074 30546 27086
rect 24770 27022 24782 27074
rect 24834 27022 24846 27074
rect 24334 27010 24386 27022
rect 30494 27010 30546 27022
rect 31166 27074 31218 27086
rect 31166 27010 31218 27022
rect 32062 27074 32114 27086
rect 32062 27010 32114 27022
rect 32622 27074 32674 27086
rect 32622 27010 32674 27022
rect 33966 27074 34018 27086
rect 33966 27010 34018 27022
rect 34414 27074 34466 27086
rect 34414 27010 34466 27022
rect 36206 27074 36258 27086
rect 36206 27010 36258 27022
rect 36430 27074 36482 27086
rect 36430 27010 36482 27022
rect 37326 27074 37378 27086
rect 37326 27010 37378 27022
rect 37774 27074 37826 27086
rect 37774 27010 37826 27022
rect 38222 27074 38274 27086
rect 38222 27010 38274 27022
rect 38782 27074 38834 27086
rect 38782 27010 38834 27022
rect 40910 27074 40962 27086
rect 40910 27010 40962 27022
rect 41358 27074 41410 27086
rect 41358 27010 41410 27022
rect 41470 27074 41522 27086
rect 41470 27010 41522 27022
rect 42590 27074 42642 27086
rect 45502 27074 45554 27086
rect 43474 27022 43486 27074
rect 43538 27022 43550 27074
rect 42590 27010 42642 27022
rect 45502 27010 45554 27022
rect 45950 27074 46002 27086
rect 45950 27010 46002 27022
rect 46398 27074 46450 27086
rect 52670 27074 52722 27086
rect 54014 27074 54066 27086
rect 47842 27022 47854 27074
rect 47906 27022 47918 27074
rect 48626 27022 48638 27074
rect 48690 27022 48702 27074
rect 51538 27022 51550 27074
rect 51602 27022 51614 27074
rect 51762 27022 51774 27074
rect 51826 27022 51838 27074
rect 53442 27022 53454 27074
rect 53506 27022 53518 27074
rect 55234 27022 55246 27074
rect 55298 27022 55310 27074
rect 46398 27010 46450 27022
rect 52670 27010 52722 27022
rect 54014 27010 54066 27022
rect 2718 26962 2770 26974
rect 5742 26962 5794 26974
rect 2034 26910 2046 26962
rect 2098 26910 2110 26962
rect 3266 26910 3278 26962
rect 3330 26910 3342 26962
rect 2718 26898 2770 26910
rect 5742 26898 5794 26910
rect 6526 26962 6578 26974
rect 6526 26898 6578 26910
rect 6750 26962 6802 26974
rect 6750 26898 6802 26910
rect 7870 26962 7922 26974
rect 7870 26898 7922 26910
rect 7982 26962 8034 26974
rect 11006 26962 11058 26974
rect 14590 26962 14642 26974
rect 8530 26910 8542 26962
rect 8594 26910 8606 26962
rect 12898 26910 12910 26962
rect 12962 26910 12974 26962
rect 7982 26898 8034 26910
rect 11006 26898 11058 26910
rect 14590 26898 14642 26910
rect 14702 26962 14754 26974
rect 19630 26962 19682 26974
rect 16034 26910 16046 26962
rect 16098 26910 16110 26962
rect 14702 26898 14754 26910
rect 19630 26898 19682 26910
rect 21534 26962 21586 26974
rect 30942 26962 30994 26974
rect 30146 26910 30158 26962
rect 30210 26910 30222 26962
rect 21534 26898 21586 26910
rect 30942 26898 30994 26910
rect 31726 26962 31778 26974
rect 31726 26898 31778 26910
rect 31838 26962 31890 26974
rect 31838 26898 31890 26910
rect 32286 26962 32338 26974
rect 32286 26898 32338 26910
rect 32958 26962 33010 26974
rect 32958 26898 33010 26910
rect 33070 26962 33122 26974
rect 33070 26898 33122 26910
rect 34750 26962 34802 26974
rect 34750 26898 34802 26910
rect 35982 26962 36034 26974
rect 35982 26898 36034 26910
rect 36878 26962 36930 26974
rect 36878 26898 36930 26910
rect 38670 26962 38722 26974
rect 38670 26898 38722 26910
rect 39342 26962 39394 26974
rect 39342 26898 39394 26910
rect 43934 26962 43986 26974
rect 43934 26898 43986 26910
rect 44046 26962 44098 26974
rect 44046 26898 44098 26910
rect 44830 26962 44882 26974
rect 44830 26898 44882 26910
rect 45726 26962 45778 26974
rect 45726 26898 45778 26910
rect 46958 26962 47010 26974
rect 52894 26962 52946 26974
rect 47506 26910 47518 26962
rect 47570 26910 47582 26962
rect 46958 26898 47010 26910
rect 52894 26898 52946 26910
rect 53006 26962 53058 26974
rect 53006 26898 53058 26910
rect 53790 26962 53842 26974
rect 53790 26898 53842 26910
rect 4062 26850 4114 26862
rect 4062 26786 4114 26798
rect 4286 26850 4338 26862
rect 4286 26786 4338 26798
rect 8206 26850 8258 26862
rect 14926 26850 14978 26862
rect 9426 26798 9438 26850
rect 9490 26798 9502 26850
rect 8206 26786 8258 26798
rect 14926 26786 14978 26798
rect 18734 26850 18786 26862
rect 18734 26786 18786 26798
rect 21758 26850 21810 26862
rect 21758 26786 21810 26798
rect 31502 26850 31554 26862
rect 31502 26786 31554 26798
rect 34638 26850 34690 26862
rect 34638 26786 34690 26798
rect 40686 26850 40738 26862
rect 40686 26786 40738 26798
rect 42030 26850 42082 26862
rect 42030 26786 42082 26798
rect 44270 26850 44322 26862
rect 44270 26786 44322 26798
rect 45054 26850 45106 26862
rect 45054 26786 45106 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 7086 26514 7138 26526
rect 7086 26450 7138 26462
rect 13358 26514 13410 26526
rect 13358 26450 13410 26462
rect 14590 26514 14642 26526
rect 14590 26450 14642 26462
rect 14814 26514 14866 26526
rect 14814 26450 14866 26462
rect 15934 26514 15986 26526
rect 15934 26450 15986 26462
rect 16382 26514 16434 26526
rect 19966 26514 20018 26526
rect 19058 26462 19070 26514
rect 19122 26462 19134 26514
rect 16382 26450 16434 26462
rect 19966 26450 20018 26462
rect 21086 26514 21138 26526
rect 21086 26450 21138 26462
rect 22766 26514 22818 26526
rect 22766 26450 22818 26462
rect 25230 26514 25282 26526
rect 25230 26450 25282 26462
rect 25342 26514 25394 26526
rect 28814 26514 28866 26526
rect 28466 26462 28478 26514
rect 28530 26462 28542 26514
rect 25342 26450 25394 26462
rect 28814 26450 28866 26462
rect 30606 26514 30658 26526
rect 33182 26514 33234 26526
rect 31266 26462 31278 26514
rect 31330 26462 31342 26514
rect 30606 26450 30658 26462
rect 33182 26450 33234 26462
rect 36206 26514 36258 26526
rect 36206 26450 36258 26462
rect 36430 26514 36482 26526
rect 36430 26450 36482 26462
rect 37214 26514 37266 26526
rect 37214 26450 37266 26462
rect 38110 26514 38162 26526
rect 38110 26450 38162 26462
rect 38446 26514 38498 26526
rect 38446 26450 38498 26462
rect 41918 26514 41970 26526
rect 41918 26450 41970 26462
rect 42814 26514 42866 26526
rect 42814 26450 42866 26462
rect 43374 26514 43426 26526
rect 43374 26450 43426 26462
rect 43710 26514 43762 26526
rect 43710 26450 43762 26462
rect 45054 26514 45106 26526
rect 45054 26450 45106 26462
rect 45502 26514 45554 26526
rect 45502 26450 45554 26462
rect 50542 26514 50594 26526
rect 50542 26450 50594 26462
rect 51438 26514 51490 26526
rect 51438 26450 51490 26462
rect 53118 26514 53170 26526
rect 53118 26450 53170 26462
rect 55246 26514 55298 26526
rect 55246 26450 55298 26462
rect 57822 26514 57874 26526
rect 57822 26450 57874 26462
rect 7982 26402 8034 26414
rect 7982 26338 8034 26350
rect 13246 26402 13298 26414
rect 13246 26338 13298 26350
rect 15038 26402 15090 26414
rect 22990 26402 23042 26414
rect 18050 26350 18062 26402
rect 18114 26350 18126 26402
rect 18386 26350 18398 26402
rect 18450 26350 18462 26402
rect 15038 26338 15090 26350
rect 22990 26338 23042 26350
rect 23102 26402 23154 26414
rect 23102 26338 23154 26350
rect 29710 26402 29762 26414
rect 29710 26338 29762 26350
rect 30158 26402 30210 26414
rect 36542 26402 36594 26414
rect 30930 26350 30942 26402
rect 30994 26350 31006 26402
rect 35746 26350 35758 26402
rect 35810 26350 35822 26402
rect 30158 26338 30210 26350
rect 36542 26338 36594 26350
rect 39902 26402 39954 26414
rect 39902 26338 39954 26350
rect 42590 26402 42642 26414
rect 42590 26338 42642 26350
rect 43150 26402 43202 26414
rect 43150 26338 43202 26350
rect 44606 26402 44658 26414
rect 44606 26338 44658 26350
rect 47854 26402 47906 26414
rect 51214 26402 51266 26414
rect 49074 26350 49086 26402
rect 49138 26350 49150 26402
rect 47854 26338 47906 26350
rect 51214 26338 51266 26350
rect 51662 26402 51714 26414
rect 51662 26338 51714 26350
rect 51774 26402 51826 26414
rect 51774 26338 51826 26350
rect 52782 26402 52834 26414
rect 52782 26338 52834 26350
rect 52894 26402 52946 26414
rect 57150 26402 57202 26414
rect 54338 26350 54350 26402
rect 54402 26350 54414 26402
rect 52894 26338 52946 26350
rect 57150 26338 57202 26350
rect 5966 26290 6018 26302
rect 1810 26238 1822 26290
rect 1874 26238 1886 26290
rect 5966 26226 6018 26238
rect 6414 26290 6466 26302
rect 6414 26226 6466 26238
rect 6638 26290 6690 26302
rect 9662 26290 9714 26302
rect 12014 26290 12066 26302
rect 8194 26238 8206 26290
rect 8258 26238 8270 26290
rect 8418 26238 8430 26290
rect 8482 26238 8494 26290
rect 9986 26238 9998 26290
rect 10050 26238 10062 26290
rect 6638 26226 6690 26238
rect 9662 26226 9714 26238
rect 12014 26226 12066 26238
rect 12238 26290 12290 26302
rect 12238 26226 12290 26238
rect 13582 26290 13634 26302
rect 13582 26226 13634 26238
rect 14366 26290 14418 26302
rect 14366 26226 14418 26238
rect 16718 26290 16770 26302
rect 16718 26226 16770 26238
rect 17502 26290 17554 26302
rect 17502 26226 17554 26238
rect 17838 26290 17890 26302
rect 21758 26290 21810 26302
rect 19282 26238 19294 26290
rect 19346 26238 19358 26290
rect 17838 26226 17890 26238
rect 21758 26226 21810 26238
rect 21982 26290 22034 26302
rect 21982 26226 22034 26238
rect 25454 26290 25506 26302
rect 25454 26226 25506 26238
rect 25902 26290 25954 26302
rect 25902 26226 25954 26238
rect 28142 26290 28194 26302
rect 28142 26226 28194 26238
rect 28926 26290 28978 26302
rect 28926 26226 28978 26238
rect 29150 26290 29202 26302
rect 29150 26226 29202 26238
rect 29486 26290 29538 26302
rect 42478 26290 42530 26302
rect 31490 26238 31502 26290
rect 31554 26238 31566 26290
rect 34402 26238 34414 26290
rect 34466 26238 34478 26290
rect 35522 26238 35534 26290
rect 35586 26238 35598 26290
rect 39218 26238 39230 26290
rect 39282 26238 39294 26290
rect 29486 26226 29538 26238
rect 42478 26226 42530 26238
rect 43038 26290 43090 26302
rect 50654 26290 50706 26302
rect 48850 26238 48862 26290
rect 48914 26238 48926 26290
rect 50306 26238 50318 26290
rect 50370 26238 50382 26290
rect 43038 26226 43090 26238
rect 50654 26226 50706 26238
rect 51102 26290 51154 26302
rect 51102 26226 51154 26238
rect 54014 26290 54066 26302
rect 54014 26226 54066 26238
rect 55134 26290 55186 26302
rect 55134 26226 55186 26238
rect 55470 26290 55522 26302
rect 55470 26226 55522 26238
rect 55582 26290 55634 26302
rect 55582 26226 55634 26238
rect 57486 26290 57538 26302
rect 58034 26238 58046 26290
rect 58098 26238 58110 26290
rect 57486 26226 57538 26238
rect 5406 26178 5458 26190
rect 2482 26126 2494 26178
rect 2546 26126 2558 26178
rect 4610 26126 4622 26178
rect 4674 26126 4686 26178
rect 5406 26114 5458 26126
rect 6190 26178 6242 26190
rect 7310 26178 7362 26190
rect 6962 26126 6974 26178
rect 7026 26126 7038 26178
rect 6190 26114 6242 26126
rect 7310 26114 7362 26126
rect 9550 26178 9602 26190
rect 20638 26178 20690 26190
rect 23550 26178 23602 26190
rect 15474 26126 15486 26178
rect 15538 26126 15550 26178
rect 22418 26126 22430 26178
rect 22482 26126 22494 26178
rect 9550 26114 9602 26126
rect 20638 26114 20690 26126
rect 23550 26114 23602 26126
rect 24110 26178 24162 26190
rect 24110 26114 24162 26126
rect 24558 26178 24610 26190
rect 24558 26114 24610 26126
rect 26238 26178 26290 26190
rect 26238 26114 26290 26126
rect 27806 26178 27858 26190
rect 27806 26114 27858 26126
rect 33742 26178 33794 26190
rect 33742 26114 33794 26126
rect 33966 26178 34018 26190
rect 33966 26114 34018 26126
rect 35086 26178 35138 26190
rect 40350 26178 40402 26190
rect 38994 26126 39006 26178
rect 39058 26126 39070 26178
rect 35086 26114 35138 26126
rect 40350 26114 40402 26126
rect 41134 26178 41186 26190
rect 41134 26114 41186 26126
rect 44158 26178 44210 26190
rect 44158 26114 44210 26126
rect 47294 26178 47346 26190
rect 53678 26178 53730 26190
rect 47954 26126 47966 26178
rect 48018 26126 48030 26178
rect 47294 26114 47346 26126
rect 53678 26114 53730 26126
rect 55358 26178 55410 26190
rect 55358 26114 55410 26126
rect 56702 26178 56754 26190
rect 56702 26114 56754 26126
rect 5070 26066 5122 26078
rect 5070 26002 5122 26014
rect 5182 26066 5234 26078
rect 5182 26002 5234 26014
rect 5630 26066 5682 26078
rect 5630 26002 5682 26014
rect 5742 26066 5794 26078
rect 14926 26066 14978 26078
rect 47630 26066 47682 26078
rect 11666 26014 11678 26066
rect 11730 26014 11742 26066
rect 47058 26014 47070 26066
rect 47122 26063 47134 26066
rect 47282 26063 47294 26066
rect 47122 26017 47294 26063
rect 47122 26014 47134 26017
rect 47282 26014 47294 26017
rect 47346 26014 47358 26066
rect 5742 26002 5794 26014
rect 14926 26002 14978 26014
rect 47630 26002 47682 26014
rect 51774 26066 51826 26078
rect 51774 26002 51826 26014
rect 56590 26066 56642 26078
rect 56590 26002 56642 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 6190 25730 6242 25742
rect 6190 25666 6242 25678
rect 13918 25730 13970 25742
rect 13918 25666 13970 25678
rect 14254 25730 14306 25742
rect 14254 25666 14306 25678
rect 19518 25730 19570 25742
rect 19518 25666 19570 25678
rect 28254 25730 28306 25742
rect 28254 25666 28306 25678
rect 48750 25730 48802 25742
rect 48750 25666 48802 25678
rect 2270 25618 2322 25630
rect 2270 25554 2322 25566
rect 3838 25618 3890 25630
rect 3838 25554 3890 25566
rect 7982 25618 8034 25630
rect 7982 25554 8034 25566
rect 15486 25618 15538 25630
rect 15486 25554 15538 25566
rect 16046 25618 16098 25630
rect 16046 25554 16098 25566
rect 18398 25618 18450 25630
rect 18398 25554 18450 25566
rect 19070 25618 19122 25630
rect 28478 25618 28530 25630
rect 21746 25566 21758 25618
rect 21810 25566 21822 25618
rect 24098 25566 24110 25618
rect 24162 25566 24174 25618
rect 19070 25554 19122 25566
rect 28478 25554 28530 25566
rect 34190 25618 34242 25630
rect 34190 25554 34242 25566
rect 38446 25618 38498 25630
rect 38446 25554 38498 25566
rect 39902 25618 39954 25630
rect 39902 25554 39954 25566
rect 42366 25618 42418 25630
rect 42366 25554 42418 25566
rect 43486 25618 43538 25630
rect 43486 25554 43538 25566
rect 43822 25618 43874 25630
rect 51998 25618 52050 25630
rect 51314 25566 51326 25618
rect 51378 25566 51390 25618
rect 43822 25554 43874 25566
rect 51998 25554 52050 25566
rect 54910 25618 54962 25630
rect 56018 25566 56030 25618
rect 56082 25566 56094 25618
rect 58146 25566 58158 25618
rect 58210 25566 58222 25618
rect 54910 25554 54962 25566
rect 1710 25506 1762 25518
rect 3726 25506 3778 25518
rect 5854 25506 5906 25518
rect 3154 25454 3166 25506
rect 3218 25454 3230 25506
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 1710 25442 1762 25454
rect 3726 25442 3778 25454
rect 5854 25442 5906 25454
rect 6078 25506 6130 25518
rect 6078 25442 6130 25454
rect 6302 25506 6354 25518
rect 7646 25506 7698 25518
rect 6962 25454 6974 25506
rect 7026 25454 7038 25506
rect 6302 25442 6354 25454
rect 7646 25442 7698 25454
rect 10334 25506 10386 25518
rect 10334 25442 10386 25454
rect 15038 25506 15090 25518
rect 15038 25442 15090 25454
rect 19294 25506 19346 25518
rect 19294 25442 19346 25454
rect 20302 25506 20354 25518
rect 24558 25506 24610 25518
rect 26798 25506 26850 25518
rect 29822 25506 29874 25518
rect 32062 25506 32114 25518
rect 37886 25506 37938 25518
rect 39790 25506 39842 25518
rect 22418 25454 22430 25506
rect 22482 25454 22494 25506
rect 26226 25454 26238 25506
rect 26290 25454 26302 25506
rect 28018 25454 28030 25506
rect 28082 25454 28094 25506
rect 30370 25454 30382 25506
rect 30434 25454 30446 25506
rect 35410 25454 35422 25506
rect 35474 25454 35486 25506
rect 39330 25454 39342 25506
rect 39394 25454 39406 25506
rect 20302 25442 20354 25454
rect 24558 25442 24610 25454
rect 26798 25442 26850 25454
rect 29822 25442 29874 25454
rect 32062 25442 32114 25454
rect 37886 25442 37938 25454
rect 39790 25442 39842 25454
rect 40574 25506 40626 25518
rect 40574 25442 40626 25454
rect 41470 25506 41522 25518
rect 48974 25506 49026 25518
rect 41906 25454 41918 25506
rect 41970 25454 41982 25506
rect 41470 25442 41522 25454
rect 48974 25442 49026 25454
rect 49198 25506 49250 25518
rect 49198 25442 49250 25454
rect 49870 25506 49922 25518
rect 49870 25442 49922 25454
rect 51662 25506 51714 25518
rect 52994 25454 53006 25506
rect 53058 25454 53070 25506
rect 55234 25454 55246 25506
rect 55298 25454 55310 25506
rect 51662 25442 51714 25454
rect 2718 25394 2770 25406
rect 2718 25330 2770 25342
rect 5630 25394 5682 25406
rect 21310 25394 21362 25406
rect 26910 25394 26962 25406
rect 6738 25342 6750 25394
rect 6802 25342 6814 25394
rect 9986 25342 9998 25394
rect 10050 25342 10062 25394
rect 22642 25342 22654 25394
rect 22706 25342 22718 25394
rect 5630 25330 5682 25342
rect 21310 25330 21362 25342
rect 26910 25330 26962 25342
rect 27246 25394 27298 25406
rect 27246 25330 27298 25342
rect 27470 25394 27522 25406
rect 28590 25394 28642 25406
rect 38558 25394 38610 25406
rect 27682 25342 27694 25394
rect 27746 25391 27758 25394
rect 28018 25391 28030 25394
rect 27746 25345 28030 25391
rect 27746 25342 27758 25345
rect 28018 25342 28030 25345
rect 28082 25342 28094 25394
rect 30594 25342 30606 25394
rect 30658 25342 30670 25394
rect 27470 25330 27522 25342
rect 28590 25330 28642 25342
rect 38558 25330 38610 25342
rect 40238 25394 40290 25406
rect 40238 25330 40290 25342
rect 40798 25394 40850 25406
rect 40798 25330 40850 25342
rect 45166 25394 45218 25406
rect 45166 25330 45218 25342
rect 49422 25394 49474 25406
rect 49422 25330 49474 25342
rect 50318 25394 50370 25406
rect 50318 25330 50370 25342
rect 50542 25394 50594 25406
rect 51326 25394 51378 25406
rect 51202 25342 51214 25394
rect 51266 25342 51278 25394
rect 50542 25330 50594 25342
rect 51326 25330 51378 25342
rect 51438 25394 51490 25406
rect 51438 25330 51490 25342
rect 52110 25394 52162 25406
rect 52110 25330 52162 25342
rect 52670 25394 52722 25406
rect 52670 25330 52722 25342
rect 52782 25394 52834 25406
rect 52782 25330 52834 25342
rect 53454 25394 53506 25406
rect 53454 25330 53506 25342
rect 3950 25282 4002 25294
rect 3378 25230 3390 25282
rect 3442 25230 3454 25282
rect 3950 25218 4002 25230
rect 4846 25282 4898 25294
rect 4846 25218 4898 25230
rect 14142 25282 14194 25294
rect 17950 25282 18002 25294
rect 25006 25282 25058 25294
rect 14690 25230 14702 25282
rect 14754 25230 14766 25282
rect 19842 25230 19854 25282
rect 19906 25230 19918 25282
rect 14142 25218 14194 25230
rect 17950 25218 18002 25230
rect 25006 25218 25058 25230
rect 27358 25282 27410 25294
rect 27358 25218 27410 25230
rect 29486 25282 29538 25294
rect 29486 25218 29538 25230
rect 31278 25282 31330 25294
rect 31278 25218 31330 25230
rect 31502 25282 31554 25294
rect 31502 25218 31554 25230
rect 33966 25282 34018 25294
rect 33966 25218 34018 25230
rect 34750 25282 34802 25294
rect 37774 25282 37826 25294
rect 35186 25230 35198 25282
rect 35250 25230 35262 25282
rect 34750 25218 34802 25230
rect 37774 25218 37826 25230
rect 38334 25282 38386 25294
rect 38334 25218 38386 25230
rect 40350 25282 40402 25294
rect 40350 25218 40402 25230
rect 40910 25282 40962 25294
rect 40910 25218 40962 25230
rect 42926 25282 42978 25294
rect 42926 25218 42978 25230
rect 44270 25282 44322 25294
rect 44270 25218 44322 25230
rect 45502 25282 45554 25294
rect 48078 25282 48130 25294
rect 47730 25230 47742 25282
rect 47794 25230 47806 25282
rect 45502 25218 45554 25230
rect 48078 25218 48130 25230
rect 48302 25282 48354 25294
rect 48302 25218 48354 25230
rect 50206 25282 50258 25294
rect 50206 25218 50258 25230
rect 53342 25282 53394 25294
rect 53342 25218 53394 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 2718 24946 2770 24958
rect 2034 24894 2046 24946
rect 2098 24894 2110 24946
rect 2718 24882 2770 24894
rect 3502 24946 3554 24958
rect 3502 24882 3554 24894
rect 4398 24946 4450 24958
rect 4398 24882 4450 24894
rect 5518 24946 5570 24958
rect 5518 24882 5570 24894
rect 7758 24946 7810 24958
rect 7758 24882 7810 24894
rect 9662 24946 9714 24958
rect 9662 24882 9714 24894
rect 10110 24946 10162 24958
rect 10110 24882 10162 24894
rect 11118 24946 11170 24958
rect 11118 24882 11170 24894
rect 18734 24946 18786 24958
rect 18734 24882 18786 24894
rect 22878 24946 22930 24958
rect 22878 24882 22930 24894
rect 25678 24946 25730 24958
rect 25678 24882 25730 24894
rect 30158 24946 30210 24958
rect 30158 24882 30210 24894
rect 35086 24946 35138 24958
rect 35086 24882 35138 24894
rect 36094 24946 36146 24958
rect 40238 24946 40290 24958
rect 38770 24894 38782 24946
rect 38834 24894 38846 24946
rect 36094 24882 36146 24894
rect 40238 24882 40290 24894
rect 41246 24946 41298 24958
rect 41246 24882 41298 24894
rect 43038 24946 43090 24958
rect 43038 24882 43090 24894
rect 54686 24946 54738 24958
rect 54686 24882 54738 24894
rect 55358 24946 55410 24958
rect 55358 24882 55410 24894
rect 56926 24946 56978 24958
rect 56926 24882 56978 24894
rect 57486 24946 57538 24958
rect 58158 24946 58210 24958
rect 57810 24894 57822 24946
rect 57874 24894 57886 24946
rect 57486 24882 57538 24894
rect 58158 24882 58210 24894
rect 5742 24834 5794 24846
rect 4722 24782 4734 24834
rect 4786 24782 4798 24834
rect 5742 24770 5794 24782
rect 6190 24834 6242 24846
rect 6190 24770 6242 24782
rect 6302 24834 6354 24846
rect 6302 24770 6354 24782
rect 14926 24834 14978 24846
rect 14926 24770 14978 24782
rect 15598 24834 15650 24846
rect 15598 24770 15650 24782
rect 15710 24834 15762 24846
rect 15710 24770 15762 24782
rect 16270 24834 16322 24846
rect 16270 24770 16322 24782
rect 16494 24834 16546 24846
rect 16494 24770 16546 24782
rect 16606 24834 16658 24846
rect 16606 24770 16658 24782
rect 23662 24834 23714 24846
rect 23662 24770 23714 24782
rect 23998 24834 24050 24846
rect 23998 24770 24050 24782
rect 26126 24834 26178 24846
rect 34750 24834 34802 24846
rect 29138 24782 29150 24834
rect 29202 24782 29214 24834
rect 26126 24770 26178 24782
rect 34750 24770 34802 24782
rect 35422 24834 35474 24846
rect 39118 24834 39170 24846
rect 35746 24782 35758 24834
rect 35810 24782 35822 24834
rect 36418 24782 36430 24834
rect 36482 24782 36494 24834
rect 35422 24770 35474 24782
rect 39118 24770 39170 24782
rect 41022 24834 41074 24846
rect 54910 24834 54962 24846
rect 45826 24782 45838 24834
rect 45890 24782 45902 24834
rect 57138 24782 57150 24834
rect 57202 24782 57214 24834
rect 41022 24770 41074 24782
rect 54910 24770 54962 24782
rect 1710 24722 1762 24734
rect 1710 24658 1762 24670
rect 2382 24722 2434 24734
rect 2382 24658 2434 24670
rect 5294 24722 5346 24734
rect 5294 24658 5346 24670
rect 7310 24722 7362 24734
rect 17502 24722 17554 24734
rect 11442 24670 11454 24722
rect 11506 24670 11518 24722
rect 7310 24658 7362 24670
rect 17502 24658 17554 24670
rect 18062 24722 18114 24734
rect 22766 24722 22818 24734
rect 19282 24670 19294 24722
rect 19346 24670 19358 24722
rect 18062 24658 18114 24670
rect 22766 24658 22818 24670
rect 25454 24722 25506 24734
rect 25454 24658 25506 24670
rect 25902 24722 25954 24734
rect 27358 24722 27410 24734
rect 26898 24670 26910 24722
rect 26962 24670 26974 24722
rect 25902 24658 25954 24670
rect 27358 24658 27410 24670
rect 27582 24722 27634 24734
rect 30046 24722 30098 24734
rect 27794 24670 27806 24722
rect 27858 24670 27870 24722
rect 28578 24670 28590 24722
rect 28642 24670 28654 24722
rect 27582 24658 27634 24670
rect 30046 24658 30098 24670
rect 30270 24722 30322 24734
rect 30270 24658 30322 24670
rect 33070 24722 33122 24734
rect 33070 24658 33122 24670
rect 33182 24722 33234 24734
rect 39342 24722 39394 24734
rect 33506 24670 33518 24722
rect 33570 24670 33582 24722
rect 33182 24658 33234 24670
rect 39342 24658 39394 24670
rect 40910 24722 40962 24734
rect 42366 24722 42418 24734
rect 42130 24670 42142 24722
rect 42194 24670 42206 24722
rect 40910 24658 40962 24670
rect 42366 24658 42418 24670
rect 42926 24722 42978 24734
rect 42926 24658 42978 24670
rect 43150 24722 43202 24734
rect 43150 24658 43202 24670
rect 43598 24722 43650 24734
rect 43598 24658 43650 24670
rect 43822 24722 43874 24734
rect 43822 24658 43874 24670
rect 44270 24722 44322 24734
rect 44270 24658 44322 24670
rect 44494 24722 44546 24734
rect 50654 24722 50706 24734
rect 45154 24670 45166 24722
rect 45218 24670 45230 24722
rect 50194 24670 50206 24722
rect 50258 24670 50270 24722
rect 44494 24658 44546 24670
rect 50654 24658 50706 24670
rect 50990 24722 51042 24734
rect 50990 24658 51042 24670
rect 51102 24722 51154 24734
rect 52446 24722 52498 24734
rect 53678 24722 53730 24734
rect 51426 24670 51438 24722
rect 51490 24670 51502 24722
rect 52770 24670 52782 24722
rect 52834 24670 52846 24722
rect 51102 24658 51154 24670
rect 52446 24658 52498 24670
rect 53678 24658 53730 24670
rect 55134 24722 55186 24734
rect 55570 24670 55582 24722
rect 55634 24670 55646 24722
rect 55134 24658 55186 24670
rect 3838 24610 3890 24622
rect 3838 24546 3890 24558
rect 5406 24610 5458 24622
rect 5406 24546 5458 24558
rect 6974 24610 7026 24622
rect 14814 24610 14866 24622
rect 23326 24610 23378 24622
rect 12226 24558 12238 24610
rect 12290 24558 12302 24610
rect 14354 24558 14366 24610
rect 14418 24558 14430 24610
rect 20066 24558 20078 24610
rect 20130 24558 20142 24610
rect 22194 24558 22206 24610
rect 22258 24558 22270 24610
rect 6974 24546 7026 24558
rect 14814 24546 14866 24558
rect 23326 24546 23378 24558
rect 24670 24610 24722 24622
rect 29822 24610 29874 24622
rect 28466 24558 28478 24610
rect 28530 24558 28542 24610
rect 24670 24546 24722 24558
rect 29822 24546 29874 24558
rect 38222 24610 38274 24622
rect 38222 24546 38274 24558
rect 44382 24610 44434 24622
rect 48974 24610 49026 24622
rect 52334 24610 52386 24622
rect 47954 24558 47966 24610
rect 48018 24558 48030 24610
rect 49746 24558 49758 24610
rect 49810 24558 49822 24610
rect 44382 24546 44434 24558
rect 48974 24546 49026 24558
rect 52334 24546 52386 24558
rect 53790 24610 53842 24622
rect 53790 24546 53842 24558
rect 55246 24610 55298 24622
rect 55246 24546 55298 24558
rect 56030 24610 56082 24622
rect 56030 24546 56082 24558
rect 6302 24498 6354 24510
rect 3826 24446 3838 24498
rect 3890 24495 3902 24498
rect 4050 24495 4062 24498
rect 3890 24449 4062 24495
rect 3890 24446 3902 24449
rect 4050 24446 4062 24449
rect 4114 24446 4126 24498
rect 6302 24434 6354 24446
rect 14702 24498 14754 24510
rect 14702 24434 14754 24446
rect 15710 24498 15762 24510
rect 15710 24434 15762 24446
rect 29598 24498 29650 24510
rect 29598 24434 29650 24446
rect 38446 24498 38498 24510
rect 38446 24434 38498 24446
rect 39566 24498 39618 24510
rect 39566 24434 39618 24446
rect 39790 24498 39842 24510
rect 55918 24498 55970 24510
rect 42466 24446 42478 24498
rect 42530 24446 42542 24498
rect 39790 24434 39842 24446
rect 55918 24434 55970 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 13806 24162 13858 24174
rect 13806 24098 13858 24110
rect 20638 24162 20690 24174
rect 20638 24098 20690 24110
rect 26686 24162 26738 24174
rect 32734 24162 32786 24174
rect 39902 24162 39954 24174
rect 30482 24110 30494 24162
rect 30546 24159 30558 24162
rect 31042 24159 31054 24162
rect 30546 24113 31054 24159
rect 30546 24110 30558 24113
rect 31042 24110 31054 24113
rect 31106 24110 31118 24162
rect 39218 24110 39230 24162
rect 39282 24159 39294 24162
rect 39778 24159 39790 24162
rect 39282 24113 39790 24159
rect 39282 24110 39294 24113
rect 39778 24110 39790 24113
rect 39842 24110 39854 24162
rect 26686 24098 26738 24110
rect 32734 24098 32786 24110
rect 39902 24098 39954 24110
rect 40574 24162 40626 24174
rect 40574 24098 40626 24110
rect 41358 24162 41410 24174
rect 41358 24098 41410 24110
rect 44942 24162 44994 24174
rect 44942 24098 44994 24110
rect 45278 24162 45330 24174
rect 45278 24098 45330 24110
rect 48078 24162 48130 24174
rect 53106 24110 53118 24162
rect 53170 24110 53182 24162
rect 48078 24098 48130 24110
rect 5070 24050 5122 24062
rect 12910 24050 12962 24062
rect 4610 23998 4622 24050
rect 4674 23998 4686 24050
rect 7074 23998 7086 24050
rect 7138 23998 7150 24050
rect 9202 23998 9214 24050
rect 9266 23998 9278 24050
rect 9538 23998 9550 24050
rect 9602 23998 9614 24050
rect 5070 23986 5122 23998
rect 12910 23986 12962 23998
rect 14254 24050 14306 24062
rect 19070 24050 19122 24062
rect 15586 23998 15598 24050
rect 15650 23998 15662 24050
rect 17714 23998 17726 24050
rect 17778 23998 17790 24050
rect 14254 23986 14306 23998
rect 19070 23986 19122 23998
rect 19966 24050 20018 24062
rect 19966 23986 20018 23998
rect 20750 24050 20802 24062
rect 29934 24050 29986 24062
rect 21410 23998 21422 24050
rect 21474 23998 21486 24050
rect 23538 23998 23550 24050
rect 23602 23998 23614 24050
rect 25666 23998 25678 24050
rect 25730 23998 25742 24050
rect 20750 23986 20802 23998
rect 29934 23986 29986 23998
rect 30606 24050 30658 24062
rect 30606 23986 30658 23998
rect 31054 24050 31106 24062
rect 31054 23986 31106 23998
rect 39790 24050 39842 24062
rect 39790 23986 39842 23998
rect 40350 24050 40402 24062
rect 54798 24050 54850 24062
rect 46610 23998 46622 24050
rect 46674 23998 46686 24050
rect 48626 23998 48638 24050
rect 48690 23998 48702 24050
rect 52882 23998 52894 24050
rect 52946 23998 52958 24050
rect 55794 23998 55806 24050
rect 55858 23998 55870 24050
rect 57922 23998 57934 24050
rect 57986 23998 57998 24050
rect 40350 23986 40402 23998
rect 54798 23986 54850 23998
rect 18062 23938 18114 23950
rect 1810 23886 1822 23938
rect 1874 23886 1886 23938
rect 5730 23886 5742 23938
rect 5794 23886 5806 23938
rect 6290 23886 6302 23938
rect 6354 23886 6366 23938
rect 12338 23886 12350 23938
rect 12402 23886 12414 23938
rect 14914 23886 14926 23938
rect 14978 23886 14990 23938
rect 18062 23874 18114 23886
rect 18622 23938 18674 23950
rect 21534 23938 21586 23950
rect 26238 23938 26290 23950
rect 19506 23886 19518 23938
rect 19570 23886 19582 23938
rect 22754 23886 22766 23938
rect 22818 23886 22830 23938
rect 18622 23874 18674 23886
rect 21534 23874 21586 23886
rect 26238 23874 26290 23886
rect 26462 23938 26514 23950
rect 26462 23874 26514 23886
rect 27358 23938 27410 23950
rect 27358 23874 27410 23886
rect 28030 23938 28082 23950
rect 28030 23874 28082 23886
rect 29486 23938 29538 23950
rect 34078 23938 34130 23950
rect 33842 23886 33854 23938
rect 33906 23886 33918 23938
rect 29486 23874 29538 23886
rect 34078 23874 34130 23886
rect 35086 23938 35138 23950
rect 37998 23938 38050 23950
rect 35522 23886 35534 23938
rect 35586 23886 35598 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 35086 23874 35138 23886
rect 37998 23874 38050 23886
rect 38894 23938 38946 23950
rect 38894 23874 38946 23886
rect 39118 23938 39170 23950
rect 39118 23874 39170 23886
rect 40798 23938 40850 23950
rect 40798 23874 40850 23886
rect 41470 23938 41522 23950
rect 41470 23874 41522 23886
rect 41694 23938 41746 23950
rect 41694 23874 41746 23886
rect 41806 23938 41858 23950
rect 41806 23874 41858 23886
rect 43710 23938 43762 23950
rect 43710 23874 43762 23886
rect 43934 23938 43986 23950
rect 47406 23938 47458 23950
rect 46946 23886 46958 23938
rect 47010 23886 47022 23938
rect 43934 23874 43986 23886
rect 47406 23874 47458 23886
rect 47630 23938 47682 23950
rect 47630 23874 47682 23886
rect 47854 23938 47906 23950
rect 47854 23874 47906 23886
rect 50654 23938 50706 23950
rect 50654 23874 50706 23886
rect 50878 23938 50930 23950
rect 50878 23874 50930 23886
rect 51102 23938 51154 23950
rect 53554 23886 53566 23938
rect 53618 23886 53630 23938
rect 55010 23886 55022 23938
rect 55074 23886 55086 23938
rect 51102 23874 51154 23886
rect 13470 23826 13522 23838
rect 2482 23774 2494 23826
rect 2546 23774 2558 23826
rect 11666 23774 11678 23826
rect 11730 23774 11742 23826
rect 13470 23762 13522 23774
rect 13694 23826 13746 23838
rect 13694 23762 13746 23774
rect 21982 23826 22034 23838
rect 21982 23762 22034 23774
rect 26014 23826 26066 23838
rect 29150 23826 29202 23838
rect 27682 23774 27694 23826
rect 27746 23774 27758 23826
rect 26014 23762 26066 23774
rect 29150 23762 29202 23774
rect 32734 23826 32786 23838
rect 32734 23762 32786 23774
rect 32846 23826 32898 23838
rect 32846 23762 32898 23774
rect 33182 23826 33234 23838
rect 33182 23762 33234 23774
rect 36990 23826 37042 23838
rect 36990 23762 37042 23774
rect 38558 23826 38610 23838
rect 38558 23762 38610 23774
rect 41022 23826 41074 23838
rect 41022 23762 41074 23774
rect 42478 23826 42530 23838
rect 50542 23826 50594 23838
rect 45602 23774 45614 23826
rect 45666 23774 45678 23826
rect 45938 23774 45950 23826
rect 46002 23774 46014 23826
rect 51426 23774 51438 23826
rect 51490 23774 51502 23826
rect 51874 23774 51886 23826
rect 51938 23774 51950 23826
rect 42478 23762 42530 23774
rect 50542 23762 50594 23774
rect 12798 23714 12850 23726
rect 5954 23662 5966 23714
rect 6018 23662 6030 23714
rect 12798 23650 12850 23662
rect 21422 23714 21474 23726
rect 21422 23650 21474 23662
rect 21758 23714 21810 23726
rect 21758 23650 21810 23662
rect 22430 23714 22482 23726
rect 22430 23650 22482 23662
rect 27134 23714 27186 23726
rect 27134 23650 27186 23662
rect 28142 23714 28194 23726
rect 28142 23650 28194 23662
rect 28366 23714 28418 23726
rect 28366 23650 28418 23662
rect 29262 23714 29314 23726
rect 29262 23650 29314 23662
rect 31950 23714 32002 23726
rect 36318 23714 36370 23726
rect 34738 23662 34750 23714
rect 34802 23662 34814 23714
rect 35746 23662 35758 23714
rect 35810 23662 35822 23714
rect 31950 23650 32002 23662
rect 36318 23650 36370 23662
rect 37326 23714 37378 23726
rect 37326 23650 37378 23662
rect 38110 23714 38162 23726
rect 38110 23650 38162 23662
rect 38222 23714 38274 23726
rect 38222 23650 38274 23662
rect 38782 23714 38834 23726
rect 38782 23650 38834 23662
rect 42590 23714 42642 23726
rect 42590 23650 42642 23662
rect 42814 23714 42866 23726
rect 42814 23650 42866 23662
rect 43262 23714 43314 23726
rect 43262 23650 43314 23662
rect 43374 23714 43426 23726
rect 43374 23650 43426 23662
rect 43486 23714 43538 23726
rect 43486 23650 43538 23662
rect 49086 23714 49138 23726
rect 49086 23650 49138 23662
rect 50318 23714 50370 23726
rect 50318 23650 50370 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 2606 23378 2658 23390
rect 2606 23314 2658 23326
rect 3726 23378 3778 23390
rect 8766 23378 8818 23390
rect 5618 23326 5630 23378
rect 5682 23326 5694 23378
rect 3726 23314 3778 23326
rect 8766 23314 8818 23326
rect 16830 23378 16882 23390
rect 16830 23314 16882 23326
rect 17390 23378 17442 23390
rect 17390 23314 17442 23326
rect 18174 23378 18226 23390
rect 18174 23314 18226 23326
rect 27694 23378 27746 23390
rect 27694 23314 27746 23326
rect 29710 23378 29762 23390
rect 29710 23314 29762 23326
rect 31278 23378 31330 23390
rect 42366 23378 42418 23390
rect 32498 23326 32510 23378
rect 32562 23326 32574 23378
rect 31278 23314 31330 23326
rect 42366 23314 42418 23326
rect 43150 23378 43202 23390
rect 43150 23314 43202 23326
rect 43486 23378 43538 23390
rect 43486 23314 43538 23326
rect 51214 23378 51266 23390
rect 57822 23378 57874 23390
rect 51986 23326 51998 23378
rect 52050 23326 52062 23378
rect 51214 23314 51266 23326
rect 57822 23314 57874 23326
rect 9662 23266 9714 23278
rect 4274 23214 4286 23266
rect 4338 23214 4350 23266
rect 5730 23214 5742 23266
rect 5794 23214 5806 23266
rect 7410 23214 7422 23266
rect 7474 23214 7486 23266
rect 9662 23202 9714 23214
rect 11678 23266 11730 23278
rect 11678 23202 11730 23214
rect 11902 23266 11954 23278
rect 27582 23266 27634 23278
rect 12338 23214 12350 23266
rect 12402 23214 12414 23266
rect 16482 23214 16494 23266
rect 16546 23214 16558 23266
rect 11902 23202 11954 23214
rect 27582 23202 27634 23214
rect 28814 23266 28866 23278
rect 28814 23202 28866 23214
rect 29038 23266 29090 23278
rect 29038 23202 29090 23214
rect 30494 23266 30546 23278
rect 30494 23202 30546 23214
rect 42814 23266 42866 23278
rect 42814 23202 42866 23214
rect 42926 23266 42978 23278
rect 48750 23266 48802 23278
rect 45602 23214 45614 23266
rect 45666 23214 45678 23266
rect 46050 23214 46062 23266
rect 46114 23214 46126 23266
rect 42926 23202 42978 23214
rect 48750 23202 48802 23214
rect 51326 23266 51378 23278
rect 51326 23202 51378 23214
rect 55582 23266 55634 23278
rect 55582 23202 55634 23214
rect 57150 23266 57202 23278
rect 57150 23202 57202 23214
rect 57486 23266 57538 23278
rect 57486 23202 57538 23214
rect 58158 23266 58210 23278
rect 58158 23202 58210 23214
rect 1710 23154 1762 23166
rect 1710 23090 1762 23102
rect 2942 23154 2994 23166
rect 2942 23090 2994 23102
rect 3278 23154 3330 23166
rect 3278 23090 3330 23102
rect 3614 23154 3666 23166
rect 3614 23090 3666 23102
rect 3950 23154 4002 23166
rect 6302 23154 6354 23166
rect 8878 23154 8930 23166
rect 4834 23102 4846 23154
rect 4898 23102 4910 23154
rect 5282 23102 5294 23154
rect 5346 23102 5358 23154
rect 7298 23102 7310 23154
rect 7362 23102 7374 23154
rect 3950 23090 4002 23102
rect 6302 23090 6354 23102
rect 8878 23090 8930 23102
rect 9550 23154 9602 23166
rect 9550 23090 9602 23102
rect 9886 23154 9938 23166
rect 9886 23090 9938 23102
rect 9998 23154 10050 23166
rect 11566 23154 11618 23166
rect 11330 23102 11342 23154
rect 11394 23102 11406 23154
rect 9998 23090 10050 23102
rect 11566 23090 11618 23102
rect 11790 23154 11842 23166
rect 11790 23090 11842 23102
rect 12686 23154 12738 23166
rect 22990 23154 23042 23166
rect 28702 23154 28754 23166
rect 17602 23102 17614 23154
rect 17666 23102 17678 23154
rect 19170 23102 19182 23154
rect 19234 23102 19246 23154
rect 23426 23102 23438 23154
rect 23490 23102 23502 23154
rect 12686 23090 12738 23102
rect 22990 23090 23042 23102
rect 28702 23090 28754 23102
rect 29486 23154 29538 23166
rect 29486 23090 29538 23102
rect 29710 23154 29762 23166
rect 29710 23090 29762 23102
rect 30046 23154 30098 23166
rect 30046 23090 30098 23102
rect 30606 23154 30658 23166
rect 30606 23090 30658 23102
rect 30830 23154 30882 23166
rect 30830 23090 30882 23102
rect 31502 23154 31554 23166
rect 33070 23154 33122 23166
rect 34638 23154 34690 23166
rect 32274 23102 32286 23154
rect 32338 23102 32350 23154
rect 33618 23102 33630 23154
rect 33682 23102 33694 23154
rect 31502 23090 31554 23102
rect 33070 23090 33122 23102
rect 34638 23090 34690 23102
rect 36878 23154 36930 23166
rect 36878 23090 36930 23102
rect 38894 23154 38946 23166
rect 40238 23154 40290 23166
rect 39330 23102 39342 23154
rect 39394 23102 39406 23154
rect 38894 23090 38946 23102
rect 40238 23090 40290 23102
rect 45278 23154 45330 23166
rect 45278 23090 45330 23102
rect 47518 23154 47570 23166
rect 50878 23154 50930 23166
rect 49410 23102 49422 23154
rect 49474 23102 49486 23154
rect 47518 23090 47570 23102
rect 50878 23090 50930 23102
rect 50990 23154 51042 23166
rect 50990 23090 51042 23102
rect 51886 23154 51938 23166
rect 55246 23154 55298 23166
rect 52210 23102 52222 23154
rect 52274 23102 52286 23154
rect 51886 23090 51938 23102
rect 55246 23090 55298 23102
rect 55358 23154 55410 23166
rect 55358 23090 55410 23102
rect 55694 23154 55746 23166
rect 55694 23090 55746 23102
rect 2270 23042 2322 23054
rect 2270 22978 2322 22990
rect 6638 23042 6690 23054
rect 6638 22978 6690 22990
rect 8430 23042 8482 23054
rect 8430 22978 8482 22990
rect 10558 23042 10610 23054
rect 10558 22978 10610 22990
rect 13134 23042 13186 23054
rect 13134 22978 13186 22990
rect 18734 23042 18786 23054
rect 22430 23042 22482 23054
rect 19842 22990 19854 23042
rect 19906 22990 19918 23042
rect 21970 22990 21982 23042
rect 22034 22990 22046 23042
rect 18734 22978 18786 22990
rect 22430 22978 22482 22990
rect 23886 23042 23938 23054
rect 23886 22978 23938 22990
rect 28366 23042 28418 23054
rect 28366 22978 28418 22990
rect 31390 23042 31442 23054
rect 34974 23042 35026 23054
rect 33954 22990 33966 23042
rect 34018 22990 34030 23042
rect 31390 22978 31442 22990
rect 34974 22978 35026 22990
rect 35758 23042 35810 23054
rect 35758 22978 35810 22990
rect 36206 23042 36258 23054
rect 39790 23042 39842 23054
rect 38098 22990 38110 23042
rect 38162 22990 38174 23042
rect 36206 22978 36258 22990
rect 39790 22978 39842 22990
rect 41134 23042 41186 23054
rect 41134 22978 41186 22990
rect 41470 23042 41522 23054
rect 41918 23042 41970 23054
rect 41682 22990 41694 23042
rect 41746 22990 41758 23042
rect 41470 22978 41522 22990
rect 8990 22930 9042 22942
rect 8990 22866 9042 22878
rect 30494 22930 30546 22942
rect 30494 22866 30546 22878
rect 34414 22930 34466 22942
rect 34414 22866 34466 22878
rect 34526 22930 34578 22942
rect 34526 22866 34578 22878
rect 35198 22930 35250 22942
rect 37102 22930 37154 22942
rect 35522 22878 35534 22930
rect 35586 22927 35598 22930
rect 36306 22927 36318 22930
rect 35586 22881 36318 22927
rect 35586 22878 35598 22881
rect 36306 22878 36318 22881
rect 36370 22878 36382 22930
rect 35198 22866 35250 22878
rect 37102 22866 37154 22878
rect 37326 22930 37378 22942
rect 37326 22866 37378 22878
rect 37550 22930 37602 22942
rect 41122 22878 41134 22930
rect 41186 22927 41198 22930
rect 41570 22927 41582 22930
rect 41186 22881 41582 22927
rect 41186 22878 41198 22881
rect 41570 22878 41582 22881
rect 41634 22878 41646 22930
rect 41697 22927 41743 22990
rect 41918 22978 41970 22990
rect 43934 23042 43986 23054
rect 43934 22978 43986 22990
rect 44382 23042 44434 23054
rect 44382 22978 44434 22990
rect 46622 23042 46674 23054
rect 46622 22978 46674 22990
rect 47070 23042 47122 23054
rect 47070 22978 47122 22990
rect 48078 23042 48130 23054
rect 55470 23042 55522 23054
rect 49634 22990 49646 23042
rect 49698 22990 49710 23042
rect 52658 22990 52670 23042
rect 52722 22990 52734 23042
rect 48078 22978 48130 22990
rect 55470 22978 55522 22990
rect 56702 23042 56754 23054
rect 56702 22978 56754 22990
rect 44942 22930 44994 22942
rect 41906 22927 41918 22930
rect 41697 22881 41918 22927
rect 41906 22878 41918 22881
rect 41970 22878 41982 22930
rect 44034 22878 44046 22930
rect 44098 22927 44110 22930
rect 44594 22927 44606 22930
rect 44098 22881 44606 22927
rect 44098 22878 44110 22881
rect 44594 22878 44606 22881
rect 44658 22878 44670 22930
rect 37550 22866 37602 22878
rect 44942 22866 44994 22878
rect 47742 22930 47794 22942
rect 47742 22866 47794 22878
rect 56590 22930 56642 22942
rect 56590 22866 56642 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 11454 22594 11506 22606
rect 20638 22594 20690 22606
rect 17042 22542 17054 22594
rect 17106 22591 17118 22594
rect 17602 22591 17614 22594
rect 17106 22545 17614 22591
rect 17106 22542 17118 22545
rect 17602 22542 17614 22545
rect 17666 22542 17678 22594
rect 11454 22530 11506 22542
rect 20638 22530 20690 22542
rect 33406 22594 33458 22606
rect 39230 22594 39282 22606
rect 37090 22542 37102 22594
rect 37154 22591 37166 22594
rect 37538 22591 37550 22594
rect 37154 22545 37550 22591
rect 37154 22542 37166 22545
rect 37538 22542 37550 22545
rect 37602 22542 37614 22594
rect 33406 22530 33458 22542
rect 39230 22530 39282 22542
rect 41694 22594 41746 22606
rect 41694 22530 41746 22542
rect 50094 22594 50146 22606
rect 50094 22530 50146 22542
rect 50990 22594 51042 22606
rect 50990 22530 51042 22542
rect 51326 22594 51378 22606
rect 51326 22530 51378 22542
rect 5070 22482 5122 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 5070 22418 5122 22430
rect 5742 22482 5794 22494
rect 5742 22418 5794 22430
rect 6190 22482 6242 22494
rect 6190 22418 6242 22430
rect 7534 22482 7586 22494
rect 7534 22418 7586 22430
rect 12014 22482 12066 22494
rect 12014 22418 12066 22430
rect 17054 22482 17106 22494
rect 17054 22418 17106 22430
rect 17950 22482 18002 22494
rect 27806 22482 27858 22494
rect 25330 22430 25342 22482
rect 25394 22430 25406 22482
rect 17950 22418 18002 22430
rect 27806 22418 27858 22430
rect 28142 22482 28194 22494
rect 31614 22482 31666 22494
rect 30930 22430 30942 22482
rect 30994 22430 31006 22482
rect 28142 22418 28194 22430
rect 31614 22418 31666 22430
rect 32622 22482 32674 22494
rect 32622 22418 32674 22430
rect 34414 22482 34466 22494
rect 34414 22418 34466 22430
rect 37550 22482 37602 22494
rect 37550 22418 37602 22430
rect 40686 22482 40738 22494
rect 40686 22418 40738 22430
rect 41246 22482 41298 22494
rect 41246 22418 41298 22430
rect 44942 22482 44994 22494
rect 44942 22418 44994 22430
rect 52782 22482 52834 22494
rect 56018 22430 56030 22482
rect 56082 22430 56094 22482
rect 58146 22430 58158 22482
rect 58210 22430 58222 22482
rect 52782 22418 52834 22430
rect 7982 22370 8034 22382
rect 11902 22370 11954 22382
rect 1810 22318 1822 22370
rect 1874 22318 1886 22370
rect 8306 22318 8318 22370
rect 8370 22318 8382 22370
rect 7982 22306 8034 22318
rect 11902 22306 11954 22318
rect 12238 22370 12290 22382
rect 12238 22306 12290 22318
rect 12350 22370 12402 22382
rect 12350 22306 12402 22318
rect 14478 22370 14530 22382
rect 14478 22306 14530 22318
rect 28030 22370 28082 22382
rect 31390 22370 31442 22382
rect 28578 22318 28590 22370
rect 28642 22318 28654 22370
rect 29138 22318 29150 22370
rect 29202 22318 29214 22370
rect 29698 22318 29710 22370
rect 29762 22318 29774 22370
rect 28030 22306 28082 22318
rect 31390 22306 31442 22318
rect 32062 22370 32114 22382
rect 32062 22306 32114 22318
rect 33182 22370 33234 22382
rect 33182 22306 33234 22318
rect 33630 22370 33682 22382
rect 33630 22306 33682 22318
rect 34526 22370 34578 22382
rect 34526 22306 34578 22318
rect 38558 22370 38610 22382
rect 38558 22306 38610 22318
rect 41806 22370 41858 22382
rect 41806 22306 41858 22318
rect 43038 22370 43090 22382
rect 43038 22306 43090 22318
rect 45502 22370 45554 22382
rect 45502 22306 45554 22318
rect 46286 22370 46338 22382
rect 54910 22370 54962 22382
rect 50418 22318 50430 22370
rect 50482 22318 50494 22370
rect 51986 22318 51998 22370
rect 52050 22318 52062 22370
rect 55234 22318 55246 22370
rect 55298 22318 55310 22370
rect 46286 22306 46338 22318
rect 54910 22306 54962 22318
rect 7870 22258 7922 22270
rect 2482 22206 2494 22258
rect 2546 22206 2558 22258
rect 7870 22194 7922 22206
rect 11342 22258 11394 22270
rect 11342 22194 11394 22206
rect 14814 22258 14866 22270
rect 14814 22194 14866 22206
rect 15262 22258 15314 22270
rect 15262 22194 15314 22206
rect 15934 22258 15986 22270
rect 15934 22194 15986 22206
rect 18734 22258 18786 22270
rect 18734 22194 18786 22206
rect 20750 22258 20802 22270
rect 20750 22194 20802 22206
rect 22318 22258 22370 22270
rect 30606 22258 30658 22270
rect 29810 22206 29822 22258
rect 29874 22206 29886 22258
rect 22318 22194 22370 22206
rect 30606 22194 30658 22206
rect 30830 22258 30882 22270
rect 30830 22194 30882 22206
rect 32958 22258 33010 22270
rect 32958 22194 33010 22206
rect 34750 22258 34802 22270
rect 34750 22194 34802 22206
rect 38334 22258 38386 22270
rect 38334 22194 38386 22206
rect 38894 22258 38946 22270
rect 38894 22194 38946 22206
rect 39118 22258 39170 22270
rect 39118 22194 39170 22206
rect 39454 22258 39506 22270
rect 39454 22194 39506 22206
rect 39790 22258 39842 22270
rect 39790 22194 39842 22206
rect 40238 22258 40290 22270
rect 40238 22194 40290 22206
rect 42366 22258 42418 22270
rect 42366 22194 42418 22206
rect 43150 22258 43202 22270
rect 43150 22194 43202 22206
rect 43598 22258 43650 22270
rect 43598 22194 43650 22206
rect 51662 22258 51714 22270
rect 51662 22194 51714 22206
rect 51774 22258 51826 22270
rect 51774 22194 51826 22206
rect 52670 22258 52722 22270
rect 52670 22194 52722 22206
rect 52894 22258 52946 22270
rect 54450 22206 54462 22258
rect 54514 22206 54526 22258
rect 52894 22194 52946 22206
rect 9214 22146 9266 22158
rect 9214 22082 9266 22094
rect 9326 22146 9378 22158
rect 9326 22082 9378 22094
rect 9438 22146 9490 22158
rect 9438 22082 9490 22094
rect 9662 22146 9714 22158
rect 9662 22082 9714 22094
rect 11454 22146 11506 22158
rect 11454 22082 11506 22094
rect 12910 22146 12962 22158
rect 12910 22082 12962 22094
rect 13470 22146 13522 22158
rect 14254 22146 14306 22158
rect 13794 22094 13806 22146
rect 13858 22094 13870 22146
rect 13470 22082 13522 22094
rect 14254 22082 14306 22094
rect 14702 22146 14754 22158
rect 14702 22082 14754 22094
rect 15150 22146 15202 22158
rect 15150 22082 15202 22094
rect 16270 22146 16322 22158
rect 16270 22082 16322 22094
rect 17502 22146 17554 22158
rect 17502 22082 17554 22094
rect 19294 22146 19346 22158
rect 19294 22082 19346 22094
rect 22430 22146 22482 22158
rect 22430 22082 22482 22094
rect 25790 22146 25842 22158
rect 25790 22082 25842 22094
rect 28254 22146 28306 22158
rect 31838 22146 31890 22158
rect 29362 22094 29374 22146
rect 29426 22094 29438 22146
rect 28254 22082 28306 22094
rect 31838 22082 31890 22094
rect 31950 22146 32002 22158
rect 31950 22082 32002 22094
rect 34078 22146 34130 22158
rect 34078 22082 34130 22094
rect 34302 22146 34354 22158
rect 34302 22082 34354 22094
rect 35534 22146 35586 22158
rect 36318 22146 36370 22158
rect 35858 22094 35870 22146
rect 35922 22094 35934 22146
rect 35534 22082 35586 22094
rect 36318 22082 36370 22094
rect 37102 22146 37154 22158
rect 37102 22082 37154 22094
rect 41694 22146 41746 22158
rect 41694 22082 41746 22094
rect 42478 22146 42530 22158
rect 42478 22082 42530 22094
rect 42590 22146 42642 22158
rect 42590 22082 42642 22094
rect 44046 22146 44098 22158
rect 44046 22082 44098 22094
rect 45838 22146 45890 22158
rect 45838 22082 45890 22094
rect 46734 22146 46786 22158
rect 46734 22082 46786 22094
rect 50206 22146 50258 22158
rect 50206 22082 50258 22094
rect 51214 22146 51266 22158
rect 51214 22082 51266 22094
rect 53454 22146 53506 22158
rect 54126 22146 54178 22158
rect 53778 22094 53790 22146
rect 53842 22094 53854 22146
rect 53454 22082 53506 22094
rect 54126 22082 54178 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 1710 21810 1762 21822
rect 1710 21746 1762 21758
rect 2942 21810 2994 21822
rect 2942 21746 2994 21758
rect 3390 21810 3442 21822
rect 3390 21746 3442 21758
rect 3838 21810 3890 21822
rect 3838 21746 3890 21758
rect 3950 21810 4002 21822
rect 3950 21746 4002 21758
rect 4734 21810 4786 21822
rect 4734 21746 4786 21758
rect 9774 21810 9826 21822
rect 13358 21810 13410 21822
rect 13010 21758 13022 21810
rect 13074 21758 13086 21810
rect 9774 21746 9826 21758
rect 13358 21746 13410 21758
rect 13694 21810 13746 21822
rect 13694 21746 13746 21758
rect 15598 21810 15650 21822
rect 15598 21746 15650 21758
rect 17614 21810 17666 21822
rect 17614 21746 17666 21758
rect 20974 21810 21026 21822
rect 20974 21746 21026 21758
rect 21086 21810 21138 21822
rect 21086 21746 21138 21758
rect 21198 21810 21250 21822
rect 21198 21746 21250 21758
rect 28702 21810 28754 21822
rect 28702 21746 28754 21758
rect 29150 21810 29202 21822
rect 29150 21746 29202 21758
rect 29598 21810 29650 21822
rect 29598 21746 29650 21758
rect 29934 21810 29986 21822
rect 29934 21746 29986 21758
rect 30942 21810 30994 21822
rect 30942 21746 30994 21758
rect 31502 21810 31554 21822
rect 34414 21810 34466 21822
rect 31502 21746 31554 21758
rect 32174 21754 32226 21766
rect 4510 21698 4562 21710
rect 4510 21634 4562 21646
rect 4846 21698 4898 21710
rect 4846 21634 4898 21646
rect 5742 21698 5794 21710
rect 5742 21634 5794 21646
rect 6414 21698 6466 21710
rect 6414 21634 6466 21646
rect 6638 21698 6690 21710
rect 6638 21634 6690 21646
rect 8990 21698 9042 21710
rect 8990 21634 9042 21646
rect 11454 21698 11506 21710
rect 11454 21634 11506 21646
rect 12686 21698 12738 21710
rect 17502 21698 17554 21710
rect 16146 21646 16158 21698
rect 16210 21646 16222 21698
rect 16706 21646 16718 21698
rect 16770 21646 16782 21698
rect 12686 21634 12738 21646
rect 17502 21634 17554 21646
rect 18174 21698 18226 21710
rect 18174 21634 18226 21646
rect 18398 21698 18450 21710
rect 18398 21634 18450 21646
rect 18510 21698 18562 21710
rect 18510 21634 18562 21646
rect 21422 21698 21474 21710
rect 26910 21698 26962 21710
rect 22530 21646 22542 21698
rect 22594 21646 22606 21698
rect 21422 21634 21474 21646
rect 26910 21634 26962 21646
rect 28478 21698 28530 21710
rect 28478 21634 28530 21646
rect 30606 21698 30658 21710
rect 30606 21634 30658 21646
rect 30718 21698 30770 21710
rect 34414 21746 34466 21758
rect 34862 21810 34914 21822
rect 34862 21746 34914 21758
rect 40014 21810 40066 21822
rect 40014 21746 40066 21758
rect 40238 21810 40290 21822
rect 40238 21746 40290 21758
rect 41022 21810 41074 21822
rect 49534 21810 49586 21822
rect 49186 21758 49198 21810
rect 49250 21758 49262 21810
rect 41022 21746 41074 21758
rect 49534 21746 49586 21758
rect 50318 21810 50370 21822
rect 52894 21810 52946 21822
rect 51090 21758 51102 21810
rect 51154 21758 51166 21810
rect 50318 21746 50370 21758
rect 52894 21746 52946 21758
rect 55246 21810 55298 21822
rect 55246 21746 55298 21758
rect 57150 21810 57202 21822
rect 57150 21746 57202 21758
rect 57598 21810 57650 21822
rect 58158 21810 58210 21822
rect 57810 21758 57822 21810
rect 57874 21758 57886 21810
rect 57598 21746 57650 21758
rect 58158 21746 58210 21758
rect 32174 21690 32226 21702
rect 32286 21698 32338 21710
rect 30718 21634 30770 21646
rect 32286 21634 32338 21646
rect 39566 21698 39618 21710
rect 39566 21634 39618 21646
rect 41470 21698 41522 21710
rect 50094 21698 50146 21710
rect 54686 21698 54738 21710
rect 46050 21646 46062 21698
rect 46114 21646 46126 21698
rect 52434 21646 52446 21698
rect 52498 21646 52510 21698
rect 41470 21634 41522 21646
rect 50094 21634 50146 21646
rect 54686 21634 54738 21646
rect 2606 21586 2658 21598
rect 2606 21522 2658 21534
rect 3726 21586 3778 21598
rect 3726 21522 3778 21534
rect 4398 21586 4450 21598
rect 4398 21522 4450 21534
rect 5294 21586 5346 21598
rect 8878 21586 8930 21598
rect 8306 21534 8318 21586
rect 8370 21534 8382 21586
rect 5294 21522 5346 21534
rect 8878 21522 8930 21534
rect 9438 21586 9490 21598
rect 9438 21522 9490 21534
rect 9886 21586 9938 21598
rect 9886 21522 9938 21534
rect 10110 21586 10162 21598
rect 12350 21586 12402 21598
rect 10770 21534 10782 21586
rect 10834 21534 10846 21586
rect 11218 21534 11230 21586
rect 11282 21534 11294 21586
rect 10110 21522 10162 21534
rect 12350 21522 12402 21534
rect 14254 21586 14306 21598
rect 14254 21522 14306 21534
rect 14590 21586 14642 21598
rect 14590 21522 14642 21534
rect 17390 21586 17442 21598
rect 17390 21522 17442 21534
rect 18062 21586 18114 21598
rect 18062 21522 18114 21534
rect 18958 21586 19010 21598
rect 20862 21586 20914 21598
rect 28030 21586 28082 21598
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 21858 21534 21870 21586
rect 21922 21534 21934 21586
rect 26002 21534 26014 21586
rect 26066 21534 26078 21586
rect 18958 21522 19010 21534
rect 20862 21522 20914 21534
rect 28030 21522 28082 21534
rect 28366 21586 28418 21598
rect 28366 21522 28418 21534
rect 29486 21586 29538 21598
rect 29486 21522 29538 21534
rect 29710 21586 29762 21598
rect 29710 21522 29762 21534
rect 31278 21586 31330 21598
rect 31278 21522 31330 21534
rect 31390 21586 31442 21598
rect 38110 21586 38162 21598
rect 31826 21534 31838 21586
rect 31890 21534 31902 21586
rect 31390 21522 31442 21534
rect 38110 21522 38162 21534
rect 38894 21586 38946 21598
rect 38894 21522 38946 21534
rect 39118 21586 39170 21598
rect 39118 21522 39170 21534
rect 39790 21586 39842 21598
rect 39790 21522 39842 21534
rect 40350 21586 40402 21598
rect 40350 21522 40402 21534
rect 41246 21586 41298 21598
rect 50430 21586 50482 21598
rect 42018 21534 42030 21586
rect 42082 21534 42094 21586
rect 45378 21534 45390 21586
rect 45442 21534 45454 21586
rect 41246 21522 41298 21534
rect 50430 21522 50482 21534
rect 50542 21586 50594 21598
rect 54910 21586 54962 21598
rect 51538 21534 51550 21586
rect 51602 21534 51614 21586
rect 52098 21534 52110 21586
rect 52162 21534 52174 21586
rect 50542 21522 50594 21534
rect 54910 21522 54962 21534
rect 55134 21586 55186 21598
rect 55134 21522 55186 21534
rect 2270 21474 2322 21486
rect 2270 21410 2322 21422
rect 15150 21474 15202 21486
rect 25342 21474 25394 21486
rect 33182 21474 33234 21486
rect 24658 21422 24670 21474
rect 24722 21422 24734 21474
rect 26674 21422 26686 21474
rect 26738 21422 26750 21474
rect 15150 21410 15202 21422
rect 25342 21410 25394 21422
rect 33182 21410 33234 21422
rect 33966 21474 34018 21486
rect 33966 21410 34018 21422
rect 35310 21474 35362 21486
rect 35310 21410 35362 21422
rect 35870 21474 35922 21486
rect 35870 21410 35922 21422
rect 36766 21474 36818 21486
rect 36766 21410 36818 21422
rect 37214 21474 37266 21486
rect 37214 21410 37266 21422
rect 37662 21474 37714 21486
rect 37662 21410 37714 21422
rect 38670 21474 38722 21486
rect 38670 21410 38722 21422
rect 39342 21474 39394 21486
rect 39342 21410 39394 21422
rect 41358 21474 41410 21486
rect 48862 21474 48914 21486
rect 53342 21474 53394 21486
rect 42690 21422 42702 21474
rect 42754 21422 42766 21474
rect 44818 21422 44830 21474
rect 44882 21422 44894 21474
rect 48178 21422 48190 21474
rect 48242 21422 48254 21474
rect 52322 21422 52334 21474
rect 52386 21422 52398 21474
rect 41358 21410 41410 21422
rect 48862 21410 48914 21422
rect 53342 21410 53394 21422
rect 53790 21474 53842 21486
rect 53790 21410 53842 21422
rect 55022 21474 55074 21486
rect 55022 21410 55074 21422
rect 55694 21474 55746 21486
rect 55694 21410 55746 21422
rect 6302 21362 6354 21374
rect 6302 21298 6354 21310
rect 15934 21362 15986 21374
rect 15934 21298 15986 21310
rect 32286 21362 32338 21374
rect 38334 21362 38386 21374
rect 55806 21362 55858 21374
rect 36754 21310 36766 21362
rect 36818 21359 36830 21362
rect 36978 21359 36990 21362
rect 36818 21313 36990 21359
rect 36818 21310 36830 21313
rect 36978 21310 36990 21313
rect 37042 21310 37054 21362
rect 53330 21310 53342 21362
rect 53394 21359 53406 21362
rect 53778 21359 53790 21362
rect 53394 21313 53790 21359
rect 53394 21310 53406 21313
rect 53778 21310 53790 21313
rect 53842 21310 53854 21362
rect 32286 21298 32338 21310
rect 38334 21298 38386 21310
rect 55806 21298 55858 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 8542 21026 8594 21038
rect 8542 20962 8594 20974
rect 37662 21026 37714 21038
rect 37662 20962 37714 20974
rect 38110 21026 38162 21038
rect 38110 20962 38162 20974
rect 45838 21026 45890 21038
rect 45838 20962 45890 20974
rect 52670 21026 52722 21038
rect 52670 20962 52722 20974
rect 53118 21026 53170 21038
rect 53118 20962 53170 20974
rect 2270 20914 2322 20926
rect 2270 20850 2322 20862
rect 4398 20914 4450 20926
rect 14926 20914 14978 20926
rect 22206 20914 22258 20926
rect 5954 20862 5966 20914
rect 6018 20862 6030 20914
rect 14466 20862 14478 20914
rect 14530 20862 14542 20914
rect 16034 20862 16046 20914
rect 16098 20862 16110 20914
rect 18162 20862 18174 20914
rect 18226 20862 18238 20914
rect 4398 20850 4450 20862
rect 14926 20850 14978 20862
rect 22206 20850 22258 20862
rect 23438 20914 23490 20926
rect 41918 20914 41970 20926
rect 26674 20862 26686 20914
rect 26738 20862 26750 20914
rect 31042 20862 31054 20914
rect 31106 20862 31118 20914
rect 33170 20862 33182 20914
rect 33234 20862 33246 20914
rect 38770 20862 38782 20914
rect 38834 20862 38846 20914
rect 40450 20862 40462 20914
rect 40514 20862 40526 20914
rect 23438 20850 23490 20862
rect 41918 20850 41970 20862
rect 43262 20914 43314 20926
rect 43262 20850 43314 20862
rect 45054 20914 45106 20926
rect 45054 20850 45106 20862
rect 50206 20914 50258 20926
rect 53230 20914 53282 20926
rect 51986 20862 51998 20914
rect 52050 20862 52062 20914
rect 50206 20850 50258 20862
rect 53230 20850 53282 20862
rect 53678 20914 53730 20926
rect 57822 20914 57874 20926
rect 54002 20862 54014 20914
rect 54066 20862 54078 20914
rect 56130 20862 56142 20914
rect 56194 20862 56206 20914
rect 53678 20850 53730 20862
rect 57822 20850 57874 20862
rect 58270 20914 58322 20926
rect 58270 20850 58322 20862
rect 3614 20802 3666 20814
rect 2706 20750 2718 20802
rect 2770 20750 2782 20802
rect 3614 20738 3666 20750
rect 4062 20802 4114 20814
rect 4062 20738 4114 20750
rect 4174 20802 4226 20814
rect 4174 20738 4226 20750
rect 4622 20802 4674 20814
rect 4622 20738 4674 20750
rect 4846 20802 4898 20814
rect 4846 20738 4898 20750
rect 7422 20802 7474 20814
rect 7422 20738 7474 20750
rect 7758 20802 7810 20814
rect 8206 20802 8258 20814
rect 7970 20750 7982 20802
rect 8034 20750 8046 20802
rect 7758 20738 7810 20750
rect 8206 20738 8258 20750
rect 8430 20802 8482 20814
rect 18510 20802 18562 20814
rect 19966 20802 20018 20814
rect 8866 20750 8878 20802
rect 8930 20750 8942 20802
rect 10882 20750 10894 20802
rect 10946 20750 10958 20802
rect 14354 20750 14366 20802
rect 14418 20750 14430 20802
rect 15250 20750 15262 20802
rect 15314 20750 15326 20802
rect 19394 20750 19406 20802
rect 19458 20750 19470 20802
rect 8430 20738 8482 20750
rect 18510 20738 18562 20750
rect 19966 20738 20018 20750
rect 20526 20802 20578 20814
rect 20526 20738 20578 20750
rect 21982 20802 22034 20814
rect 21982 20738 22034 20750
rect 22094 20802 22146 20814
rect 28478 20802 28530 20814
rect 23874 20750 23886 20802
rect 23938 20750 23950 20802
rect 27906 20750 27918 20802
rect 27970 20750 27982 20802
rect 22094 20738 22146 20750
rect 28478 20738 28530 20750
rect 30046 20802 30098 20814
rect 30046 20738 30098 20750
rect 30494 20802 30546 20814
rect 34414 20802 34466 20814
rect 35086 20802 35138 20814
rect 33954 20750 33966 20802
rect 34018 20750 34030 20802
rect 34738 20750 34750 20802
rect 34802 20750 34814 20802
rect 30494 20738 30546 20750
rect 34414 20738 34466 20750
rect 35086 20738 35138 20750
rect 35646 20802 35698 20814
rect 35646 20738 35698 20750
rect 35870 20802 35922 20814
rect 35870 20738 35922 20750
rect 36094 20802 36146 20814
rect 36094 20738 36146 20750
rect 37214 20802 37266 20814
rect 37214 20738 37266 20750
rect 37438 20802 37490 20814
rect 41806 20802 41858 20814
rect 38994 20750 39006 20802
rect 39058 20750 39070 20802
rect 40562 20750 40574 20802
rect 40626 20750 40638 20802
rect 37438 20738 37490 20750
rect 41806 20738 41858 20750
rect 42030 20802 42082 20814
rect 42030 20738 42082 20750
rect 42366 20802 42418 20814
rect 42366 20738 42418 20750
rect 44270 20802 44322 20814
rect 50318 20802 50370 20814
rect 51550 20802 51602 20814
rect 46274 20750 46286 20802
rect 46338 20750 46350 20802
rect 50866 20750 50878 20802
rect 50930 20750 50942 20802
rect 56802 20750 56814 20802
rect 56866 20750 56878 20802
rect 44270 20738 44322 20750
rect 50318 20738 50370 20750
rect 51550 20738 51602 20750
rect 6190 20690 6242 20702
rect 12014 20690 12066 20702
rect 2930 20638 2942 20690
rect 2994 20638 3006 20690
rect 8978 20638 8990 20690
rect 9042 20638 9054 20690
rect 6190 20626 6242 20638
rect 12014 20626 12066 20638
rect 18846 20690 18898 20702
rect 18846 20626 18898 20638
rect 19630 20690 19682 20702
rect 19630 20626 19682 20638
rect 22318 20690 22370 20702
rect 22318 20626 22370 20638
rect 22542 20690 22594 20702
rect 27022 20690 27074 20702
rect 29934 20690 29986 20702
rect 24546 20638 24558 20690
rect 24610 20638 24622 20690
rect 28130 20638 28142 20690
rect 28194 20638 28206 20690
rect 29138 20638 29150 20690
rect 29202 20638 29214 20690
rect 22542 20626 22594 20638
rect 27022 20626 27074 20638
rect 29934 20626 29986 20638
rect 36990 20690 37042 20702
rect 36990 20626 37042 20638
rect 39566 20690 39618 20702
rect 39566 20626 39618 20638
rect 39902 20690 39954 20702
rect 39902 20626 39954 20638
rect 40350 20690 40402 20702
rect 40350 20626 40402 20638
rect 40910 20690 40962 20702
rect 40910 20626 40962 20638
rect 45502 20690 45554 20702
rect 47070 20690 47122 20702
rect 46386 20638 46398 20690
rect 46450 20638 46462 20690
rect 45502 20626 45554 20638
rect 47070 20626 47122 20638
rect 52782 20690 52834 20702
rect 52782 20626 52834 20638
rect 1710 20578 1762 20590
rect 1710 20514 1762 20526
rect 3390 20578 3442 20590
rect 3390 20514 3442 20526
rect 3502 20578 3554 20590
rect 3502 20514 3554 20526
rect 5966 20578 6018 20590
rect 5966 20514 6018 20526
rect 6974 20578 7026 20590
rect 6974 20514 7026 20526
rect 7534 20578 7586 20590
rect 27134 20578 27186 20590
rect 10322 20526 10334 20578
rect 10386 20526 10398 20578
rect 7534 20514 7586 20526
rect 27134 20514 27186 20526
rect 28590 20578 28642 20590
rect 28590 20514 28642 20526
rect 29486 20578 29538 20590
rect 29486 20514 29538 20526
rect 29822 20578 29874 20590
rect 29822 20514 29874 20526
rect 35198 20578 35250 20590
rect 35198 20514 35250 20526
rect 35310 20578 35362 20590
rect 35310 20514 35362 20526
rect 36542 20578 36594 20590
rect 36542 20514 36594 20526
rect 40126 20578 40178 20590
rect 40126 20514 40178 20526
rect 41022 20578 41074 20590
rect 41022 20514 41074 20526
rect 41134 20578 41186 20590
rect 41134 20514 41186 20526
rect 42702 20578 42754 20590
rect 42702 20514 42754 20526
rect 43710 20578 43762 20590
rect 43710 20514 43762 20526
rect 47406 20578 47458 20590
rect 47406 20514 47458 20526
rect 47854 20578 47906 20590
rect 47854 20514 47906 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 4846 20242 4898 20254
rect 4846 20178 4898 20190
rect 11230 20242 11282 20254
rect 11230 20178 11282 20190
rect 11678 20242 11730 20254
rect 11678 20178 11730 20190
rect 14478 20242 14530 20254
rect 14478 20178 14530 20190
rect 19406 20242 19458 20254
rect 19406 20178 19458 20190
rect 19742 20242 19794 20254
rect 19742 20178 19794 20190
rect 38558 20242 38610 20254
rect 38558 20178 38610 20190
rect 38894 20242 38946 20254
rect 38894 20178 38946 20190
rect 39006 20242 39058 20254
rect 39006 20178 39058 20190
rect 41022 20242 41074 20254
rect 41022 20178 41074 20190
rect 5070 20130 5122 20142
rect 2482 20078 2494 20130
rect 2546 20078 2558 20130
rect 5070 20066 5122 20078
rect 5182 20130 5234 20142
rect 5182 20066 5234 20078
rect 6078 20130 6130 20142
rect 6078 20066 6130 20078
rect 6414 20130 6466 20142
rect 6414 20066 6466 20078
rect 6750 20130 6802 20142
rect 6750 20066 6802 20078
rect 7310 20130 7362 20142
rect 7310 20066 7362 20078
rect 7422 20130 7474 20142
rect 7422 20066 7474 20078
rect 8654 20130 8706 20142
rect 8654 20066 8706 20078
rect 8878 20130 8930 20142
rect 13582 20130 13634 20142
rect 12002 20078 12014 20130
rect 12066 20078 12078 20130
rect 12450 20078 12462 20130
rect 12514 20078 12526 20130
rect 13234 20078 13246 20130
rect 13298 20078 13310 20130
rect 8878 20066 8930 20078
rect 13582 20066 13634 20078
rect 17950 20130 18002 20142
rect 17950 20066 18002 20078
rect 18398 20130 18450 20142
rect 18398 20066 18450 20078
rect 24110 20130 24162 20142
rect 24110 20066 24162 20078
rect 26686 20130 26738 20142
rect 31950 20130 32002 20142
rect 28242 20078 28254 20130
rect 28306 20078 28318 20130
rect 26686 20066 26738 20078
rect 31950 20066 32002 20078
rect 32062 20130 32114 20142
rect 32062 20066 32114 20078
rect 34974 20130 35026 20142
rect 34974 20066 35026 20078
rect 39790 20130 39842 20142
rect 39790 20066 39842 20078
rect 39902 20130 39954 20142
rect 48862 20130 48914 20142
rect 46274 20078 46286 20130
rect 46338 20078 46350 20130
rect 46610 20078 46622 20130
rect 46674 20078 46686 20130
rect 39902 20066 39954 20078
rect 48862 20066 48914 20078
rect 50206 20130 50258 20142
rect 50206 20066 50258 20078
rect 51550 20130 51602 20142
rect 51550 20066 51602 20078
rect 7086 20018 7138 20030
rect 7982 20018 8034 20030
rect 1810 19966 1822 20018
rect 1874 19966 1886 20018
rect 7746 19966 7758 20018
rect 7810 19966 7822 20018
rect 7086 19954 7138 19966
rect 7982 19954 8034 19966
rect 8990 20018 9042 20030
rect 8990 19954 9042 19966
rect 9550 20018 9602 20030
rect 9550 19954 9602 19966
rect 9774 20018 9826 20030
rect 26462 20018 26514 20030
rect 34862 20018 34914 20030
rect 10098 19966 10110 20018
rect 10162 19966 10174 20018
rect 10994 19966 11006 20018
rect 11058 19966 11070 20018
rect 12674 19966 12686 20018
rect 12738 19966 12750 20018
rect 14690 19966 14702 20018
rect 14754 19966 14766 20018
rect 21186 19966 21198 20018
rect 21250 19966 21262 20018
rect 25778 19966 25790 20018
rect 25842 19966 25854 20018
rect 28130 19966 28142 20018
rect 28194 19966 28206 20018
rect 29698 19966 29710 20018
rect 29762 19966 29774 20018
rect 31042 19966 31054 20018
rect 31106 19966 31118 20018
rect 9774 19954 9826 19966
rect 26462 19954 26514 19966
rect 34862 19954 34914 19966
rect 35870 20018 35922 20030
rect 38782 20018 38834 20030
rect 36306 19966 36318 20018
rect 36370 19966 36382 20018
rect 35870 19954 35922 19966
rect 38782 19954 38834 19966
rect 39230 20018 39282 20030
rect 47294 20018 47346 20030
rect 39554 19966 39566 20018
rect 39618 19966 39630 20018
rect 43138 19966 43150 20018
rect 43202 19966 43214 20018
rect 39230 19954 39282 19966
rect 47294 19954 47346 19966
rect 47854 20018 47906 20030
rect 51102 20018 51154 20030
rect 52446 20018 52498 20030
rect 50866 19966 50878 20018
rect 50930 19966 50942 20018
rect 52210 19966 52222 20018
rect 52274 19966 52286 20018
rect 47854 19954 47906 19966
rect 51102 19954 51154 19966
rect 52446 19954 52498 19966
rect 5630 19906 5682 19918
rect 20302 19906 20354 19918
rect 23662 19906 23714 19918
rect 36766 19906 36818 19918
rect 4610 19854 4622 19906
rect 4674 19854 4686 19906
rect 18946 19854 18958 19906
rect 19010 19854 19022 19906
rect 21858 19854 21870 19906
rect 21922 19854 21934 19906
rect 29362 19854 29374 19906
rect 29426 19854 29438 19906
rect 5630 19842 5682 19854
rect 20302 19842 20354 19854
rect 23662 19842 23714 19854
rect 36766 19842 36818 19854
rect 37214 19906 37266 19918
rect 37214 19842 37266 19854
rect 37662 19906 37714 19918
rect 37662 19842 37714 19854
rect 38110 19906 38162 19918
rect 38110 19842 38162 19854
rect 40238 19906 40290 19918
rect 40238 19842 40290 19854
rect 41470 19906 41522 19918
rect 41470 19842 41522 19854
rect 42254 19906 42306 19918
rect 53902 19906 53954 19918
rect 44930 19854 44942 19906
rect 44994 19854 45006 19906
rect 42254 19842 42306 19854
rect 53902 19842 53954 19854
rect 8094 19794 8146 19806
rect 5506 19742 5518 19794
rect 5570 19791 5582 19794
rect 6178 19791 6190 19794
rect 5570 19745 6190 19791
rect 5570 19742 5582 19745
rect 6178 19742 6190 19745
rect 6242 19742 6254 19794
rect 8094 19730 8146 19742
rect 11342 19794 11394 19806
rect 11342 19730 11394 19742
rect 14366 19794 14418 19806
rect 14366 19730 14418 19742
rect 23550 19794 23602 19806
rect 23550 19730 23602 19742
rect 32062 19794 32114 19806
rect 32062 19730 32114 19742
rect 34974 19794 35026 19806
rect 42142 19794 42194 19806
rect 37202 19742 37214 19794
rect 37266 19791 37278 19794
rect 37650 19791 37662 19794
rect 37266 19745 37662 19791
rect 37266 19742 37278 19745
rect 37650 19742 37662 19745
rect 37714 19742 37726 19794
rect 34974 19730 35026 19742
rect 42142 19730 42194 19742
rect 45614 19794 45666 19806
rect 45614 19730 45666 19742
rect 45950 19794 46002 19806
rect 45950 19730 46002 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 10558 19458 10610 19470
rect 10558 19394 10610 19406
rect 15374 19458 15426 19470
rect 15374 19394 15426 19406
rect 26350 19458 26402 19470
rect 39330 19406 39342 19458
rect 39394 19455 39406 19458
rect 40002 19455 40014 19458
rect 39394 19409 40014 19455
rect 39394 19406 39406 19409
rect 40002 19406 40014 19409
rect 40066 19406 40078 19458
rect 41458 19406 41470 19458
rect 41522 19455 41534 19458
rect 41906 19455 41918 19458
rect 41522 19409 41918 19455
rect 41522 19406 41534 19409
rect 41906 19406 41918 19409
rect 41970 19406 41982 19458
rect 26350 19394 26402 19406
rect 4062 19346 4114 19358
rect 10670 19346 10722 19358
rect 6514 19294 6526 19346
rect 6578 19294 6590 19346
rect 8418 19294 8430 19346
rect 8482 19294 8494 19346
rect 4062 19282 4114 19294
rect 10670 19282 10722 19294
rect 12910 19346 12962 19358
rect 26910 19346 26962 19358
rect 17602 19294 17614 19346
rect 17666 19294 17678 19346
rect 22306 19294 22318 19346
rect 22370 19294 22382 19346
rect 24434 19294 24446 19346
rect 24498 19294 24510 19346
rect 25218 19294 25230 19346
rect 25282 19294 25294 19346
rect 26002 19294 26014 19346
rect 26066 19294 26078 19346
rect 12910 19282 12962 19294
rect 26910 19282 26962 19294
rect 28366 19346 28418 19358
rect 31278 19346 31330 19358
rect 38558 19346 38610 19358
rect 29474 19294 29486 19346
rect 29538 19294 29550 19346
rect 35298 19294 35310 19346
rect 35362 19294 35374 19346
rect 28366 19282 28418 19294
rect 31278 19282 31330 19294
rect 38558 19282 38610 19294
rect 39118 19346 39170 19358
rect 39118 19282 39170 19294
rect 41022 19346 41074 19358
rect 41022 19282 41074 19294
rect 41470 19346 41522 19358
rect 41470 19282 41522 19294
rect 43150 19346 43202 19358
rect 43150 19282 43202 19294
rect 43710 19346 43762 19358
rect 43710 19282 43762 19294
rect 44046 19346 44098 19358
rect 44046 19282 44098 19294
rect 46174 19346 46226 19358
rect 47842 19294 47854 19346
rect 47906 19294 47918 19346
rect 49970 19294 49982 19346
rect 50034 19294 50046 19346
rect 46174 19282 46226 19294
rect 1710 19234 1762 19246
rect 3838 19234 3890 19246
rect 3378 19182 3390 19234
rect 3442 19182 3454 19234
rect 1710 19170 1762 19182
rect 3838 19170 3890 19182
rect 4174 19234 4226 19246
rect 4174 19170 4226 19182
rect 5070 19234 5122 19246
rect 9886 19234 9938 19246
rect 6066 19182 6078 19234
rect 6130 19182 6142 19234
rect 7522 19182 7534 19234
rect 7586 19182 7598 19234
rect 5070 19170 5122 19182
rect 9886 19170 9938 19182
rect 13582 19234 13634 19246
rect 13582 19170 13634 19182
rect 16046 19234 16098 19246
rect 16046 19170 16098 19182
rect 17950 19234 18002 19246
rect 17950 19170 18002 19182
rect 18174 19234 18226 19246
rect 18174 19170 18226 19182
rect 18622 19234 18674 19246
rect 25678 19234 25730 19246
rect 28590 19234 28642 19246
rect 19954 19182 19966 19234
rect 20018 19182 20030 19234
rect 21634 19182 21646 19234
rect 21698 19182 21710 19234
rect 28018 19182 28030 19234
rect 28082 19182 28094 19234
rect 18622 19170 18674 19182
rect 25678 19170 25730 19182
rect 28590 19170 28642 19182
rect 29374 19234 29426 19246
rect 32286 19234 32338 19246
rect 29698 19182 29710 19234
rect 29762 19182 29774 19234
rect 31602 19182 31614 19234
rect 31666 19182 31678 19234
rect 29374 19170 29426 19182
rect 32286 19170 32338 19182
rect 32846 19234 32898 19246
rect 37438 19234 37490 19246
rect 33282 19182 33294 19234
rect 33346 19182 33358 19234
rect 33506 19182 33518 19234
rect 33570 19182 33582 19234
rect 35746 19182 35758 19234
rect 35810 19182 35822 19234
rect 32846 19170 32898 19182
rect 37438 19170 37490 19182
rect 37886 19234 37938 19246
rect 37886 19170 37938 19182
rect 38110 19234 38162 19246
rect 38110 19170 38162 19182
rect 42142 19234 42194 19246
rect 42142 19170 42194 19182
rect 43486 19234 43538 19246
rect 53678 19234 53730 19246
rect 45154 19182 45166 19234
rect 45218 19182 45230 19234
rect 47058 19182 47070 19234
rect 47122 19182 47134 19234
rect 53890 19182 53902 19234
rect 53954 19182 53966 19234
rect 43486 19170 43538 19182
rect 53678 19170 53730 19182
rect 2382 19122 2434 19134
rect 2382 19058 2434 19070
rect 2718 19122 2770 19134
rect 2718 19058 2770 19070
rect 4510 19122 4562 19134
rect 4510 19058 4562 19070
rect 5630 19122 5682 19134
rect 5630 19058 5682 19070
rect 13694 19122 13746 19134
rect 13694 19058 13746 19070
rect 14142 19122 14194 19134
rect 14142 19058 14194 19070
rect 14478 19122 14530 19134
rect 14478 19058 14530 19070
rect 14590 19122 14642 19134
rect 14590 19058 14642 19070
rect 15710 19122 15762 19134
rect 15710 19058 15762 19070
rect 17278 19122 17330 19134
rect 26126 19122 26178 19134
rect 20738 19070 20750 19122
rect 20802 19070 20814 19122
rect 17278 19058 17330 19070
rect 26126 19058 26178 19070
rect 32398 19122 32450 19134
rect 32398 19058 32450 19070
rect 36206 19122 36258 19134
rect 36206 19058 36258 19070
rect 42702 19122 42754 19134
rect 42702 19058 42754 19070
rect 53454 19122 53506 19134
rect 54562 19070 54574 19122
rect 54626 19070 54638 19122
rect 53454 19058 53506 19070
rect 2046 19010 2098 19022
rect 4734 19010 4786 19022
rect 3602 18958 3614 19010
rect 3666 18958 3678 19010
rect 2046 18946 2098 18958
rect 4734 18946 4786 18958
rect 4958 19010 5010 19022
rect 11118 19010 11170 19022
rect 10210 18958 10222 19010
rect 10274 18958 10286 19010
rect 4958 18946 5010 18958
rect 11118 18946 11170 18958
rect 13806 19010 13858 19022
rect 13806 18946 13858 18958
rect 13918 19010 13970 19022
rect 13918 18946 13970 18958
rect 15486 19010 15538 19022
rect 15486 18946 15538 18958
rect 16158 19010 16210 19022
rect 16158 18946 16210 18958
rect 16382 19010 16434 19022
rect 16382 18946 16434 18958
rect 17502 19010 17554 19022
rect 17502 18946 17554 18958
rect 18398 19010 18450 19022
rect 18398 18946 18450 18958
rect 18958 19010 19010 19022
rect 18958 18946 19010 18958
rect 19406 19010 19458 19022
rect 20414 19010 20466 19022
rect 19730 18958 19742 19010
rect 19794 18958 19806 19010
rect 19406 18946 19458 18958
rect 20414 18946 20466 18958
rect 27246 19010 27298 19022
rect 27246 18946 27298 18958
rect 29038 19010 29090 19022
rect 32510 19010 32562 19022
rect 31826 18958 31838 19010
rect 31890 18958 31902 19010
rect 29038 18946 29090 18958
rect 32510 18946 32562 18958
rect 32958 19010 33010 19022
rect 32958 18946 33010 18958
rect 33070 19010 33122 19022
rect 33070 18946 33122 18958
rect 37102 19010 37154 19022
rect 37102 18946 37154 18958
rect 37998 19010 38050 19022
rect 37998 18946 38050 18958
rect 39566 19010 39618 19022
rect 39566 18946 39618 18958
rect 40014 19010 40066 19022
rect 40014 18946 40066 18958
rect 40462 19010 40514 19022
rect 40462 18946 40514 18958
rect 43934 19010 43986 19022
rect 43934 18946 43986 18958
rect 44158 19010 44210 19022
rect 44158 18946 44210 18958
rect 45390 19010 45442 19022
rect 45390 18946 45442 18958
rect 50430 19010 50482 19022
rect 50430 18946 50482 18958
rect 53342 19010 53394 19022
rect 53342 18946 53394 18958
rect 53566 19010 53618 19022
rect 53566 18946 53618 18958
rect 54238 19010 54290 19022
rect 54238 18946 54290 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 2718 18674 2770 18686
rect 2718 18610 2770 18622
rect 3166 18674 3218 18686
rect 3166 18610 3218 18622
rect 3614 18674 3666 18686
rect 3614 18610 3666 18622
rect 5182 18674 5234 18686
rect 5182 18610 5234 18622
rect 7870 18674 7922 18686
rect 7870 18610 7922 18622
rect 8878 18674 8930 18686
rect 8878 18610 8930 18622
rect 9998 18674 10050 18686
rect 9998 18610 10050 18622
rect 15038 18674 15090 18686
rect 15038 18610 15090 18622
rect 18958 18674 19010 18686
rect 18958 18610 19010 18622
rect 19182 18674 19234 18686
rect 19182 18610 19234 18622
rect 20862 18674 20914 18686
rect 20862 18610 20914 18622
rect 21086 18674 21138 18686
rect 21086 18610 21138 18622
rect 22094 18674 22146 18686
rect 22094 18610 22146 18622
rect 22318 18674 22370 18686
rect 22318 18610 22370 18622
rect 26798 18674 26850 18686
rect 26798 18610 26850 18622
rect 36654 18674 36706 18686
rect 36654 18610 36706 18622
rect 39902 18674 39954 18686
rect 39902 18610 39954 18622
rect 42366 18674 42418 18686
rect 42366 18610 42418 18622
rect 43038 18674 43090 18686
rect 43038 18610 43090 18622
rect 43934 18674 43986 18686
rect 43934 18610 43986 18622
rect 2046 18562 2098 18574
rect 2046 18498 2098 18510
rect 5854 18562 5906 18574
rect 5854 18498 5906 18510
rect 6078 18562 6130 18574
rect 6078 18498 6130 18510
rect 8990 18562 9042 18574
rect 25790 18562 25842 18574
rect 32062 18562 32114 18574
rect 10322 18510 10334 18562
rect 10386 18510 10398 18562
rect 21410 18510 21422 18562
rect 21474 18510 21486 18562
rect 28466 18510 28478 18562
rect 28530 18510 28542 18562
rect 31602 18510 31614 18562
rect 31666 18510 31678 18562
rect 8990 18498 9042 18510
rect 25790 18498 25842 18510
rect 32062 18498 32114 18510
rect 32286 18562 32338 18574
rect 32286 18498 32338 18510
rect 36766 18562 36818 18574
rect 38222 18562 38274 18574
rect 37874 18510 37886 18562
rect 37938 18510 37950 18562
rect 36766 18498 36818 18510
rect 38222 18498 38274 18510
rect 38334 18562 38386 18574
rect 38334 18498 38386 18510
rect 44158 18562 44210 18574
rect 44158 18498 44210 18510
rect 44270 18562 44322 18574
rect 44270 18498 44322 18510
rect 44718 18562 44770 18574
rect 46050 18510 46062 18562
rect 46114 18510 46126 18562
rect 44718 18498 44770 18510
rect 1710 18450 1762 18462
rect 1710 18386 1762 18398
rect 3838 18450 3890 18462
rect 3838 18386 3890 18398
rect 4286 18450 4338 18462
rect 4286 18386 4338 18398
rect 4398 18450 4450 18462
rect 8094 18450 8146 18462
rect 11342 18450 11394 18462
rect 14926 18450 14978 18462
rect 16382 18450 16434 18462
rect 6962 18398 6974 18450
rect 7026 18398 7038 18450
rect 8418 18398 8430 18450
rect 8482 18398 8494 18450
rect 11666 18398 11678 18450
rect 11730 18398 11742 18450
rect 12450 18398 12462 18450
rect 12514 18398 12526 18450
rect 15810 18398 15822 18450
rect 15874 18398 15886 18450
rect 4398 18386 4450 18398
rect 8094 18386 8146 18398
rect 11342 18386 11394 18398
rect 14926 18386 14978 18398
rect 16382 18386 16434 18398
rect 16494 18450 16546 18462
rect 16494 18386 16546 18398
rect 17278 18450 17330 18462
rect 19630 18450 19682 18462
rect 18050 18398 18062 18450
rect 18114 18398 18126 18450
rect 18274 18398 18286 18450
rect 18338 18398 18350 18450
rect 17278 18386 17330 18398
rect 19630 18386 19682 18398
rect 21982 18450 22034 18462
rect 21982 18386 22034 18398
rect 22206 18450 22258 18462
rect 22206 18386 22258 18398
rect 22430 18450 22482 18462
rect 22430 18386 22482 18398
rect 24222 18450 24274 18462
rect 24222 18386 24274 18398
rect 24670 18450 24722 18462
rect 24670 18386 24722 18398
rect 25230 18450 25282 18462
rect 25230 18386 25282 18398
rect 25454 18450 25506 18462
rect 26574 18450 26626 18462
rect 26338 18398 26350 18450
rect 26402 18398 26414 18450
rect 25454 18386 25506 18398
rect 26574 18386 26626 18398
rect 26686 18450 26738 18462
rect 29934 18450 29986 18462
rect 27010 18398 27022 18450
rect 27074 18398 27086 18450
rect 29362 18398 29374 18450
rect 29426 18398 29438 18450
rect 26686 18386 26738 18398
rect 29934 18386 29986 18398
rect 30942 18450 30994 18462
rect 33070 18450 33122 18462
rect 31378 18398 31390 18450
rect 31442 18398 31454 18450
rect 30942 18386 30994 18398
rect 33070 18386 33122 18398
rect 33294 18450 33346 18462
rect 36430 18450 36482 18462
rect 33618 18398 33630 18450
rect 33682 18398 33694 18450
rect 33294 18386 33346 18398
rect 36430 18386 36482 18398
rect 36878 18450 36930 18462
rect 36878 18386 36930 18398
rect 37326 18450 37378 18462
rect 37326 18386 37378 18398
rect 37550 18450 37602 18462
rect 37550 18386 37602 18398
rect 38558 18450 38610 18462
rect 38558 18386 38610 18398
rect 39230 18450 39282 18462
rect 39230 18386 39282 18398
rect 39678 18450 39730 18462
rect 39678 18386 39730 18398
rect 40350 18450 40402 18462
rect 40350 18386 40402 18398
rect 42478 18450 42530 18462
rect 48862 18450 48914 18462
rect 45378 18398 45390 18450
rect 45442 18398 45454 18450
rect 42478 18386 42530 18398
rect 48862 18386 48914 18398
rect 51998 18450 52050 18462
rect 55234 18398 55246 18450
rect 55298 18398 55310 18450
rect 51998 18386 52050 18398
rect 4062 18338 4114 18350
rect 6526 18338 6578 18350
rect 7982 18338 8034 18350
rect 19070 18338 19122 18350
rect 5058 18286 5070 18338
rect 5122 18286 5134 18338
rect 5730 18286 5742 18338
rect 5794 18286 5806 18338
rect 7410 18286 7422 18338
rect 7474 18286 7486 18338
rect 14578 18286 14590 18338
rect 14642 18286 14654 18338
rect 18386 18286 18398 18338
rect 18450 18286 18462 18338
rect 4062 18274 4114 18286
rect 6526 18274 6578 18286
rect 7982 18274 8034 18286
rect 19070 18274 19122 18286
rect 23886 18338 23938 18350
rect 23886 18274 23938 18286
rect 25342 18338 25394 18350
rect 25342 18274 25394 18286
rect 27470 18338 27522 18350
rect 27470 18274 27522 18286
rect 28030 18338 28082 18350
rect 28030 18274 28082 18286
rect 29822 18338 29874 18350
rect 33182 18338 33234 18350
rect 31938 18286 31950 18338
rect 32002 18286 32014 18338
rect 29822 18274 29874 18286
rect 33182 18274 33234 18286
rect 39790 18338 39842 18350
rect 39790 18274 39842 18286
rect 43486 18338 43538 18350
rect 48178 18286 48190 18338
rect 48242 18286 48254 18338
rect 52322 18286 52334 18338
rect 52386 18286 52398 18338
rect 54450 18286 54462 18338
rect 54514 18286 54526 18338
rect 43486 18274 43538 18286
rect 5406 18226 5458 18238
rect 5406 18162 5458 18174
rect 8878 18226 8930 18238
rect 8878 18162 8930 18174
rect 15038 18226 15090 18238
rect 42366 18226 42418 18238
rect 28018 18174 28030 18226
rect 28082 18223 28094 18226
rect 28242 18223 28254 18226
rect 28082 18177 28254 18223
rect 28082 18174 28094 18177
rect 28242 18174 28254 18177
rect 28306 18174 28318 18226
rect 28914 18174 28926 18226
rect 28978 18174 28990 18226
rect 15038 18162 15090 18174
rect 42366 18162 42418 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 6862 17890 6914 17902
rect 5506 17838 5518 17890
rect 5570 17887 5582 17890
rect 6514 17887 6526 17890
rect 5570 17841 6526 17887
rect 5570 17838 5582 17841
rect 6514 17838 6526 17841
rect 6578 17838 6590 17890
rect 6862 17826 6914 17838
rect 33518 17890 33570 17902
rect 33518 17826 33570 17838
rect 37438 17890 37490 17902
rect 37438 17826 37490 17838
rect 42814 17890 42866 17902
rect 42814 17826 42866 17838
rect 53566 17890 53618 17902
rect 53566 17826 53618 17838
rect 5070 17778 5122 17790
rect 4610 17726 4622 17778
rect 4674 17726 4686 17778
rect 5070 17714 5122 17726
rect 5854 17778 5906 17790
rect 5854 17714 5906 17726
rect 7646 17778 7698 17790
rect 7646 17714 7698 17726
rect 11342 17778 11394 17790
rect 15262 17778 15314 17790
rect 13682 17726 13694 17778
rect 13746 17726 13758 17778
rect 11342 17714 11394 17726
rect 15262 17714 15314 17726
rect 16494 17778 16546 17790
rect 20862 17778 20914 17790
rect 27022 17778 27074 17790
rect 43598 17778 43650 17790
rect 17378 17726 17390 17778
rect 17442 17726 17454 17778
rect 19506 17726 19518 17778
rect 19570 17726 19582 17778
rect 22082 17726 22094 17778
rect 22146 17726 22158 17778
rect 24210 17726 24222 17778
rect 24274 17726 24286 17778
rect 32610 17726 32622 17778
rect 32674 17726 32686 17778
rect 40338 17726 40350 17778
rect 40402 17726 40414 17778
rect 42466 17726 42478 17778
rect 42530 17726 42542 17778
rect 16494 17714 16546 17726
rect 20862 17714 20914 17726
rect 27022 17714 27074 17726
rect 43598 17714 43650 17726
rect 44046 17778 44098 17790
rect 49758 17778 49810 17790
rect 51662 17778 51714 17790
rect 47618 17726 47630 17778
rect 47682 17726 47694 17778
rect 51202 17726 51214 17778
rect 51266 17726 51278 17778
rect 44046 17714 44098 17726
rect 49758 17714 49810 17726
rect 51662 17714 51714 17726
rect 53454 17778 53506 17790
rect 53454 17714 53506 17726
rect 6190 17666 6242 17678
rect 14590 17666 14642 17678
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 8306 17614 8318 17666
rect 8370 17614 8382 17666
rect 8866 17614 8878 17666
rect 8930 17614 8942 17666
rect 9314 17614 9326 17666
rect 9378 17614 9390 17666
rect 14018 17614 14030 17666
rect 14082 17614 14094 17666
rect 6190 17602 6242 17614
rect 14590 17602 14642 17614
rect 15934 17666 15986 17678
rect 25566 17666 25618 17678
rect 20290 17614 20302 17666
rect 20354 17614 20366 17666
rect 21410 17614 21422 17666
rect 21474 17614 21486 17666
rect 25218 17614 25230 17666
rect 25282 17614 25294 17666
rect 15934 17602 15986 17614
rect 25566 17602 25618 17614
rect 25678 17666 25730 17678
rect 25678 17602 25730 17614
rect 26126 17666 26178 17678
rect 27582 17666 27634 17678
rect 26562 17614 26574 17666
rect 26626 17614 26638 17666
rect 26126 17602 26178 17614
rect 27582 17602 27634 17614
rect 28142 17666 28194 17678
rect 28142 17602 28194 17614
rect 28366 17666 28418 17678
rect 28366 17602 28418 17614
rect 29374 17666 29426 17678
rect 29374 17602 29426 17614
rect 29822 17666 29874 17678
rect 29822 17602 29874 17614
rect 30158 17666 30210 17678
rect 30158 17602 30210 17614
rect 30270 17666 30322 17678
rect 33070 17666 33122 17678
rect 31042 17614 31054 17666
rect 31106 17614 31118 17666
rect 32386 17614 32398 17666
rect 32450 17614 32462 17666
rect 30270 17602 30322 17614
rect 33070 17602 33122 17614
rect 33294 17666 33346 17678
rect 33294 17602 33346 17614
rect 37886 17666 37938 17678
rect 37886 17602 37938 17614
rect 38222 17666 38274 17678
rect 38222 17602 38274 17614
rect 38558 17666 38610 17678
rect 38558 17602 38610 17614
rect 39230 17666 39282 17678
rect 45614 17666 45666 17678
rect 50766 17666 50818 17678
rect 39666 17614 39678 17666
rect 39730 17614 39742 17666
rect 46498 17614 46510 17666
rect 46562 17614 46574 17666
rect 39230 17602 39282 17614
rect 45614 17602 45666 17614
rect 50766 17602 50818 17614
rect 6974 17554 7026 17566
rect 2482 17502 2494 17554
rect 2546 17502 2558 17554
rect 6974 17490 7026 17502
rect 7310 17554 7362 17566
rect 7310 17490 7362 17502
rect 7534 17554 7586 17566
rect 7534 17490 7586 17502
rect 7758 17554 7810 17566
rect 10782 17554 10834 17566
rect 27246 17554 27298 17566
rect 8082 17502 8094 17554
rect 8146 17502 8158 17554
rect 17042 17502 17054 17554
rect 17106 17502 17118 17554
rect 7758 17490 7810 17502
rect 10782 17490 10834 17502
rect 27246 17490 27298 17502
rect 28590 17554 28642 17566
rect 28590 17490 28642 17502
rect 29150 17554 29202 17566
rect 29150 17490 29202 17502
rect 31726 17554 31778 17566
rect 31726 17490 31778 17502
rect 37550 17554 37602 17566
rect 37550 17490 37602 17502
rect 42926 17554 42978 17566
rect 42926 17490 42978 17502
rect 43150 17554 43202 17566
rect 43150 17490 43202 17502
rect 45278 17554 45330 17566
rect 45278 17490 45330 17502
rect 45950 17554 46002 17566
rect 45950 17490 46002 17502
rect 46174 17554 46226 17566
rect 46174 17490 46226 17502
rect 51214 17554 51266 17566
rect 51214 17490 51266 17502
rect 6862 17442 6914 17454
rect 6862 17378 6914 17390
rect 9438 17442 9490 17454
rect 10222 17442 10274 17454
rect 9874 17390 9886 17442
rect 9938 17390 9950 17442
rect 9438 17378 9490 17390
rect 10222 17378 10274 17390
rect 15598 17442 15650 17454
rect 15598 17378 15650 17390
rect 16718 17442 16770 17454
rect 16718 17378 16770 17390
rect 27470 17442 27522 17454
rect 27470 17378 27522 17390
rect 28478 17442 28530 17454
rect 28478 17378 28530 17390
rect 29262 17442 29314 17454
rect 29262 17378 29314 17390
rect 30046 17442 30098 17454
rect 30046 17378 30098 17390
rect 30494 17442 30546 17454
rect 33966 17442 34018 17454
rect 31266 17390 31278 17442
rect 31330 17390 31342 17442
rect 30494 17378 30546 17390
rect 33966 17378 34018 17390
rect 34750 17442 34802 17454
rect 36430 17442 36482 17454
rect 35074 17390 35086 17442
rect 35138 17390 35150 17442
rect 34750 17378 34802 17390
rect 36430 17378 36482 17390
rect 37438 17442 37490 17454
rect 37438 17378 37490 17390
rect 37998 17442 38050 17454
rect 37998 17378 38050 17390
rect 39006 17442 39058 17454
rect 39006 17378 39058 17390
rect 39118 17442 39170 17454
rect 39118 17378 39170 17390
rect 45166 17442 45218 17454
rect 45166 17378 45218 17390
rect 45726 17442 45778 17454
rect 45726 17378 45778 17390
rect 50878 17442 50930 17454
rect 50878 17378 50930 17390
rect 51102 17442 51154 17454
rect 51102 17378 51154 17390
rect 51774 17442 51826 17454
rect 51774 17378 51826 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 1710 17106 1762 17118
rect 1710 17042 1762 17054
rect 3166 17106 3218 17118
rect 3166 17042 3218 17054
rect 3614 17106 3666 17118
rect 11342 17106 11394 17118
rect 4274 17054 4286 17106
rect 4338 17054 4350 17106
rect 3614 17042 3666 17054
rect 11342 17042 11394 17054
rect 13358 17106 13410 17118
rect 13358 17042 13410 17054
rect 19070 17106 19122 17118
rect 19070 17042 19122 17054
rect 20078 17106 20130 17118
rect 20078 17042 20130 17054
rect 20414 17106 20466 17118
rect 26686 17106 26738 17118
rect 20738 17054 20750 17106
rect 20802 17054 20814 17106
rect 25778 17054 25790 17106
rect 25842 17054 25854 17106
rect 20414 17042 20466 17054
rect 26686 17042 26738 17054
rect 26798 17106 26850 17118
rect 26798 17042 26850 17054
rect 28254 17106 28306 17118
rect 28254 17042 28306 17054
rect 37774 17106 37826 17118
rect 37774 17042 37826 17054
rect 41694 17106 41746 17118
rect 41694 17042 41746 17054
rect 42366 17106 42418 17118
rect 42366 17042 42418 17054
rect 43486 17106 43538 17118
rect 43486 17042 43538 17054
rect 46062 17106 46114 17118
rect 46062 17042 46114 17054
rect 47070 17106 47122 17118
rect 47070 17042 47122 17054
rect 47294 17106 47346 17118
rect 47294 17042 47346 17054
rect 47966 17106 48018 17118
rect 47966 17042 48018 17054
rect 2718 16994 2770 17006
rect 13022 16994 13074 17006
rect 2034 16942 2046 16994
rect 2098 16942 2110 16994
rect 4162 16942 4174 16994
rect 4226 16942 4238 16994
rect 5618 16942 5630 16994
rect 5682 16942 5694 16994
rect 9874 16942 9886 16994
rect 9938 16942 9950 16994
rect 11666 16942 11678 16994
rect 11730 16942 11742 16994
rect 2718 16930 2770 16942
rect 13022 16930 13074 16942
rect 13134 16994 13186 17006
rect 13134 16930 13186 16942
rect 15038 16994 15090 17006
rect 15038 16930 15090 16942
rect 16270 16994 16322 17006
rect 16270 16930 16322 16942
rect 18846 16994 18898 17006
rect 30270 16994 30322 17006
rect 22866 16942 22878 16994
rect 22930 16942 22942 16994
rect 24658 16942 24670 16994
rect 24722 16942 24734 16994
rect 29474 16942 29486 16994
rect 29538 16942 29550 16994
rect 18846 16930 18898 16942
rect 30270 16930 30322 16942
rect 31054 16994 31106 17006
rect 31054 16930 31106 16942
rect 39454 16994 39506 17006
rect 39454 16930 39506 16942
rect 42142 16994 42194 17006
rect 42142 16930 42194 16942
rect 42814 16994 42866 17006
rect 42814 16930 42866 16942
rect 44046 16994 44098 17006
rect 44046 16930 44098 16942
rect 44606 16994 44658 17006
rect 44606 16930 44658 16942
rect 47742 16994 47794 17006
rect 47742 16930 47794 16942
rect 48750 16994 48802 17006
rect 52210 16942 52222 16994
rect 52274 16942 52286 16994
rect 48750 16930 48802 16942
rect 2382 16882 2434 16894
rect 2382 16818 2434 16830
rect 3278 16882 3330 16894
rect 3278 16818 3330 16830
rect 3390 16882 3442 16894
rect 14366 16882 14418 16894
rect 4050 16830 4062 16882
rect 4114 16830 4126 16882
rect 5058 16830 5070 16882
rect 5122 16830 5134 16882
rect 8642 16830 8654 16882
rect 8706 16830 8718 16882
rect 10098 16830 10110 16882
rect 10162 16830 10174 16882
rect 3390 16818 3442 16830
rect 14366 16818 14418 16830
rect 14814 16882 14866 16894
rect 14814 16818 14866 16830
rect 16158 16882 16210 16894
rect 16158 16818 16210 16830
rect 18734 16882 18786 16894
rect 24334 16882 24386 16894
rect 26910 16882 26962 16894
rect 28926 16882 28978 16894
rect 42030 16882 42082 16894
rect 45950 16882 46002 16894
rect 21186 16830 21198 16882
rect 21250 16830 21262 16882
rect 25554 16830 25566 16882
rect 25618 16830 25630 16882
rect 27234 16830 27246 16882
rect 27298 16830 27310 16882
rect 29362 16830 29374 16882
rect 29426 16830 29438 16882
rect 34402 16830 34414 16882
rect 34466 16830 34478 16882
rect 35186 16830 35198 16882
rect 35250 16830 35262 16882
rect 45154 16830 45166 16882
rect 45218 16830 45230 16882
rect 18734 16818 18786 16830
rect 24334 16818 24386 16830
rect 26910 16818 26962 16830
rect 28926 16818 28978 16830
rect 42030 16818 42082 16830
rect 45950 16818 46002 16830
rect 46734 16882 46786 16894
rect 46734 16818 46786 16830
rect 47630 16882 47682 16894
rect 49410 16830 49422 16882
rect 49474 16830 49486 16882
rect 52994 16830 53006 16882
rect 53058 16830 53070 16882
rect 47630 16818 47682 16830
rect 14926 16770 14978 16782
rect 43262 16770 43314 16782
rect 6626 16718 6638 16770
rect 6690 16718 6702 16770
rect 37314 16718 37326 16770
rect 37378 16718 37390 16770
rect 42914 16718 42926 16770
rect 42978 16718 42990 16770
rect 44930 16718 44942 16770
rect 44994 16718 45006 16770
rect 47170 16718 47182 16770
rect 47234 16718 47246 16770
rect 49186 16718 49198 16770
rect 49250 16718 49262 16770
rect 50082 16718 50094 16770
rect 50146 16718 50158 16770
rect 14926 16706 14978 16718
rect 43262 16706 43314 16718
rect 16270 16658 16322 16670
rect 16270 16594 16322 16606
rect 28590 16658 28642 16670
rect 28590 16594 28642 16606
rect 42590 16658 42642 16670
rect 42590 16594 42642 16606
rect 43598 16658 43650 16670
rect 43598 16594 43650 16606
rect 46062 16658 46114 16670
rect 46062 16594 46114 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 8766 16322 8818 16334
rect 8766 16258 8818 16270
rect 9102 16322 9154 16334
rect 9102 16258 9154 16270
rect 10782 16322 10834 16334
rect 10782 16258 10834 16270
rect 17166 16322 17218 16334
rect 25790 16322 25842 16334
rect 24658 16270 24670 16322
rect 24722 16319 24734 16322
rect 25106 16319 25118 16322
rect 24722 16273 25118 16319
rect 24722 16270 24734 16273
rect 25106 16270 25118 16273
rect 25170 16270 25182 16322
rect 17166 16258 17218 16270
rect 25790 16258 25842 16270
rect 26798 16322 26850 16334
rect 26798 16258 26850 16270
rect 33070 16322 33122 16334
rect 33070 16258 33122 16270
rect 43710 16322 43762 16334
rect 43710 16258 43762 16270
rect 46510 16322 46562 16334
rect 46510 16258 46562 16270
rect 48750 16322 48802 16334
rect 48750 16258 48802 16270
rect 49086 16322 49138 16334
rect 49086 16258 49138 16270
rect 5070 16210 5122 16222
rect 4610 16158 4622 16210
rect 4674 16158 4686 16210
rect 5070 16146 5122 16158
rect 9662 16210 9714 16222
rect 14702 16210 14754 16222
rect 25118 16210 25170 16222
rect 11106 16158 11118 16210
rect 11170 16158 11182 16210
rect 12674 16158 12686 16210
rect 12738 16158 12750 16210
rect 15026 16158 15038 16210
rect 15090 16158 15102 16210
rect 24322 16158 24334 16210
rect 24386 16158 24398 16210
rect 9662 16146 9714 16158
rect 14702 16146 14754 16158
rect 25118 16146 25170 16158
rect 25678 16210 25730 16222
rect 28366 16210 28418 16222
rect 27346 16158 27358 16210
rect 27410 16158 27422 16210
rect 25678 16146 25730 16158
rect 28366 16146 28418 16158
rect 35646 16210 35698 16222
rect 35646 16146 35698 16158
rect 38222 16210 38274 16222
rect 45054 16210 45106 16222
rect 39778 16158 39790 16210
rect 39842 16158 39854 16210
rect 41906 16158 41918 16210
rect 41970 16158 41982 16210
rect 38222 16146 38274 16158
rect 45054 16146 45106 16158
rect 46734 16210 46786 16222
rect 46734 16146 46786 16158
rect 47070 16210 47122 16222
rect 49646 16210 49698 16222
rect 48402 16158 48414 16210
rect 48466 16158 48478 16210
rect 47070 16146 47122 16158
rect 49646 16146 49698 16158
rect 50094 16210 50146 16222
rect 50094 16146 50146 16158
rect 7870 16098 7922 16110
rect 1810 16046 1822 16098
rect 1874 16046 1886 16098
rect 6738 16046 6750 16098
rect 6802 16046 6814 16098
rect 6962 16046 6974 16098
rect 7026 16046 7038 16098
rect 7870 16034 7922 16046
rect 8094 16098 8146 16110
rect 8094 16034 8146 16046
rect 11790 16098 11842 16110
rect 11790 16034 11842 16046
rect 12126 16098 12178 16110
rect 12126 16034 12178 16046
rect 12350 16098 12402 16110
rect 12350 16034 12402 16046
rect 14590 16098 14642 16110
rect 16718 16098 16770 16110
rect 15250 16046 15262 16098
rect 15314 16046 15326 16098
rect 14590 16034 14642 16046
rect 16718 16034 16770 16046
rect 17614 16098 17666 16110
rect 17614 16034 17666 16046
rect 17838 16098 17890 16110
rect 17838 16034 17890 16046
rect 18062 16098 18114 16110
rect 18062 16034 18114 16046
rect 21982 16098 22034 16110
rect 21982 16034 22034 16046
rect 22206 16098 22258 16110
rect 26350 16098 26402 16110
rect 22978 16046 22990 16098
rect 23042 16046 23054 16098
rect 23650 16046 23662 16098
rect 23714 16046 23726 16098
rect 22206 16034 22258 16046
rect 26350 16034 26402 16046
rect 26574 16098 26626 16110
rect 26574 16034 26626 16046
rect 31838 16098 31890 16110
rect 31838 16034 31890 16046
rect 32062 16098 32114 16110
rect 32062 16034 32114 16046
rect 32286 16098 32338 16110
rect 32286 16034 32338 16046
rect 33182 16098 33234 16110
rect 33182 16034 33234 16046
rect 34750 16098 34802 16110
rect 34750 16034 34802 16046
rect 35534 16098 35586 16110
rect 35534 16034 35586 16046
rect 35758 16098 35810 16110
rect 43262 16098 43314 16110
rect 39106 16046 39118 16098
rect 39170 16046 39182 16098
rect 42914 16046 42926 16098
rect 42978 16046 42990 16098
rect 35758 16034 35810 16046
rect 43262 16034 43314 16046
rect 45390 16098 45442 16110
rect 45390 16034 45442 16046
rect 47182 16098 47234 16110
rect 49198 16098 49250 16110
rect 47506 16046 47518 16098
rect 47570 16046 47582 16098
rect 47182 16034 47234 16046
rect 49198 16034 49250 16046
rect 50654 16098 50706 16110
rect 50654 16034 50706 16046
rect 50766 16098 50818 16110
rect 50766 16034 50818 16046
rect 6190 15986 6242 15998
rect 2482 15934 2494 15986
rect 2546 15934 2558 15986
rect 6190 15922 6242 15934
rect 6526 15986 6578 15998
rect 6526 15922 6578 15934
rect 11454 15986 11506 15998
rect 15934 15986 15986 15998
rect 13682 15934 13694 15986
rect 13746 15934 13758 15986
rect 14018 15934 14030 15986
rect 14082 15934 14094 15986
rect 11454 15922 11506 15934
rect 15934 15922 15986 15934
rect 16830 15986 16882 15998
rect 16830 15922 16882 15934
rect 22430 15986 22482 15998
rect 24558 15986 24610 15998
rect 22754 15934 22766 15986
rect 22818 15934 22830 15986
rect 22430 15922 22482 15934
rect 24558 15922 24610 15934
rect 26126 15986 26178 15998
rect 26126 15922 26178 15934
rect 27694 15986 27746 15998
rect 27694 15922 27746 15934
rect 27806 15986 27858 15998
rect 27806 15922 27858 15934
rect 32734 15986 32786 15998
rect 32734 15922 32786 15934
rect 33070 15986 33122 15998
rect 33070 15922 33122 15934
rect 33854 15986 33906 15998
rect 33854 15922 33906 15934
rect 35198 15986 35250 15998
rect 35198 15922 35250 15934
rect 36990 15986 37042 15998
rect 36990 15922 37042 15934
rect 37550 15986 37602 15998
rect 37550 15922 37602 15934
rect 37886 15986 37938 15998
rect 37886 15922 37938 15934
rect 43374 15986 43426 15998
rect 43374 15922 43426 15934
rect 43934 15986 43986 15998
rect 43934 15922 43986 15934
rect 50990 15986 51042 15998
rect 50990 15922 51042 15934
rect 51550 15986 51602 15998
rect 53442 15934 53454 15986
rect 53506 15934 53518 15986
rect 51550 15922 51602 15934
rect 5966 15874 6018 15886
rect 5966 15810 6018 15822
rect 6078 15874 6130 15886
rect 6078 15810 6130 15822
rect 7982 15874 8034 15886
rect 7982 15810 8034 15822
rect 8318 15874 8370 15886
rect 8318 15810 8370 15822
rect 8990 15874 9042 15886
rect 8990 15810 9042 15822
rect 11006 15874 11058 15886
rect 11006 15810 11058 15822
rect 11790 15874 11842 15886
rect 11790 15810 11842 15822
rect 12574 15874 12626 15886
rect 12574 15810 12626 15822
rect 17054 15874 17106 15886
rect 17054 15810 17106 15822
rect 21870 15874 21922 15886
rect 21870 15810 21922 15822
rect 22094 15874 22146 15886
rect 22094 15810 22146 15822
rect 28030 15874 28082 15886
rect 28030 15810 28082 15822
rect 34078 15874 34130 15886
rect 34078 15810 34130 15822
rect 34190 15874 34242 15886
rect 34190 15810 34242 15822
rect 34302 15874 34354 15886
rect 34302 15810 34354 15822
rect 35982 15874 36034 15886
rect 35982 15810 36034 15822
rect 37102 15874 37154 15886
rect 37102 15810 37154 15822
rect 37326 15874 37378 15886
rect 37326 15810 37378 15822
rect 37662 15874 37714 15886
rect 37662 15810 37714 15822
rect 43822 15874 43874 15886
rect 43822 15810 43874 15822
rect 45502 15874 45554 15886
rect 45502 15810 45554 15822
rect 45726 15874 45778 15886
rect 48526 15874 48578 15886
rect 46162 15822 46174 15874
rect 46226 15822 46238 15874
rect 45726 15810 45778 15822
rect 48526 15810 48578 15822
rect 49534 15874 49586 15886
rect 49534 15810 49586 15822
rect 50878 15874 50930 15886
rect 50878 15810 50930 15822
rect 51102 15874 51154 15886
rect 51102 15810 51154 15822
rect 51662 15874 51714 15886
rect 51662 15810 51714 15822
rect 52782 15874 52834 15886
rect 52782 15810 52834 15822
rect 53118 15874 53170 15886
rect 53118 15810 53170 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 2718 15538 2770 15550
rect 2718 15474 2770 15486
rect 3166 15538 3218 15550
rect 3166 15474 3218 15486
rect 3278 15538 3330 15550
rect 3278 15474 3330 15486
rect 4734 15538 4786 15550
rect 4734 15474 4786 15486
rect 4958 15538 5010 15550
rect 4958 15474 5010 15486
rect 5518 15538 5570 15550
rect 5518 15474 5570 15486
rect 8990 15538 9042 15550
rect 16830 15538 16882 15550
rect 10434 15486 10446 15538
rect 10498 15486 10510 15538
rect 8990 15474 9042 15486
rect 16830 15474 16882 15486
rect 24446 15538 24498 15550
rect 24446 15474 24498 15486
rect 32510 15538 32562 15550
rect 32510 15474 32562 15486
rect 35982 15538 36034 15550
rect 35982 15474 36034 15486
rect 38222 15538 38274 15550
rect 38222 15474 38274 15486
rect 38334 15538 38386 15550
rect 38334 15474 38386 15486
rect 39230 15538 39282 15550
rect 39230 15474 39282 15486
rect 41246 15538 41298 15550
rect 41246 15474 41298 15486
rect 42030 15538 42082 15550
rect 44718 15538 44770 15550
rect 44146 15486 44158 15538
rect 44210 15486 44222 15538
rect 42030 15474 42082 15486
rect 44718 15474 44770 15486
rect 45614 15538 45666 15550
rect 45614 15474 45666 15486
rect 45838 15538 45890 15550
rect 45838 15474 45890 15486
rect 47966 15538 48018 15550
rect 47966 15474 48018 15486
rect 1710 15426 1762 15438
rect 1710 15362 1762 15374
rect 2046 15426 2098 15438
rect 2046 15362 2098 15374
rect 2382 15426 2434 15438
rect 2382 15362 2434 15374
rect 8094 15426 8146 15438
rect 8094 15362 8146 15374
rect 8206 15426 8258 15438
rect 13470 15426 13522 15438
rect 8642 15374 8654 15426
rect 8706 15374 8718 15426
rect 8206 15362 8258 15374
rect 13470 15362 13522 15374
rect 19294 15426 19346 15438
rect 19294 15362 19346 15374
rect 19630 15426 19682 15438
rect 19630 15362 19682 15374
rect 23662 15426 23714 15438
rect 23662 15362 23714 15374
rect 23998 15426 24050 15438
rect 23998 15362 24050 15374
rect 27582 15426 27634 15438
rect 27582 15362 27634 15374
rect 28814 15426 28866 15438
rect 28814 15362 28866 15374
rect 29038 15426 29090 15438
rect 29038 15362 29090 15374
rect 32286 15426 32338 15438
rect 32286 15362 32338 15374
rect 33070 15426 33122 15438
rect 33070 15362 33122 15374
rect 38446 15426 38498 15438
rect 38446 15362 38498 15374
rect 39006 15426 39058 15438
rect 39006 15362 39058 15374
rect 42254 15426 42306 15438
rect 42254 15362 42306 15374
rect 46958 15426 47010 15438
rect 47742 15426 47794 15438
rect 47170 15374 47182 15426
rect 47234 15374 47246 15426
rect 46958 15362 47010 15374
rect 47742 15362 47794 15374
rect 48078 15426 48130 15438
rect 48078 15362 48130 15374
rect 49422 15426 49474 15438
rect 49422 15362 49474 15374
rect 49646 15426 49698 15438
rect 52546 15374 52558 15426
rect 52610 15374 52622 15426
rect 49646 15362 49698 15374
rect 3054 15314 3106 15326
rect 3054 15250 3106 15262
rect 3726 15314 3778 15326
rect 3726 15250 3778 15262
rect 3838 15314 3890 15326
rect 3838 15250 3890 15262
rect 4062 15314 4114 15326
rect 4062 15250 4114 15262
rect 4174 15314 4226 15326
rect 4174 15250 4226 15262
rect 4510 15314 4562 15326
rect 4510 15250 4562 15262
rect 5070 15314 5122 15326
rect 7534 15314 7586 15326
rect 7074 15262 7086 15314
rect 7138 15262 7150 15314
rect 5070 15250 5122 15262
rect 7534 15250 7586 15262
rect 9438 15314 9490 15326
rect 9438 15250 9490 15262
rect 9886 15314 9938 15326
rect 9886 15250 9938 15262
rect 10110 15314 10162 15326
rect 12798 15314 12850 15326
rect 10658 15262 10670 15314
rect 10722 15262 10734 15314
rect 11330 15262 11342 15314
rect 11394 15262 11406 15314
rect 11666 15262 11678 15314
rect 11730 15262 11742 15314
rect 10110 15250 10162 15262
rect 12798 15250 12850 15262
rect 13022 15314 13074 15326
rect 13022 15250 13074 15262
rect 13134 15314 13186 15326
rect 13134 15250 13186 15262
rect 13806 15314 13858 15326
rect 13806 15250 13858 15262
rect 14030 15314 14082 15326
rect 14030 15250 14082 15262
rect 14366 15314 14418 15326
rect 14366 15250 14418 15262
rect 14702 15314 14754 15326
rect 14702 15250 14754 15262
rect 14926 15314 14978 15326
rect 14926 15250 14978 15262
rect 15150 15314 15202 15326
rect 15150 15250 15202 15262
rect 16158 15314 16210 15326
rect 16158 15250 16210 15262
rect 16606 15314 16658 15326
rect 19070 15314 19122 15326
rect 27918 15314 27970 15326
rect 17826 15262 17838 15314
rect 17890 15262 17902 15314
rect 20514 15262 20526 15314
rect 20578 15262 20590 15314
rect 26898 15262 26910 15314
rect 26962 15262 26974 15314
rect 16606 15250 16658 15262
rect 19070 15250 19122 15262
rect 27918 15250 27970 15262
rect 28478 15314 28530 15326
rect 31838 15314 31890 15326
rect 31042 15262 31054 15314
rect 31106 15262 31118 15314
rect 28478 15250 28530 15262
rect 31838 15250 31890 15262
rect 33294 15314 33346 15326
rect 33294 15250 33346 15262
rect 33518 15314 33570 15326
rect 33518 15250 33570 15262
rect 34526 15314 34578 15326
rect 35870 15314 35922 15326
rect 34962 15262 34974 15314
rect 35026 15262 35038 15314
rect 34526 15250 34578 15262
rect 35870 15250 35922 15262
rect 36206 15314 36258 15326
rect 37326 15314 37378 15326
rect 36978 15262 36990 15314
rect 37042 15262 37054 15314
rect 36206 15250 36258 15262
rect 37326 15250 37378 15262
rect 38894 15314 38946 15326
rect 38894 15250 38946 15262
rect 39342 15314 39394 15326
rect 43150 15314 43202 15326
rect 42914 15262 42926 15314
rect 42978 15262 42990 15314
rect 39342 15250 39394 15262
rect 43150 15250 43202 15262
rect 43598 15314 43650 15326
rect 43598 15250 43650 15262
rect 43822 15314 43874 15326
rect 43822 15250 43874 15262
rect 44494 15314 44546 15326
rect 44494 15250 44546 15262
rect 44606 15314 44658 15326
rect 44606 15250 44658 15262
rect 45166 15314 45218 15326
rect 45166 15250 45218 15262
rect 45390 15314 45442 15326
rect 45390 15250 45442 15262
rect 46510 15314 46562 15326
rect 46510 15250 46562 15262
rect 46622 15314 46674 15326
rect 46622 15250 46674 15262
rect 47294 15314 47346 15326
rect 49870 15314 49922 15326
rect 47506 15262 47518 15314
rect 47570 15262 47582 15314
rect 50082 15262 50094 15314
rect 50146 15262 50158 15314
rect 53218 15262 53230 15314
rect 53282 15262 53294 15314
rect 47294 15250 47346 15262
rect 49870 15250 49922 15262
rect 5966 15202 6018 15214
rect 5966 15138 6018 15150
rect 6638 15202 6690 15214
rect 6638 15138 6690 15150
rect 9998 15202 10050 15214
rect 9998 15138 10050 15150
rect 11118 15202 11170 15214
rect 11118 15138 11170 15150
rect 14254 15202 14306 15214
rect 14254 15138 14306 15150
rect 15598 15202 15650 15214
rect 15598 15138 15650 15150
rect 16718 15202 16770 15214
rect 18510 15202 18562 15214
rect 17602 15150 17614 15202
rect 17666 15150 17678 15202
rect 16718 15138 16770 15150
rect 18510 15138 18562 15150
rect 19518 15202 19570 15214
rect 32398 15202 32450 15214
rect 21186 15150 21198 15202
rect 21250 15150 21262 15202
rect 23314 15150 23326 15202
rect 23378 15150 23390 15202
rect 26786 15150 26798 15202
rect 26850 15150 26862 15202
rect 29138 15150 29150 15202
rect 29202 15150 29214 15202
rect 31154 15150 31166 15202
rect 31218 15150 31230 15202
rect 19518 15138 19570 15150
rect 32398 15138 32450 15150
rect 35422 15202 35474 15214
rect 35422 15138 35474 15150
rect 37438 15202 37490 15214
rect 37438 15138 37490 15150
rect 45502 15202 45554 15214
rect 45502 15138 45554 15150
rect 49758 15202 49810 15214
rect 50418 15150 50430 15202
rect 50482 15150 50494 15202
rect 49758 15138 49810 15150
rect 8094 15090 8146 15102
rect 33742 15090 33794 15102
rect 30594 15038 30606 15090
rect 30658 15038 30670 15090
rect 8094 15026 8146 15038
rect 33742 15026 33794 15038
rect 34190 15090 34242 15102
rect 34190 15026 34242 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 6302 14754 6354 14766
rect 4386 14702 4398 14754
rect 4450 14751 4462 14754
rect 4946 14751 4958 14754
rect 4450 14705 4958 14751
rect 4450 14702 4462 14705
rect 4946 14702 4958 14705
rect 5010 14702 5022 14754
rect 6302 14690 6354 14702
rect 8430 14754 8482 14766
rect 19070 14754 19122 14766
rect 9762 14702 9774 14754
rect 9826 14702 9838 14754
rect 8430 14690 8482 14702
rect 19070 14690 19122 14702
rect 21534 14754 21586 14766
rect 21534 14690 21586 14702
rect 27694 14754 27746 14766
rect 27694 14690 27746 14702
rect 28030 14754 28082 14766
rect 28030 14690 28082 14702
rect 34302 14754 34354 14766
rect 34302 14690 34354 14702
rect 45614 14754 45666 14766
rect 45614 14690 45666 14702
rect 46846 14754 46898 14766
rect 46846 14690 46898 14702
rect 47182 14754 47234 14766
rect 47182 14690 47234 14702
rect 3166 14642 3218 14654
rect 3166 14578 3218 14590
rect 3614 14642 3666 14654
rect 3614 14578 3666 14590
rect 4622 14642 4674 14654
rect 7534 14642 7586 14654
rect 14926 14642 14978 14654
rect 21646 14642 21698 14654
rect 25902 14642 25954 14654
rect 32622 14642 32674 14654
rect 40798 14642 40850 14654
rect 43822 14642 43874 14654
rect 5954 14590 5966 14642
rect 6018 14590 6030 14642
rect 10098 14590 10110 14642
rect 10162 14590 10174 14642
rect 11778 14590 11790 14642
rect 11842 14590 11854 14642
rect 13794 14590 13806 14642
rect 13858 14590 13870 14642
rect 16258 14590 16270 14642
rect 16322 14590 16334 14642
rect 17490 14590 17502 14642
rect 17554 14590 17566 14642
rect 23202 14590 23214 14642
rect 23266 14590 23278 14642
rect 25330 14590 25342 14642
rect 25394 14590 25406 14642
rect 31602 14590 31614 14642
rect 31666 14590 31678 14642
rect 33170 14590 33182 14642
rect 33234 14590 33246 14642
rect 38658 14590 38670 14642
rect 38722 14590 38734 14642
rect 42018 14590 42030 14642
rect 42082 14590 42094 14642
rect 42914 14590 42926 14642
rect 42978 14590 42990 14642
rect 4622 14578 4674 14590
rect 7534 14578 7586 14590
rect 14926 14578 14978 14590
rect 21646 14578 21698 14590
rect 25902 14578 25954 14590
rect 32622 14578 32674 14590
rect 40798 14578 40850 14590
rect 43822 14578 43874 14590
rect 45054 14642 45106 14654
rect 45054 14578 45106 14590
rect 45278 14642 45330 14654
rect 45278 14578 45330 14590
rect 48526 14642 48578 14654
rect 48850 14590 48862 14642
rect 48914 14590 48926 14642
rect 48526 14578 48578 14590
rect 1710 14530 1762 14542
rect 4174 14530 4226 14542
rect 2482 14478 2494 14530
rect 2546 14478 2558 14530
rect 1710 14466 1762 14478
rect 4174 14466 4226 14478
rect 5070 14530 5122 14542
rect 5070 14466 5122 14478
rect 6638 14530 6690 14542
rect 6638 14466 6690 14478
rect 7310 14530 7362 14542
rect 7310 14466 7362 14478
rect 7758 14530 7810 14542
rect 7758 14466 7810 14478
rect 7982 14530 8034 14542
rect 11006 14530 11058 14542
rect 14814 14530 14866 14542
rect 18734 14530 18786 14542
rect 26574 14530 26626 14542
rect 9426 14478 9438 14530
rect 9490 14478 9502 14530
rect 9762 14478 9774 14530
rect 9826 14478 9838 14530
rect 11890 14478 11902 14530
rect 11954 14478 11966 14530
rect 13906 14478 13918 14530
rect 13970 14478 13982 14530
rect 16370 14478 16382 14530
rect 16434 14478 16446 14530
rect 17938 14478 17950 14530
rect 18002 14478 18014 14530
rect 19730 14478 19742 14530
rect 19794 14478 19806 14530
rect 22418 14478 22430 14530
rect 22482 14478 22494 14530
rect 26338 14478 26350 14530
rect 26402 14478 26414 14530
rect 7982 14466 8034 14478
rect 11006 14466 11058 14478
rect 14814 14466 14866 14478
rect 18734 14466 18786 14478
rect 26574 14466 26626 14478
rect 26686 14530 26738 14542
rect 26686 14466 26738 14478
rect 26910 14530 26962 14542
rect 34750 14530 34802 14542
rect 31154 14478 31166 14530
rect 31218 14478 31230 14530
rect 33282 14478 33294 14530
rect 33346 14478 33358 14530
rect 26910 14466 26962 14478
rect 34750 14466 34802 14478
rect 34974 14530 35026 14542
rect 34974 14466 35026 14478
rect 35198 14530 35250 14542
rect 35198 14466 35250 14478
rect 35758 14530 35810 14542
rect 35758 14466 35810 14478
rect 37214 14530 37266 14542
rect 37214 14466 37266 14478
rect 37662 14530 37714 14542
rect 37874 14478 37886 14530
rect 37938 14478 37950 14530
rect 41346 14478 41358 14530
rect 41410 14478 41422 14530
rect 42242 14478 42254 14530
rect 42306 14478 42318 14530
rect 43362 14478 43374 14530
rect 43426 14478 43438 14530
rect 45602 14478 45614 14530
rect 45666 14478 45678 14530
rect 51650 14478 51662 14530
rect 51714 14478 51726 14530
rect 37662 14466 37714 14478
rect 2718 14418 2770 14430
rect 2034 14366 2046 14418
rect 2098 14366 2110 14418
rect 2718 14354 2770 14366
rect 4062 14418 4114 14430
rect 4062 14354 4114 14366
rect 6078 14418 6130 14430
rect 6078 14354 6130 14366
rect 12574 14418 12626 14430
rect 12574 14354 12626 14366
rect 13470 14418 13522 14430
rect 13470 14354 13522 14366
rect 17054 14418 17106 14430
rect 17054 14354 17106 14366
rect 18398 14418 18450 14430
rect 18398 14354 18450 14366
rect 18958 14418 19010 14430
rect 18958 14354 19010 14366
rect 19406 14418 19458 14430
rect 19406 14354 19458 14366
rect 26014 14418 26066 14430
rect 26014 14354 26066 14366
rect 26798 14418 26850 14430
rect 26798 14354 26850 14366
rect 27806 14418 27858 14430
rect 27806 14354 27858 14366
rect 30718 14418 30770 14430
rect 30718 14354 30770 14366
rect 32846 14418 32898 14430
rect 32846 14354 32898 14366
rect 35422 14418 35474 14430
rect 35422 14354 35474 14366
rect 36206 14418 36258 14430
rect 46622 14418 46674 14430
rect 41458 14366 41470 14418
rect 41522 14366 41534 14418
rect 50978 14366 50990 14418
rect 51042 14366 51054 14418
rect 36206 14354 36258 14366
rect 46622 14354 46674 14366
rect 3838 14306 3890 14318
rect 3838 14242 3890 14254
rect 6750 14306 6802 14318
rect 6750 14242 6802 14254
rect 6862 14306 6914 14318
rect 6862 14242 6914 14254
rect 11118 14306 11170 14318
rect 11118 14242 11170 14254
rect 11342 14306 11394 14318
rect 11342 14242 11394 14254
rect 15038 14306 15090 14318
rect 15038 14242 15090 14254
rect 19518 14306 19570 14318
rect 19518 14242 19570 14254
rect 22094 14306 22146 14318
rect 22094 14242 22146 14254
rect 35870 14306 35922 14318
rect 35870 14242 35922 14254
rect 35982 14306 36034 14318
rect 35982 14242 36034 14254
rect 36990 14306 37042 14318
rect 36990 14242 37042 14254
rect 37102 14306 37154 14318
rect 37102 14242 37154 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 13022 13970 13074 13982
rect 13022 13906 13074 13918
rect 18510 13970 18562 13982
rect 18510 13906 18562 13918
rect 24670 13970 24722 13982
rect 24670 13906 24722 13918
rect 25566 13970 25618 13982
rect 25566 13906 25618 13918
rect 26014 13970 26066 13982
rect 26014 13906 26066 13918
rect 28926 13970 28978 13982
rect 28926 13906 28978 13918
rect 30942 13970 30994 13982
rect 30942 13906 30994 13918
rect 33406 13970 33458 13982
rect 33406 13906 33458 13918
rect 34974 13970 35026 13982
rect 34974 13906 35026 13918
rect 37662 13970 37714 13982
rect 37662 13906 37714 13918
rect 37774 13970 37826 13982
rect 37774 13906 37826 13918
rect 37886 13970 37938 13982
rect 37886 13906 37938 13918
rect 38782 13970 38834 13982
rect 38782 13906 38834 13918
rect 39454 13970 39506 13982
rect 39454 13906 39506 13918
rect 40014 13970 40066 13982
rect 44830 13970 44882 13982
rect 43474 13918 43486 13970
rect 43538 13918 43550 13970
rect 40014 13906 40066 13918
rect 44830 13906 44882 13918
rect 45950 13970 46002 13982
rect 45950 13906 46002 13918
rect 46174 13970 46226 13982
rect 46174 13906 46226 13918
rect 47070 13970 47122 13982
rect 47070 13906 47122 13918
rect 49422 13970 49474 13982
rect 50878 13970 50930 13982
rect 49746 13918 49758 13970
rect 49810 13918 49822 13970
rect 49422 13906 49474 13918
rect 50878 13906 50930 13918
rect 5294 13858 5346 13870
rect 5294 13794 5346 13806
rect 5518 13858 5570 13870
rect 5518 13794 5570 13806
rect 7646 13858 7698 13870
rect 7646 13794 7698 13806
rect 13134 13858 13186 13870
rect 13134 13794 13186 13806
rect 18286 13858 18338 13870
rect 18286 13794 18338 13806
rect 27134 13858 27186 13870
rect 27134 13794 27186 13806
rect 27694 13858 27746 13870
rect 27694 13794 27746 13806
rect 28366 13858 28418 13870
rect 28366 13794 28418 13806
rect 29374 13858 29426 13870
rect 29374 13794 29426 13806
rect 33294 13858 33346 13870
rect 33294 13794 33346 13806
rect 39566 13858 39618 13870
rect 47294 13858 47346 13870
rect 41122 13806 41134 13858
rect 41186 13806 41198 13858
rect 41570 13806 41582 13858
rect 41634 13806 41646 13858
rect 42690 13806 42702 13858
rect 42754 13806 42766 13858
rect 46498 13806 46510 13858
rect 46562 13806 46574 13858
rect 39566 13794 39618 13806
rect 47294 13794 47346 13806
rect 47518 13858 47570 13870
rect 50766 13858 50818 13870
rect 50082 13806 50094 13858
rect 50146 13806 50158 13858
rect 47518 13794 47570 13806
rect 50766 13794 50818 13806
rect 4958 13746 5010 13758
rect 7198 13746 7250 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 6962 13694 6974 13746
rect 7026 13694 7038 13746
rect 4958 13682 5010 13694
rect 7198 13682 7250 13694
rect 7870 13746 7922 13758
rect 7870 13682 7922 13694
rect 8430 13746 8482 13758
rect 26462 13746 26514 13758
rect 9986 13694 9998 13746
rect 10050 13694 10062 13746
rect 13794 13694 13806 13746
rect 13858 13694 13870 13746
rect 14242 13694 14254 13746
rect 14306 13694 14318 13746
rect 22194 13694 22206 13746
rect 22258 13694 22270 13746
rect 26002 13694 26014 13746
rect 26066 13694 26078 13746
rect 8430 13682 8482 13694
rect 26462 13682 26514 13694
rect 26798 13746 26850 13758
rect 31166 13746 31218 13758
rect 27458 13694 27470 13746
rect 27522 13694 27534 13746
rect 26798 13682 26850 13694
rect 31166 13682 31218 13694
rect 31726 13746 31778 13758
rect 31726 13682 31778 13694
rect 34078 13746 34130 13758
rect 34078 13682 34130 13694
rect 34526 13746 34578 13758
rect 36654 13746 36706 13758
rect 36194 13694 36206 13746
rect 36258 13694 36270 13746
rect 34526 13682 34578 13694
rect 36654 13682 36706 13694
rect 36766 13746 36818 13758
rect 36766 13682 36818 13694
rect 37326 13746 37378 13758
rect 37326 13682 37378 13694
rect 38334 13746 38386 13758
rect 38334 13682 38386 13694
rect 38558 13746 38610 13758
rect 38558 13682 38610 13694
rect 38894 13746 38946 13758
rect 44046 13746 44098 13758
rect 42578 13694 42590 13746
rect 42642 13694 42654 13746
rect 43474 13694 43486 13746
rect 43538 13694 43550 13746
rect 44258 13694 44270 13746
rect 44322 13694 44334 13746
rect 44594 13694 44606 13746
rect 44658 13694 44670 13746
rect 46834 13694 46846 13746
rect 46898 13694 46910 13746
rect 50306 13694 50318 13746
rect 50370 13694 50382 13746
rect 38894 13682 38946 13694
rect 44046 13682 44098 13694
rect 5070 13634 5122 13646
rect 2482 13582 2494 13634
rect 2546 13582 2558 13634
rect 4610 13582 4622 13634
rect 4674 13582 4686 13634
rect 5070 13570 5122 13582
rect 6302 13634 6354 13646
rect 9550 13634 9602 13646
rect 14478 13634 14530 13646
rect 7970 13582 7982 13634
rect 8034 13582 8046 13634
rect 10322 13582 10334 13634
rect 10386 13582 10398 13634
rect 6302 13570 6354 13582
rect 9550 13570 9602 13582
rect 14478 13570 14530 13582
rect 17390 13634 17442 13646
rect 17390 13570 17442 13582
rect 17950 13634 18002 13646
rect 17950 13570 18002 13582
rect 18398 13634 18450 13646
rect 22766 13634 22818 13646
rect 19394 13582 19406 13634
rect 19458 13582 19470 13634
rect 21522 13582 21534 13634
rect 21586 13582 21598 13634
rect 18398 13570 18450 13582
rect 22766 13570 22818 13582
rect 26686 13634 26738 13646
rect 26686 13570 26738 13582
rect 28254 13634 28306 13646
rect 28254 13570 28306 13582
rect 38110 13634 38162 13646
rect 38110 13570 38162 13582
rect 47182 13634 47234 13646
rect 47182 13570 47234 13582
rect 49086 13634 49138 13646
rect 49086 13570 49138 13582
rect 8206 13522 8258 13534
rect 8206 13458 8258 13470
rect 13022 13522 13074 13534
rect 13022 13458 13074 13470
rect 17614 13522 17666 13534
rect 17614 13458 17666 13470
rect 27806 13522 27858 13534
rect 27806 13458 27858 13470
rect 28142 13522 28194 13534
rect 28142 13458 28194 13470
rect 33406 13522 33458 13534
rect 33406 13458 33458 13470
rect 34302 13522 34354 13534
rect 34302 13458 34354 13470
rect 39454 13522 39506 13534
rect 39454 13458 39506 13470
rect 41806 13522 41858 13534
rect 41806 13458 41858 13470
rect 42142 13522 42194 13534
rect 44594 13470 44606 13522
rect 44658 13470 44670 13522
rect 42142 13458 42194 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 13470 13186 13522 13198
rect 13470 13122 13522 13134
rect 25006 13186 25058 13198
rect 25006 13122 25058 13134
rect 26238 13186 26290 13198
rect 26238 13122 26290 13134
rect 27582 13186 27634 13198
rect 27582 13122 27634 13134
rect 27806 13186 27858 13198
rect 27806 13122 27858 13134
rect 41134 13186 41186 13198
rect 41134 13122 41186 13134
rect 44270 13186 44322 13198
rect 44270 13122 44322 13134
rect 3390 13074 3442 13086
rect 16830 13074 16882 13086
rect 6626 13022 6638 13074
rect 6690 13022 6702 13074
rect 7970 13022 7982 13074
rect 8034 13022 8046 13074
rect 3390 13010 3442 13022
rect 16830 13010 16882 13022
rect 20190 13074 20242 13086
rect 20190 13010 20242 13022
rect 23886 13074 23938 13086
rect 23886 13010 23938 13022
rect 26126 13074 26178 13086
rect 26126 13010 26178 13022
rect 29934 13074 29986 13086
rect 29934 13010 29986 13022
rect 37438 13074 37490 13086
rect 37438 13010 37490 13022
rect 40686 13074 40738 13086
rect 40686 13010 40738 13022
rect 41806 13074 41858 13086
rect 41806 13010 41858 13022
rect 46958 13074 47010 13086
rect 46958 13010 47010 13022
rect 1710 12962 1762 12974
rect 1710 12898 1762 12910
rect 2382 12962 2434 12974
rect 2382 12898 2434 12910
rect 3278 12962 3330 12974
rect 4398 12962 4450 12974
rect 3826 12910 3838 12962
rect 3890 12910 3902 12962
rect 3278 12898 3330 12910
rect 4398 12898 4450 12910
rect 5742 12962 5794 12974
rect 18846 12962 18898 12974
rect 6402 12910 6414 12962
rect 6466 12910 6478 12962
rect 7746 12910 7758 12962
rect 7810 12910 7822 12962
rect 10882 12910 10894 12962
rect 10946 12910 10958 12962
rect 5742 12898 5794 12910
rect 18846 12898 18898 12910
rect 19406 12962 19458 12974
rect 19406 12898 19458 12910
rect 19630 12962 19682 12974
rect 19630 12898 19682 12910
rect 20302 12962 20354 12974
rect 20302 12898 20354 12910
rect 24334 12962 24386 12974
rect 26686 12962 26738 12974
rect 25330 12910 25342 12962
rect 25394 12910 25406 12962
rect 24334 12898 24386 12910
rect 26686 12898 26738 12910
rect 26910 12962 26962 12974
rect 26910 12898 26962 12910
rect 27022 12962 27074 12974
rect 28366 12962 28418 12974
rect 27234 12910 27246 12962
rect 27298 12910 27310 12962
rect 28130 12910 28142 12962
rect 28194 12910 28206 12962
rect 27022 12898 27074 12910
rect 28366 12898 28418 12910
rect 29150 12962 29202 12974
rect 30942 12962 30994 12974
rect 29362 12910 29374 12962
rect 29426 12910 29438 12962
rect 29150 12898 29202 12910
rect 30942 12898 30994 12910
rect 31614 12962 31666 12974
rect 31614 12898 31666 12910
rect 33854 12962 33906 12974
rect 42142 12962 42194 12974
rect 38770 12910 38782 12962
rect 38834 12910 38846 12962
rect 33854 12898 33906 12910
rect 42142 12898 42194 12910
rect 42366 12962 42418 12974
rect 42366 12898 42418 12910
rect 42590 12962 42642 12974
rect 42590 12898 42642 12910
rect 43038 12962 43090 12974
rect 43038 12898 43090 12910
rect 43374 12962 43426 12974
rect 43374 12898 43426 12910
rect 2718 12850 2770 12862
rect 2718 12786 2770 12798
rect 4286 12850 4338 12862
rect 4286 12786 4338 12798
rect 4846 12850 4898 12862
rect 4846 12786 4898 12798
rect 7086 12850 7138 12862
rect 7086 12786 7138 12798
rect 8430 12850 8482 12862
rect 8430 12786 8482 12798
rect 19182 12850 19234 12862
rect 19182 12786 19234 12798
rect 24110 12850 24162 12862
rect 24110 12786 24162 12798
rect 24670 12850 24722 12862
rect 24670 12786 24722 12798
rect 25118 12850 25170 12862
rect 25118 12786 25170 12798
rect 31390 12850 31442 12862
rect 31390 12786 31442 12798
rect 31950 12850 32002 12862
rect 31950 12786 32002 12798
rect 32062 12850 32114 12862
rect 32062 12786 32114 12798
rect 33182 12850 33234 12862
rect 33182 12786 33234 12798
rect 33406 12850 33458 12862
rect 33406 12786 33458 12798
rect 41022 12850 41074 12862
rect 41022 12786 41074 12798
rect 41134 12850 41186 12862
rect 41134 12786 41186 12798
rect 44158 12850 44210 12862
rect 44158 12786 44210 12798
rect 3502 12738 3554 12750
rect 2034 12686 2046 12738
rect 2098 12686 2110 12738
rect 3502 12674 3554 12686
rect 4062 12738 4114 12750
rect 4062 12674 4114 12686
rect 10670 12738 10722 12750
rect 10670 12674 10722 12686
rect 13582 12738 13634 12750
rect 13582 12674 13634 12686
rect 13694 12738 13746 12750
rect 13694 12674 13746 12686
rect 19070 12738 19122 12750
rect 19070 12674 19122 12686
rect 20078 12738 20130 12750
rect 20078 12674 20130 12686
rect 24222 12738 24274 12750
rect 24222 12674 24274 12686
rect 26014 12738 26066 12750
rect 26014 12674 26066 12686
rect 26798 12738 26850 12750
rect 26798 12674 26850 12686
rect 28254 12738 28306 12750
rect 28254 12674 28306 12686
rect 28478 12738 28530 12750
rect 28478 12674 28530 12686
rect 31502 12738 31554 12750
rect 31502 12674 31554 12686
rect 32286 12738 32338 12750
rect 32286 12674 32338 12686
rect 33294 12738 33346 12750
rect 33294 12674 33346 12686
rect 34302 12738 34354 12750
rect 42366 12738 42418 12750
rect 38546 12686 38558 12738
rect 38610 12686 38622 12738
rect 34302 12674 34354 12686
rect 42366 12674 42418 12686
rect 43150 12738 43202 12750
rect 43150 12674 43202 12686
rect 44046 12738 44098 12750
rect 44046 12674 44098 12686
rect 47070 12738 47122 12750
rect 47070 12674 47122 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 2046 12402 2098 12414
rect 3390 12402 3442 12414
rect 2818 12350 2830 12402
rect 2882 12350 2894 12402
rect 2046 12338 2098 12350
rect 3390 12338 3442 12350
rect 4174 12402 4226 12414
rect 4174 12338 4226 12350
rect 4510 12402 4562 12414
rect 4510 12338 4562 12350
rect 5854 12402 5906 12414
rect 5854 12338 5906 12350
rect 9774 12402 9826 12414
rect 9774 12338 9826 12350
rect 13134 12402 13186 12414
rect 13134 12338 13186 12350
rect 14702 12402 14754 12414
rect 14702 12338 14754 12350
rect 17614 12402 17666 12414
rect 19742 12402 19794 12414
rect 18610 12350 18622 12402
rect 18674 12350 18686 12402
rect 17614 12338 17666 12350
rect 19742 12338 19794 12350
rect 19966 12402 20018 12414
rect 19966 12338 20018 12350
rect 26686 12402 26738 12414
rect 26686 12338 26738 12350
rect 26798 12402 26850 12414
rect 26798 12338 26850 12350
rect 26910 12402 26962 12414
rect 26910 12338 26962 12350
rect 29822 12402 29874 12414
rect 29822 12338 29874 12350
rect 30382 12402 30434 12414
rect 30382 12338 30434 12350
rect 33182 12402 33234 12414
rect 33182 12338 33234 12350
rect 33854 12402 33906 12414
rect 33854 12338 33906 12350
rect 34750 12402 34802 12414
rect 34750 12338 34802 12350
rect 38782 12402 38834 12414
rect 38782 12338 38834 12350
rect 40350 12402 40402 12414
rect 40350 12338 40402 12350
rect 6414 12290 6466 12302
rect 4834 12238 4846 12290
rect 4898 12238 4910 12290
rect 6414 12226 6466 12238
rect 6862 12290 6914 12302
rect 6862 12226 6914 12238
rect 7086 12290 7138 12302
rect 7086 12226 7138 12238
rect 8430 12290 8482 12302
rect 8430 12226 8482 12238
rect 8766 12290 8818 12302
rect 8766 12226 8818 12238
rect 9998 12290 10050 12302
rect 9998 12226 10050 12238
rect 11790 12290 11842 12302
rect 11790 12226 11842 12238
rect 12686 12290 12738 12302
rect 12686 12226 12738 12238
rect 13918 12290 13970 12302
rect 13918 12226 13970 12238
rect 14478 12290 14530 12302
rect 14478 12226 14530 12238
rect 15822 12290 15874 12302
rect 17950 12290 18002 12302
rect 16594 12238 16606 12290
rect 16658 12238 16670 12290
rect 15822 12226 15874 12238
rect 17950 12226 18002 12238
rect 19182 12290 19234 12302
rect 19182 12226 19234 12238
rect 19294 12290 19346 12302
rect 19294 12226 19346 12238
rect 19518 12290 19570 12302
rect 19518 12226 19570 12238
rect 20638 12290 20690 12302
rect 20638 12226 20690 12238
rect 20750 12290 20802 12302
rect 26238 12290 26290 12302
rect 29598 12290 29650 12302
rect 22530 12238 22542 12290
rect 22594 12238 22606 12290
rect 28802 12238 28814 12290
rect 28866 12238 28878 12290
rect 20750 12226 20802 12238
rect 26238 12226 26290 12238
rect 29598 12226 29650 12238
rect 30718 12290 30770 12302
rect 30718 12226 30770 12238
rect 32510 12290 32562 12302
rect 32510 12226 32562 12238
rect 33294 12290 33346 12302
rect 33294 12226 33346 12238
rect 33966 12290 34018 12302
rect 33966 12226 34018 12238
rect 34974 12290 35026 12302
rect 34974 12226 35026 12238
rect 35198 12290 35250 12302
rect 35198 12226 35250 12238
rect 37102 12290 37154 12302
rect 37102 12226 37154 12238
rect 37774 12290 37826 12302
rect 37774 12226 37826 12238
rect 38670 12290 38722 12302
rect 38670 12226 38722 12238
rect 39230 12290 39282 12302
rect 39230 12226 39282 12238
rect 40910 12290 40962 12302
rect 40910 12226 40962 12238
rect 42142 12290 42194 12302
rect 42142 12226 42194 12238
rect 42366 12290 42418 12302
rect 46174 12290 46226 12302
rect 43586 12238 43598 12290
rect 43650 12238 43662 12290
rect 42366 12226 42418 12238
rect 46174 12226 46226 12238
rect 1710 12178 1762 12190
rect 1710 12114 1762 12126
rect 2494 12178 2546 12190
rect 2494 12114 2546 12126
rect 3166 12178 3218 12190
rect 3166 12114 3218 12126
rect 3838 12178 3890 12190
rect 3838 12114 3890 12126
rect 5294 12178 5346 12190
rect 8990 12178 9042 12190
rect 12126 12178 12178 12190
rect 6066 12126 6078 12178
rect 6130 12126 6142 12178
rect 10322 12126 10334 12178
rect 10386 12126 10398 12178
rect 5294 12114 5346 12126
rect 8990 12114 9042 12126
rect 12126 12114 12178 12126
rect 12238 12178 12290 12190
rect 12238 12114 12290 12126
rect 12910 12178 12962 12190
rect 12910 12114 12962 12126
rect 13246 12178 13298 12190
rect 13246 12114 13298 12126
rect 13582 12178 13634 12190
rect 13582 12114 13634 12126
rect 14142 12178 14194 12190
rect 17390 12178 17442 12190
rect 15474 12126 15486 12178
rect 15538 12126 15550 12178
rect 16370 12126 16382 12178
rect 16434 12126 16446 12178
rect 14142 12114 14194 12126
rect 17390 12114 17442 12126
rect 17726 12178 17778 12190
rect 20414 12178 20466 12190
rect 25342 12178 25394 12190
rect 27358 12178 27410 12190
rect 29486 12178 29538 12190
rect 18386 12126 18398 12178
rect 18450 12126 18462 12178
rect 21858 12126 21870 12178
rect 21922 12126 21934 12178
rect 25778 12126 25790 12178
rect 25842 12126 25854 12178
rect 27570 12126 27582 12178
rect 27634 12126 27646 12178
rect 27906 12126 27918 12178
rect 27970 12126 27982 12178
rect 29138 12126 29150 12178
rect 29202 12126 29214 12178
rect 17726 12114 17778 12126
rect 20414 12114 20466 12126
rect 25342 12114 25394 12126
rect 27358 12114 27410 12126
rect 29486 12114 29538 12126
rect 30270 12178 30322 12190
rect 30270 12114 30322 12126
rect 30494 12178 30546 12190
rect 32958 12178 33010 12190
rect 31602 12126 31614 12178
rect 31666 12126 31678 12178
rect 30494 12114 30546 12126
rect 32958 12114 33010 12126
rect 33742 12178 33794 12190
rect 33742 12114 33794 12126
rect 34414 12178 34466 12190
rect 34414 12114 34466 12126
rect 34526 12178 34578 12190
rect 34526 12114 34578 12126
rect 36206 12178 36258 12190
rect 36206 12114 36258 12126
rect 36766 12178 36818 12190
rect 41470 12178 41522 12190
rect 38210 12126 38222 12178
rect 38274 12126 38286 12178
rect 38434 12126 38446 12178
rect 38498 12126 38510 12178
rect 42802 12126 42814 12178
rect 42866 12126 42878 12178
rect 36766 12114 36818 12126
rect 41470 12114 41522 12126
rect 3278 12066 3330 12078
rect 3278 12002 3330 12014
rect 8542 12066 8594 12078
rect 8542 12002 8594 12014
rect 10110 12066 10162 12078
rect 10110 12002 10162 12014
rect 11902 12066 11954 12078
rect 11902 12002 11954 12014
rect 13694 12066 13746 12078
rect 13694 12002 13746 12014
rect 14590 12066 14642 12078
rect 19854 12066 19906 12078
rect 32062 12066 32114 12078
rect 15586 12014 15598 12066
rect 15650 12014 15662 12066
rect 24658 12014 24670 12066
rect 24722 12014 24734 12066
rect 29026 12014 29038 12066
rect 29090 12014 29102 12066
rect 14590 12002 14642 12014
rect 19854 12002 19906 12014
rect 32062 12002 32114 12014
rect 39118 12066 39170 12078
rect 42466 12014 42478 12066
rect 42530 12014 42542 12066
rect 45714 12014 45726 12066
rect 45778 12014 45790 12066
rect 39118 12002 39170 12014
rect 6078 11954 6130 11966
rect 6078 11890 6130 11902
rect 6750 11954 6802 11966
rect 6750 11890 6802 11902
rect 20750 11954 20802 11966
rect 20750 11890 20802 11902
rect 37214 11954 37266 11966
rect 37214 11890 37266 11902
rect 37886 11954 37938 11966
rect 37886 11890 37938 11902
rect 39006 11954 39058 11966
rect 39006 11890 39058 11902
rect 41022 11954 41074 11966
rect 41022 11890 41074 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 9102 11618 9154 11630
rect 38222 11618 38274 11630
rect 43038 11618 43090 11630
rect 14802 11566 14814 11618
rect 14866 11566 14878 11618
rect 27346 11566 27358 11618
rect 27410 11566 27422 11618
rect 41794 11566 41806 11618
rect 41858 11566 41870 11618
rect 9102 11554 9154 11566
rect 38222 11554 38274 11566
rect 43038 11554 43090 11566
rect 5070 11506 5122 11518
rect 2482 11454 2494 11506
rect 2546 11454 2558 11506
rect 4610 11454 4622 11506
rect 4674 11454 4686 11506
rect 5070 11442 5122 11454
rect 5742 11506 5794 11518
rect 5742 11442 5794 11454
rect 9214 11506 9266 11518
rect 9214 11442 9266 11454
rect 9998 11506 10050 11518
rect 9998 11442 10050 11454
rect 11342 11506 11394 11518
rect 28366 11506 28418 11518
rect 27122 11454 27134 11506
rect 27186 11454 27198 11506
rect 11342 11442 11394 11454
rect 28366 11442 28418 11454
rect 34302 11506 34354 11518
rect 36094 11506 36146 11518
rect 35186 11454 35198 11506
rect 35250 11454 35262 11506
rect 34302 11442 34354 11454
rect 36094 11442 36146 11454
rect 41246 11506 41298 11518
rect 49310 11506 49362 11518
rect 45826 11454 45838 11506
rect 45890 11454 45902 11506
rect 41246 11442 41298 11454
rect 49310 11442 49362 11454
rect 6078 11394 6130 11406
rect 11678 11394 11730 11406
rect 13582 11394 13634 11406
rect 1810 11342 1822 11394
rect 1874 11342 1886 11394
rect 9426 11342 9438 11394
rect 9490 11342 9502 11394
rect 12226 11342 12238 11394
rect 12290 11342 12302 11394
rect 12786 11342 12798 11394
rect 12850 11342 12862 11394
rect 6078 11330 6130 11342
rect 11678 11330 11730 11342
rect 13582 11330 13634 11342
rect 13694 11394 13746 11406
rect 13694 11330 13746 11342
rect 14030 11394 14082 11406
rect 25902 11394 25954 11406
rect 14690 11342 14702 11394
rect 14754 11342 14766 11394
rect 15026 11342 15038 11394
rect 15090 11342 15102 11394
rect 15698 11342 15710 11394
rect 15762 11342 15774 11394
rect 16930 11342 16942 11394
rect 16994 11342 17006 11394
rect 20738 11342 20750 11394
rect 20802 11342 20814 11394
rect 25330 11342 25342 11394
rect 25394 11342 25406 11394
rect 14030 11330 14082 11342
rect 25902 11330 25954 11342
rect 26014 11394 26066 11406
rect 26014 11330 26066 11342
rect 26574 11394 26626 11406
rect 30270 11394 30322 11406
rect 27458 11342 27470 11394
rect 27522 11342 27534 11394
rect 26574 11330 26626 11342
rect 30270 11330 30322 11342
rect 30942 11394 30994 11406
rect 30942 11330 30994 11342
rect 31278 11394 31330 11406
rect 32174 11394 32226 11406
rect 31826 11342 31838 11394
rect 31890 11342 31902 11394
rect 31278 11330 31330 11342
rect 32174 11330 32226 11342
rect 32846 11394 32898 11406
rect 32846 11330 32898 11342
rect 33630 11394 33682 11406
rect 33630 11330 33682 11342
rect 34078 11394 34130 11406
rect 34078 11330 34130 11342
rect 34526 11394 34578 11406
rect 34526 11330 34578 11342
rect 34638 11394 34690 11406
rect 38782 11394 38834 11406
rect 35410 11342 35422 11394
rect 35474 11342 35486 11394
rect 37090 11342 37102 11394
rect 37154 11342 37166 11394
rect 37762 11342 37774 11394
rect 37826 11342 37838 11394
rect 38210 11342 38222 11394
rect 38274 11342 38286 11394
rect 34638 11330 34690 11342
rect 38782 11330 38834 11342
rect 39118 11394 39170 11406
rect 39790 11394 39842 11406
rect 39330 11342 39342 11394
rect 39394 11342 39406 11394
rect 39118 11330 39170 11342
rect 39790 11330 39842 11342
rect 40350 11394 40402 11406
rect 40786 11342 40798 11394
rect 40850 11342 40862 11394
rect 41570 11342 41582 11394
rect 41634 11342 41646 11394
rect 43362 11342 43374 11394
rect 43426 11342 43438 11394
rect 47954 11342 47966 11394
rect 48018 11342 48030 11394
rect 48738 11342 48750 11394
rect 48802 11342 48814 11394
rect 40350 11330 40402 11342
rect 5630 11282 5682 11294
rect 5630 11218 5682 11230
rect 5966 11282 6018 11294
rect 19518 11282 19570 11294
rect 29934 11282 29986 11294
rect 15810 11230 15822 11282
rect 15874 11230 15886 11282
rect 17042 11230 17054 11282
rect 17106 11230 17118 11282
rect 25554 11230 25566 11282
rect 25618 11230 25630 11282
rect 5966 11218 6018 11230
rect 19518 11218 19570 11230
rect 29934 11218 29986 11230
rect 30046 11282 30098 11294
rect 30046 11218 30098 11230
rect 30718 11282 30770 11294
rect 30718 11218 30770 11230
rect 31502 11282 31554 11294
rect 31502 11218 31554 11230
rect 37214 11282 37266 11294
rect 37214 11218 37266 11230
rect 38894 11282 38946 11294
rect 38894 11218 38946 11230
rect 39678 11282 39730 11294
rect 42254 11282 42306 11294
rect 42130 11230 42142 11282
rect 42194 11230 42206 11282
rect 39678 11218 39730 11230
rect 42254 11218 42306 11230
rect 42366 11282 42418 11294
rect 42366 11218 42418 11230
rect 42702 11282 42754 11294
rect 42702 11218 42754 11230
rect 11790 11170 11842 11182
rect 11790 11106 11842 11118
rect 11902 11170 11954 11182
rect 11902 11106 11954 11118
rect 12014 11170 12066 11182
rect 13806 11170 13858 11182
rect 12562 11118 12574 11170
rect 12626 11118 12638 11170
rect 12014 11106 12066 11118
rect 13806 11106 13858 11118
rect 13918 11170 13970 11182
rect 24894 11170 24946 11182
rect 17154 11118 17166 11170
rect 17218 11118 17230 11170
rect 13918 11106 13970 11118
rect 24894 11106 24946 11118
rect 26126 11170 26178 11182
rect 26126 11106 26178 11118
rect 30606 11170 30658 11182
rect 30606 11106 30658 11118
rect 31390 11170 31442 11182
rect 31390 11106 31442 11118
rect 32286 11170 32338 11182
rect 32286 11106 32338 11118
rect 32398 11170 32450 11182
rect 32398 11106 32450 11118
rect 33070 11170 33122 11182
rect 33070 11106 33122 11118
rect 39902 11170 39954 11182
rect 39902 11106 39954 11118
rect 42926 11170 42978 11182
rect 42926 11106 42978 11118
rect 43486 11170 43538 11182
rect 43486 11106 43538 11118
rect 44158 11170 44210 11182
rect 44158 11106 44210 11118
rect 44942 11170 44994 11182
rect 44942 11106 44994 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 2046 10834 2098 10846
rect 2046 10770 2098 10782
rect 2718 10834 2770 10846
rect 3950 10834 4002 10846
rect 5518 10834 5570 10846
rect 3378 10782 3390 10834
rect 3442 10782 3454 10834
rect 4834 10782 4846 10834
rect 4898 10782 4910 10834
rect 2718 10770 2770 10782
rect 3950 10770 4002 10782
rect 5518 10770 5570 10782
rect 7310 10834 7362 10846
rect 7310 10770 7362 10782
rect 8654 10834 8706 10846
rect 17950 10834 18002 10846
rect 13234 10782 13246 10834
rect 13298 10782 13310 10834
rect 8654 10770 8706 10782
rect 17950 10770 18002 10782
rect 26798 10834 26850 10846
rect 26798 10770 26850 10782
rect 33742 10834 33794 10846
rect 33742 10770 33794 10782
rect 34638 10834 34690 10846
rect 34638 10770 34690 10782
rect 36206 10834 36258 10846
rect 36206 10770 36258 10782
rect 37326 10834 37378 10846
rect 37326 10770 37378 10782
rect 38558 10834 38610 10846
rect 38558 10770 38610 10782
rect 39006 10834 39058 10846
rect 39006 10770 39058 10782
rect 39566 10834 39618 10846
rect 39566 10770 39618 10782
rect 42254 10834 42306 10846
rect 42254 10770 42306 10782
rect 43598 10834 43650 10846
rect 43598 10770 43650 10782
rect 1710 10722 1762 10734
rect 1710 10658 1762 10670
rect 2382 10722 2434 10734
rect 2382 10658 2434 10670
rect 4286 10722 4338 10734
rect 4286 10658 4338 10670
rect 4398 10722 4450 10734
rect 6750 10722 6802 10734
rect 12126 10722 12178 10734
rect 16830 10722 16882 10734
rect 34526 10722 34578 10734
rect 5842 10670 5854 10722
rect 5906 10670 5918 10722
rect 9650 10670 9662 10722
rect 9714 10670 9726 10722
rect 13794 10670 13806 10722
rect 13858 10670 13870 10722
rect 15362 10670 15374 10722
rect 15426 10670 15438 10722
rect 19954 10670 19966 10722
rect 20018 10670 20030 10722
rect 27234 10670 27246 10722
rect 27298 10670 27310 10722
rect 4398 10658 4450 10670
rect 6750 10658 6802 10670
rect 12126 10658 12178 10670
rect 16830 10658 16882 10670
rect 34526 10658 34578 10670
rect 36990 10722 37042 10734
rect 36990 10658 37042 10670
rect 37102 10722 37154 10734
rect 37102 10658 37154 10670
rect 37886 10722 37938 10734
rect 42590 10722 42642 10734
rect 41458 10670 41470 10722
rect 41522 10670 41534 10722
rect 37886 10658 37938 10670
rect 42590 10658 42642 10670
rect 42814 10722 42866 10734
rect 43250 10670 43262 10722
rect 43314 10670 43326 10722
rect 42814 10658 42866 10670
rect 3054 10610 3106 10622
rect 3054 10546 3106 10558
rect 5182 10610 5234 10622
rect 5182 10546 5234 10558
rect 6190 10610 6242 10622
rect 6190 10546 6242 10558
rect 6526 10610 6578 10622
rect 6526 10546 6578 10558
rect 8430 10610 8482 10622
rect 8430 10546 8482 10558
rect 8766 10610 8818 10622
rect 8766 10546 8818 10558
rect 8990 10610 9042 10622
rect 16270 10610 16322 10622
rect 9538 10558 9550 10610
rect 9602 10558 9614 10610
rect 11554 10558 11566 10610
rect 11618 10558 11630 10610
rect 14466 10558 14478 10610
rect 14530 10558 14542 10610
rect 14802 10558 14814 10610
rect 14866 10558 14878 10610
rect 8990 10546 9042 10558
rect 16270 10546 16322 10558
rect 16606 10610 16658 10622
rect 16606 10546 16658 10558
rect 18174 10610 18226 10622
rect 27582 10610 27634 10622
rect 18498 10558 18510 10610
rect 18562 10558 18574 10610
rect 19282 10558 19294 10610
rect 19346 10558 19358 10610
rect 18174 10546 18226 10558
rect 27582 10546 27634 10558
rect 33182 10610 33234 10622
rect 35758 10610 35810 10622
rect 34850 10558 34862 10610
rect 34914 10558 34926 10610
rect 33182 10546 33234 10558
rect 35758 10546 35810 10558
rect 35982 10610 36034 10622
rect 35982 10546 36034 10558
rect 36094 10610 36146 10622
rect 36094 10546 36146 10558
rect 38222 10610 38274 10622
rect 39778 10558 39790 10610
rect 39842 10558 39854 10610
rect 41234 10558 41246 10610
rect 41298 10558 41310 10610
rect 44706 10558 44718 10610
rect 44770 10558 44782 10610
rect 45154 10558 45166 10610
rect 45218 10558 45230 10610
rect 38222 10546 38274 10558
rect 6302 10498 6354 10510
rect 16718 10498 16770 10510
rect 15026 10446 15038 10498
rect 15090 10446 15102 10498
rect 6302 10434 6354 10446
rect 16718 10434 16770 10446
rect 18062 10498 18114 10510
rect 22542 10498 22594 10510
rect 22082 10446 22094 10498
rect 22146 10446 22158 10498
rect 18062 10434 18114 10446
rect 22542 10434 22594 10446
rect 23550 10498 23602 10510
rect 23550 10434 23602 10446
rect 31278 10498 31330 10510
rect 31278 10434 31330 10446
rect 33854 10498 33906 10510
rect 33854 10434 33906 10446
rect 39118 10498 39170 10510
rect 42914 10446 42926 10498
rect 42978 10446 42990 10498
rect 44034 10446 44046 10498
rect 44098 10446 44110 10498
rect 39118 10434 39170 10446
rect 4398 10386 4450 10398
rect 4398 10322 4450 10334
rect 23438 10386 23490 10398
rect 35534 10386 35586 10398
rect 30930 10334 30942 10386
rect 30994 10383 31006 10386
rect 31266 10383 31278 10386
rect 30994 10337 31278 10383
rect 30994 10334 31006 10337
rect 31266 10334 31278 10337
rect 31330 10334 31342 10386
rect 23438 10322 23490 10334
rect 35534 10322 35586 10334
rect 37662 10386 37714 10398
rect 37662 10322 37714 10334
rect 38446 10386 38498 10398
rect 38446 10322 38498 10334
rect 39454 10386 39506 10398
rect 39454 10322 39506 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 7086 10050 7138 10062
rect 7086 9986 7138 9998
rect 11902 10050 11954 10062
rect 11902 9986 11954 9998
rect 14366 10050 14418 10062
rect 14366 9986 14418 9998
rect 18510 10050 18562 10062
rect 18510 9986 18562 9998
rect 35870 10050 35922 10062
rect 35870 9986 35922 9998
rect 37550 10050 37602 10062
rect 37550 9986 37602 9998
rect 13582 9938 13634 9950
rect 4834 9886 4846 9938
rect 4898 9886 4910 9938
rect 8530 9886 8542 9938
rect 8594 9886 8606 9938
rect 10658 9886 10670 9938
rect 10722 9886 10734 9938
rect 13582 9874 13634 9886
rect 16830 9938 16882 9950
rect 34190 9938 34242 9950
rect 22978 9886 22990 9938
rect 23042 9886 23054 9938
rect 25106 9886 25118 9938
rect 25170 9886 25182 9938
rect 26674 9886 26686 9938
rect 26738 9886 26750 9938
rect 29698 9886 29710 9938
rect 29762 9886 29774 9938
rect 16830 9874 16882 9886
rect 34190 9874 34242 9886
rect 34638 9938 34690 9950
rect 34638 9874 34690 9886
rect 34862 9938 34914 9950
rect 34862 9874 34914 9886
rect 36542 9938 36594 9950
rect 36542 9874 36594 9886
rect 37214 9938 37266 9950
rect 37214 9874 37266 9886
rect 38782 9938 38834 9950
rect 41234 9886 41246 9938
rect 41298 9886 41310 9938
rect 38782 9874 38834 9886
rect 5518 9826 5570 9838
rect 2034 9774 2046 9826
rect 2098 9774 2110 9826
rect 5518 9762 5570 9774
rect 5966 9826 6018 9838
rect 5966 9762 6018 9774
rect 6190 9826 6242 9838
rect 11790 9826 11842 9838
rect 7522 9774 7534 9826
rect 7586 9774 7598 9826
rect 11330 9774 11342 9826
rect 11394 9774 11406 9826
rect 6190 9762 6242 9774
rect 11790 9762 11842 9774
rect 12350 9826 12402 9838
rect 12350 9762 12402 9774
rect 12910 9826 12962 9838
rect 12910 9762 12962 9774
rect 13358 9826 13410 9838
rect 13358 9762 13410 9774
rect 13918 9826 13970 9838
rect 13918 9762 13970 9774
rect 16270 9826 16322 9838
rect 16270 9762 16322 9774
rect 17054 9826 17106 9838
rect 17054 9762 17106 9774
rect 17726 9826 17778 9838
rect 17726 9762 17778 9774
rect 18622 9826 18674 9838
rect 18622 9762 18674 9774
rect 19070 9826 19122 9838
rect 19070 9762 19122 9774
rect 19854 9826 19906 9838
rect 27022 9826 27074 9838
rect 27806 9826 27858 9838
rect 22194 9774 22206 9826
rect 22258 9774 22270 9826
rect 27234 9774 27246 9826
rect 27298 9774 27310 9826
rect 19854 9762 19906 9774
rect 27022 9762 27074 9774
rect 27806 9762 27858 9774
rect 28030 9826 28082 9838
rect 35422 9826 35474 9838
rect 43374 9826 43426 9838
rect 32610 9774 32622 9826
rect 32674 9774 32686 9826
rect 39106 9774 39118 9826
rect 39170 9774 39182 9826
rect 41122 9774 41134 9826
rect 41186 9774 41198 9826
rect 28030 9762 28082 9774
rect 35422 9762 35474 9774
rect 43374 9762 43426 9774
rect 43486 9826 43538 9838
rect 43922 9774 43934 9826
rect 43986 9774 43998 9826
rect 43486 9762 43538 9774
rect 6078 9714 6130 9726
rect 12686 9714 12738 9726
rect 2706 9662 2718 9714
rect 2770 9662 2782 9714
rect 7746 9662 7758 9714
rect 7810 9662 7822 9714
rect 6078 9650 6130 9662
rect 12686 9650 12738 9662
rect 13806 9714 13858 9726
rect 13806 9650 13858 9662
rect 14478 9714 14530 9726
rect 14478 9650 14530 9662
rect 17502 9714 17554 9726
rect 17502 9650 17554 9662
rect 18510 9714 18562 9726
rect 28254 9714 28306 9726
rect 35758 9714 35810 9726
rect 19394 9662 19406 9714
rect 19458 9662 19470 9714
rect 31826 9662 31838 9714
rect 31890 9662 31902 9714
rect 37550 9714 37602 9726
rect 18510 9650 18562 9662
rect 28254 9650 28306 9662
rect 35758 9650 35810 9662
rect 37438 9658 37490 9670
rect 6750 9602 6802 9614
rect 6750 9538 6802 9550
rect 12462 9602 12514 9614
rect 12462 9538 12514 9550
rect 17614 9602 17666 9614
rect 17614 9538 17666 9550
rect 21870 9602 21922 9614
rect 21870 9538 21922 9550
rect 26686 9602 26738 9614
rect 26686 9538 26738 9550
rect 26798 9602 26850 9614
rect 26798 9538 26850 9550
rect 27694 9602 27746 9614
rect 27694 9538 27746 9550
rect 27918 9602 27970 9614
rect 27918 9538 27970 9550
rect 33070 9602 33122 9614
rect 39218 9662 39230 9714
rect 39282 9662 39294 9714
rect 42802 9662 42814 9714
rect 42866 9662 42878 9714
rect 37550 9650 37602 9662
rect 37438 9594 37490 9606
rect 43598 9602 43650 9614
rect 33070 9538 33122 9550
rect 43598 9538 43650 9550
rect 43710 9602 43762 9614
rect 45166 9602 45218 9614
rect 44818 9550 44830 9602
rect 44882 9550 44894 9602
rect 43710 9538 43762 9550
rect 45166 9538 45218 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 2158 9266 2210 9278
rect 2158 9202 2210 9214
rect 2494 9266 2546 9278
rect 2494 9202 2546 9214
rect 3838 9266 3890 9278
rect 3838 9202 3890 9214
rect 8430 9266 8482 9278
rect 8430 9202 8482 9214
rect 9550 9266 9602 9278
rect 9550 9202 9602 9214
rect 9774 9266 9826 9278
rect 9774 9202 9826 9214
rect 10446 9266 10498 9278
rect 10446 9202 10498 9214
rect 12574 9266 12626 9278
rect 12574 9202 12626 9214
rect 16046 9266 16098 9278
rect 16046 9202 16098 9214
rect 16270 9266 16322 9278
rect 16270 9202 16322 9214
rect 22430 9266 22482 9278
rect 22430 9202 22482 9214
rect 22654 9266 22706 9278
rect 23662 9266 23714 9278
rect 22978 9214 22990 9266
rect 23042 9214 23054 9266
rect 22654 9202 22706 9214
rect 23662 9202 23714 9214
rect 23774 9266 23826 9278
rect 23774 9202 23826 9214
rect 23886 9266 23938 9278
rect 23886 9202 23938 9214
rect 24670 9266 24722 9278
rect 33742 9266 33794 9278
rect 29138 9214 29150 9266
rect 29202 9214 29214 9266
rect 24670 9202 24722 9214
rect 33742 9202 33794 9214
rect 34526 9266 34578 9278
rect 34526 9202 34578 9214
rect 34974 9266 35026 9278
rect 34974 9202 35026 9214
rect 35086 9266 35138 9278
rect 40014 9266 40066 9278
rect 35858 9214 35870 9266
rect 35922 9214 35934 9266
rect 35086 9202 35138 9214
rect 40014 9202 40066 9214
rect 40126 9266 40178 9278
rect 40126 9202 40178 9214
rect 42366 9266 42418 9278
rect 42366 9202 42418 9214
rect 46062 9266 46114 9278
rect 46062 9202 46114 9214
rect 24110 9154 24162 9166
rect 10770 9102 10782 9154
rect 10834 9102 10846 9154
rect 19506 9102 19518 9154
rect 19570 9102 19582 9154
rect 24110 9090 24162 9102
rect 28590 9154 28642 9166
rect 28590 9090 28642 9102
rect 33966 9154 34018 9166
rect 33966 9090 34018 9102
rect 35310 9154 35362 9166
rect 35310 9090 35362 9102
rect 35534 9154 35586 9166
rect 39790 9154 39842 9166
rect 39106 9102 39118 9154
rect 39170 9102 39182 9154
rect 35534 9090 35586 9102
rect 39790 9090 39842 9102
rect 40910 9154 40962 9166
rect 40910 9090 40962 9102
rect 4622 9042 4674 9054
rect 10222 9042 10274 9054
rect 5058 8990 5070 9042
rect 5122 8990 5134 9042
rect 4622 8978 4674 8990
rect 10222 8978 10274 8990
rect 12686 9042 12738 9054
rect 12686 8978 12738 8990
rect 15934 9042 15986 9054
rect 20750 9042 20802 9054
rect 29486 9042 29538 9054
rect 37214 9042 37266 9054
rect 41022 9042 41074 9054
rect 20178 8990 20190 9042
rect 20242 8990 20254 9042
rect 23426 8990 23438 9042
rect 23490 8990 23502 9042
rect 25218 8990 25230 9042
rect 25282 8990 25294 9042
rect 30258 8990 30270 9042
rect 30322 8990 30334 9042
rect 36082 8990 36094 9042
rect 36146 8990 36158 9042
rect 37650 8990 37662 9042
rect 37714 8990 37726 9042
rect 38210 8990 38222 9042
rect 38274 8990 38286 9042
rect 39554 8990 39566 9042
rect 39618 8990 39630 9042
rect 41346 8990 41358 9042
rect 41410 8990 41422 9042
rect 42690 8990 42702 9042
rect 42754 8990 42766 9042
rect 15934 8978 15986 8990
rect 20750 8978 20802 8990
rect 29486 8978 29538 8990
rect 37214 8978 37266 8990
rect 41022 8978 41074 8990
rect 8766 8930 8818 8942
rect 5730 8878 5742 8930
rect 5794 8878 5806 8930
rect 7858 8878 7870 8930
rect 7922 8878 7934 8930
rect 8766 8866 8818 8878
rect 9662 8930 9714 8942
rect 30830 8930 30882 8942
rect 39902 8930 39954 8942
rect 17378 8878 17390 8930
rect 17442 8878 17454 8930
rect 26002 8878 26014 8930
rect 26066 8878 26078 8930
rect 28130 8878 28142 8930
rect 28194 8878 28206 8930
rect 30034 8878 30046 8930
rect 30098 8878 30110 8930
rect 35074 8878 35086 8930
rect 35138 8878 35150 8930
rect 43474 8878 43486 8930
rect 43538 8878 43550 8930
rect 45602 8878 45614 8930
rect 45666 8878 45678 8930
rect 9662 8866 9714 8878
rect 30830 8866 30882 8878
rect 39902 8866 39954 8878
rect 12574 8818 12626 8830
rect 12574 8754 12626 8766
rect 28478 8818 28530 8830
rect 28478 8754 28530 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 26126 8482 26178 8494
rect 26126 8418 26178 8430
rect 43486 8482 43538 8494
rect 43486 8418 43538 8430
rect 11230 8370 11282 8382
rect 26238 8370 26290 8382
rect 38334 8370 38386 8382
rect 43598 8370 43650 8382
rect 8082 8318 8094 8370
rect 8146 8318 8158 8370
rect 10210 8318 10222 8370
rect 10274 8318 10286 8370
rect 15586 8318 15598 8370
rect 15650 8318 15662 8370
rect 17714 8318 17726 8370
rect 17778 8318 17790 8370
rect 32162 8318 32174 8370
rect 32226 8318 32238 8370
rect 34290 8318 34302 8370
rect 34354 8318 34366 8370
rect 39666 8318 39678 8370
rect 39730 8318 39742 8370
rect 11230 8306 11282 8318
rect 26238 8306 26290 8318
rect 38334 8306 38386 8318
rect 43598 8306 43650 8318
rect 6302 8258 6354 8270
rect 10446 8258 10498 8270
rect 7298 8206 7310 8258
rect 7362 8206 7374 8258
rect 6302 8194 6354 8206
rect 10446 8194 10498 8206
rect 10782 8258 10834 8270
rect 10782 8194 10834 8206
rect 12014 8258 12066 8270
rect 12014 8194 12066 8206
rect 12238 8258 12290 8270
rect 13470 8258 13522 8270
rect 12562 8206 12574 8258
rect 12626 8206 12638 8258
rect 12238 8194 12290 8206
rect 13470 8194 13522 8206
rect 13694 8258 13746 8270
rect 14254 8258 14306 8270
rect 14018 8206 14030 8258
rect 14082 8206 14094 8258
rect 13694 8194 13746 8206
rect 14254 8194 14306 8206
rect 14590 8258 14642 8270
rect 18958 8258 19010 8270
rect 18498 8206 18510 8258
rect 18562 8206 18574 8258
rect 31490 8206 31502 8258
rect 31554 8206 31566 8258
rect 35410 8206 35422 8258
rect 35474 8206 35486 8258
rect 35970 8206 35982 8258
rect 36034 8206 36046 8258
rect 38882 8206 38894 8258
rect 38946 8206 38958 8258
rect 42578 8206 42590 8258
rect 42642 8206 42654 8258
rect 14590 8194 14642 8206
rect 18958 8194 19010 8206
rect 5966 8146 6018 8158
rect 5966 8082 6018 8094
rect 10670 8146 10722 8158
rect 42926 8146 42978 8158
rect 34738 8094 34750 8146
rect 34802 8094 34814 8146
rect 38658 8094 38670 8146
rect 38722 8094 38734 8146
rect 41794 8094 41806 8146
rect 41858 8094 41870 8146
rect 10670 8082 10722 8094
rect 42926 8082 42978 8094
rect 43038 8146 43090 8158
rect 43038 8082 43090 8094
rect 12126 8034 12178 8046
rect 12126 7970 12178 7982
rect 13582 8034 13634 8046
rect 13582 7970 13634 7982
rect 14478 8034 14530 8046
rect 14478 7970 14530 7982
rect 38222 8034 38274 8046
rect 38222 7970 38274 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 8094 7698 8146 7710
rect 8094 7634 8146 7646
rect 8990 7698 9042 7710
rect 8990 7634 9042 7646
rect 27022 7698 27074 7710
rect 27022 7634 27074 7646
rect 36430 7698 36482 7710
rect 36430 7634 36482 7646
rect 40126 7698 40178 7710
rect 40126 7634 40178 7646
rect 41134 7698 41186 7710
rect 41134 7634 41186 7646
rect 41246 7698 41298 7710
rect 41246 7634 41298 7646
rect 41358 7698 41410 7710
rect 41358 7634 41410 7646
rect 41470 7698 41522 7710
rect 41470 7634 41522 7646
rect 42814 7698 42866 7710
rect 42814 7634 42866 7646
rect 41694 7586 41746 7598
rect 10546 7534 10558 7586
rect 10610 7534 10622 7586
rect 15138 7534 15150 7586
rect 15202 7534 15214 7586
rect 28130 7534 28142 7586
rect 28194 7534 28206 7586
rect 37538 7534 37550 7586
rect 37602 7534 37614 7586
rect 41694 7522 41746 7534
rect 16382 7474 16434 7486
rect 9762 7422 9774 7474
rect 9826 7422 9838 7474
rect 15922 7422 15934 7474
rect 15986 7422 15998 7474
rect 27346 7422 27358 7474
rect 27410 7422 27422 7474
rect 33170 7422 33182 7474
rect 33234 7422 33246 7474
rect 36866 7422 36878 7474
rect 36930 7422 36942 7474
rect 16382 7410 16434 7422
rect 12674 7310 12686 7362
rect 12738 7310 12750 7362
rect 13010 7310 13022 7362
rect 13074 7310 13086 7362
rect 30258 7310 30270 7362
rect 30322 7310 30334 7362
rect 33842 7310 33854 7362
rect 33906 7310 33918 7362
rect 35970 7310 35982 7362
rect 36034 7310 36046 7362
rect 39666 7310 39678 7362
rect 39730 7310 39742 7362
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 34638 6914 34690 6926
rect 34638 6850 34690 6862
rect 35310 6802 35362 6814
rect 35310 6738 35362 6750
rect 34850 6638 34862 6690
rect 34914 6687 34926 6690
rect 35074 6687 35086 6690
rect 34914 6641 35086 6687
rect 34914 6638 34926 6641
rect 35074 6638 35086 6641
rect 35138 6638 35150 6690
rect 34750 6578 34802 6590
rect 34750 6514 34802 6526
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 11454 6130 11506 6142
rect 11454 6066 11506 6078
rect 12562 5966 12574 6018
rect 12626 5966 12638 6018
rect 11778 5854 11790 5906
rect 11842 5854 11854 5906
rect 14690 5742 14702 5794
rect 14754 5742 14766 5794
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 38546 4510 38558 4562
rect 38610 4510 38622 4562
rect 38770 4286 38782 4338
rect 38834 4286 38846 4338
rect 17614 4226 17666 4238
rect 17614 4162 17666 4174
rect 18174 4226 18226 4238
rect 18174 4162 18226 4174
rect 30942 4226 30994 4238
rect 30942 4162 30994 4174
rect 31950 4226 32002 4238
rect 31950 4162 32002 4174
rect 32622 4226 32674 4238
rect 32622 4162 32674 4174
rect 33294 4226 33346 4238
rect 33294 4162 33346 4174
rect 34190 4226 34242 4238
rect 34190 4162 34242 4174
rect 34862 4226 34914 4238
rect 34862 4162 34914 4174
rect 35758 4226 35810 4238
rect 35758 4162 35810 4174
rect 36430 4226 36482 4238
rect 36430 4162 36482 4174
rect 37102 4226 37154 4238
rect 37102 4162 37154 4174
rect 37774 4226 37826 4238
rect 37774 4162 37826 4174
rect 38334 4226 38386 4238
rect 38334 4162 38386 4174
rect 39342 4226 39394 4238
rect 39342 4162 39394 4174
rect 39790 4226 39842 4238
rect 39790 4162 39842 4174
rect 40350 4226 40402 4238
rect 40350 4162 40402 4174
rect 37762 4062 37774 4114
rect 37826 4111 37838 4114
rect 38210 4111 38222 4114
rect 37826 4065 38222 4111
rect 37826 4062 37838 4065
rect 38210 4062 38222 4065
rect 38274 4062 38286 4114
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 24994 3614 25006 3666
rect 25058 3614 25070 3666
rect 33954 3614 33966 3666
rect 34018 3614 34030 3666
rect 29150 3554 29202 3566
rect 18610 3502 18622 3554
rect 18674 3502 18686 3554
rect 29150 3490 29202 3502
rect 31166 3554 31218 3566
rect 31166 3490 31218 3502
rect 32174 3554 32226 3566
rect 32174 3490 32226 3502
rect 32846 3554 32898 3566
rect 32846 3490 32898 3502
rect 33518 3554 33570 3566
rect 33518 3490 33570 3502
rect 34414 3554 34466 3566
rect 39006 3554 39058 3566
rect 36194 3502 36206 3554
rect 36258 3502 36270 3554
rect 36866 3502 36878 3554
rect 36930 3502 36942 3554
rect 37538 3502 37550 3554
rect 37602 3502 37614 3554
rect 38210 3502 38222 3554
rect 38274 3502 38286 3554
rect 34414 3490 34466 3502
rect 39006 3490 39058 3502
rect 39790 3554 39842 3566
rect 40674 3502 40686 3554
rect 40738 3502 40750 3554
rect 39790 3490 39842 3502
rect 16494 3442 16546 3454
rect 16494 3378 16546 3390
rect 17054 3442 17106 3454
rect 17054 3378 17106 3390
rect 17390 3442 17442 3454
rect 17390 3378 17442 3390
rect 17726 3442 17778 3454
rect 18398 3442 18450 3454
rect 18050 3390 18062 3442
rect 18114 3390 18126 3442
rect 17726 3378 17778 3390
rect 18398 3378 18450 3390
rect 24110 3442 24162 3454
rect 24110 3378 24162 3390
rect 24558 3442 24610 3454
rect 24558 3378 24610 3390
rect 29822 3442 29874 3454
rect 29822 3378 29874 3390
rect 30158 3442 30210 3454
rect 30158 3378 30210 3390
rect 30494 3442 30546 3454
rect 31502 3442 31554 3454
rect 33182 3442 33234 3454
rect 35086 3442 35138 3454
rect 36654 3442 36706 3454
rect 30818 3390 30830 3442
rect 30882 3390 30894 3442
rect 32498 3390 32510 3442
rect 32562 3390 32574 3442
rect 34738 3390 34750 3442
rect 34802 3390 34814 3442
rect 35410 3390 35422 3442
rect 35474 3390 35486 3442
rect 35970 3390 35982 3442
rect 36034 3390 36046 3442
rect 30494 3378 30546 3390
rect 31502 3378 31554 3390
rect 33182 3378 33234 3390
rect 35086 3378 35138 3390
rect 36654 3378 36706 3390
rect 37326 3442 37378 3454
rect 40462 3442 40514 3454
rect 37986 3390 37998 3442
rect 38050 3390 38062 3442
rect 38658 3390 38670 3442
rect 38722 3390 38734 3442
rect 40114 3390 40126 3442
rect 40178 3390 40190 3442
rect 37326 3378 37378 3390
rect 40462 3378 40514 3390
rect 29598 3330 29650 3342
rect 29598 3266 29650 3278
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
rect 35634 2494 35646 2546
rect 35698 2543 35710 2546
rect 36418 2543 36430 2546
rect 35698 2497 36430 2543
rect 35698 2494 35710 2497
rect 36418 2494 36430 2497
rect 36482 2543 36494 2546
rect 36866 2543 36878 2546
rect 36482 2497 36878 2543
rect 36482 2494 36494 2497
rect 36866 2494 36878 2497
rect 36930 2494 36942 2546
rect 36978 2382 36990 2434
rect 37042 2431 37054 2434
rect 38210 2431 38222 2434
rect 37042 2385 38222 2431
rect 37042 2382 37054 2385
rect 38210 2382 38222 2385
rect 38274 2382 38286 2434
<< via1 >>
rect 19182 56590 19234 56642
rect 20078 56590 20130 56642
rect 23998 56590 24050 56642
rect 25006 56590 25058 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 19182 56254 19234 56306
rect 33182 56254 33234 56306
rect 20190 56030 20242 56082
rect 23998 56030 24050 56082
rect 27358 56030 27410 56082
rect 29486 56030 29538 56082
rect 32398 56030 32450 56082
rect 35982 56030 36034 56082
rect 42814 56030 42866 56082
rect 46174 56030 46226 56082
rect 46622 56030 46674 56082
rect 49534 56030 49586 56082
rect 50430 56030 50482 56082
rect 24670 55918 24722 55970
rect 30942 55918 30994 55970
rect 35310 55918 35362 55970
rect 36766 55918 36818 55970
rect 39006 55918 39058 55970
rect 40014 55918 40066 55970
rect 42142 55918 42194 55970
rect 47630 55918 47682 55970
rect 22990 55806 23042 55858
rect 24558 55806 24610 55858
rect 26798 55806 26850 55858
rect 43822 55806 43874 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 35758 55470 35810 55522
rect 14590 55358 14642 55410
rect 20750 55358 20802 55410
rect 24222 55358 24274 55410
rect 26350 55358 26402 55410
rect 33742 55358 33794 55410
rect 37102 55358 37154 55410
rect 40574 55358 40626 55410
rect 42142 55358 42194 55410
rect 45502 55358 45554 55410
rect 51662 55358 51714 55410
rect 17502 55246 17554 55298
rect 17950 55246 18002 55298
rect 23550 55246 23602 55298
rect 30942 55246 30994 55298
rect 37662 55246 37714 55298
rect 40910 55246 40962 55298
rect 48414 55246 48466 55298
rect 48750 55246 48802 55298
rect 16718 55134 16770 55186
rect 18622 55134 18674 55186
rect 28478 55134 28530 55186
rect 31614 55134 31666 55186
rect 35646 55134 35698 55186
rect 36318 55134 36370 55186
rect 38446 55134 38498 55186
rect 43934 55134 43986 55186
rect 47630 55134 47682 55186
rect 49534 55134 49586 55186
rect 28366 55022 28418 55074
rect 34190 55022 34242 55074
rect 34638 55022 34690 55074
rect 35086 55022 35138 55074
rect 36206 55022 36258 55074
rect 43822 55022 43874 55074
rect 44942 55022 44994 55074
rect 52110 55022 52162 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 16718 54686 16770 54738
rect 17726 54686 17778 54738
rect 18510 54686 18562 54738
rect 23662 54686 23714 54738
rect 25678 54686 25730 54738
rect 31390 54686 31442 54738
rect 34190 54686 34242 54738
rect 38334 54686 38386 54738
rect 39006 54686 39058 54738
rect 39790 54686 39842 54738
rect 41246 54686 41298 54738
rect 42030 54686 42082 54738
rect 46286 54686 46338 54738
rect 46398 54686 46450 54738
rect 48078 54686 48130 54738
rect 48862 54686 48914 54738
rect 49422 54686 49474 54738
rect 16830 54574 16882 54626
rect 25566 54574 25618 54626
rect 27022 54574 27074 54626
rect 28366 54574 28418 54626
rect 32174 54574 32226 54626
rect 33630 54574 33682 54626
rect 35534 54574 35586 54626
rect 38222 54574 38274 54626
rect 39118 54574 39170 54626
rect 40126 54574 40178 54626
rect 41918 54574 41970 54626
rect 43374 54574 43426 54626
rect 17502 54462 17554 54514
rect 17614 54462 17666 54514
rect 17838 54462 17890 54514
rect 18062 54462 18114 54514
rect 18958 54462 19010 54514
rect 24670 54462 24722 54514
rect 25454 54462 25506 54514
rect 26574 54462 26626 54514
rect 27694 54462 27746 54514
rect 32510 54462 32562 54514
rect 33182 54462 33234 54514
rect 33294 54462 33346 54514
rect 34750 54462 34802 54514
rect 37998 54462 38050 54514
rect 38446 54462 38498 54514
rect 38558 54462 38610 54514
rect 39566 54462 39618 54514
rect 39678 54462 39730 54514
rect 39902 54462 39954 54514
rect 40910 54462 40962 54514
rect 41134 54462 41186 54514
rect 41358 54462 41410 54514
rect 41582 54462 41634 54514
rect 42590 54462 42642 54514
rect 46062 54462 46114 54514
rect 46510 54462 46562 54514
rect 46622 54462 46674 54514
rect 47070 54462 47122 54514
rect 47294 54462 47346 54514
rect 47518 54462 47570 54514
rect 47742 54462 47794 54514
rect 53006 54462 53058 54514
rect 53566 54462 53618 54514
rect 18398 54350 18450 54402
rect 19630 54350 19682 54402
rect 21758 54350 21810 54402
rect 30494 54350 30546 54402
rect 30942 54350 30994 54402
rect 31390 54350 31442 54402
rect 33518 54350 33570 54402
rect 33966 54350 34018 54402
rect 34190 54350 34242 54402
rect 37662 54350 37714 54402
rect 45502 54350 45554 54402
rect 47406 54350 47458 54402
rect 48190 54350 48242 54402
rect 49310 54350 49362 54402
rect 49870 54350 49922 54402
rect 50206 54350 50258 54402
rect 52334 54350 52386 54402
rect 31614 54238 31666 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 16718 53790 16770 53842
rect 17390 53790 17442 53842
rect 19854 53790 19906 53842
rect 26574 53790 26626 53842
rect 27246 53790 27298 53842
rect 27806 53790 27858 53842
rect 29262 53790 29314 53842
rect 31390 53790 31442 53842
rect 33518 53790 33570 53842
rect 37662 53790 37714 53842
rect 41918 53790 41970 53842
rect 44158 53790 44210 53842
rect 44942 53790 44994 53842
rect 45614 53790 45666 53842
rect 48974 53790 49026 53842
rect 49534 53790 49586 53842
rect 50766 53790 50818 53842
rect 51438 53790 51490 53842
rect 13806 53678 13858 53730
rect 17614 53678 17666 53730
rect 18846 53678 18898 53730
rect 19294 53678 19346 53730
rect 19742 53678 19794 53730
rect 23214 53678 23266 53730
rect 23774 53678 23826 53730
rect 28366 53678 28418 53730
rect 29150 53678 29202 53730
rect 29374 53678 29426 53730
rect 29822 53678 29874 53730
rect 30718 53678 30770 53730
rect 33854 53678 33906 53730
rect 37774 53678 37826 53730
rect 39118 53678 39170 53730
rect 43150 53678 43202 53730
rect 43598 53678 43650 53730
rect 43822 53678 43874 53730
rect 48414 53678 48466 53730
rect 49646 53678 49698 53730
rect 50430 53678 50482 53730
rect 51550 53678 51602 53730
rect 14590 53566 14642 53618
rect 17054 53566 17106 53618
rect 18398 53566 18450 53618
rect 18958 53566 19010 53618
rect 19182 53566 19234 53618
rect 20190 53566 20242 53618
rect 20414 53566 20466 53618
rect 22654 53566 22706 53618
rect 24446 53566 24498 53618
rect 27806 53566 27858 53618
rect 35422 53566 35474 53618
rect 38222 53566 38274 53618
rect 39790 53566 39842 53618
rect 42254 53566 42306 53618
rect 42926 53566 42978 53618
rect 44158 53566 44210 53618
rect 47742 53566 47794 53618
rect 50094 53566 50146 53618
rect 50878 53566 50930 53618
rect 51102 53566 51154 53618
rect 17278 53454 17330 53506
rect 17502 53454 17554 53506
rect 18062 53454 18114 53506
rect 19070 53454 19122 53506
rect 19966 53454 20018 53506
rect 21646 53454 21698 53506
rect 22094 53454 22146 53506
rect 22318 53454 22370 53506
rect 22990 53454 23042 53506
rect 27358 53454 27410 53506
rect 27918 53454 27970 53506
rect 28142 53454 28194 53506
rect 29598 53454 29650 53506
rect 37214 53454 37266 53506
rect 37662 53454 37714 53506
rect 37998 53454 38050 53506
rect 38670 53454 38722 53506
rect 42590 53454 42642 53506
rect 44046 53454 44098 53506
rect 44830 53454 44882 53506
rect 49534 53454 49586 53506
rect 49870 53454 49922 53506
rect 50654 53454 50706 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 15486 53118 15538 53170
rect 19630 53118 19682 53170
rect 24110 53118 24162 53170
rect 24334 53118 24386 53170
rect 25342 53118 25394 53170
rect 30158 53118 30210 53170
rect 30718 53118 30770 53170
rect 31614 53118 31666 53170
rect 32510 53118 32562 53170
rect 34078 53118 34130 53170
rect 36990 53118 37042 53170
rect 41022 53118 41074 53170
rect 41470 53118 41522 53170
rect 41918 53118 41970 53170
rect 45614 53118 45666 53170
rect 46174 53118 46226 53170
rect 46286 53118 46338 53170
rect 46510 53118 46562 53170
rect 46958 53118 47010 53170
rect 47742 53118 47794 53170
rect 49086 53118 49138 53170
rect 15598 53006 15650 53058
rect 17390 53006 17442 53058
rect 17726 53006 17778 53058
rect 18174 53006 18226 53058
rect 24446 53006 24498 53058
rect 25678 53006 25730 53058
rect 25902 53006 25954 53058
rect 27582 53006 27634 53058
rect 31838 53006 31890 53058
rect 40238 53006 40290 53058
rect 44158 53006 44210 53058
rect 47630 53006 47682 53058
rect 19742 52894 19794 52946
rect 20750 52894 20802 52946
rect 24222 52894 24274 52946
rect 24670 52894 24722 52946
rect 25454 52894 25506 52946
rect 26910 52894 26962 52946
rect 31502 52894 31554 52946
rect 31950 52894 32002 52946
rect 33518 52894 33570 52946
rect 35982 52894 36034 52946
rect 39230 52894 39282 52946
rect 39566 52894 39618 52946
rect 39790 52894 39842 52946
rect 44942 52894 44994 52946
rect 45390 52894 45442 52946
rect 46062 52894 46114 52946
rect 46398 52894 46450 52946
rect 47182 52894 47234 52946
rect 48750 52894 48802 52946
rect 50878 52894 50930 52946
rect 51326 52894 51378 52946
rect 51662 52894 51714 52946
rect 52446 52894 52498 52946
rect 18622 52782 18674 52834
rect 21422 52782 21474 52834
rect 23550 52782 23602 52834
rect 25342 52782 25394 52834
rect 29710 52782 29762 52834
rect 30606 52782 30658 52834
rect 39342 52782 39394 52834
rect 39902 52782 39954 52834
rect 40126 52782 40178 52834
rect 48190 52782 48242 52834
rect 49534 52782 49586 52834
rect 50430 52782 50482 52834
rect 51214 52782 51266 52834
rect 54574 52782 54626 52834
rect 30494 52670 30546 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 18174 52334 18226 52386
rect 18398 52334 18450 52386
rect 24558 52334 24610 52386
rect 26798 52334 26850 52386
rect 31390 52334 31442 52386
rect 48750 52334 48802 52386
rect 49534 52334 49586 52386
rect 16382 52222 16434 52274
rect 18958 52222 19010 52274
rect 20638 52222 20690 52274
rect 24222 52222 24274 52274
rect 24670 52222 24722 52274
rect 46622 52222 46674 52274
rect 48750 52222 48802 52274
rect 51214 52222 51266 52274
rect 13582 52110 13634 52162
rect 16830 52110 16882 52162
rect 17838 52110 17890 52162
rect 17950 52110 18002 52162
rect 19182 52110 19234 52162
rect 20414 52110 20466 52162
rect 20750 52110 20802 52162
rect 21982 52110 22034 52162
rect 22094 52110 22146 52162
rect 22430 52110 22482 52162
rect 25230 52110 25282 52162
rect 26238 52110 26290 52162
rect 29374 52110 29426 52162
rect 29598 52110 29650 52162
rect 29822 52110 29874 52162
rect 30382 52110 30434 52162
rect 33294 52110 33346 52162
rect 37326 52110 37378 52162
rect 39566 52110 39618 52162
rect 40014 52110 40066 52162
rect 45166 52110 45218 52162
rect 49310 52110 49362 52162
rect 49758 52110 49810 52162
rect 50318 52110 50370 52162
rect 50766 52110 50818 52162
rect 51326 52110 51378 52162
rect 14254 51998 14306 52050
rect 18846 51998 18898 52050
rect 21870 51998 21922 52050
rect 30046 51998 30098 52050
rect 34078 51998 34130 52050
rect 37662 51998 37714 52050
rect 38558 51998 38610 52050
rect 41806 51998 41858 52050
rect 51214 51998 51266 52050
rect 17838 51886 17890 51938
rect 25454 51886 25506 51938
rect 36318 51886 36370 51938
rect 40238 51886 40290 51938
rect 49982 51886 50034 51938
rect 50094 51886 50146 51938
rect 50206 51886 50258 51938
rect 50990 51886 51042 51938
rect 52782 51886 52834 51938
rect 53230 51886 53282 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 14478 51550 14530 51602
rect 16046 51550 16098 51602
rect 29150 51550 29202 51602
rect 33070 51550 33122 51602
rect 34638 51550 34690 51602
rect 39006 51550 39058 51602
rect 44158 51550 44210 51602
rect 16494 51438 16546 51490
rect 18398 51438 18450 51490
rect 23662 51438 23714 51490
rect 30382 51438 30434 51490
rect 33854 51438 33906 51490
rect 34974 51438 35026 51490
rect 39118 51438 39170 51490
rect 39454 51438 39506 51490
rect 39790 51438 39842 51490
rect 42478 51438 42530 51490
rect 45390 51438 45442 51490
rect 46062 51438 46114 51490
rect 47182 51438 47234 51490
rect 47854 51438 47906 51490
rect 52446 51438 52498 51490
rect 15822 51326 15874 51378
rect 16270 51326 16322 51378
rect 17614 51326 17666 51378
rect 21870 51326 21922 51378
rect 22206 51326 22258 51378
rect 22542 51326 22594 51378
rect 23438 51326 23490 51378
rect 25678 51326 25730 51378
rect 29710 51326 29762 51378
rect 33294 51326 33346 51378
rect 33966 51326 34018 51378
rect 34302 51326 34354 51378
rect 34526 51326 34578 51378
rect 34750 51326 34802 51378
rect 35422 51326 35474 51378
rect 38782 51326 38834 51378
rect 40014 51326 40066 51378
rect 40910 51326 40962 51378
rect 43822 51326 43874 51378
rect 45054 51326 45106 51378
rect 46622 51326 46674 51378
rect 46958 51326 47010 51378
rect 51998 51326 52050 51378
rect 52670 51326 52722 51378
rect 53118 51326 53170 51378
rect 53342 51326 53394 51378
rect 53566 51326 53618 51378
rect 53902 51326 53954 51378
rect 14590 51214 14642 51266
rect 16158 51214 16210 51266
rect 20526 51214 20578 51266
rect 22094 51214 22146 51266
rect 22990 51214 23042 51266
rect 26350 51214 26402 51266
rect 28590 51214 28642 51266
rect 32510 51214 32562 51266
rect 36094 51214 36146 51266
rect 38334 51214 38386 51266
rect 39566 51214 39618 51266
rect 46062 51214 46114 51266
rect 46734 51214 46786 51266
rect 47966 51214 48018 51266
rect 49198 51214 49250 51266
rect 51326 51214 51378 51266
rect 52894 51214 52946 51266
rect 53790 51214 53842 51266
rect 46286 51102 46338 51154
rect 48078 51102 48130 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 41134 50766 41186 50818
rect 51886 50766 51938 50818
rect 1934 50654 1986 50706
rect 13694 50654 13746 50706
rect 15822 50654 15874 50706
rect 17054 50654 17106 50706
rect 18622 50654 18674 50706
rect 24222 50654 24274 50706
rect 27582 50654 27634 50706
rect 32062 50654 32114 50706
rect 50430 50654 50482 50706
rect 51998 50654 52050 50706
rect 55582 50654 55634 50706
rect 3838 50542 3890 50594
rect 15374 50542 15426 50594
rect 15710 50542 15762 50594
rect 16158 50542 16210 50594
rect 17166 50542 17218 50594
rect 17502 50542 17554 50594
rect 17838 50542 17890 50594
rect 18734 50542 18786 50594
rect 19070 50542 19122 50594
rect 21422 50542 21474 50594
rect 24558 50542 24610 50594
rect 29150 50542 29202 50594
rect 32622 50542 32674 50594
rect 36430 50542 36482 50594
rect 36990 50542 37042 50594
rect 39118 50542 39170 50594
rect 41918 50542 41970 50594
rect 46398 50542 46450 50594
rect 46846 50542 46898 50594
rect 49534 50542 49586 50594
rect 52670 50542 52722 50594
rect 13582 50430 13634 50482
rect 14926 50430 14978 50482
rect 15822 50430 15874 50482
rect 18062 50430 18114 50482
rect 18510 50430 18562 50482
rect 19742 50430 19794 50482
rect 22094 50430 22146 50482
rect 25342 50430 25394 50482
rect 28366 50430 28418 50482
rect 28478 50430 28530 50482
rect 28590 50430 28642 50482
rect 29934 50430 29986 50482
rect 32734 50430 32786 50482
rect 35310 50430 35362 50482
rect 37102 50430 37154 50482
rect 40798 50430 40850 50482
rect 41246 50430 41298 50482
rect 41358 50430 41410 50482
rect 42254 50430 42306 50482
rect 42590 50430 42642 50482
rect 43038 50430 43090 50482
rect 44942 50430 44994 50482
rect 47406 50430 47458 50482
rect 53454 50430 53506 50482
rect 16046 50318 16098 50370
rect 16942 50318 16994 50370
rect 19406 50318 19458 50370
rect 34862 50318 34914 50370
rect 39790 50318 39842 50370
rect 45054 50318 45106 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 18398 49982 18450 50034
rect 20638 49982 20690 50034
rect 21758 49982 21810 50034
rect 23214 49982 23266 50034
rect 25342 49982 25394 50034
rect 26462 49982 26514 50034
rect 27246 49982 27298 50034
rect 27358 49982 27410 50034
rect 30494 49982 30546 50034
rect 34414 49982 34466 50034
rect 34750 49982 34802 50034
rect 35982 49982 36034 50034
rect 36318 49982 36370 50034
rect 36878 49982 36930 50034
rect 48862 49982 48914 50034
rect 50766 49982 50818 50034
rect 54014 49982 54066 50034
rect 54126 49982 54178 50034
rect 54798 49982 54850 50034
rect 2046 49870 2098 49922
rect 12910 49870 12962 49922
rect 15710 49870 15762 49922
rect 16830 49870 16882 49922
rect 17390 49870 17442 49922
rect 21982 49870 22034 49922
rect 24670 49870 24722 49922
rect 26574 49870 26626 49922
rect 27582 49870 27634 49922
rect 29486 49870 29538 49922
rect 30158 49870 30210 49922
rect 32510 49870 32562 49922
rect 38222 49870 38274 49922
rect 46062 49870 46114 49922
rect 48750 49870 48802 49922
rect 49086 49870 49138 49922
rect 49758 49870 49810 49922
rect 52334 49870 52386 49922
rect 53902 49870 53954 49922
rect 54574 49870 54626 49922
rect 1710 49758 1762 49810
rect 12238 49758 12290 49810
rect 15374 49758 15426 49810
rect 16494 49758 16546 49810
rect 17502 49758 17554 49810
rect 17950 49758 18002 49810
rect 19518 49758 19570 49810
rect 19742 49758 19794 49810
rect 20078 49758 20130 49810
rect 23438 49758 23490 49810
rect 25790 49758 25842 49810
rect 26126 49758 26178 49810
rect 26350 49758 26402 49810
rect 26798 49758 26850 49810
rect 27694 49758 27746 49810
rect 28814 49758 28866 49810
rect 29262 49758 29314 49810
rect 32174 49758 32226 49810
rect 33630 49758 33682 49810
rect 36094 49758 36146 49810
rect 36542 49758 36594 49810
rect 37438 49758 37490 49810
rect 41694 49758 41746 49810
rect 44942 49758 44994 49810
rect 45390 49758 45442 49810
rect 49198 49758 49250 49810
rect 51438 49758 51490 49810
rect 51886 49758 51938 49810
rect 2494 49646 2546 49698
rect 11566 49646 11618 49698
rect 15038 49646 15090 49698
rect 16158 49646 16210 49698
rect 19070 49646 19122 49698
rect 19630 49646 19682 49698
rect 20414 49646 20466 49698
rect 20526 49646 20578 49698
rect 21646 49646 21698 49698
rect 25230 49646 25282 49698
rect 25678 49646 25730 49698
rect 27470 49646 27522 49698
rect 28254 49646 28306 49698
rect 29038 49646 29090 49698
rect 31838 49646 31890 49698
rect 33294 49646 33346 49698
rect 34078 49646 34130 49698
rect 35198 49646 35250 49698
rect 36206 49646 36258 49698
rect 36990 49646 37042 49698
rect 40350 49646 40402 49698
rect 42366 49646 42418 49698
rect 44494 49646 44546 49698
rect 48190 49646 48242 49698
rect 54798 49646 54850 49698
rect 11454 49534 11506 49586
rect 17726 49534 17778 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 42366 49198 42418 49250
rect 10782 49086 10834 49138
rect 12910 49086 12962 49138
rect 27022 49086 27074 49138
rect 27582 49086 27634 49138
rect 33742 49086 33794 49138
rect 37214 49086 37266 49138
rect 37550 49086 37602 49138
rect 42702 49086 42754 49138
rect 43150 49086 43202 49138
rect 47070 49086 47122 49138
rect 48078 49086 48130 49138
rect 50206 49086 50258 49138
rect 52670 49086 52722 49138
rect 54798 49086 54850 49138
rect 10110 48974 10162 49026
rect 14702 48974 14754 49026
rect 14814 48974 14866 49026
rect 15150 48974 15202 49026
rect 15822 48974 15874 49026
rect 17054 48974 17106 49026
rect 17390 48974 17442 49026
rect 22766 48974 22818 49026
rect 24110 48974 24162 49026
rect 30718 48974 30770 49026
rect 32958 48974 33010 49026
rect 38110 48974 38162 49026
rect 39790 48974 39842 49026
rect 41470 48974 41522 49026
rect 43374 48974 43426 49026
rect 44830 48974 44882 49026
rect 47294 48974 47346 49026
rect 55470 48974 55522 49026
rect 1710 48862 1762 48914
rect 16830 48862 16882 48914
rect 22542 48862 22594 48914
rect 24894 48862 24946 48914
rect 30942 48862 30994 48914
rect 39902 48862 39954 48914
rect 40574 48862 40626 48914
rect 43038 48862 43090 48914
rect 43598 48862 43650 48914
rect 50878 48862 50930 48914
rect 2046 48750 2098 48802
rect 2494 48750 2546 48802
rect 13918 48750 13970 48802
rect 17166 48750 17218 48802
rect 29374 48750 29426 48802
rect 30382 48750 30434 48802
rect 31390 48750 31442 48802
rect 35534 48750 35586 48802
rect 36318 48750 36370 48802
rect 42478 48750 42530 48802
rect 45166 48750 45218 48802
rect 50542 48750 50594 48802
rect 51326 48750 51378 48802
rect 51774 48750 51826 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 12126 48414 12178 48466
rect 12238 48414 12290 48466
rect 13358 48414 13410 48466
rect 25454 48414 25506 48466
rect 30718 48414 30770 48466
rect 36542 48414 36594 48466
rect 38782 48414 38834 48466
rect 41134 48414 41186 48466
rect 42814 48414 42866 48466
rect 45726 48414 45778 48466
rect 51886 48414 51938 48466
rect 2046 48302 2098 48354
rect 17838 48302 17890 48354
rect 20302 48302 20354 48354
rect 25790 48302 25842 48354
rect 31502 48302 31554 48354
rect 42142 48302 42194 48354
rect 43038 48302 43090 48354
rect 43598 48302 43650 48354
rect 45838 48302 45890 48354
rect 46846 48302 46898 48354
rect 47742 48302 47794 48354
rect 1710 48190 1762 48242
rect 11790 48190 11842 48242
rect 12014 48190 12066 48242
rect 12462 48190 12514 48242
rect 14030 48190 14082 48242
rect 19518 48190 19570 48242
rect 25230 48190 25282 48242
rect 25566 48190 25618 48242
rect 30046 48190 30098 48242
rect 30382 48190 30434 48242
rect 30830 48190 30882 48242
rect 30942 48190 30994 48242
rect 31726 48190 31778 48242
rect 31950 48190 32002 48242
rect 33182 48190 33234 48242
rect 36878 48190 36930 48242
rect 37102 48190 37154 48242
rect 37438 48190 37490 48242
rect 37662 48190 37714 48242
rect 37998 48190 38050 48242
rect 38334 48190 38386 48242
rect 41358 48190 41410 48242
rect 41806 48190 41858 48242
rect 42590 48190 42642 48242
rect 42814 48190 42866 48242
rect 43934 48190 43986 48242
rect 45390 48190 45442 48242
rect 46062 48190 46114 48242
rect 46398 48190 46450 48242
rect 47070 48190 47122 48242
rect 47406 48190 47458 48242
rect 48750 48190 48802 48242
rect 52670 48190 52722 48242
rect 2494 48078 2546 48130
rect 12910 48078 12962 48130
rect 14702 48078 14754 48130
rect 16830 48078 16882 48130
rect 17838 48078 17890 48130
rect 22430 48078 22482 48130
rect 24670 48078 24722 48130
rect 27246 48078 27298 48130
rect 29374 48078 29426 48130
rect 33966 48078 34018 48130
rect 36094 48078 36146 48130
rect 36990 48078 37042 48130
rect 37886 48078 37938 48130
rect 40014 48078 40066 48130
rect 40350 48078 40402 48130
rect 42030 48078 42082 48130
rect 46622 48078 46674 48130
rect 48190 48078 48242 48130
rect 49870 48078 49922 48130
rect 53118 48078 53170 48130
rect 17614 47966 17666 48018
rect 32174 47966 32226 48018
rect 32622 47966 32674 48018
rect 51662 47966 51714 48018
rect 51998 47966 52050 48018
rect 52334 47966 52386 48018
rect 52670 47966 52722 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 16382 47630 16434 47682
rect 16718 47630 16770 47682
rect 26798 47630 26850 47682
rect 29262 47630 29314 47682
rect 33294 47630 33346 47682
rect 36430 47630 36482 47682
rect 45838 47630 45890 47682
rect 12462 47518 12514 47570
rect 12910 47518 12962 47570
rect 17838 47518 17890 47570
rect 19966 47518 20018 47570
rect 26910 47518 26962 47570
rect 27806 47518 27858 47570
rect 30718 47518 30770 47570
rect 32846 47518 32898 47570
rect 39902 47518 39954 47570
rect 40350 47518 40402 47570
rect 42142 47518 42194 47570
rect 44270 47518 44322 47570
rect 46846 47518 46898 47570
rect 50206 47518 50258 47570
rect 51102 47518 51154 47570
rect 57934 47518 57986 47570
rect 9662 47406 9714 47458
rect 17166 47406 17218 47458
rect 20302 47406 20354 47458
rect 24334 47406 24386 47458
rect 24894 47406 24946 47458
rect 28366 47406 28418 47458
rect 30046 47406 30098 47458
rect 33182 47406 33234 47458
rect 34078 47406 34130 47458
rect 35198 47406 35250 47458
rect 36094 47406 36146 47458
rect 36990 47406 37042 47458
rect 40126 47406 40178 47458
rect 41470 47406 41522 47458
rect 48974 47406 49026 47458
rect 49646 47406 49698 47458
rect 50990 47406 51042 47458
rect 51214 47406 51266 47458
rect 51438 47406 51490 47458
rect 51886 47406 51938 47458
rect 55582 47406 55634 47458
rect 1710 47294 1762 47346
rect 10334 47294 10386 47346
rect 16494 47294 16546 47346
rect 21310 47294 21362 47346
rect 22766 47294 22818 47346
rect 25342 47294 25394 47346
rect 27022 47294 27074 47346
rect 29150 47294 29202 47346
rect 29262 47294 29314 47346
rect 34974 47294 35026 47346
rect 36318 47294 36370 47346
rect 37774 47294 37826 47346
rect 50654 47294 50706 47346
rect 52110 47294 52162 47346
rect 2046 47182 2098 47234
rect 2494 47182 2546 47234
rect 20638 47182 20690 47234
rect 21646 47182 21698 47234
rect 26350 47182 26402 47234
rect 27694 47182 27746 47234
rect 27918 47182 27970 47234
rect 33294 47182 33346 47234
rect 34190 47182 34242 47234
rect 34302 47182 34354 47234
rect 34526 47182 34578 47234
rect 35758 47182 35810 47234
rect 40462 47182 40514 47234
rect 40686 47182 40738 47234
rect 44942 47182 44994 47234
rect 45950 47182 46002 47234
rect 46062 47182 46114 47234
rect 51774 47182 51826 47234
rect 55246 47182 55298 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 10894 46846 10946 46898
rect 11902 46846 11954 46898
rect 17614 46846 17666 46898
rect 31838 46846 31890 46898
rect 33742 46846 33794 46898
rect 35534 46846 35586 46898
rect 36542 46846 36594 46898
rect 44270 46846 44322 46898
rect 48750 46846 48802 46898
rect 49534 46846 49586 46898
rect 50206 46846 50258 46898
rect 53902 46846 53954 46898
rect 2046 46734 2098 46786
rect 11006 46734 11058 46786
rect 11790 46734 11842 46786
rect 16718 46734 16770 46786
rect 17390 46734 17442 46786
rect 21086 46734 21138 46786
rect 26238 46734 26290 46786
rect 32174 46734 32226 46786
rect 32286 46734 32338 46786
rect 34078 46734 34130 46786
rect 36766 46734 36818 46786
rect 41246 46734 41298 46786
rect 42366 46734 42418 46786
rect 45838 46734 45890 46786
rect 49422 46734 49474 46786
rect 52670 46734 52722 46786
rect 1710 46622 1762 46674
rect 11566 46622 11618 46674
rect 11678 46622 11730 46674
rect 12014 46622 12066 46674
rect 13246 46622 13298 46674
rect 16382 46622 16434 46674
rect 17614 46622 17666 46674
rect 17950 46622 18002 46674
rect 19854 46622 19906 46674
rect 20078 46622 20130 46674
rect 20526 46622 20578 46674
rect 23662 46622 23714 46674
rect 25678 46622 25730 46674
rect 26574 46622 26626 46674
rect 26798 46622 26850 46674
rect 27022 46622 27074 46674
rect 27582 46622 27634 46674
rect 30942 46622 30994 46674
rect 33966 46622 34018 46674
rect 35198 46622 35250 46674
rect 36654 46622 36706 46674
rect 37102 46622 37154 46674
rect 37886 46622 37938 46674
rect 40910 46622 40962 46674
rect 41134 46622 41186 46674
rect 41694 46622 41746 46674
rect 42254 46622 42306 46674
rect 45054 46622 45106 46674
rect 48974 46622 49026 46674
rect 49758 46622 49810 46674
rect 53342 46622 53394 46674
rect 2494 46510 2546 46562
rect 2942 46510 2994 46562
rect 9886 46510 9938 46562
rect 12686 46510 12738 46562
rect 13918 46510 13970 46562
rect 16046 46510 16098 46562
rect 21870 46510 21922 46562
rect 24446 46510 24498 46562
rect 25342 46510 25394 46562
rect 26686 46510 26738 46562
rect 28254 46510 28306 46562
rect 30382 46510 30434 46562
rect 33182 46510 33234 46562
rect 34862 46510 34914 46562
rect 36206 46510 36258 46562
rect 40014 46510 40066 46562
rect 44382 46510 44434 46562
rect 47966 46510 48018 46562
rect 50542 46510 50594 46562
rect 2270 46398 2322 46450
rect 3054 46398 3106 46450
rect 9774 46398 9826 46450
rect 20302 46398 20354 46450
rect 32286 46398 32338 46450
rect 41918 46398 41970 46450
rect 42142 46398 42194 46450
rect 44494 46398 44546 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 13582 46062 13634 46114
rect 14590 46062 14642 46114
rect 20190 46062 20242 46114
rect 26686 46062 26738 46114
rect 48302 46062 48354 46114
rect 48526 46062 48578 46114
rect 9102 45950 9154 46002
rect 11230 45950 11282 46002
rect 11790 45950 11842 46002
rect 13022 45950 13074 46002
rect 14142 45950 14194 46002
rect 14702 45950 14754 46002
rect 15150 45950 15202 46002
rect 19630 45950 19682 46002
rect 20750 45950 20802 46002
rect 23886 45950 23938 46002
rect 26014 45950 26066 46002
rect 26462 45950 26514 46002
rect 31726 45950 31778 46002
rect 33966 45950 34018 46002
rect 37998 45950 38050 46002
rect 40238 45950 40290 46002
rect 40798 45950 40850 46002
rect 42142 45950 42194 46002
rect 48078 45950 48130 46002
rect 49198 45950 49250 46002
rect 50430 45950 50482 46002
rect 54910 45950 54962 46002
rect 57710 45950 57762 46002
rect 1822 45838 1874 45890
rect 8430 45838 8482 45890
rect 11566 45838 11618 45890
rect 13694 45838 13746 45890
rect 13918 45838 13970 45890
rect 15262 45838 15314 45890
rect 15710 45838 15762 45890
rect 19966 45838 20018 45890
rect 20414 45838 20466 45890
rect 20526 45838 20578 45890
rect 21870 45838 21922 45890
rect 22094 45838 22146 45890
rect 23214 45838 23266 45890
rect 26350 45838 26402 45890
rect 28142 45838 28194 45890
rect 28702 45838 28754 45890
rect 32286 45838 32338 45890
rect 33406 45838 33458 45890
rect 40126 45838 40178 45890
rect 41022 45838 41074 45890
rect 43710 45838 43762 45890
rect 45166 45838 45218 45890
rect 45278 45838 45330 45890
rect 47518 45838 47570 45890
rect 48638 45838 48690 45890
rect 52670 45838 52722 45890
rect 55806 45838 55858 45890
rect 2382 45726 2434 45778
rect 3166 45726 3218 45778
rect 11790 45726 11842 45778
rect 12238 45726 12290 45778
rect 14254 45726 14306 45778
rect 18062 45726 18114 45778
rect 18286 45726 18338 45778
rect 22766 45726 22818 45778
rect 32062 45726 32114 45778
rect 41694 45726 41746 45778
rect 45390 45726 45442 45778
rect 47294 45726 47346 45778
rect 47966 45726 48018 45778
rect 51886 45726 51938 45778
rect 2046 45614 2098 45666
rect 2718 45614 2770 45666
rect 12014 45614 12066 45666
rect 15150 45614 15202 45666
rect 15486 45614 15538 45666
rect 18174 45614 18226 45666
rect 21422 45614 21474 45666
rect 27134 45614 27186 45666
rect 28030 45614 28082 45666
rect 28254 45614 28306 45666
rect 29262 45614 29314 45666
rect 32398 45614 32450 45666
rect 32510 45614 32562 45666
rect 35870 45614 35922 45666
rect 39566 45614 39618 45666
rect 39902 45614 39954 45666
rect 40350 45614 40402 45666
rect 43486 45614 43538 45666
rect 45838 45614 45890 45666
rect 51998 45614 52050 45666
rect 52222 45614 52274 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 10670 45278 10722 45330
rect 16606 45278 16658 45330
rect 20638 45278 20690 45330
rect 21422 45278 21474 45330
rect 25342 45278 25394 45330
rect 27022 45278 27074 45330
rect 38334 45278 38386 45330
rect 50878 45278 50930 45330
rect 54686 45278 54738 45330
rect 2046 45166 2098 45218
rect 11230 45166 11282 45218
rect 14926 45166 14978 45218
rect 18174 45166 18226 45218
rect 20974 45166 21026 45218
rect 21758 45166 21810 45218
rect 26238 45166 26290 45218
rect 30606 45166 30658 45218
rect 31390 45166 31442 45218
rect 34414 45166 34466 45218
rect 34526 45166 34578 45218
rect 45054 45166 45106 45218
rect 45166 45166 45218 45218
rect 47182 45166 47234 45218
rect 53342 45166 53394 45218
rect 1710 45054 1762 45106
rect 10782 45054 10834 45106
rect 11006 45054 11058 45106
rect 12126 45054 12178 45106
rect 14366 45054 14418 45106
rect 14702 45054 14754 45106
rect 15262 45054 15314 45106
rect 16270 45054 16322 45106
rect 17502 45054 17554 45106
rect 22094 45054 22146 45106
rect 26014 45054 26066 45106
rect 26798 45054 26850 45106
rect 27470 45054 27522 45106
rect 29486 45054 29538 45106
rect 30382 45054 30434 45106
rect 31166 45054 31218 45106
rect 31726 45054 31778 45106
rect 31950 45054 32002 45106
rect 33406 45054 33458 45106
rect 33854 45054 33906 45106
rect 34750 45054 34802 45106
rect 35086 45054 35138 45106
rect 35758 45054 35810 45106
rect 36318 45054 36370 45106
rect 37326 45054 37378 45106
rect 37886 45054 37938 45106
rect 38670 45054 38722 45106
rect 41582 45054 41634 45106
rect 42814 45054 42866 45106
rect 43150 45054 43202 45106
rect 43486 45054 43538 45106
rect 44270 45054 44322 45106
rect 47630 45054 47682 45106
rect 54014 45054 54066 45106
rect 54462 45054 54514 45106
rect 55134 45054 55186 45106
rect 55470 45054 55522 45106
rect 2494 44942 2546 44994
rect 9774 44942 9826 44994
rect 10894 44942 10946 44994
rect 13246 44942 13298 44994
rect 14814 44942 14866 44994
rect 15374 44942 15426 44994
rect 15822 44942 15874 44994
rect 20302 44942 20354 44994
rect 23214 44942 23266 44994
rect 26910 44942 26962 44994
rect 29934 44942 29986 44994
rect 31502 44942 31554 44994
rect 34078 44942 34130 44994
rect 37998 44942 38050 44994
rect 38894 44942 38946 44994
rect 41806 44942 41858 44994
rect 42254 44942 42306 44994
rect 43262 44942 43314 44994
rect 43822 44942 43874 44994
rect 44718 44942 44770 44994
rect 47406 44942 47458 44994
rect 51214 44942 51266 44994
rect 54574 44942 54626 44994
rect 9662 44830 9714 44882
rect 45166 44830 45218 44882
rect 47854 44830 47906 44882
rect 48302 44830 48354 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 24334 44494 24386 44546
rect 24558 44494 24610 44546
rect 25902 44494 25954 44546
rect 38110 44494 38162 44546
rect 38782 44494 38834 44546
rect 43710 44494 43762 44546
rect 46286 44494 46338 44546
rect 46510 44494 46562 44546
rect 49422 44494 49474 44546
rect 51662 44494 51714 44546
rect 1934 44382 1986 44434
rect 8878 44382 8930 44434
rect 11006 44382 11058 44434
rect 15598 44382 15650 44434
rect 18510 44382 18562 44434
rect 20750 44382 20802 44434
rect 23662 44382 23714 44434
rect 24558 44382 24610 44434
rect 25006 44382 25058 44434
rect 25678 44382 25730 44434
rect 27246 44382 27298 44434
rect 27918 44382 27970 44434
rect 32062 44382 32114 44434
rect 32958 44382 33010 44434
rect 39006 44382 39058 44434
rect 43822 44382 43874 44434
rect 45390 44382 45442 44434
rect 45726 44382 45778 44434
rect 49086 44382 49138 44434
rect 50878 44382 50930 44434
rect 51886 44382 51938 44434
rect 52110 44382 52162 44434
rect 55022 44382 55074 44434
rect 57822 44382 57874 44434
rect 4286 44270 4338 44322
rect 8206 44270 8258 44322
rect 12462 44270 12514 44322
rect 12574 44270 12626 44322
rect 13022 44270 13074 44322
rect 13918 44270 13970 44322
rect 14254 44270 14306 44322
rect 17614 44270 17666 44322
rect 18622 44270 18674 44322
rect 21422 44270 21474 44322
rect 21870 44270 21922 44322
rect 23102 44270 23154 44322
rect 24222 44270 24274 44322
rect 26126 44270 26178 44322
rect 27134 44270 27186 44322
rect 29150 44270 29202 44322
rect 32510 44270 32562 44322
rect 33182 44270 33234 44322
rect 35310 44270 35362 44322
rect 35646 44270 35698 44322
rect 38558 44270 38610 44322
rect 39566 44270 39618 44322
rect 40014 44270 40066 44322
rect 41470 44270 41522 44322
rect 41806 44270 41858 44322
rect 42926 44270 42978 44322
rect 43038 44270 43090 44322
rect 45950 44270 46002 44322
rect 47070 44270 47122 44322
rect 47518 44270 47570 44322
rect 48974 44270 49026 44322
rect 52670 44270 52722 44322
rect 55694 44270 55746 44322
rect 13582 44158 13634 44210
rect 14478 44158 14530 44210
rect 14926 44158 14978 44210
rect 15262 44158 15314 44210
rect 15486 44158 15538 44210
rect 16270 44158 16322 44210
rect 18398 44158 18450 44210
rect 18958 44158 19010 44210
rect 19406 44158 19458 44210
rect 22318 44158 22370 44210
rect 22654 44158 22706 44210
rect 23550 44158 23602 44210
rect 23774 44158 23826 44210
rect 29934 44158 29986 44210
rect 33854 44158 33906 44210
rect 34190 44158 34242 44210
rect 34414 44158 34466 44210
rect 34750 44158 34802 44210
rect 35086 44158 35138 44210
rect 39342 44158 39394 44210
rect 43262 44158 43314 44210
rect 47966 44158 48018 44210
rect 50766 44158 50818 44210
rect 50990 44158 51042 44210
rect 51214 44158 51266 44210
rect 11454 44046 11506 44098
rect 12798 44046 12850 44098
rect 14030 44046 14082 44098
rect 15934 44046 15986 44098
rect 17278 44046 17330 44098
rect 18062 44046 18114 44098
rect 20414 44046 20466 44098
rect 26574 44046 26626 44098
rect 34638 44046 34690 44098
rect 35198 44046 35250 44098
rect 39454 44046 39506 44098
rect 41582 44046 41634 44098
rect 42814 44046 42866 44098
rect 46622 44046 46674 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 10222 43710 10274 43762
rect 27470 43710 27522 43762
rect 29710 43710 29762 43762
rect 33630 43710 33682 43762
rect 42926 43710 42978 43762
rect 49086 43710 49138 43762
rect 2046 43598 2098 43650
rect 4846 43598 4898 43650
rect 5294 43598 5346 43650
rect 17502 43598 17554 43650
rect 19630 43598 19682 43650
rect 19854 43598 19906 43650
rect 19966 43598 20018 43650
rect 20078 43598 20130 43650
rect 22318 43598 22370 43650
rect 23214 43598 23266 43650
rect 23438 43598 23490 43650
rect 23662 43598 23714 43650
rect 24334 43598 24386 43650
rect 27022 43598 27074 43650
rect 29038 43598 29090 43650
rect 29150 43598 29202 43650
rect 33406 43598 33458 43650
rect 33518 43598 33570 43650
rect 35198 43598 35250 43650
rect 37774 43598 37826 43650
rect 40126 43598 40178 43650
rect 40238 43598 40290 43650
rect 43374 43598 43426 43650
rect 48750 43598 48802 43650
rect 48862 43598 48914 43650
rect 49870 43598 49922 43650
rect 49982 43598 50034 43650
rect 53006 43598 53058 43650
rect 53118 43598 53170 43650
rect 1710 43486 1762 43538
rect 8654 43486 8706 43538
rect 9998 43486 10050 43538
rect 10558 43486 10610 43538
rect 13918 43486 13970 43538
rect 17838 43486 17890 43538
rect 20750 43486 20802 43538
rect 23998 43486 24050 43538
rect 25790 43486 25842 43538
rect 27246 43486 27298 43538
rect 29598 43486 29650 43538
rect 29822 43486 29874 43538
rect 30158 43486 30210 43538
rect 32958 43486 33010 43538
rect 34526 43486 34578 43538
rect 37662 43486 37714 43538
rect 39006 43486 39058 43538
rect 42142 43486 42194 43538
rect 42590 43486 42642 43538
rect 42814 43486 42866 43538
rect 46062 43486 46114 43538
rect 47406 43486 47458 43538
rect 50878 43486 50930 43538
rect 51214 43486 51266 43538
rect 51774 43486 51826 43538
rect 52110 43486 52162 43538
rect 53454 43486 53506 43538
rect 2494 43374 2546 43426
rect 5742 43374 5794 43426
rect 7870 43374 7922 43426
rect 11342 43374 11394 43426
rect 13470 43374 13522 43426
rect 14702 43374 14754 43426
rect 16830 43374 16882 43426
rect 20526 43374 20578 43426
rect 21422 43374 21474 43426
rect 22878 43374 22930 43426
rect 23550 43374 23602 43426
rect 26462 43374 26514 43426
rect 27134 43374 27186 43426
rect 28702 43374 28754 43426
rect 37326 43374 37378 43426
rect 38222 43374 38274 43426
rect 39342 43374 39394 43426
rect 41022 43374 41074 43426
rect 43822 43374 43874 43426
rect 46286 43374 46338 43426
rect 46734 43374 46786 43426
rect 47518 43374 47570 43426
rect 51326 43374 51378 43426
rect 51662 43374 51714 43426
rect 4622 43262 4674 43314
rect 4958 43262 5010 43314
rect 5406 43262 5458 43314
rect 22542 43262 22594 43314
rect 26574 43262 26626 43314
rect 29150 43262 29202 43314
rect 39006 43262 39058 43314
rect 40126 43262 40178 43314
rect 42030 43262 42082 43314
rect 43262 43262 43314 43314
rect 48078 43262 48130 43314
rect 49870 43262 49922 43314
rect 55358 43262 55410 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 4062 42926 4114 42978
rect 11230 42926 11282 42978
rect 12014 42926 12066 42978
rect 13470 42926 13522 42978
rect 14366 42926 14418 42978
rect 14702 42926 14754 42978
rect 17950 42926 18002 42978
rect 18174 42926 18226 42978
rect 20526 42926 20578 42978
rect 46286 42926 46338 42978
rect 6078 42814 6130 42866
rect 8878 42814 8930 42866
rect 10446 42814 10498 42866
rect 13582 42814 13634 42866
rect 18286 42814 18338 42866
rect 20078 42814 20130 42866
rect 47518 42814 47570 42866
rect 51214 42814 51266 42866
rect 3390 42702 3442 42754
rect 3726 42702 3778 42754
rect 5630 42702 5682 42754
rect 5854 42702 5906 42754
rect 6750 42702 6802 42754
rect 8318 42702 8370 42754
rect 14702 42702 14754 42754
rect 15486 42702 15538 42754
rect 22542 42702 22594 42754
rect 22766 42702 22818 42754
rect 23326 42702 23378 42754
rect 23886 42702 23938 42754
rect 24334 42702 24386 42754
rect 24558 42702 24610 42754
rect 25118 42702 25170 42754
rect 25678 42702 25730 42754
rect 26910 42702 26962 42754
rect 28142 42702 28194 42754
rect 32510 42702 32562 42754
rect 35422 42702 35474 42754
rect 35534 42702 35586 42754
rect 39006 42702 39058 42754
rect 39678 42702 39730 42754
rect 40126 42702 40178 42754
rect 42142 42702 42194 42754
rect 42590 42702 42642 42754
rect 42814 42702 42866 42754
rect 46398 42702 46450 42754
rect 47406 42702 47458 42754
rect 47630 42702 47682 42754
rect 49422 42702 49474 42754
rect 50430 42702 50482 42754
rect 50766 42702 50818 42754
rect 51438 42702 51490 42754
rect 54798 42702 54850 42754
rect 55582 42702 55634 42754
rect 1710 42590 1762 42642
rect 2046 42590 2098 42642
rect 6190 42590 6242 42642
rect 6862 42590 6914 42642
rect 7534 42590 7586 42642
rect 8094 42590 8146 42642
rect 8766 42590 8818 42642
rect 11342 42590 11394 42642
rect 11566 42590 11618 42642
rect 11902 42590 11954 42642
rect 17838 42590 17890 42642
rect 19070 42590 19122 42642
rect 19406 42590 19458 42642
rect 2494 42478 2546 42530
rect 3950 42478 4002 42530
rect 7646 42478 7698 42530
rect 13694 42478 13746 42530
rect 15150 42478 15202 42530
rect 18734 42478 18786 42530
rect 19518 42478 19570 42530
rect 20414 42534 20466 42586
rect 20526 42590 20578 42642
rect 23774 42590 23826 42642
rect 25342 42590 25394 42642
rect 26350 42590 26402 42642
rect 26574 42590 26626 42642
rect 28254 42590 28306 42642
rect 29262 42590 29314 42642
rect 30382 42590 30434 42642
rect 30718 42590 30770 42642
rect 31278 42590 31330 42642
rect 32734 42590 32786 42642
rect 33742 42590 33794 42642
rect 34078 42590 34130 42642
rect 34414 42590 34466 42642
rect 35870 42590 35922 42642
rect 40350 42590 40402 42642
rect 42366 42590 42418 42642
rect 46286 42590 46338 42642
rect 47854 42590 47906 42642
rect 50654 42590 50706 42642
rect 52110 42590 52162 42642
rect 53678 42590 53730 42642
rect 57374 42590 57426 42642
rect 21870 42478 21922 42530
rect 22318 42478 22370 42530
rect 22990 42478 23042 42530
rect 23102 42478 23154 42530
rect 23662 42478 23714 42530
rect 24782 42478 24834 42530
rect 24894 42478 24946 42530
rect 25566 42478 25618 42530
rect 26686 42478 26738 42530
rect 28478 42478 28530 42530
rect 34750 42478 34802 42530
rect 35758 42478 35810 42530
rect 38446 42478 38498 42530
rect 38670 42478 38722 42530
rect 38894 42478 38946 42530
rect 42478 42478 42530 42530
rect 43486 42478 43538 42530
rect 45054 42478 45106 42530
rect 48862 42478 48914 42530
rect 49086 42478 49138 42530
rect 49310 42478 49362 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 2046 42142 2098 42194
rect 3950 42142 4002 42194
rect 5854 42142 5906 42194
rect 12126 42142 12178 42194
rect 25902 42142 25954 42194
rect 26126 42142 26178 42194
rect 29374 42142 29426 42194
rect 31950 42142 32002 42194
rect 33742 42142 33794 42194
rect 34750 42142 34802 42194
rect 41582 42142 41634 42194
rect 45726 42142 45778 42194
rect 49534 42142 49586 42194
rect 51214 42142 51266 42194
rect 51326 42142 51378 42194
rect 51438 42142 51490 42194
rect 4398 42030 4450 42082
rect 5966 42030 6018 42082
rect 6190 42030 6242 42082
rect 6526 42030 6578 42082
rect 7086 42030 7138 42082
rect 8206 42030 8258 42082
rect 10334 42030 10386 42082
rect 11454 42030 11506 42082
rect 12574 42030 12626 42082
rect 12686 42030 12738 42082
rect 13806 42030 13858 42082
rect 21310 42030 21362 42082
rect 21646 42030 21698 42082
rect 23214 42030 23266 42082
rect 23550 42030 23602 42082
rect 23662 42030 23714 42082
rect 26350 42030 26402 42082
rect 26798 42030 26850 42082
rect 30718 42030 30770 42082
rect 35870 42030 35922 42082
rect 39678 42030 39730 42082
rect 43150 42030 43202 42082
rect 47966 42030 48018 42082
rect 48078 42030 48130 42082
rect 49310 42030 49362 42082
rect 1710 41918 1762 41970
rect 3838 41918 3890 41970
rect 4286 41918 4338 41970
rect 5406 41918 5458 41970
rect 6302 41918 6354 41970
rect 8094 41918 8146 41970
rect 10558 41918 10610 41970
rect 11118 41918 11170 41970
rect 12014 41918 12066 41970
rect 12350 41918 12402 41970
rect 12910 41918 12962 41970
rect 13470 41918 13522 41970
rect 17390 41918 17442 41970
rect 18174 41918 18226 41970
rect 20750 41918 20802 41970
rect 21086 41918 21138 41970
rect 22542 41918 22594 41970
rect 22990 41918 23042 41970
rect 26686 41918 26738 41970
rect 29038 41918 29090 41970
rect 30270 41918 30322 41970
rect 30494 41918 30546 41970
rect 30942 41918 30994 41970
rect 35086 41918 35138 41970
rect 39230 41918 39282 41970
rect 39902 41918 39954 41970
rect 41246 41918 41298 41970
rect 42366 41918 42418 41970
rect 46062 41918 46114 41970
rect 47518 41918 47570 41970
rect 49086 41918 49138 41970
rect 51886 41918 51938 41970
rect 52558 41918 52610 41970
rect 53006 41918 53058 41970
rect 53454 41918 53506 41970
rect 2494 41806 2546 41858
rect 2942 41806 2994 41858
rect 8654 41806 8706 41858
rect 14254 41806 14306 41858
rect 14926 41806 14978 41858
rect 16942 41806 16994 41858
rect 20302 41806 20354 41858
rect 22766 41806 22818 41858
rect 24222 41806 24274 41858
rect 24670 41806 24722 41858
rect 27358 41806 27410 41858
rect 30830 41806 30882 41858
rect 31390 41806 31442 41858
rect 37998 41806 38050 41858
rect 38446 41806 38498 41858
rect 38894 41806 38946 41858
rect 39790 41806 39842 41858
rect 40350 41806 40402 41858
rect 45278 41806 45330 41858
rect 46510 41806 46562 41858
rect 49198 41806 49250 41858
rect 50878 41806 50930 41858
rect 53118 41806 53170 41858
rect 55246 41806 55298 41858
rect 8206 41694 8258 41746
rect 8766 41694 8818 41746
rect 23662 41694 23714 41746
rect 26238 41694 26290 41746
rect 26798 41694 26850 41746
rect 47966 41694 48018 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 13582 41358 13634 41410
rect 12686 41246 12738 41298
rect 20190 41246 20242 41298
rect 22094 41246 22146 41298
rect 28590 41246 28642 41298
rect 31390 41246 31442 41298
rect 33518 41246 33570 41298
rect 36430 41246 36482 41298
rect 37438 41246 37490 41298
rect 39566 41246 39618 41298
rect 41694 41246 41746 41298
rect 42142 41246 42194 41298
rect 43598 41246 43650 41298
rect 51214 41246 51266 41298
rect 55022 41246 55074 41298
rect 57934 41246 57986 41298
rect 1822 41134 1874 41186
rect 7646 41134 7698 41186
rect 8206 41134 8258 41186
rect 10894 41134 10946 41186
rect 13694 41134 13746 41186
rect 14030 41134 14082 41186
rect 14366 41134 14418 41186
rect 15038 41134 15090 41186
rect 15150 41134 15202 41186
rect 15822 41134 15874 41186
rect 19182 41134 19234 41186
rect 19518 41134 19570 41186
rect 22430 41134 22482 41186
rect 22542 41134 22594 41186
rect 23326 41134 23378 41186
rect 23550 41134 23602 41186
rect 23774 41134 23826 41186
rect 23998 41134 24050 41186
rect 24334 41134 24386 41186
rect 25790 41134 25842 41186
rect 30046 41134 30098 41186
rect 30718 41134 30770 41186
rect 34190 41134 34242 41186
rect 38222 41134 38274 41186
rect 38782 41134 38834 41186
rect 42254 41134 42306 41186
rect 42814 41134 42866 41186
rect 43934 41134 43986 41186
rect 45166 41134 45218 41186
rect 47630 41134 47682 41186
rect 47966 41134 48018 41186
rect 48414 41134 48466 41186
rect 52670 41134 52722 41186
rect 55918 41134 55970 41186
rect 2046 41022 2098 41074
rect 2382 41022 2434 41074
rect 2718 41022 2770 41074
rect 3166 41022 3218 41074
rect 6190 41022 6242 41074
rect 8654 41022 8706 41074
rect 13582 41022 13634 41074
rect 14590 41022 14642 41074
rect 14926 41022 14978 41074
rect 15486 41022 15538 41074
rect 16046 41022 16098 41074
rect 19630 41022 19682 41074
rect 19854 41022 19906 41074
rect 24670 41022 24722 41074
rect 25006 41022 25058 41074
rect 26462 41022 26514 41074
rect 38446 41022 38498 41074
rect 45278 41022 45330 41074
rect 46734 41022 46786 41074
rect 47518 41022 47570 41074
rect 49086 41022 49138 41074
rect 6302 40910 6354 40962
rect 14142 40910 14194 40962
rect 15934 40910 15986 40962
rect 16606 40910 16658 40962
rect 18398 40910 18450 40962
rect 18734 40910 18786 40962
rect 18958 40910 19010 40962
rect 19070 40910 19122 40962
rect 21646 40910 21698 40962
rect 22654 40910 22706 40962
rect 22766 40910 22818 40962
rect 23438 40910 23490 40962
rect 24446 40910 24498 40962
rect 29486 40910 29538 40962
rect 34750 40910 34802 40962
rect 35646 40910 35698 40962
rect 36990 40910 37042 40962
rect 45502 40910 45554 40962
rect 45950 40910 46002 40962
rect 46398 40910 46450 40962
rect 47406 40910 47458 40962
rect 51662 40910 51714 40962
rect 52110 40910 52162 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 8654 40574 8706 40626
rect 13358 40574 13410 40626
rect 21422 40574 21474 40626
rect 25342 40574 25394 40626
rect 26686 40574 26738 40626
rect 26798 40574 26850 40626
rect 26910 40574 26962 40626
rect 27918 40574 27970 40626
rect 28814 40574 28866 40626
rect 29934 40574 29986 40626
rect 30942 40574 30994 40626
rect 31614 40574 31666 40626
rect 31950 40574 32002 40626
rect 38110 40574 38162 40626
rect 38670 40574 38722 40626
rect 41470 40574 41522 40626
rect 41694 40574 41746 40626
rect 42030 40574 42082 40626
rect 56590 40574 56642 40626
rect 2046 40462 2098 40514
rect 10334 40462 10386 40514
rect 12798 40462 12850 40514
rect 13582 40462 13634 40514
rect 14702 40462 14754 40514
rect 22542 40462 22594 40514
rect 25678 40462 25730 40514
rect 25790 40462 25842 40514
rect 29822 40462 29874 40514
rect 30718 40462 30770 40514
rect 39566 40462 39618 40514
rect 41022 40462 41074 40514
rect 41358 40462 41410 40514
rect 42590 40462 42642 40514
rect 50094 40462 50146 40514
rect 1710 40350 1762 40402
rect 2494 40350 2546 40402
rect 4622 40350 4674 40402
rect 7870 40350 7922 40402
rect 9550 40350 9602 40402
rect 14030 40350 14082 40402
rect 18846 40350 18898 40402
rect 19406 40350 19458 40402
rect 21198 40350 21250 40402
rect 21870 40350 21922 40402
rect 30046 40350 30098 40402
rect 30382 40350 30434 40402
rect 31278 40350 31330 40402
rect 32510 40350 32562 40402
rect 33854 40350 33906 40402
rect 37774 40350 37826 40402
rect 39902 40350 39954 40402
rect 42814 40350 42866 40402
rect 43262 40350 43314 40402
rect 43486 40350 43538 40402
rect 44382 40350 44434 40402
rect 45278 40350 45330 40402
rect 48862 40350 48914 40402
rect 49310 40350 49362 40402
rect 52782 40350 52834 40402
rect 53454 40350 53506 40402
rect 56814 40350 56866 40402
rect 57150 40350 57202 40402
rect 5294 40238 5346 40290
rect 7422 40238 7474 40290
rect 12462 40238 12514 40290
rect 12910 40238 12962 40290
rect 13470 40238 13522 40290
rect 16830 40238 16882 40290
rect 19518 40238 19570 40290
rect 24670 40238 24722 40290
rect 26238 40238 26290 40290
rect 26462 40238 26514 40290
rect 34526 40238 34578 40290
rect 36654 40238 36706 40290
rect 37438 40238 37490 40290
rect 39118 40238 39170 40290
rect 43374 40238 43426 40290
rect 43934 40238 43986 40290
rect 44830 40238 44882 40290
rect 45950 40238 46002 40290
rect 48078 40238 48130 40290
rect 52222 40238 52274 40290
rect 55582 40238 55634 40290
rect 56030 40238 56082 40290
rect 56702 40238 56754 40290
rect 7758 40126 7810 40178
rect 8318 40126 8370 40178
rect 8542 40126 8594 40178
rect 25790 40126 25842 40178
rect 31054 40126 31106 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 10334 39790 10386 39842
rect 10670 39790 10722 39842
rect 12126 39790 12178 39842
rect 32398 39790 32450 39842
rect 1934 39678 1986 39730
rect 6526 39678 6578 39730
rect 7086 39678 7138 39730
rect 9214 39678 9266 39730
rect 10894 39678 10946 39730
rect 11566 39678 11618 39730
rect 14254 39678 14306 39730
rect 16382 39678 16434 39730
rect 22094 39678 22146 39730
rect 24222 39678 24274 39730
rect 24782 39678 24834 39730
rect 29262 39678 29314 39730
rect 30606 39678 30658 39730
rect 34078 39678 34130 39730
rect 44270 39678 44322 39730
rect 44942 39678 44994 39730
rect 45726 39678 45778 39730
rect 48974 39678 49026 39730
rect 51214 39678 51266 39730
rect 51662 39678 51714 39730
rect 52782 39678 52834 39730
rect 53230 39678 53282 39730
rect 55358 39678 55410 39730
rect 4286 39566 4338 39618
rect 6078 39566 6130 39618
rect 9998 39566 10050 39618
rect 11902 39566 11954 39618
rect 12910 39566 12962 39618
rect 13582 39566 13634 39618
rect 18398 39566 18450 39618
rect 18958 39566 19010 39618
rect 21310 39566 21362 39618
rect 27694 39566 27746 39618
rect 28254 39566 28306 39618
rect 28590 39566 28642 39618
rect 32286 39566 32338 39618
rect 34526 39566 34578 39618
rect 35086 39566 35138 39618
rect 35870 39566 35922 39618
rect 37214 39566 37266 39618
rect 38446 39566 38498 39618
rect 41470 39566 41522 39618
rect 45278 39566 45330 39618
rect 45838 39566 45890 39618
rect 51550 39566 51602 39618
rect 52222 39566 52274 39618
rect 56030 39566 56082 39618
rect 5966 39454 6018 39506
rect 19070 39454 19122 39506
rect 26910 39454 26962 39506
rect 31614 39454 31666 39506
rect 31950 39454 32002 39506
rect 33966 39454 34018 39506
rect 37550 39454 37602 39506
rect 42142 39454 42194 39506
rect 5742 39342 5794 39394
rect 6414 39342 6466 39394
rect 12462 39342 12514 39394
rect 28030 39342 28082 39394
rect 28142 39342 28194 39394
rect 31390 39342 31442 39394
rect 32398 39342 32450 39394
rect 33742 39342 33794 39394
rect 34190 39342 34242 39394
rect 34862 39342 34914 39394
rect 36206 39342 36258 39394
rect 37998 39342 38050 39394
rect 38894 39342 38946 39394
rect 45614 39342 45666 39394
rect 50318 39342 50370 39394
rect 50766 39342 50818 39394
rect 51774 39342 51826 39394
rect 56590 39342 56642 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 7646 39006 7698 39058
rect 8990 39006 9042 39058
rect 10222 39006 10274 39058
rect 11118 39006 11170 39058
rect 13022 39006 13074 39058
rect 13582 39006 13634 39058
rect 14142 39006 14194 39058
rect 15598 39006 15650 39058
rect 24446 39006 24498 39058
rect 25678 39006 25730 39058
rect 25902 39006 25954 39058
rect 33182 39006 33234 39058
rect 33966 39006 34018 39058
rect 34302 39006 34354 39058
rect 34526 39006 34578 39058
rect 35758 39006 35810 39058
rect 41806 39006 41858 39058
rect 41918 39006 41970 39058
rect 43822 39006 43874 39058
rect 52222 39006 52274 39058
rect 53230 39006 53282 39058
rect 2046 38894 2098 38946
rect 4622 38894 4674 38946
rect 6414 38894 6466 38946
rect 12686 38894 12738 38946
rect 13358 38894 13410 38946
rect 15934 38894 15986 38946
rect 21422 38894 21474 38946
rect 27134 38894 27186 38946
rect 35422 38894 35474 38946
rect 35982 38894 36034 38946
rect 36654 38894 36706 38946
rect 36990 38894 37042 38946
rect 42590 38894 42642 38946
rect 42814 38894 42866 38946
rect 45502 38894 45554 38946
rect 52446 38894 52498 38946
rect 53006 38894 53058 38946
rect 56702 38894 56754 38946
rect 1710 38782 1762 38834
rect 4734 38782 4786 38834
rect 5966 38782 6018 38834
rect 6862 38782 6914 38834
rect 20862 38782 20914 38834
rect 21198 38782 21250 38834
rect 21870 38782 21922 38834
rect 22430 38782 22482 38834
rect 25230 38782 25282 38834
rect 25790 38782 25842 38834
rect 26462 38782 26514 38834
rect 29598 38770 29650 38822
rect 34190 38782 34242 38834
rect 35534 38782 35586 38834
rect 36094 38782 36146 38834
rect 36878 38782 36930 38834
rect 37438 38782 37490 38834
rect 41582 38782 41634 38834
rect 42030 38782 42082 38834
rect 42478 38782 42530 38834
rect 42926 38782 42978 38834
rect 45838 38782 45890 38834
rect 48862 38782 48914 38834
rect 52558 38782 52610 38834
rect 52894 38782 52946 38834
rect 53454 38782 53506 38834
rect 2494 38670 2546 38722
rect 5070 38670 5122 38722
rect 6750 38670 6802 38722
rect 25454 38670 25506 38722
rect 29262 38670 29314 38722
rect 30382 38670 30434 38722
rect 32510 38670 32562 38722
rect 35086 38670 35138 38722
rect 38222 38670 38274 38722
rect 40350 38670 40402 38722
rect 44158 38670 44210 38722
rect 46510 38670 46562 38722
rect 49534 38670 49586 38722
rect 51662 38670 51714 38722
rect 5182 38558 5234 38610
rect 5518 38558 5570 38610
rect 5630 38558 5682 38610
rect 5854 38558 5906 38610
rect 6526 38558 6578 38610
rect 13694 38558 13746 38610
rect 13918 38558 13970 38610
rect 14254 38558 14306 38610
rect 35422 38558 35474 38610
rect 36990 38558 37042 38610
rect 46622 38558 46674 38610
rect 55358 38558 55410 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 5854 38222 5906 38274
rect 6190 38222 6242 38274
rect 12574 38222 12626 38274
rect 36542 38222 36594 38274
rect 37326 38222 37378 38274
rect 39678 38222 39730 38274
rect 40014 38222 40066 38274
rect 10894 38110 10946 38162
rect 14814 38110 14866 38162
rect 18734 38110 18786 38162
rect 23774 38110 23826 38162
rect 29486 38110 29538 38162
rect 30270 38110 30322 38162
rect 30830 38110 30882 38162
rect 31838 38110 31890 38162
rect 37886 38110 37938 38162
rect 44158 38110 44210 38162
rect 45054 38110 45106 38162
rect 47182 38110 47234 38162
rect 51662 38110 51714 38162
rect 55918 38110 55970 38162
rect 5966 37998 6018 38050
rect 6414 37998 6466 38050
rect 8094 37998 8146 38050
rect 12014 37998 12066 38050
rect 12238 37998 12290 38050
rect 13806 37998 13858 38050
rect 14366 37998 14418 38050
rect 15262 37998 15314 38050
rect 15822 37998 15874 38050
rect 19966 37998 20018 38050
rect 21870 37998 21922 38050
rect 22318 37998 22370 38050
rect 29710 37998 29762 38050
rect 30158 37998 30210 38050
rect 32174 37998 32226 38050
rect 35646 37998 35698 38050
rect 37550 37998 37602 38050
rect 37774 37998 37826 38050
rect 37998 37998 38050 38050
rect 40238 37998 40290 38050
rect 40686 37998 40738 38050
rect 40910 37998 40962 38050
rect 41358 37998 41410 38050
rect 46622 37998 46674 38050
rect 46958 37998 47010 38050
rect 47070 37998 47122 38050
rect 47294 37998 47346 38050
rect 48750 37998 48802 38050
rect 53006 37998 53058 38050
rect 1710 37886 1762 37938
rect 2046 37886 2098 37938
rect 6526 37886 6578 37938
rect 7310 37886 7362 37938
rect 7646 37886 7698 37938
rect 8766 37886 8818 37938
rect 11342 37886 11394 37938
rect 11566 37886 11618 37938
rect 14030 37886 14082 37938
rect 15486 37886 15538 37938
rect 16606 37886 16658 37938
rect 20190 37886 20242 37938
rect 20862 37886 20914 37938
rect 34302 37886 34354 37938
rect 34974 37886 35026 37938
rect 35982 37886 36034 37938
rect 36430 37886 36482 37938
rect 40574 37886 40626 37938
rect 42030 37886 42082 37938
rect 46286 37886 46338 37938
rect 47518 37886 47570 37938
rect 49534 37886 49586 37938
rect 53790 37886 53842 37938
rect 2494 37774 2546 37826
rect 11454 37774 11506 37826
rect 14254 37774 14306 37826
rect 19630 37774 19682 37826
rect 21310 37774 21362 37826
rect 22542 37774 22594 37826
rect 23214 37774 23266 37826
rect 27806 37774 27858 37826
rect 28590 37774 28642 37826
rect 30382 37774 30434 37826
rect 32510 37774 32562 37826
rect 33182 37774 33234 37826
rect 33630 37774 33682 37826
rect 33966 37774 34018 37826
rect 34638 37774 34690 37826
rect 35310 37774 35362 37826
rect 36206 37774 36258 37826
rect 40014 37774 40066 37826
rect 40462 37774 40514 37826
rect 46398 37774 46450 37826
rect 52222 37774 52274 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 2046 37438 2098 37490
rect 6302 37438 6354 37490
rect 15374 37438 15426 37490
rect 28366 37438 28418 37490
rect 28926 37438 28978 37490
rect 29038 37438 29090 37490
rect 30382 37438 30434 37490
rect 30718 37438 30770 37490
rect 31390 37438 31442 37490
rect 33406 37438 33458 37490
rect 34414 37438 34466 37490
rect 37326 37438 37378 37490
rect 39454 37438 39506 37490
rect 40126 37438 40178 37490
rect 41358 37438 41410 37490
rect 45838 37438 45890 37490
rect 46174 37438 46226 37490
rect 50430 37438 50482 37490
rect 50878 37438 50930 37490
rect 51438 37438 51490 37490
rect 52446 37438 52498 37490
rect 6974 37326 7026 37378
rect 7310 37326 7362 37378
rect 11230 37326 11282 37378
rect 12462 37326 12514 37378
rect 14814 37326 14866 37378
rect 15934 37326 15986 37378
rect 16494 37326 16546 37378
rect 24334 37326 24386 37378
rect 25230 37326 25282 37378
rect 26910 37326 26962 37378
rect 29262 37326 29314 37378
rect 34750 37326 34802 37378
rect 37102 37326 37154 37378
rect 37438 37326 37490 37378
rect 39902 37326 39954 37378
rect 41134 37326 41186 37378
rect 42142 37326 42194 37378
rect 46286 37326 46338 37378
rect 47630 37326 47682 37378
rect 51214 37326 51266 37378
rect 52222 37326 52274 37378
rect 1710 37214 1762 37266
rect 5854 37214 5906 37266
rect 5966 37214 6018 37266
rect 6190 37214 6242 37266
rect 11566 37214 11618 37266
rect 13358 37214 13410 37266
rect 13806 37214 13858 37266
rect 14366 37214 14418 37266
rect 20974 37214 21026 37266
rect 21310 37214 21362 37266
rect 21422 37214 21474 37266
rect 21646 37214 21698 37266
rect 21870 37214 21922 37266
rect 22318 37214 22370 37266
rect 23662 37214 23714 37266
rect 25678 37214 25730 37266
rect 26686 37214 26738 37266
rect 27022 37214 27074 37266
rect 27582 37214 27634 37266
rect 27918 37214 27970 37266
rect 28030 37214 28082 37266
rect 28142 37214 28194 37266
rect 28814 37214 28866 37266
rect 36878 37214 36930 37266
rect 37774 37214 37826 37266
rect 38222 37214 38274 37266
rect 39790 37214 39842 37266
rect 40910 37214 40962 37266
rect 41806 37214 41858 37266
rect 46062 37214 46114 37266
rect 47070 37214 47122 37266
rect 48078 37214 48130 37266
rect 48862 37214 48914 37266
rect 51550 37214 51602 37266
rect 51662 37214 51714 37266
rect 51774 37214 51826 37266
rect 52670 37214 52722 37266
rect 52782 37214 52834 37266
rect 56030 37214 56082 37266
rect 2494 37102 2546 37154
rect 2942 37102 2994 37154
rect 12574 37102 12626 37154
rect 12910 37102 12962 37154
rect 17502 37102 17554 37154
rect 18062 37102 18114 37154
rect 20190 37102 20242 37154
rect 23998 37102 24050 37154
rect 25566 37102 25618 37154
rect 31838 37102 31890 37154
rect 33854 37102 33906 37154
rect 35310 37102 35362 37154
rect 35758 37102 35810 37154
rect 36094 37102 36146 37154
rect 36542 37102 36594 37154
rect 39342 37102 39394 37154
rect 41022 37102 41074 37154
rect 45390 37102 45442 37154
rect 46846 37102 46898 37154
rect 52558 37102 52610 37154
rect 6414 36990 6466 37042
rect 12238 36990 12290 37042
rect 15710 36990 15762 37042
rect 36094 36990 36146 37042
rect 36430 36990 36482 37042
rect 36766 36990 36818 37042
rect 55022 36990 55074 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 23102 36654 23154 36706
rect 23550 36654 23602 36706
rect 25566 36654 25618 36706
rect 51326 36654 51378 36706
rect 8430 36542 8482 36594
rect 10558 36542 10610 36594
rect 17838 36542 17890 36594
rect 20078 36542 20130 36594
rect 20638 36542 20690 36594
rect 21422 36542 21474 36594
rect 24782 36542 24834 36594
rect 26238 36542 26290 36594
rect 28478 36542 28530 36594
rect 30942 36542 30994 36594
rect 32734 36542 32786 36594
rect 35086 36542 35138 36594
rect 37102 36542 37154 36594
rect 39790 36542 39842 36594
rect 42590 36542 42642 36594
rect 47070 36542 47122 36594
rect 47854 36542 47906 36594
rect 49534 36542 49586 36594
rect 49982 36542 50034 36594
rect 50430 36542 50482 36594
rect 52782 36542 52834 36594
rect 54462 36542 54514 36594
rect 56590 36542 56642 36594
rect 7758 36430 7810 36482
rect 11790 36430 11842 36482
rect 12686 36430 12738 36482
rect 13806 36430 13858 36482
rect 16718 36430 16770 36482
rect 17166 36430 17218 36482
rect 19518 36430 19570 36482
rect 19966 36430 20018 36482
rect 20190 36430 20242 36482
rect 22206 36430 22258 36482
rect 23102 36430 23154 36482
rect 23774 36430 23826 36482
rect 24334 36430 24386 36482
rect 26462 36430 26514 36482
rect 26798 36430 26850 36482
rect 28702 36430 28754 36482
rect 30382 36430 30434 36482
rect 30830 36430 30882 36482
rect 33294 36430 33346 36482
rect 34638 36430 34690 36482
rect 34750 36430 34802 36482
rect 36094 36430 36146 36482
rect 39118 36430 39170 36482
rect 39566 36430 39618 36482
rect 40238 36430 40290 36482
rect 41694 36430 41746 36482
rect 42254 36430 42306 36482
rect 42702 36430 42754 36482
rect 42814 36430 42866 36482
rect 45278 36430 45330 36482
rect 45502 36430 45554 36482
rect 45726 36430 45778 36482
rect 47518 36430 47570 36482
rect 47742 36430 47794 36482
rect 50654 36430 50706 36482
rect 50990 36430 51042 36482
rect 51438 36430 51490 36482
rect 53118 36430 53170 36482
rect 53790 36430 53842 36482
rect 1710 36318 1762 36370
rect 2382 36318 2434 36370
rect 2718 36318 2770 36370
rect 3166 36318 3218 36370
rect 12910 36318 12962 36370
rect 16382 36318 16434 36370
rect 17390 36318 17442 36370
rect 22654 36318 22706 36370
rect 22990 36318 23042 36370
rect 25454 36318 25506 36370
rect 27806 36318 27858 36370
rect 28030 36318 28082 36370
rect 28254 36318 28306 36370
rect 30046 36318 30098 36370
rect 33070 36318 33122 36370
rect 33966 36318 34018 36370
rect 34078 36318 34130 36370
rect 34302 36318 34354 36370
rect 35534 36318 35586 36370
rect 35870 36318 35922 36370
rect 41918 36318 41970 36370
rect 46734 36318 46786 36370
rect 48526 36318 48578 36370
rect 48862 36318 48914 36370
rect 49086 36318 49138 36370
rect 51886 36318 51938 36370
rect 52110 36318 52162 36370
rect 52670 36318 52722 36370
rect 53006 36318 53058 36370
rect 2046 36206 2098 36258
rect 11006 36206 11058 36258
rect 12238 36206 12290 36258
rect 13470 36206 13522 36258
rect 16046 36206 16098 36258
rect 19742 36206 19794 36258
rect 25566 36206 25618 36258
rect 29710 36206 29762 36258
rect 30270 36206 30322 36258
rect 30494 36206 30546 36258
rect 31054 36206 31106 36258
rect 31278 36206 31330 36258
rect 31838 36206 31890 36258
rect 34974 36206 35026 36258
rect 35086 36206 35138 36258
rect 35646 36206 35698 36258
rect 40126 36206 40178 36258
rect 40350 36206 40402 36258
rect 40574 36206 40626 36258
rect 41134 36206 41186 36258
rect 42478 36206 42530 36258
rect 43486 36206 43538 36258
rect 44942 36206 44994 36258
rect 46174 36206 46226 36258
rect 46958 36206 47010 36258
rect 47182 36206 47234 36258
rect 47966 36206 48018 36258
rect 48078 36206 48130 36258
rect 48638 36206 48690 36258
rect 51214 36206 51266 36258
rect 51774 36206 51826 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 13470 35870 13522 35922
rect 15598 35870 15650 35922
rect 18510 35870 18562 35922
rect 18734 35870 18786 35922
rect 23326 35870 23378 35922
rect 23774 35870 23826 35922
rect 24110 35870 24162 35922
rect 24670 35870 24722 35922
rect 26686 35870 26738 35922
rect 28702 35870 28754 35922
rect 30830 35870 30882 35922
rect 32174 35870 32226 35922
rect 34526 35870 34578 35922
rect 39678 35870 39730 35922
rect 39902 35870 39954 35922
rect 40238 35870 40290 35922
rect 41246 35870 41298 35922
rect 41918 35870 41970 35922
rect 51326 35870 51378 35922
rect 51662 35870 51714 35922
rect 52222 35870 52274 35922
rect 52670 35870 52722 35922
rect 5854 35758 5906 35810
rect 19070 35758 19122 35810
rect 25230 35758 25282 35810
rect 27246 35758 27298 35810
rect 30270 35758 30322 35810
rect 30606 35758 30658 35810
rect 31166 35758 31218 35810
rect 31614 35758 31666 35810
rect 33070 35758 33122 35810
rect 33406 35758 33458 35810
rect 34414 35758 34466 35810
rect 35534 35758 35586 35810
rect 41470 35758 41522 35810
rect 42254 35758 42306 35810
rect 43374 35758 43426 35810
rect 47854 35758 47906 35810
rect 47966 35758 48018 35810
rect 48750 35758 48802 35810
rect 50094 35758 50146 35810
rect 51550 35758 51602 35810
rect 52894 35758 52946 35810
rect 4286 35646 4338 35698
rect 5182 35646 5234 35698
rect 9550 35646 9602 35698
rect 14142 35646 14194 35698
rect 14366 35646 14418 35698
rect 14590 35646 14642 35698
rect 23662 35646 23714 35698
rect 23886 35646 23938 35698
rect 25902 35646 25954 35698
rect 26126 35646 26178 35698
rect 26462 35646 26514 35698
rect 26798 35646 26850 35698
rect 27918 35646 27970 35698
rect 28142 35646 28194 35698
rect 28478 35646 28530 35698
rect 28814 35646 28866 35698
rect 29822 35646 29874 35698
rect 30046 35646 30098 35698
rect 30830 35646 30882 35698
rect 32510 35646 32562 35698
rect 33966 35646 34018 35698
rect 34190 35646 34242 35698
rect 34862 35646 34914 35698
rect 39566 35646 39618 35698
rect 41134 35646 41186 35698
rect 41582 35646 41634 35698
rect 42030 35646 42082 35698
rect 42702 35646 42754 35698
rect 47182 35646 47234 35698
rect 48862 35646 48914 35698
rect 49198 35646 49250 35698
rect 50318 35646 50370 35698
rect 50990 35646 51042 35698
rect 51774 35646 51826 35698
rect 52446 35646 52498 35698
rect 53006 35646 53058 35698
rect 53454 35646 53506 35698
rect 7982 35534 8034 35586
rect 8430 35534 8482 35586
rect 10334 35534 10386 35586
rect 12462 35534 12514 35586
rect 12910 35534 12962 35586
rect 14254 35534 14306 35586
rect 15150 35534 15202 35586
rect 16158 35534 16210 35586
rect 37662 35534 37714 35586
rect 38110 35534 38162 35586
rect 45502 35534 45554 35586
rect 45950 35534 46002 35586
rect 46398 35534 46450 35586
rect 46734 35534 46786 35586
rect 52334 35534 52386 35586
rect 1934 35422 1986 35474
rect 16046 35422 16098 35474
rect 45726 35422 45778 35474
rect 46398 35422 46450 35474
rect 46958 35422 47010 35474
rect 47630 35422 47682 35474
rect 47966 35422 48018 35474
rect 55358 35422 55410 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 10894 35086 10946 35138
rect 22990 35086 23042 35138
rect 23438 35086 23490 35138
rect 26798 35086 26850 35138
rect 29038 35086 29090 35138
rect 41806 35086 41858 35138
rect 11006 34974 11058 35026
rect 15822 34974 15874 35026
rect 17950 34974 18002 35026
rect 25118 34974 25170 35026
rect 29934 34974 29986 35026
rect 30382 34974 30434 35026
rect 30942 34974 30994 35026
rect 15150 34862 15202 34914
rect 22206 34862 22258 34914
rect 23214 34862 23266 34914
rect 24110 34862 24162 34914
rect 26462 34862 26514 34914
rect 28142 34862 28194 34914
rect 29486 34862 29538 34914
rect 29710 34862 29762 34914
rect 32958 34974 33010 35026
rect 33630 34974 33682 35026
rect 36094 34974 36146 35026
rect 37102 34974 37154 35026
rect 39678 34974 39730 35026
rect 40910 34974 40962 35026
rect 44942 34974 44994 35026
rect 48190 34974 48242 35026
rect 52670 34974 52722 35026
rect 54126 34974 54178 35026
rect 57934 34974 57986 35026
rect 30942 34862 30994 34914
rect 31166 34862 31218 34914
rect 31726 34862 31778 34914
rect 32062 34862 32114 34914
rect 32286 34862 32338 34914
rect 34638 34862 34690 34914
rect 35198 34862 35250 34914
rect 35646 34862 35698 34914
rect 39230 34862 39282 34914
rect 39454 34862 39506 34914
rect 40126 34862 40178 34914
rect 41134 34862 41186 34914
rect 41470 34862 41522 34914
rect 42254 34862 42306 34914
rect 42702 34862 42754 34914
rect 42926 34862 42978 34914
rect 43486 34862 43538 34914
rect 46958 34862 47010 34914
rect 50654 34862 50706 34914
rect 50990 34862 51042 34914
rect 51326 34862 51378 34914
rect 51662 34862 51714 34914
rect 51774 34862 51826 34914
rect 52110 34862 52162 34914
rect 52782 34862 52834 34914
rect 53342 34862 53394 34914
rect 55582 34862 55634 34914
rect 5854 34750 5906 34802
rect 14254 34750 14306 34802
rect 21646 34750 21698 34802
rect 22766 34750 22818 34802
rect 23886 34750 23938 34802
rect 26238 34750 26290 34802
rect 31390 34750 31442 34802
rect 31502 34750 31554 34802
rect 38558 34750 38610 34802
rect 49982 34750 50034 34802
rect 5518 34638 5570 34690
rect 5742 34638 5794 34690
rect 14142 34638 14194 34690
rect 14702 34638 14754 34690
rect 21310 34638 21362 34690
rect 22430 34638 22482 34690
rect 24446 34638 24498 34690
rect 25902 34638 25954 34690
rect 27246 34638 27298 34690
rect 27694 34638 27746 34690
rect 30270 34638 30322 34690
rect 30494 34638 30546 34690
rect 34302 34638 34354 34690
rect 34526 34638 34578 34690
rect 34750 34638 34802 34690
rect 37662 34638 37714 34690
rect 38222 34638 38274 34690
rect 38782 34638 38834 34690
rect 40350 34638 40402 34690
rect 41694 34638 41746 34690
rect 42030 34638 42082 34690
rect 42142 34638 42194 34690
rect 44046 34638 44098 34690
rect 45950 34638 46002 34690
rect 46286 34638 46338 34690
rect 46622 34638 46674 34690
rect 49870 34638 49922 34690
rect 50542 34638 50594 34690
rect 51102 34638 51154 34690
rect 51550 34638 51602 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 7982 34302 8034 34354
rect 12238 34302 12290 34354
rect 16270 34302 16322 34354
rect 16494 34302 16546 34354
rect 18398 34302 18450 34354
rect 22878 34302 22930 34354
rect 24782 34302 24834 34354
rect 25230 34302 25282 34354
rect 31166 34302 31218 34354
rect 37102 34302 37154 34354
rect 43262 34302 43314 34354
rect 46958 34302 47010 34354
rect 48078 34302 48130 34354
rect 48302 34302 48354 34354
rect 48862 34302 48914 34354
rect 50206 34302 50258 34354
rect 51326 34302 51378 34354
rect 8542 34190 8594 34242
rect 10558 34190 10610 34242
rect 13358 34190 13410 34242
rect 16158 34190 16210 34242
rect 20190 34190 20242 34242
rect 23550 34190 23602 34242
rect 23774 34190 23826 34242
rect 25566 34190 25618 34242
rect 29934 34190 29986 34242
rect 38222 34190 38274 34242
rect 42590 34190 42642 34242
rect 45390 34190 45442 34242
rect 45838 34190 45890 34242
rect 47182 34190 47234 34242
rect 47630 34190 47682 34242
rect 47966 34190 48018 34242
rect 48750 34190 48802 34242
rect 52782 34190 52834 34242
rect 4286 34078 4338 34130
rect 4734 34078 4786 34130
rect 8318 34078 8370 34130
rect 8654 34078 8706 34130
rect 10222 34078 10274 34130
rect 12686 34078 12738 34130
rect 15934 34078 15986 34130
rect 16382 34078 16434 34130
rect 18286 34078 18338 34130
rect 18622 34078 18674 34130
rect 18846 34078 18898 34130
rect 19518 34078 19570 34130
rect 29598 34078 29650 34130
rect 35534 34078 35586 34130
rect 35982 34078 36034 34130
rect 36206 34078 36258 34130
rect 37550 34078 37602 34130
rect 42030 34078 42082 34130
rect 43038 34078 43090 34130
rect 47406 34078 47458 34130
rect 48974 34078 49026 34130
rect 49422 34078 49474 34130
rect 50654 34078 50706 34130
rect 50878 34078 50930 34130
rect 51998 34078 52050 34130
rect 52894 34078 52946 34130
rect 53230 34078 53282 34130
rect 1822 33966 1874 34018
rect 5406 33966 5458 34018
rect 7534 33966 7586 34018
rect 11006 33966 11058 34018
rect 15486 33966 15538 34018
rect 17726 33966 17778 34018
rect 18510 33966 18562 34018
rect 22318 33966 22370 34018
rect 26462 33966 26514 34018
rect 31614 33966 31666 34018
rect 33742 33966 33794 34018
rect 34190 33966 34242 34018
rect 34750 33966 34802 34018
rect 36094 33966 36146 34018
rect 36542 33966 36594 34018
rect 40350 33966 40402 34018
rect 42142 33966 42194 34018
rect 43710 33966 43762 34018
rect 47518 33966 47570 34018
rect 49870 33966 49922 34018
rect 51102 33966 51154 34018
rect 52222 33966 52274 34018
rect 17838 33854 17890 33906
rect 23214 33854 23266 33906
rect 34974 33854 35026 33906
rect 35310 33854 35362 33906
rect 36766 33854 36818 33906
rect 44830 33854 44882 33906
rect 45166 33854 45218 33906
rect 51774 33854 51826 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 5518 33518 5570 33570
rect 5854 33518 5906 33570
rect 34302 33518 34354 33570
rect 38558 33518 38610 33570
rect 42702 33518 42754 33570
rect 43038 33518 43090 33570
rect 52782 33518 52834 33570
rect 57934 33518 57986 33570
rect 4734 33406 4786 33458
rect 6190 33406 6242 33458
rect 10446 33406 10498 33458
rect 10894 33406 10946 33458
rect 15486 33406 15538 33458
rect 15934 33406 15986 33458
rect 16606 33406 16658 33458
rect 18174 33406 18226 33458
rect 20302 33406 20354 33458
rect 24110 33406 24162 33458
rect 27806 33406 27858 33458
rect 29150 33406 29202 33458
rect 34862 33406 34914 33458
rect 35758 33406 35810 33458
rect 37662 33406 37714 33458
rect 42702 33406 42754 33458
rect 47742 33406 47794 33458
rect 50990 33406 51042 33458
rect 51438 33406 51490 33458
rect 1934 33294 1986 33346
rect 6638 33294 6690 33346
rect 6862 33294 6914 33346
rect 7198 33294 7250 33346
rect 7646 33294 7698 33346
rect 11566 33294 11618 33346
rect 12350 33294 12402 33346
rect 12910 33294 12962 33346
rect 15374 33294 15426 33346
rect 17054 33294 17106 33346
rect 17390 33294 17442 33346
rect 21870 33294 21922 33346
rect 22318 33294 22370 33346
rect 22990 33294 23042 33346
rect 24894 33294 24946 33346
rect 32062 33294 32114 33346
rect 35310 33294 35362 33346
rect 38894 33294 38946 33346
rect 39454 33294 39506 33346
rect 43038 33294 43090 33346
rect 44046 33294 44098 33346
rect 44942 33294 44994 33346
rect 48190 33294 48242 33346
rect 52670 33294 52722 33346
rect 55582 33294 55634 33346
rect 2606 33182 2658 33234
rect 8318 33182 8370 33234
rect 14254 33182 14306 33234
rect 14926 33182 14978 33234
rect 15486 33182 15538 33234
rect 22542 33182 22594 33234
rect 24446 33182 24498 33234
rect 24558 33182 24610 33234
rect 25678 33182 25730 33234
rect 28478 33182 28530 33234
rect 28590 33182 28642 33234
rect 31278 33182 31330 33234
rect 32510 33182 32562 33234
rect 34414 33182 34466 33234
rect 36094 33182 36146 33234
rect 36430 33182 36482 33234
rect 39678 33182 39730 33234
rect 44270 33182 44322 33234
rect 45614 33182 45666 33234
rect 48862 33182 48914 33234
rect 51326 33182 51378 33234
rect 54462 33182 54514 33234
rect 5854 33070 5906 33122
rect 6078 33070 6130 33122
rect 6302 33070 6354 33122
rect 7086 33070 7138 33122
rect 11678 33070 11730 33122
rect 11902 33070 11954 33122
rect 13470 33070 13522 33122
rect 13806 33070 13858 33122
rect 15150 33070 15202 33122
rect 16046 33070 16098 33122
rect 32398 33070 32450 33122
rect 32958 33070 33010 33122
rect 33854 33070 33906 33122
rect 34302 33070 34354 33122
rect 37102 33070 37154 33122
rect 37998 33070 38050 33122
rect 51886 33070 51938 33122
rect 53230 33070 53282 33122
rect 54574 33070 54626 33122
rect 55358 33070 55410 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 8094 32734 8146 32786
rect 8430 32734 8482 32786
rect 14366 32734 14418 32786
rect 15822 32734 15874 32786
rect 16494 32734 16546 32786
rect 16830 32734 16882 32786
rect 20862 32734 20914 32786
rect 25566 32734 25618 32786
rect 25678 32734 25730 32786
rect 29822 32734 29874 32786
rect 31726 32734 31778 32786
rect 38894 32734 38946 32786
rect 39342 32734 39394 32786
rect 50542 32734 50594 32786
rect 52558 32734 52610 32786
rect 5406 32622 5458 32674
rect 6862 32622 6914 32674
rect 9774 32622 9826 32674
rect 15710 32622 15762 32674
rect 25230 32622 25282 32674
rect 26462 32622 26514 32674
rect 29486 32622 29538 32674
rect 30046 32622 30098 32674
rect 51774 32622 51826 32674
rect 55246 32622 55298 32674
rect 1822 32510 1874 32562
rect 5294 32510 5346 32562
rect 6974 32510 7026 32562
rect 8318 32510 8370 32562
rect 8542 32510 8594 32562
rect 9550 32510 9602 32562
rect 9998 32510 10050 32562
rect 10222 32510 10274 32562
rect 10558 32510 10610 32562
rect 14702 32510 14754 32562
rect 15038 32510 15090 32562
rect 15374 32510 15426 32562
rect 19742 32510 19794 32562
rect 21086 32510 21138 32562
rect 25454 32510 25506 32562
rect 25902 32510 25954 32562
rect 26798 32510 26850 32562
rect 29710 32510 29762 32562
rect 29934 32510 29986 32562
rect 31390 32510 31442 32562
rect 31614 32510 31666 32562
rect 31838 32510 31890 32562
rect 31950 32510 32002 32562
rect 34750 32510 34802 32562
rect 35310 32510 35362 32562
rect 35982 32510 36034 32562
rect 36206 32510 36258 32562
rect 38782 32510 38834 32562
rect 41694 32510 41746 32562
rect 45054 32510 45106 32562
rect 47966 32510 48018 32562
rect 51886 32510 51938 32562
rect 52222 32510 52274 32562
rect 55918 32510 55970 32562
rect 2494 32398 2546 32450
rect 4622 32398 4674 32450
rect 5854 32398 5906 32450
rect 7646 32398 7698 32450
rect 9102 32398 9154 32450
rect 11230 32398 11282 32450
rect 13358 32398 13410 32450
rect 13918 32398 13970 32450
rect 14926 32398 14978 32450
rect 27246 32398 27298 32450
rect 29150 32398 29202 32450
rect 31054 32398 31106 32450
rect 33966 32398 34018 32450
rect 36766 32398 36818 32450
rect 37214 32398 37266 32450
rect 39454 32398 39506 32450
rect 42478 32398 42530 32450
rect 44606 32398 44658 32450
rect 53118 32398 53170 32450
rect 14142 32286 14194 32338
rect 14478 32286 14530 32338
rect 15822 32286 15874 32338
rect 19742 32286 19794 32338
rect 20078 32286 20130 32338
rect 34638 32286 34690 32338
rect 35086 32286 35138 32338
rect 38894 32286 38946 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 15150 31950 15202 32002
rect 42142 31950 42194 32002
rect 51886 31950 51938 32002
rect 2830 31838 2882 31890
rect 6078 31838 6130 31890
rect 7646 31838 7698 31890
rect 8878 31838 8930 31890
rect 9438 31838 9490 31890
rect 11230 31838 11282 31890
rect 12910 31838 12962 31890
rect 15822 31838 15874 31890
rect 22542 31838 22594 31890
rect 23998 31838 24050 31890
rect 25454 31838 25506 31890
rect 26462 31838 26514 31890
rect 28590 31838 28642 31890
rect 29710 31838 29762 31890
rect 39006 31838 39058 31890
rect 40686 31838 40738 31890
rect 41582 31838 41634 31890
rect 42030 31838 42082 31890
rect 43598 31838 43650 31890
rect 50318 31838 50370 31890
rect 51550 31838 51602 31890
rect 54350 31838 54402 31890
rect 1710 31726 1762 31778
rect 4622 31726 4674 31778
rect 4846 31726 4898 31778
rect 6190 31726 6242 31778
rect 6526 31726 6578 31778
rect 8542 31726 8594 31778
rect 11678 31726 11730 31778
rect 14142 31726 14194 31778
rect 14590 31726 14642 31778
rect 15598 31726 15650 31778
rect 16270 31726 16322 31778
rect 19182 31726 19234 31778
rect 19630 31726 19682 31778
rect 19854 31726 19906 31778
rect 22654 31726 22706 31778
rect 23214 31726 23266 31778
rect 24222 31726 24274 31778
rect 25678 31726 25730 31778
rect 29486 31726 29538 31778
rect 30158 31726 30210 31778
rect 38558 31726 38610 31778
rect 39902 31726 39954 31778
rect 41246 31726 41298 31778
rect 41470 31726 41522 31778
rect 47518 31726 47570 31778
rect 50878 31726 50930 31778
rect 52558 31726 52610 31778
rect 53230 31726 53282 31778
rect 53790 31726 53842 31778
rect 55022 31726 55074 31778
rect 2942 31614 2994 31666
rect 3614 31614 3666 31666
rect 3838 31614 3890 31666
rect 4062 31614 4114 31666
rect 4510 31614 4562 31666
rect 5070 31614 5122 31666
rect 5966 31614 6018 31666
rect 7758 31614 7810 31666
rect 8094 31614 8146 31666
rect 9774 31614 9826 31666
rect 10110 31614 10162 31666
rect 10334 31614 10386 31666
rect 11342 31614 11394 31666
rect 14702 31614 14754 31666
rect 15038 31614 15090 31666
rect 15262 31614 15314 31666
rect 16606 31614 16658 31666
rect 16830 31614 16882 31666
rect 17054 31614 17106 31666
rect 17390 31614 17442 31666
rect 18622 31614 18674 31666
rect 18734 31614 18786 31666
rect 18958 31614 19010 31666
rect 20526 31614 20578 31666
rect 22990 31614 23042 31666
rect 23550 31614 23602 31666
rect 23886 31614 23938 31666
rect 24782 31614 24834 31666
rect 32174 31614 32226 31666
rect 38110 31614 38162 31666
rect 39678 31614 39730 31666
rect 41022 31614 41074 31666
rect 48190 31614 48242 31666
rect 52110 31614 52162 31666
rect 2046 31502 2098 31554
rect 2718 31502 2770 31554
rect 3166 31502 3218 31554
rect 3726 31502 3778 31554
rect 7198 31502 7250 31554
rect 7534 31502 7586 31554
rect 9550 31502 9602 31554
rect 10222 31502 10274 31554
rect 11118 31502 11170 31554
rect 12126 31502 12178 31554
rect 16382 31502 16434 31554
rect 17166 31502 17218 31554
rect 17726 31502 17778 31554
rect 18062 31502 18114 31554
rect 23214 31502 23266 31554
rect 24446 31502 24498 31554
rect 24670 31502 24722 31554
rect 29822 31502 29874 31554
rect 36206 31502 36258 31554
rect 41582 31502 41634 31554
rect 42702 31502 42754 31554
rect 43150 31502 43202 31554
rect 44158 31502 44210 31554
rect 50990 31502 51042 31554
rect 53006 31502 53058 31554
rect 53118 31502 53170 31554
rect 54014 31502 54066 31554
rect 54238 31502 54290 31554
rect 54350 31502 54402 31554
rect 54798 31502 54850 31554
rect 55694 31502 55746 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 4734 31166 4786 31218
rect 4958 31166 5010 31218
rect 5630 31166 5682 31218
rect 5966 31166 6018 31218
rect 12574 31166 12626 31218
rect 14926 31166 14978 31218
rect 18846 31166 18898 31218
rect 19406 31166 19458 31218
rect 19966 31166 20018 31218
rect 20302 31166 20354 31218
rect 21534 31166 21586 31218
rect 25454 31166 25506 31218
rect 26798 31166 26850 31218
rect 34302 31166 34354 31218
rect 34974 31166 35026 31218
rect 49422 31166 49474 31218
rect 54910 31166 54962 31218
rect 56702 31166 56754 31218
rect 2046 31054 2098 31106
rect 2718 31054 2770 31106
rect 3390 31054 3442 31106
rect 4510 31054 4562 31106
rect 8990 31054 9042 31106
rect 9550 31054 9602 31106
rect 16494 31054 16546 31106
rect 18734 31054 18786 31106
rect 19518 31054 19570 31106
rect 22206 31054 22258 31106
rect 25230 31054 25282 31106
rect 27806 31054 27858 31106
rect 29710 31054 29762 31106
rect 31726 31054 31778 31106
rect 33182 31054 33234 31106
rect 36654 31054 36706 31106
rect 39342 31054 39394 31106
rect 39678 31054 39730 31106
rect 44606 31054 44658 31106
rect 45726 31054 45778 31106
rect 54350 31054 54402 31106
rect 1822 30942 1874 30994
rect 2382 30942 2434 30994
rect 3054 30942 3106 30994
rect 4174 30942 4226 30994
rect 5070 30942 5122 30994
rect 8430 30942 8482 30994
rect 9998 30942 10050 30994
rect 11342 30942 11394 30994
rect 11902 30942 11954 30994
rect 12238 30942 12290 30994
rect 12462 30942 12514 30994
rect 12798 30942 12850 30994
rect 16046 30942 16098 30994
rect 17726 30942 17778 30994
rect 19854 30942 19906 30994
rect 20078 30942 20130 30994
rect 21870 30942 21922 30994
rect 22990 30942 23042 30994
rect 23774 30942 23826 30994
rect 24222 30942 24274 30994
rect 24446 30942 24498 30994
rect 27918 30942 27970 30994
rect 29486 30942 29538 30994
rect 29822 30942 29874 30994
rect 30718 30942 30770 30994
rect 31502 30942 31554 30994
rect 31838 30942 31890 30994
rect 31950 30942 32002 30994
rect 32174 30942 32226 30994
rect 33518 30942 33570 30994
rect 34190 30942 34242 30994
rect 35422 30942 35474 30994
rect 38110 30942 38162 30994
rect 43822 30942 43874 30994
rect 44382 30942 44434 30994
rect 45054 30942 45106 30994
rect 49758 30942 49810 30994
rect 53006 30942 53058 30994
rect 53678 30942 53730 30994
rect 54574 30942 54626 30994
rect 54686 30942 54738 30994
rect 54798 30942 54850 30994
rect 55582 30942 55634 30994
rect 3838 30830 3890 30882
rect 6414 30830 6466 30882
rect 8206 30830 8258 30882
rect 9886 30830 9938 30882
rect 11118 30830 11170 30882
rect 13246 30830 13298 30882
rect 15598 30830 15650 30882
rect 17502 30830 17554 30882
rect 18398 30830 18450 30882
rect 22542 30830 22594 30882
rect 23326 30830 23378 30882
rect 24334 30830 24386 30882
rect 25342 30830 25394 30882
rect 30382 30830 30434 30882
rect 31166 30830 31218 30882
rect 33854 30830 33906 30882
rect 35870 30830 35922 30882
rect 37214 30830 37266 30882
rect 37662 30830 37714 30882
rect 38558 30830 38610 30882
rect 40910 30803 40962 30855
rect 43038 30830 43090 30882
rect 47854 30830 47906 30882
rect 48862 30830 48914 30882
rect 51998 30830 52050 30882
rect 53118 30830 53170 30882
rect 11566 30718 11618 30770
rect 18846 30718 18898 30770
rect 27134 30718 27186 30770
rect 33070 30718 33122 30770
rect 33518 30718 33570 30770
rect 34302 30718 34354 30770
rect 35646 30718 35698 30770
rect 36542 30718 36594 30770
rect 39902 30718 39954 30770
rect 40238 30718 40290 30770
rect 53006 30718 53058 30770
rect 55694 30718 55746 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 8878 30382 8930 30434
rect 9102 30382 9154 30434
rect 9326 30382 9378 30434
rect 10782 30382 10834 30434
rect 11006 30382 11058 30434
rect 18734 30382 18786 30434
rect 22430 30382 22482 30434
rect 22878 30382 22930 30434
rect 37102 30382 37154 30434
rect 39678 30382 39730 30434
rect 44942 30382 44994 30434
rect 4622 30270 4674 30322
rect 10222 30270 10274 30322
rect 16158 30270 16210 30322
rect 17054 30270 17106 30322
rect 18958 30270 19010 30322
rect 23102 30270 23154 30322
rect 23550 30270 23602 30322
rect 23774 30270 23826 30322
rect 24110 30270 24162 30322
rect 30158 30270 30210 30322
rect 34414 30270 34466 30322
rect 37214 30270 37266 30322
rect 39342 30270 39394 30322
rect 44046 30270 44098 30322
rect 49086 30270 49138 30322
rect 49646 30270 49698 30322
rect 56030 30270 56082 30322
rect 58158 30270 58210 30322
rect 1822 30158 1874 30210
rect 5518 30158 5570 30210
rect 5742 30158 5794 30210
rect 6078 30158 6130 30210
rect 7982 30158 8034 30210
rect 8654 30158 8706 30210
rect 10558 30158 10610 30210
rect 16942 30158 16994 30210
rect 17166 30158 17218 30210
rect 17838 30158 17890 30210
rect 18062 30158 18114 30210
rect 22542 30158 22594 30210
rect 27134 30158 27186 30210
rect 30046 30158 30098 30210
rect 30830 30158 30882 30210
rect 31614 30158 31666 30210
rect 32286 30158 32338 30210
rect 34862 30158 34914 30210
rect 35870 30158 35922 30210
rect 37438 30158 37490 30210
rect 37886 30158 37938 30210
rect 38222 30158 38274 30210
rect 38670 30158 38722 30210
rect 39006 30158 39058 30210
rect 40126 30158 40178 30210
rect 40686 30158 40738 30210
rect 45278 30158 45330 30210
rect 48750 30158 48802 30210
rect 50094 30158 50146 30210
rect 51550 30158 51602 30210
rect 52670 30158 52722 30210
rect 53230 30158 53282 30210
rect 53566 30158 53618 30210
rect 54462 30158 54514 30210
rect 54910 30158 54962 30210
rect 55246 30158 55298 30210
rect 2494 30046 2546 30098
rect 5966 30046 6018 30098
rect 10446 30046 10498 30098
rect 11678 30046 11730 30098
rect 13806 30046 13858 30098
rect 16270 30046 16322 30098
rect 16606 30046 16658 30098
rect 21646 30046 21698 30098
rect 22430 30046 22482 30098
rect 23102 30046 23154 30098
rect 30270 30046 30322 30098
rect 30382 30046 30434 30098
rect 35422 30046 35474 30098
rect 36318 30046 36370 30098
rect 36430 30046 36482 30098
rect 38446 30046 38498 30098
rect 41022 30046 41074 30098
rect 45502 30046 45554 30098
rect 46062 30046 46114 30098
rect 48190 30046 48242 30098
rect 50542 30046 50594 30098
rect 51998 30046 52050 30098
rect 53006 30046 53058 30098
rect 53342 30046 53394 30098
rect 54126 30046 54178 30098
rect 5070 29934 5122 29986
rect 8318 29934 8370 29986
rect 9774 29934 9826 29986
rect 12014 29934 12066 29986
rect 12574 29934 12626 29986
rect 13470 29934 13522 29986
rect 17614 29934 17666 29986
rect 17950 29934 18002 29986
rect 18398 29934 18450 29986
rect 19518 29934 19570 29986
rect 21310 29934 21362 29986
rect 23998 29934 24050 29986
rect 24222 29934 24274 29986
rect 24894 29934 24946 29986
rect 27358 29934 27410 29986
rect 34862 29934 34914 29986
rect 36094 29934 36146 29986
rect 37998 29934 38050 29986
rect 38558 29934 38610 29986
rect 39454 29934 39506 29986
rect 40014 29934 40066 29986
rect 51438 29934 51490 29986
rect 52782 29934 52834 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 2046 29598 2098 29650
rect 3166 29598 3218 29650
rect 3614 29598 3666 29650
rect 3726 29598 3778 29650
rect 6078 29598 6130 29650
rect 7982 29598 8034 29650
rect 8654 29598 8706 29650
rect 8878 29598 8930 29650
rect 9998 29598 10050 29650
rect 10110 29598 10162 29650
rect 17502 29598 17554 29650
rect 22430 29598 22482 29650
rect 25342 29598 25394 29650
rect 34078 29598 34130 29650
rect 34302 29598 34354 29650
rect 37438 29598 37490 29650
rect 39006 29598 39058 29650
rect 39230 29598 39282 29650
rect 45278 29598 45330 29650
rect 45950 29598 46002 29650
rect 47966 29598 48018 29650
rect 50990 29598 51042 29650
rect 52446 29598 52498 29650
rect 52558 29598 52610 29650
rect 53118 29598 53170 29650
rect 54014 29598 54066 29650
rect 54238 29598 54290 29650
rect 55806 29598 55858 29650
rect 57150 29598 57202 29650
rect 58158 29598 58210 29650
rect 2718 29486 2770 29538
rect 4286 29486 4338 29538
rect 4510 29486 4562 29538
rect 5966 29486 6018 29538
rect 9662 29486 9714 29538
rect 13022 29486 13074 29538
rect 18062 29486 18114 29538
rect 18622 29486 18674 29538
rect 21198 29486 21250 29538
rect 23326 29486 23378 29538
rect 27358 29486 27410 29538
rect 33294 29486 33346 29538
rect 35086 29486 35138 29538
rect 35422 29486 35474 29538
rect 35646 29486 35698 29538
rect 36542 29486 36594 29538
rect 38110 29486 38162 29538
rect 43262 29486 43314 29538
rect 43710 29486 43762 29538
rect 44382 29486 44434 29538
rect 47182 29486 47234 29538
rect 47854 29486 47906 29538
rect 51214 29486 51266 29538
rect 53790 29486 53842 29538
rect 54686 29486 54738 29538
rect 55134 29486 55186 29538
rect 55246 29486 55298 29538
rect 55582 29486 55634 29538
rect 55918 29486 55970 29538
rect 57822 29486 57874 29538
rect 1710 29374 1762 29426
rect 2382 29374 2434 29426
rect 3502 29374 3554 29426
rect 4174 29374 4226 29426
rect 4622 29374 4674 29426
rect 6974 29374 7026 29426
rect 7422 29374 7474 29426
rect 7758 29374 7810 29426
rect 8094 29374 8146 29426
rect 8990 29374 9042 29426
rect 9886 29374 9938 29426
rect 12238 29374 12290 29426
rect 21982 29374 22034 29426
rect 23438 29374 23490 29426
rect 26574 29374 26626 29426
rect 30382 29374 30434 29426
rect 30942 29374 30994 29426
rect 31838 29374 31890 29426
rect 33182 29374 33234 29426
rect 33406 29374 33458 29426
rect 33518 29374 33570 29426
rect 33854 29374 33906 29426
rect 34414 29374 34466 29426
rect 35198 29374 35250 29426
rect 36318 29374 36370 29426
rect 36654 29374 36706 29426
rect 36990 29374 37042 29426
rect 37214 29374 37266 29426
rect 37550 29374 37602 29426
rect 38446 29374 38498 29426
rect 38782 29374 38834 29426
rect 39454 29374 39506 29426
rect 42702 29374 42754 29426
rect 43038 29374 43090 29426
rect 43374 29374 43426 29426
rect 44158 29374 44210 29426
rect 47406 29374 47458 29426
rect 48078 29374 48130 29426
rect 49758 29374 49810 29426
rect 49982 29374 50034 29426
rect 50878 29374 50930 29426
rect 51326 29374 51378 29426
rect 51998 29374 52050 29426
rect 52222 29374 52274 29426
rect 53230 29374 53282 29426
rect 54126 29374 54178 29426
rect 54798 29374 54850 29426
rect 57486 29374 57538 29426
rect 5070 29262 5122 29314
rect 5518 29262 5570 29314
rect 6190 29262 6242 29314
rect 6526 29262 6578 29314
rect 10670 29262 10722 29314
rect 11902 29262 11954 29314
rect 15150 29262 15202 29314
rect 19070 29262 19122 29314
rect 26350 29262 26402 29314
rect 29486 29262 29538 29314
rect 31054 29262 31106 29314
rect 31614 29262 31666 29314
rect 32398 29262 32450 29314
rect 36430 29262 36482 29314
rect 38558 29262 38610 29314
rect 41470 29262 41522 29314
rect 42478 29262 42530 29314
rect 49086 29262 49138 29314
rect 52558 29262 52610 29314
rect 56926 29262 56978 29314
rect 17838 29150 17890 29202
rect 22766 29150 22818 29202
rect 38894 29150 38946 29202
rect 44942 29150 44994 29202
rect 53118 29150 53170 29202
rect 54686 29150 54738 29202
rect 55246 29150 55298 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 18062 28814 18114 28866
rect 25678 28814 25730 28866
rect 27246 28814 27298 28866
rect 32510 28814 32562 28866
rect 37214 28814 37266 28866
rect 37774 28814 37826 28866
rect 4622 28702 4674 28754
rect 5966 28702 6018 28754
rect 7534 28702 7586 28754
rect 8094 28702 8146 28754
rect 13918 28702 13970 28754
rect 18286 28702 18338 28754
rect 18622 28702 18674 28754
rect 19294 28702 19346 28754
rect 22206 28702 22258 28754
rect 25118 28702 25170 28754
rect 30830 28702 30882 28754
rect 31614 28702 31666 28754
rect 32398 28702 32450 28754
rect 33294 28702 33346 28754
rect 33406 28702 33458 28754
rect 33854 28702 33906 28754
rect 34750 28702 34802 28754
rect 35646 28702 35698 28754
rect 37214 28702 37266 28754
rect 37998 28702 38050 28754
rect 40686 28702 40738 28754
rect 42254 28702 42306 28754
rect 44270 28702 44322 28754
rect 47966 28702 48018 28754
rect 48526 28702 48578 28754
rect 49870 28702 49922 28754
rect 51326 28702 51378 28754
rect 55246 28702 55298 28754
rect 55806 28702 55858 28754
rect 56366 28702 56418 28754
rect 57598 28702 57650 28754
rect 1822 28590 1874 28642
rect 6302 28590 6354 28642
rect 6638 28590 6690 28642
rect 7310 28590 7362 28642
rect 7982 28590 8034 28642
rect 8206 28590 8258 28642
rect 8654 28590 8706 28642
rect 9438 28590 9490 28642
rect 12462 28590 12514 28642
rect 13358 28590 13410 28642
rect 18510 28590 18562 28642
rect 26462 28590 26514 28642
rect 27582 28590 27634 28642
rect 28030 28590 28082 28642
rect 29934 28590 29986 28642
rect 30382 28590 30434 28642
rect 31502 28590 31554 28642
rect 31726 28590 31778 28642
rect 32062 28590 32114 28642
rect 35198 28590 35250 28642
rect 35534 28590 35586 28642
rect 35870 28590 35922 28642
rect 36542 28590 36594 28642
rect 40798 28590 40850 28642
rect 41134 28590 41186 28642
rect 41918 28590 41970 28642
rect 42590 28590 42642 28642
rect 43262 28590 43314 28642
rect 43486 28590 43538 28642
rect 45950 28590 46002 28642
rect 46174 28590 46226 28642
rect 47406 28590 47458 28642
rect 50430 28590 50482 28642
rect 50766 28590 50818 28642
rect 51886 28590 51938 28642
rect 53342 28590 53394 28642
rect 53902 28590 53954 28642
rect 54126 28590 54178 28642
rect 54686 28590 54738 28642
rect 55134 28590 55186 28642
rect 57150 28590 57202 28642
rect 58158 28590 58210 28642
rect 2494 28478 2546 28530
rect 6078 28478 6130 28530
rect 9102 28478 9154 28530
rect 12798 28478 12850 28530
rect 18734 28478 18786 28530
rect 25902 28478 25954 28530
rect 28366 28478 28418 28530
rect 29598 28478 29650 28530
rect 33182 28478 33234 28530
rect 34862 28478 34914 28530
rect 35086 28478 35138 28530
rect 36206 28478 36258 28530
rect 36318 28478 36370 28530
rect 43710 28478 43762 28530
rect 43822 28478 43874 28530
rect 46622 28478 46674 28530
rect 51438 28478 51490 28530
rect 52894 28478 52946 28530
rect 5070 28366 5122 28418
rect 12686 28366 12738 28418
rect 13806 28366 13858 28418
rect 14030 28366 14082 28418
rect 17838 28366 17890 28418
rect 19854 28366 19906 28418
rect 20302 28366 20354 28418
rect 23662 28366 23714 28418
rect 23998 28366 24050 28418
rect 24670 28366 24722 28418
rect 25790 28366 25842 28418
rect 37550 28366 37602 28418
rect 38558 28366 38610 28418
rect 39006 28366 39058 28418
rect 40574 28366 40626 28418
rect 45278 28366 45330 28418
rect 45390 28366 45442 28418
rect 45502 28366 45554 28418
rect 46734 28366 46786 28418
rect 46846 28366 46898 28418
rect 47854 28366 47906 28418
rect 48078 28366 48130 28418
rect 51214 28366 51266 28418
rect 52670 28366 52722 28418
rect 52782 28366 52834 28418
rect 53566 28366 53618 28418
rect 54910 28366 54962 28418
rect 55246 28366 55298 28418
rect 55918 28366 55970 28418
rect 57822 28366 57874 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 2718 28030 2770 28082
rect 3166 28030 3218 28082
rect 3614 28030 3666 28082
rect 3726 28030 3778 28082
rect 4622 28030 4674 28082
rect 13022 28030 13074 28082
rect 13582 28030 13634 28082
rect 14254 28030 14306 28082
rect 18062 28030 18114 28082
rect 22094 28030 22146 28082
rect 26686 28030 26738 28082
rect 28366 28030 28418 28082
rect 29262 28030 29314 28082
rect 30270 28030 30322 28082
rect 31838 28030 31890 28082
rect 39006 28030 39058 28082
rect 42254 28030 42306 28082
rect 42366 28030 42418 28082
rect 43150 28030 43202 28082
rect 44158 28030 44210 28082
rect 44270 28030 44322 28082
rect 48862 28030 48914 28082
rect 49982 28030 50034 28082
rect 55358 28030 55410 28082
rect 1710 27918 1762 27970
rect 2046 27918 2098 27970
rect 5070 27918 5122 27970
rect 5518 27918 5570 27970
rect 5630 27918 5682 27970
rect 8430 27918 8482 27970
rect 11566 27918 11618 27970
rect 12798 27918 12850 27970
rect 13246 27918 13298 27970
rect 13806 27918 13858 27970
rect 13918 27918 13970 27970
rect 14590 27918 14642 27970
rect 17390 27918 17442 27970
rect 19182 27918 19234 27970
rect 22990 27918 23042 27970
rect 23662 27918 23714 27970
rect 28590 27918 28642 27970
rect 29710 27918 29762 27970
rect 33294 27918 33346 27970
rect 35870 27918 35922 27970
rect 40238 27918 40290 27970
rect 42590 27918 42642 27970
rect 44046 27918 44098 27970
rect 46062 27918 46114 27970
rect 50430 27918 50482 27970
rect 53006 27918 53058 27970
rect 57822 27918 57874 27970
rect 2494 27806 2546 27858
rect 3502 27806 3554 27858
rect 4174 27806 4226 27858
rect 4398 27806 4450 27858
rect 4846 27806 4898 27858
rect 5294 27806 5346 27858
rect 7646 27806 7698 27858
rect 9550 27806 9602 27858
rect 9774 27806 9826 27858
rect 10222 27806 10274 27858
rect 11790 27806 11842 27858
rect 12462 27806 12514 27858
rect 13358 27806 13410 27858
rect 18286 27806 18338 27858
rect 18622 27806 18674 27858
rect 19630 27806 19682 27858
rect 21086 27806 21138 27858
rect 21646 27806 21698 27858
rect 22430 27806 22482 27858
rect 23214 27806 23266 27858
rect 24110 27806 24162 27858
rect 25566 27806 25618 27858
rect 25902 27806 25954 27858
rect 26014 27806 26066 27858
rect 28702 27806 28754 27858
rect 28814 27806 28866 27858
rect 29038 27806 29090 27858
rect 29374 27806 29426 27858
rect 31950 27806 32002 27858
rect 32062 27806 32114 27858
rect 33966 27806 34018 27858
rect 36094 27806 36146 27858
rect 36318 27806 36370 27858
rect 37662 27806 37714 27858
rect 38558 27806 38610 27858
rect 39230 27806 39282 27858
rect 40126 27806 40178 27858
rect 40462 27806 40514 27858
rect 41358 27806 41410 27858
rect 41582 27806 41634 27858
rect 41806 27806 41858 27858
rect 42142 27806 42194 27858
rect 43486 27806 43538 27858
rect 43822 27806 43874 27858
rect 45390 27806 45442 27858
rect 51550 27806 51602 27858
rect 51998 27806 52050 27858
rect 54238 27806 54290 27858
rect 54686 27806 54738 27858
rect 55694 27806 55746 27858
rect 58158 27806 58210 27858
rect 7422 27694 7474 27746
rect 9662 27694 9714 27746
rect 17726 27694 17778 27746
rect 18174 27694 18226 27746
rect 20078 27694 20130 27746
rect 21198 27694 21250 27746
rect 24558 27694 24610 27746
rect 25678 27694 25730 27746
rect 31054 27694 31106 27746
rect 32286 27694 32338 27746
rect 34190 27694 34242 27746
rect 34750 27694 34802 27746
rect 35198 27694 35250 27746
rect 37326 27694 37378 27746
rect 38222 27694 38274 27746
rect 38782 27694 38834 27746
rect 39118 27694 39170 27746
rect 44718 27694 44770 27746
rect 48190 27694 48242 27746
rect 54014 27694 54066 27746
rect 57150 27694 57202 27746
rect 57598 27694 57650 27746
rect 7982 27582 8034 27634
rect 8654 27582 8706 27634
rect 8990 27582 9042 27634
rect 12126 27582 12178 27634
rect 32510 27582 32562 27634
rect 40910 27582 40962 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 18622 27246 18674 27298
rect 19742 27246 19794 27298
rect 20190 27246 20242 27298
rect 24110 27246 24162 27298
rect 33070 27246 33122 27298
rect 38670 27246 38722 27298
rect 51214 27246 51266 27298
rect 54350 27246 54402 27298
rect 54574 27246 54626 27298
rect 55022 27246 55074 27298
rect 6414 27134 6466 27186
rect 14142 27134 14194 27186
rect 18174 27134 18226 27186
rect 21422 27134 21474 27186
rect 22430 27134 22482 27186
rect 23214 27134 23266 27186
rect 25454 27134 25506 27186
rect 27582 27134 27634 27186
rect 32510 27134 32562 27186
rect 33630 27134 33682 27186
rect 34190 27134 34242 27186
rect 35310 27134 35362 27186
rect 36318 27134 36370 27186
rect 37550 27134 37602 27186
rect 40238 27134 40290 27186
rect 41134 27134 41186 27186
rect 43038 27134 43090 27186
rect 43934 27134 43986 27186
rect 44942 27134 44994 27186
rect 46174 27134 46226 27186
rect 47742 27134 47794 27186
rect 51102 27134 51154 27186
rect 52782 27134 52834 27186
rect 54910 27134 54962 27186
rect 56030 27134 56082 27186
rect 58158 27134 58210 27186
rect 1710 27022 1762 27074
rect 2494 27022 2546 27074
rect 3502 27022 3554 27074
rect 3950 27022 4002 27074
rect 4398 27022 4450 27074
rect 4622 27022 4674 27074
rect 4734 27022 4786 27074
rect 5070 27022 5122 27074
rect 8430 27022 8482 27074
rect 10446 27022 10498 27074
rect 12574 27022 12626 27074
rect 13806 27022 13858 27074
rect 14030 27022 14082 27074
rect 14366 27022 14418 27074
rect 15262 27022 15314 27074
rect 18958 27022 19010 27074
rect 19294 27022 19346 27074
rect 19854 27022 19906 27074
rect 20414 27022 20466 27074
rect 21310 27022 21362 27074
rect 22766 27022 22818 27074
rect 23438 27022 23490 27074
rect 23886 27022 23938 27074
rect 24334 27022 24386 27074
rect 24782 27022 24834 27074
rect 30494 27022 30546 27074
rect 31166 27022 31218 27074
rect 32062 27022 32114 27074
rect 32622 27022 32674 27074
rect 33966 27022 34018 27074
rect 34414 27022 34466 27074
rect 36206 27022 36258 27074
rect 36430 27022 36482 27074
rect 37326 27022 37378 27074
rect 37774 27022 37826 27074
rect 38222 27022 38274 27074
rect 38782 27022 38834 27074
rect 40910 27022 40962 27074
rect 41358 27022 41410 27074
rect 41470 27022 41522 27074
rect 42590 27022 42642 27074
rect 43486 27022 43538 27074
rect 45502 27022 45554 27074
rect 45950 27022 46002 27074
rect 46398 27022 46450 27074
rect 47854 27022 47906 27074
rect 48638 27022 48690 27074
rect 51550 27022 51602 27074
rect 51774 27022 51826 27074
rect 52670 27022 52722 27074
rect 53454 27022 53506 27074
rect 54014 27022 54066 27074
rect 55246 27022 55298 27074
rect 2046 26910 2098 26962
rect 2718 26910 2770 26962
rect 3278 26910 3330 26962
rect 5742 26910 5794 26962
rect 6526 26910 6578 26962
rect 6750 26910 6802 26962
rect 7870 26910 7922 26962
rect 7982 26910 8034 26962
rect 8542 26910 8594 26962
rect 11006 26910 11058 26962
rect 12910 26910 12962 26962
rect 14590 26910 14642 26962
rect 14702 26910 14754 26962
rect 16046 26910 16098 26962
rect 19630 26910 19682 26962
rect 21534 26910 21586 26962
rect 30158 26910 30210 26962
rect 30942 26910 30994 26962
rect 31726 26910 31778 26962
rect 31838 26910 31890 26962
rect 32286 26910 32338 26962
rect 32958 26910 33010 26962
rect 33070 26910 33122 26962
rect 34750 26910 34802 26962
rect 35982 26910 36034 26962
rect 36878 26910 36930 26962
rect 38670 26910 38722 26962
rect 39342 26910 39394 26962
rect 43934 26910 43986 26962
rect 44046 26910 44098 26962
rect 44830 26910 44882 26962
rect 45726 26910 45778 26962
rect 46958 26910 47010 26962
rect 47518 26910 47570 26962
rect 52894 26910 52946 26962
rect 53006 26910 53058 26962
rect 53790 26910 53842 26962
rect 4062 26798 4114 26850
rect 4286 26798 4338 26850
rect 8206 26798 8258 26850
rect 9438 26798 9490 26850
rect 14926 26798 14978 26850
rect 18734 26798 18786 26850
rect 21758 26798 21810 26850
rect 31502 26798 31554 26850
rect 34638 26798 34690 26850
rect 40686 26798 40738 26850
rect 42030 26798 42082 26850
rect 44270 26798 44322 26850
rect 45054 26798 45106 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 7086 26462 7138 26514
rect 13358 26462 13410 26514
rect 14590 26462 14642 26514
rect 14814 26462 14866 26514
rect 15934 26462 15986 26514
rect 16382 26462 16434 26514
rect 19070 26462 19122 26514
rect 19966 26462 20018 26514
rect 21086 26462 21138 26514
rect 22766 26462 22818 26514
rect 25230 26462 25282 26514
rect 25342 26462 25394 26514
rect 28478 26462 28530 26514
rect 28814 26462 28866 26514
rect 30606 26462 30658 26514
rect 31278 26462 31330 26514
rect 33182 26462 33234 26514
rect 36206 26462 36258 26514
rect 36430 26462 36482 26514
rect 37214 26462 37266 26514
rect 38110 26462 38162 26514
rect 38446 26462 38498 26514
rect 41918 26462 41970 26514
rect 42814 26462 42866 26514
rect 43374 26462 43426 26514
rect 43710 26462 43762 26514
rect 45054 26462 45106 26514
rect 45502 26462 45554 26514
rect 50542 26462 50594 26514
rect 51438 26462 51490 26514
rect 53118 26462 53170 26514
rect 55246 26462 55298 26514
rect 57822 26462 57874 26514
rect 7982 26350 8034 26402
rect 13246 26350 13298 26402
rect 15038 26350 15090 26402
rect 18062 26350 18114 26402
rect 18398 26350 18450 26402
rect 22990 26350 23042 26402
rect 23102 26350 23154 26402
rect 29710 26350 29762 26402
rect 30158 26350 30210 26402
rect 30942 26350 30994 26402
rect 35758 26350 35810 26402
rect 36542 26350 36594 26402
rect 39902 26350 39954 26402
rect 42590 26350 42642 26402
rect 43150 26350 43202 26402
rect 44606 26350 44658 26402
rect 47854 26350 47906 26402
rect 49086 26350 49138 26402
rect 51214 26350 51266 26402
rect 51662 26350 51714 26402
rect 51774 26350 51826 26402
rect 52782 26350 52834 26402
rect 52894 26350 52946 26402
rect 54350 26350 54402 26402
rect 57150 26350 57202 26402
rect 1822 26238 1874 26290
rect 5966 26238 6018 26290
rect 6414 26238 6466 26290
rect 6638 26238 6690 26290
rect 8206 26238 8258 26290
rect 8430 26238 8482 26290
rect 9662 26238 9714 26290
rect 9998 26238 10050 26290
rect 12014 26238 12066 26290
rect 12238 26238 12290 26290
rect 13582 26238 13634 26290
rect 14366 26238 14418 26290
rect 16718 26238 16770 26290
rect 17502 26238 17554 26290
rect 17838 26238 17890 26290
rect 19294 26238 19346 26290
rect 21758 26238 21810 26290
rect 21982 26238 22034 26290
rect 25454 26238 25506 26290
rect 25902 26238 25954 26290
rect 28142 26238 28194 26290
rect 28926 26238 28978 26290
rect 29150 26238 29202 26290
rect 29486 26238 29538 26290
rect 31502 26238 31554 26290
rect 34414 26238 34466 26290
rect 35534 26238 35586 26290
rect 39230 26238 39282 26290
rect 42478 26238 42530 26290
rect 43038 26238 43090 26290
rect 48862 26238 48914 26290
rect 50318 26238 50370 26290
rect 50654 26238 50706 26290
rect 51102 26238 51154 26290
rect 54014 26238 54066 26290
rect 55134 26238 55186 26290
rect 55470 26238 55522 26290
rect 55582 26238 55634 26290
rect 57486 26238 57538 26290
rect 58046 26238 58098 26290
rect 2494 26126 2546 26178
rect 4622 26126 4674 26178
rect 5406 26126 5458 26178
rect 6190 26126 6242 26178
rect 6974 26126 7026 26178
rect 7310 26126 7362 26178
rect 9550 26126 9602 26178
rect 15486 26126 15538 26178
rect 20638 26126 20690 26178
rect 22430 26126 22482 26178
rect 23550 26126 23602 26178
rect 24110 26126 24162 26178
rect 24558 26126 24610 26178
rect 26238 26126 26290 26178
rect 27806 26126 27858 26178
rect 33742 26126 33794 26178
rect 33966 26126 34018 26178
rect 35086 26126 35138 26178
rect 39006 26126 39058 26178
rect 40350 26126 40402 26178
rect 41134 26126 41186 26178
rect 44158 26126 44210 26178
rect 47294 26126 47346 26178
rect 47966 26126 48018 26178
rect 53678 26126 53730 26178
rect 55358 26126 55410 26178
rect 56702 26126 56754 26178
rect 5070 26014 5122 26066
rect 5182 26014 5234 26066
rect 5630 26014 5682 26066
rect 5742 26014 5794 26066
rect 11678 26014 11730 26066
rect 14926 26014 14978 26066
rect 47070 26014 47122 26066
rect 47294 26014 47346 26066
rect 47630 26014 47682 26066
rect 51774 26014 51826 26066
rect 56590 26014 56642 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 6190 25678 6242 25730
rect 13918 25678 13970 25730
rect 14254 25678 14306 25730
rect 19518 25678 19570 25730
rect 28254 25678 28306 25730
rect 48750 25678 48802 25730
rect 2270 25566 2322 25618
rect 3838 25566 3890 25618
rect 7982 25566 8034 25618
rect 15486 25566 15538 25618
rect 16046 25566 16098 25618
rect 18398 25566 18450 25618
rect 19070 25566 19122 25618
rect 21758 25566 21810 25618
rect 24110 25566 24162 25618
rect 28478 25566 28530 25618
rect 34190 25566 34242 25618
rect 38446 25566 38498 25618
rect 39902 25566 39954 25618
rect 42366 25566 42418 25618
rect 43486 25566 43538 25618
rect 43822 25566 43874 25618
rect 51326 25566 51378 25618
rect 51998 25566 52050 25618
rect 54910 25566 54962 25618
rect 56030 25566 56082 25618
rect 58158 25566 58210 25618
rect 1710 25454 1762 25506
rect 3166 25454 3218 25506
rect 3726 25454 3778 25506
rect 4286 25454 4338 25506
rect 5854 25454 5906 25506
rect 6078 25454 6130 25506
rect 6302 25454 6354 25506
rect 6974 25454 7026 25506
rect 7646 25454 7698 25506
rect 10334 25454 10386 25506
rect 15038 25454 15090 25506
rect 19294 25454 19346 25506
rect 20302 25454 20354 25506
rect 22430 25454 22482 25506
rect 24558 25454 24610 25506
rect 26238 25454 26290 25506
rect 26798 25454 26850 25506
rect 28030 25454 28082 25506
rect 29822 25454 29874 25506
rect 30382 25454 30434 25506
rect 32062 25454 32114 25506
rect 35422 25454 35474 25506
rect 37886 25454 37938 25506
rect 39342 25454 39394 25506
rect 39790 25454 39842 25506
rect 40574 25454 40626 25506
rect 41470 25454 41522 25506
rect 41918 25454 41970 25506
rect 48974 25454 49026 25506
rect 49198 25454 49250 25506
rect 49870 25454 49922 25506
rect 51662 25454 51714 25506
rect 53006 25454 53058 25506
rect 55246 25454 55298 25506
rect 2718 25342 2770 25394
rect 5630 25342 5682 25394
rect 6750 25342 6802 25394
rect 9998 25342 10050 25394
rect 21310 25342 21362 25394
rect 22654 25342 22706 25394
rect 26910 25342 26962 25394
rect 27246 25342 27298 25394
rect 27470 25342 27522 25394
rect 27694 25342 27746 25394
rect 28030 25342 28082 25394
rect 28590 25342 28642 25394
rect 30606 25342 30658 25394
rect 38558 25342 38610 25394
rect 40238 25342 40290 25394
rect 40798 25342 40850 25394
rect 45166 25342 45218 25394
rect 49422 25342 49474 25394
rect 50318 25342 50370 25394
rect 50542 25342 50594 25394
rect 51214 25342 51266 25394
rect 51326 25342 51378 25394
rect 51438 25342 51490 25394
rect 52110 25342 52162 25394
rect 52670 25342 52722 25394
rect 52782 25342 52834 25394
rect 53454 25342 53506 25394
rect 3390 25230 3442 25282
rect 3950 25230 4002 25282
rect 4846 25230 4898 25282
rect 14142 25230 14194 25282
rect 14702 25230 14754 25282
rect 17950 25230 18002 25282
rect 19854 25230 19906 25282
rect 25006 25230 25058 25282
rect 27358 25230 27410 25282
rect 29486 25230 29538 25282
rect 31278 25230 31330 25282
rect 31502 25230 31554 25282
rect 33966 25230 34018 25282
rect 34750 25230 34802 25282
rect 35198 25230 35250 25282
rect 37774 25230 37826 25282
rect 38334 25230 38386 25282
rect 40350 25230 40402 25282
rect 40910 25230 40962 25282
rect 42926 25230 42978 25282
rect 44270 25230 44322 25282
rect 45502 25230 45554 25282
rect 47742 25230 47794 25282
rect 48078 25230 48130 25282
rect 48302 25230 48354 25282
rect 50206 25230 50258 25282
rect 53342 25230 53394 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 2046 24894 2098 24946
rect 2718 24894 2770 24946
rect 3502 24894 3554 24946
rect 4398 24894 4450 24946
rect 5518 24894 5570 24946
rect 7758 24894 7810 24946
rect 9662 24894 9714 24946
rect 10110 24894 10162 24946
rect 11118 24894 11170 24946
rect 18734 24894 18786 24946
rect 22878 24894 22930 24946
rect 25678 24894 25730 24946
rect 30158 24894 30210 24946
rect 35086 24894 35138 24946
rect 36094 24894 36146 24946
rect 38782 24894 38834 24946
rect 40238 24894 40290 24946
rect 41246 24894 41298 24946
rect 43038 24894 43090 24946
rect 54686 24894 54738 24946
rect 55358 24894 55410 24946
rect 56926 24894 56978 24946
rect 57486 24894 57538 24946
rect 57822 24894 57874 24946
rect 58158 24894 58210 24946
rect 4734 24782 4786 24834
rect 5742 24782 5794 24834
rect 6190 24782 6242 24834
rect 6302 24782 6354 24834
rect 14926 24782 14978 24834
rect 15598 24782 15650 24834
rect 15710 24782 15762 24834
rect 16270 24782 16322 24834
rect 16494 24782 16546 24834
rect 16606 24782 16658 24834
rect 23662 24782 23714 24834
rect 23998 24782 24050 24834
rect 26126 24782 26178 24834
rect 29150 24782 29202 24834
rect 34750 24782 34802 24834
rect 35422 24782 35474 24834
rect 35758 24782 35810 24834
rect 36430 24782 36482 24834
rect 39118 24782 39170 24834
rect 41022 24782 41074 24834
rect 45838 24782 45890 24834
rect 54910 24782 54962 24834
rect 57150 24782 57202 24834
rect 1710 24670 1762 24722
rect 2382 24670 2434 24722
rect 5294 24670 5346 24722
rect 7310 24670 7362 24722
rect 11454 24670 11506 24722
rect 17502 24670 17554 24722
rect 18062 24670 18114 24722
rect 19294 24670 19346 24722
rect 22766 24670 22818 24722
rect 25454 24670 25506 24722
rect 25902 24670 25954 24722
rect 26910 24670 26962 24722
rect 27358 24670 27410 24722
rect 27582 24670 27634 24722
rect 27806 24670 27858 24722
rect 28590 24670 28642 24722
rect 30046 24670 30098 24722
rect 30270 24670 30322 24722
rect 33070 24670 33122 24722
rect 33182 24670 33234 24722
rect 33518 24670 33570 24722
rect 39342 24670 39394 24722
rect 40910 24670 40962 24722
rect 42142 24670 42194 24722
rect 42366 24670 42418 24722
rect 42926 24670 42978 24722
rect 43150 24670 43202 24722
rect 43598 24670 43650 24722
rect 43822 24670 43874 24722
rect 44270 24670 44322 24722
rect 44494 24670 44546 24722
rect 45166 24670 45218 24722
rect 50206 24670 50258 24722
rect 50654 24670 50706 24722
rect 50990 24670 51042 24722
rect 51102 24670 51154 24722
rect 51438 24670 51490 24722
rect 52446 24670 52498 24722
rect 52782 24670 52834 24722
rect 53678 24670 53730 24722
rect 55134 24670 55186 24722
rect 55582 24670 55634 24722
rect 3838 24558 3890 24610
rect 5406 24558 5458 24610
rect 6974 24558 7026 24610
rect 12238 24558 12290 24610
rect 14366 24558 14418 24610
rect 14814 24558 14866 24610
rect 20078 24558 20130 24610
rect 22206 24558 22258 24610
rect 23326 24558 23378 24610
rect 24670 24558 24722 24610
rect 28478 24558 28530 24610
rect 29822 24558 29874 24610
rect 38222 24558 38274 24610
rect 44382 24558 44434 24610
rect 47966 24558 48018 24610
rect 48974 24558 49026 24610
rect 49758 24558 49810 24610
rect 52334 24558 52386 24610
rect 53790 24558 53842 24610
rect 55246 24558 55298 24610
rect 56030 24558 56082 24610
rect 3838 24446 3890 24498
rect 4062 24446 4114 24498
rect 6302 24446 6354 24498
rect 14702 24446 14754 24498
rect 15710 24446 15762 24498
rect 29598 24446 29650 24498
rect 38446 24446 38498 24498
rect 39566 24446 39618 24498
rect 39790 24446 39842 24498
rect 42478 24446 42530 24498
rect 55918 24446 55970 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 13806 24110 13858 24162
rect 20638 24110 20690 24162
rect 26686 24110 26738 24162
rect 30494 24110 30546 24162
rect 31054 24110 31106 24162
rect 32734 24110 32786 24162
rect 39230 24110 39282 24162
rect 39790 24110 39842 24162
rect 39902 24110 39954 24162
rect 40574 24110 40626 24162
rect 41358 24110 41410 24162
rect 44942 24110 44994 24162
rect 45278 24110 45330 24162
rect 48078 24110 48130 24162
rect 53118 24110 53170 24162
rect 4622 23998 4674 24050
rect 5070 23998 5122 24050
rect 7086 23998 7138 24050
rect 9214 23998 9266 24050
rect 9550 23998 9602 24050
rect 12910 23998 12962 24050
rect 14254 23998 14306 24050
rect 15598 23998 15650 24050
rect 17726 23998 17778 24050
rect 19070 23998 19122 24050
rect 19966 23998 20018 24050
rect 20750 23998 20802 24050
rect 21422 23998 21474 24050
rect 23550 23998 23602 24050
rect 25678 23998 25730 24050
rect 29934 23998 29986 24050
rect 30606 23998 30658 24050
rect 31054 23998 31106 24050
rect 39790 23998 39842 24050
rect 40350 23998 40402 24050
rect 46622 23998 46674 24050
rect 48638 23998 48690 24050
rect 52894 23998 52946 24050
rect 54798 23998 54850 24050
rect 55806 23998 55858 24050
rect 57934 23998 57986 24050
rect 1822 23886 1874 23938
rect 5742 23886 5794 23938
rect 6302 23886 6354 23938
rect 12350 23886 12402 23938
rect 14926 23886 14978 23938
rect 18062 23886 18114 23938
rect 18622 23886 18674 23938
rect 19518 23886 19570 23938
rect 21534 23886 21586 23938
rect 22766 23886 22818 23938
rect 26238 23886 26290 23938
rect 26462 23886 26514 23938
rect 27358 23886 27410 23938
rect 28030 23886 28082 23938
rect 29486 23886 29538 23938
rect 33854 23886 33906 23938
rect 34078 23886 34130 23938
rect 35086 23886 35138 23938
rect 35534 23886 35586 23938
rect 37662 23886 37714 23938
rect 37998 23886 38050 23938
rect 38894 23886 38946 23938
rect 39118 23886 39170 23938
rect 40798 23886 40850 23938
rect 41470 23886 41522 23938
rect 41694 23886 41746 23938
rect 41806 23886 41858 23938
rect 43710 23886 43762 23938
rect 43934 23886 43986 23938
rect 46958 23886 47010 23938
rect 47406 23886 47458 23938
rect 47630 23886 47682 23938
rect 47854 23886 47906 23938
rect 50654 23886 50706 23938
rect 50878 23886 50930 23938
rect 51102 23886 51154 23938
rect 53566 23886 53618 23938
rect 55022 23886 55074 23938
rect 2494 23774 2546 23826
rect 11678 23774 11730 23826
rect 13470 23774 13522 23826
rect 13694 23774 13746 23826
rect 21982 23774 22034 23826
rect 26014 23774 26066 23826
rect 27694 23774 27746 23826
rect 29150 23774 29202 23826
rect 32734 23774 32786 23826
rect 32846 23774 32898 23826
rect 33182 23774 33234 23826
rect 36990 23774 37042 23826
rect 38558 23774 38610 23826
rect 41022 23774 41074 23826
rect 42478 23774 42530 23826
rect 45614 23774 45666 23826
rect 45950 23774 46002 23826
rect 50542 23774 50594 23826
rect 51438 23774 51490 23826
rect 51886 23774 51938 23826
rect 5966 23662 6018 23714
rect 12798 23662 12850 23714
rect 21422 23662 21474 23714
rect 21758 23662 21810 23714
rect 22430 23662 22482 23714
rect 27134 23662 27186 23714
rect 28142 23662 28194 23714
rect 28366 23662 28418 23714
rect 29262 23662 29314 23714
rect 31950 23662 32002 23714
rect 34750 23662 34802 23714
rect 35758 23662 35810 23714
rect 36318 23662 36370 23714
rect 37326 23662 37378 23714
rect 38110 23662 38162 23714
rect 38222 23662 38274 23714
rect 38782 23662 38834 23714
rect 42590 23662 42642 23714
rect 42814 23662 42866 23714
rect 43262 23662 43314 23714
rect 43374 23662 43426 23714
rect 43486 23662 43538 23714
rect 49086 23662 49138 23714
rect 50318 23662 50370 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 2606 23326 2658 23378
rect 3726 23326 3778 23378
rect 5630 23326 5682 23378
rect 8766 23326 8818 23378
rect 16830 23326 16882 23378
rect 17390 23326 17442 23378
rect 18174 23326 18226 23378
rect 27694 23326 27746 23378
rect 29710 23326 29762 23378
rect 31278 23326 31330 23378
rect 32510 23326 32562 23378
rect 42366 23326 42418 23378
rect 43150 23326 43202 23378
rect 43486 23326 43538 23378
rect 51214 23326 51266 23378
rect 51998 23326 52050 23378
rect 57822 23326 57874 23378
rect 4286 23214 4338 23266
rect 5742 23214 5794 23266
rect 7422 23214 7474 23266
rect 9662 23214 9714 23266
rect 11678 23214 11730 23266
rect 11902 23214 11954 23266
rect 12350 23214 12402 23266
rect 16494 23214 16546 23266
rect 27582 23214 27634 23266
rect 28814 23214 28866 23266
rect 29038 23214 29090 23266
rect 30494 23214 30546 23266
rect 42814 23214 42866 23266
rect 42926 23214 42978 23266
rect 45614 23214 45666 23266
rect 46062 23214 46114 23266
rect 48750 23214 48802 23266
rect 51326 23214 51378 23266
rect 55582 23214 55634 23266
rect 57150 23214 57202 23266
rect 57486 23214 57538 23266
rect 58158 23214 58210 23266
rect 1710 23102 1762 23154
rect 2942 23102 2994 23154
rect 3278 23102 3330 23154
rect 3614 23102 3666 23154
rect 3950 23102 4002 23154
rect 4846 23102 4898 23154
rect 5294 23102 5346 23154
rect 6302 23102 6354 23154
rect 7310 23102 7362 23154
rect 8878 23102 8930 23154
rect 9550 23102 9602 23154
rect 9886 23102 9938 23154
rect 9998 23102 10050 23154
rect 11342 23102 11394 23154
rect 11566 23102 11618 23154
rect 11790 23102 11842 23154
rect 12686 23102 12738 23154
rect 17614 23102 17666 23154
rect 19182 23102 19234 23154
rect 22990 23102 23042 23154
rect 23438 23102 23490 23154
rect 28702 23102 28754 23154
rect 29486 23102 29538 23154
rect 29710 23102 29762 23154
rect 30046 23102 30098 23154
rect 30606 23102 30658 23154
rect 30830 23102 30882 23154
rect 31502 23102 31554 23154
rect 32286 23102 32338 23154
rect 33070 23102 33122 23154
rect 33630 23102 33682 23154
rect 34638 23102 34690 23154
rect 36878 23102 36930 23154
rect 38894 23102 38946 23154
rect 39342 23102 39394 23154
rect 40238 23102 40290 23154
rect 45278 23102 45330 23154
rect 47518 23102 47570 23154
rect 49422 23102 49474 23154
rect 50878 23102 50930 23154
rect 50990 23102 51042 23154
rect 51886 23102 51938 23154
rect 52222 23102 52274 23154
rect 55246 23102 55298 23154
rect 55358 23102 55410 23154
rect 55694 23102 55746 23154
rect 2270 22990 2322 23042
rect 6638 22990 6690 23042
rect 8430 22990 8482 23042
rect 10558 22990 10610 23042
rect 13134 22990 13186 23042
rect 18734 22990 18786 23042
rect 19854 22990 19906 23042
rect 21982 22990 22034 23042
rect 22430 22990 22482 23042
rect 23886 22990 23938 23042
rect 28366 22990 28418 23042
rect 31390 22990 31442 23042
rect 33966 22990 34018 23042
rect 34974 22990 35026 23042
rect 35758 22990 35810 23042
rect 36206 22990 36258 23042
rect 38110 22990 38162 23042
rect 39790 22990 39842 23042
rect 41134 22990 41186 23042
rect 41470 22990 41522 23042
rect 41694 22990 41746 23042
rect 41918 22990 41970 23042
rect 8990 22878 9042 22930
rect 30494 22878 30546 22930
rect 34414 22878 34466 22930
rect 34526 22878 34578 22930
rect 35198 22878 35250 22930
rect 35534 22878 35586 22930
rect 36318 22878 36370 22930
rect 37102 22878 37154 22930
rect 37326 22878 37378 22930
rect 37550 22878 37602 22930
rect 41134 22878 41186 22930
rect 41582 22878 41634 22930
rect 43934 22990 43986 23042
rect 44382 22990 44434 23042
rect 46622 22990 46674 23042
rect 47070 22990 47122 23042
rect 48078 22990 48130 23042
rect 49646 22990 49698 23042
rect 52670 22990 52722 23042
rect 55470 22990 55522 23042
rect 56702 22990 56754 23042
rect 41918 22878 41970 22930
rect 44046 22878 44098 22930
rect 44606 22878 44658 22930
rect 44942 22878 44994 22930
rect 47742 22878 47794 22930
rect 56590 22878 56642 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 11454 22542 11506 22594
rect 17054 22542 17106 22594
rect 17614 22542 17666 22594
rect 20638 22542 20690 22594
rect 33406 22542 33458 22594
rect 37102 22542 37154 22594
rect 37550 22542 37602 22594
rect 39230 22542 39282 22594
rect 41694 22542 41746 22594
rect 50094 22542 50146 22594
rect 50990 22542 51042 22594
rect 51326 22542 51378 22594
rect 4622 22430 4674 22482
rect 5070 22430 5122 22482
rect 5742 22430 5794 22482
rect 6190 22430 6242 22482
rect 7534 22430 7586 22482
rect 12014 22430 12066 22482
rect 17054 22430 17106 22482
rect 17950 22430 18002 22482
rect 25342 22430 25394 22482
rect 27806 22430 27858 22482
rect 28142 22430 28194 22482
rect 30942 22430 30994 22482
rect 31614 22430 31666 22482
rect 32622 22430 32674 22482
rect 34414 22430 34466 22482
rect 37550 22430 37602 22482
rect 40686 22430 40738 22482
rect 41246 22430 41298 22482
rect 44942 22430 44994 22482
rect 52782 22430 52834 22482
rect 56030 22430 56082 22482
rect 58158 22430 58210 22482
rect 1822 22318 1874 22370
rect 7982 22318 8034 22370
rect 8318 22318 8370 22370
rect 11902 22318 11954 22370
rect 12238 22318 12290 22370
rect 12350 22318 12402 22370
rect 14478 22318 14530 22370
rect 28030 22318 28082 22370
rect 28590 22318 28642 22370
rect 29150 22318 29202 22370
rect 29710 22318 29762 22370
rect 31390 22318 31442 22370
rect 32062 22318 32114 22370
rect 33182 22318 33234 22370
rect 33630 22318 33682 22370
rect 34526 22318 34578 22370
rect 38558 22318 38610 22370
rect 41806 22318 41858 22370
rect 43038 22318 43090 22370
rect 45502 22318 45554 22370
rect 46286 22318 46338 22370
rect 50430 22318 50482 22370
rect 51998 22318 52050 22370
rect 54910 22318 54962 22370
rect 55246 22318 55298 22370
rect 2494 22206 2546 22258
rect 7870 22206 7922 22258
rect 11342 22206 11394 22258
rect 14814 22206 14866 22258
rect 15262 22206 15314 22258
rect 15934 22206 15986 22258
rect 18734 22206 18786 22258
rect 20750 22206 20802 22258
rect 22318 22206 22370 22258
rect 29822 22206 29874 22258
rect 30606 22206 30658 22258
rect 30830 22206 30882 22258
rect 32958 22206 33010 22258
rect 34750 22206 34802 22258
rect 38334 22206 38386 22258
rect 38894 22206 38946 22258
rect 39118 22206 39170 22258
rect 39454 22206 39506 22258
rect 39790 22206 39842 22258
rect 40238 22206 40290 22258
rect 42366 22206 42418 22258
rect 43150 22206 43202 22258
rect 43598 22206 43650 22258
rect 51662 22206 51714 22258
rect 51774 22206 51826 22258
rect 52670 22206 52722 22258
rect 52894 22206 52946 22258
rect 54462 22206 54514 22258
rect 9214 22094 9266 22146
rect 9326 22094 9378 22146
rect 9438 22094 9490 22146
rect 9662 22094 9714 22146
rect 11454 22094 11506 22146
rect 12910 22094 12962 22146
rect 13470 22094 13522 22146
rect 13806 22094 13858 22146
rect 14254 22094 14306 22146
rect 14702 22094 14754 22146
rect 15150 22094 15202 22146
rect 16270 22094 16322 22146
rect 17502 22094 17554 22146
rect 19294 22094 19346 22146
rect 22430 22094 22482 22146
rect 25790 22094 25842 22146
rect 28254 22094 28306 22146
rect 29374 22094 29426 22146
rect 31838 22094 31890 22146
rect 31950 22094 32002 22146
rect 34078 22094 34130 22146
rect 34302 22094 34354 22146
rect 35534 22094 35586 22146
rect 35870 22094 35922 22146
rect 36318 22094 36370 22146
rect 37102 22094 37154 22146
rect 41694 22094 41746 22146
rect 42478 22094 42530 22146
rect 42590 22094 42642 22146
rect 44046 22094 44098 22146
rect 45838 22094 45890 22146
rect 46734 22094 46786 22146
rect 50206 22094 50258 22146
rect 51214 22094 51266 22146
rect 53454 22094 53506 22146
rect 53790 22094 53842 22146
rect 54126 22094 54178 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 1710 21758 1762 21810
rect 2942 21758 2994 21810
rect 3390 21758 3442 21810
rect 3838 21758 3890 21810
rect 3950 21758 4002 21810
rect 4734 21758 4786 21810
rect 9774 21758 9826 21810
rect 13022 21758 13074 21810
rect 13358 21758 13410 21810
rect 13694 21758 13746 21810
rect 15598 21758 15650 21810
rect 17614 21758 17666 21810
rect 20974 21758 21026 21810
rect 21086 21758 21138 21810
rect 21198 21758 21250 21810
rect 28702 21758 28754 21810
rect 29150 21758 29202 21810
rect 29598 21758 29650 21810
rect 29934 21758 29986 21810
rect 30942 21758 30994 21810
rect 31502 21758 31554 21810
rect 4510 21646 4562 21698
rect 4846 21646 4898 21698
rect 5742 21646 5794 21698
rect 6414 21646 6466 21698
rect 6638 21646 6690 21698
rect 8990 21646 9042 21698
rect 11454 21646 11506 21698
rect 12686 21646 12738 21698
rect 16158 21646 16210 21698
rect 16718 21646 16770 21698
rect 17502 21646 17554 21698
rect 18174 21646 18226 21698
rect 18398 21646 18450 21698
rect 18510 21646 18562 21698
rect 21422 21646 21474 21698
rect 22542 21646 22594 21698
rect 26910 21646 26962 21698
rect 28478 21646 28530 21698
rect 30606 21646 30658 21698
rect 30718 21646 30770 21698
rect 32174 21702 32226 21754
rect 34414 21758 34466 21810
rect 34862 21758 34914 21810
rect 40014 21758 40066 21810
rect 40238 21758 40290 21810
rect 41022 21758 41074 21810
rect 49198 21758 49250 21810
rect 49534 21758 49586 21810
rect 50318 21758 50370 21810
rect 51102 21758 51154 21810
rect 52894 21758 52946 21810
rect 55246 21758 55298 21810
rect 57150 21758 57202 21810
rect 57598 21758 57650 21810
rect 57822 21758 57874 21810
rect 58158 21758 58210 21810
rect 32286 21646 32338 21698
rect 39566 21646 39618 21698
rect 41470 21646 41522 21698
rect 46062 21646 46114 21698
rect 50094 21646 50146 21698
rect 52446 21646 52498 21698
rect 54686 21646 54738 21698
rect 2606 21534 2658 21586
rect 3726 21534 3778 21586
rect 4398 21534 4450 21586
rect 5294 21534 5346 21586
rect 8318 21534 8370 21586
rect 8878 21534 8930 21586
rect 9438 21534 9490 21586
rect 9886 21534 9938 21586
rect 10110 21534 10162 21586
rect 10782 21534 10834 21586
rect 11230 21534 11282 21586
rect 12350 21534 12402 21586
rect 14254 21534 14306 21586
rect 14590 21534 14642 21586
rect 17390 21534 17442 21586
rect 18062 21534 18114 21586
rect 18958 21534 19010 21586
rect 19406 21534 19458 21586
rect 20862 21534 20914 21586
rect 21870 21534 21922 21586
rect 26014 21534 26066 21586
rect 28030 21534 28082 21586
rect 28366 21534 28418 21586
rect 29486 21534 29538 21586
rect 29710 21534 29762 21586
rect 31278 21534 31330 21586
rect 31390 21534 31442 21586
rect 31838 21534 31890 21586
rect 38110 21534 38162 21586
rect 38894 21534 38946 21586
rect 39118 21534 39170 21586
rect 39790 21534 39842 21586
rect 40350 21534 40402 21586
rect 41246 21534 41298 21586
rect 42030 21534 42082 21586
rect 45390 21534 45442 21586
rect 50430 21534 50482 21586
rect 50542 21534 50594 21586
rect 51550 21534 51602 21586
rect 52110 21534 52162 21586
rect 54910 21534 54962 21586
rect 55134 21534 55186 21586
rect 2270 21422 2322 21474
rect 15150 21422 15202 21474
rect 24670 21422 24722 21474
rect 25342 21422 25394 21474
rect 26686 21422 26738 21474
rect 33182 21422 33234 21474
rect 33966 21422 34018 21474
rect 35310 21422 35362 21474
rect 35870 21422 35922 21474
rect 36766 21422 36818 21474
rect 37214 21422 37266 21474
rect 37662 21422 37714 21474
rect 38670 21422 38722 21474
rect 39342 21422 39394 21474
rect 41358 21422 41410 21474
rect 42702 21422 42754 21474
rect 44830 21422 44882 21474
rect 48190 21422 48242 21474
rect 48862 21422 48914 21474
rect 52334 21422 52386 21474
rect 53342 21422 53394 21474
rect 53790 21422 53842 21474
rect 55022 21422 55074 21474
rect 55694 21422 55746 21474
rect 6302 21310 6354 21362
rect 15934 21310 15986 21362
rect 32286 21310 32338 21362
rect 36766 21310 36818 21362
rect 36990 21310 37042 21362
rect 38334 21310 38386 21362
rect 53342 21310 53394 21362
rect 53790 21310 53842 21362
rect 55806 21310 55858 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 8542 20974 8594 21026
rect 37662 20974 37714 21026
rect 38110 20974 38162 21026
rect 45838 20974 45890 21026
rect 52670 20974 52722 21026
rect 53118 20974 53170 21026
rect 2270 20862 2322 20914
rect 4398 20862 4450 20914
rect 5966 20862 6018 20914
rect 14478 20862 14530 20914
rect 14926 20862 14978 20914
rect 16046 20862 16098 20914
rect 18174 20862 18226 20914
rect 22206 20862 22258 20914
rect 23438 20862 23490 20914
rect 26686 20862 26738 20914
rect 31054 20862 31106 20914
rect 33182 20862 33234 20914
rect 38782 20862 38834 20914
rect 40462 20862 40514 20914
rect 41918 20862 41970 20914
rect 43262 20862 43314 20914
rect 45054 20862 45106 20914
rect 50206 20862 50258 20914
rect 51998 20862 52050 20914
rect 53230 20862 53282 20914
rect 53678 20862 53730 20914
rect 54014 20862 54066 20914
rect 56142 20862 56194 20914
rect 57822 20862 57874 20914
rect 58270 20862 58322 20914
rect 2718 20750 2770 20802
rect 3614 20750 3666 20802
rect 4062 20750 4114 20802
rect 4174 20750 4226 20802
rect 4622 20750 4674 20802
rect 4846 20750 4898 20802
rect 7422 20750 7474 20802
rect 7758 20750 7810 20802
rect 7982 20750 8034 20802
rect 8206 20750 8258 20802
rect 8430 20750 8482 20802
rect 8878 20750 8930 20802
rect 10894 20750 10946 20802
rect 14366 20750 14418 20802
rect 15262 20750 15314 20802
rect 18510 20750 18562 20802
rect 19406 20750 19458 20802
rect 19966 20750 20018 20802
rect 20526 20750 20578 20802
rect 21982 20750 22034 20802
rect 22094 20750 22146 20802
rect 23886 20750 23938 20802
rect 27918 20750 27970 20802
rect 28478 20750 28530 20802
rect 30046 20750 30098 20802
rect 30494 20750 30546 20802
rect 33966 20750 34018 20802
rect 34414 20750 34466 20802
rect 34750 20750 34802 20802
rect 35086 20750 35138 20802
rect 35646 20750 35698 20802
rect 35870 20750 35922 20802
rect 36094 20750 36146 20802
rect 37214 20750 37266 20802
rect 37438 20750 37490 20802
rect 39006 20750 39058 20802
rect 40574 20750 40626 20802
rect 41806 20750 41858 20802
rect 42030 20750 42082 20802
rect 42366 20750 42418 20802
rect 44270 20750 44322 20802
rect 46286 20750 46338 20802
rect 50318 20750 50370 20802
rect 50878 20750 50930 20802
rect 51550 20750 51602 20802
rect 56814 20750 56866 20802
rect 2942 20638 2994 20690
rect 6190 20638 6242 20690
rect 8990 20638 9042 20690
rect 12014 20638 12066 20690
rect 18846 20638 18898 20690
rect 19630 20638 19682 20690
rect 22318 20638 22370 20690
rect 22542 20638 22594 20690
rect 24558 20638 24610 20690
rect 27022 20638 27074 20690
rect 28142 20638 28194 20690
rect 29150 20638 29202 20690
rect 29934 20638 29986 20690
rect 36990 20638 37042 20690
rect 39566 20638 39618 20690
rect 39902 20638 39954 20690
rect 40350 20638 40402 20690
rect 40910 20638 40962 20690
rect 45502 20638 45554 20690
rect 46398 20638 46450 20690
rect 47070 20638 47122 20690
rect 52782 20638 52834 20690
rect 1710 20526 1762 20578
rect 3390 20526 3442 20578
rect 3502 20526 3554 20578
rect 5966 20526 6018 20578
rect 6974 20526 7026 20578
rect 7534 20526 7586 20578
rect 10334 20526 10386 20578
rect 27134 20526 27186 20578
rect 28590 20526 28642 20578
rect 29486 20526 29538 20578
rect 29822 20526 29874 20578
rect 35198 20526 35250 20578
rect 35310 20526 35362 20578
rect 36542 20526 36594 20578
rect 40126 20526 40178 20578
rect 41022 20526 41074 20578
rect 41134 20526 41186 20578
rect 42702 20526 42754 20578
rect 43710 20526 43762 20578
rect 47406 20526 47458 20578
rect 47854 20526 47906 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 4846 20190 4898 20242
rect 11230 20190 11282 20242
rect 11678 20190 11730 20242
rect 14478 20190 14530 20242
rect 19406 20190 19458 20242
rect 19742 20190 19794 20242
rect 38558 20190 38610 20242
rect 38894 20190 38946 20242
rect 39006 20190 39058 20242
rect 41022 20190 41074 20242
rect 2494 20078 2546 20130
rect 5070 20078 5122 20130
rect 5182 20078 5234 20130
rect 6078 20078 6130 20130
rect 6414 20078 6466 20130
rect 6750 20078 6802 20130
rect 7310 20078 7362 20130
rect 7422 20078 7474 20130
rect 8654 20078 8706 20130
rect 8878 20078 8930 20130
rect 12014 20078 12066 20130
rect 12462 20078 12514 20130
rect 13246 20078 13298 20130
rect 13582 20078 13634 20130
rect 17950 20078 18002 20130
rect 18398 20078 18450 20130
rect 24110 20078 24162 20130
rect 26686 20078 26738 20130
rect 28254 20078 28306 20130
rect 31950 20078 32002 20130
rect 32062 20078 32114 20130
rect 34974 20078 35026 20130
rect 39790 20078 39842 20130
rect 39902 20078 39954 20130
rect 46286 20078 46338 20130
rect 46622 20078 46674 20130
rect 48862 20078 48914 20130
rect 50206 20078 50258 20130
rect 51550 20078 51602 20130
rect 1822 19966 1874 20018
rect 7086 19966 7138 20018
rect 7758 19966 7810 20018
rect 7982 19966 8034 20018
rect 8990 19966 9042 20018
rect 9550 19966 9602 20018
rect 9774 19966 9826 20018
rect 10110 19966 10162 20018
rect 11006 19966 11058 20018
rect 12686 19966 12738 20018
rect 14702 19966 14754 20018
rect 21198 19966 21250 20018
rect 25790 19966 25842 20018
rect 26462 19966 26514 20018
rect 28142 19966 28194 20018
rect 29710 19966 29762 20018
rect 31054 19966 31106 20018
rect 34862 19966 34914 20018
rect 35870 19966 35922 20018
rect 36318 19966 36370 20018
rect 38782 19966 38834 20018
rect 39230 19966 39282 20018
rect 39566 19966 39618 20018
rect 43150 19966 43202 20018
rect 47294 19966 47346 20018
rect 47854 19966 47906 20018
rect 50878 19966 50930 20018
rect 51102 19966 51154 20018
rect 52222 19966 52274 20018
rect 52446 19966 52498 20018
rect 4622 19854 4674 19906
rect 5630 19854 5682 19906
rect 18958 19854 19010 19906
rect 20302 19854 20354 19906
rect 21870 19854 21922 19906
rect 23662 19854 23714 19906
rect 29374 19854 29426 19906
rect 36766 19854 36818 19906
rect 37214 19854 37266 19906
rect 37662 19854 37714 19906
rect 38110 19854 38162 19906
rect 40238 19854 40290 19906
rect 41470 19854 41522 19906
rect 42254 19854 42306 19906
rect 44942 19854 44994 19906
rect 53902 19854 53954 19906
rect 5518 19742 5570 19794
rect 6190 19742 6242 19794
rect 8094 19742 8146 19794
rect 11342 19742 11394 19794
rect 14366 19742 14418 19794
rect 23550 19742 23602 19794
rect 32062 19742 32114 19794
rect 34974 19742 35026 19794
rect 37214 19742 37266 19794
rect 37662 19742 37714 19794
rect 42142 19742 42194 19794
rect 45614 19742 45666 19794
rect 45950 19742 46002 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 10558 19406 10610 19458
rect 15374 19406 15426 19458
rect 26350 19406 26402 19458
rect 39342 19406 39394 19458
rect 40014 19406 40066 19458
rect 41470 19406 41522 19458
rect 41918 19406 41970 19458
rect 4062 19294 4114 19346
rect 6526 19294 6578 19346
rect 8430 19294 8482 19346
rect 10670 19294 10722 19346
rect 12910 19294 12962 19346
rect 17614 19294 17666 19346
rect 22318 19294 22370 19346
rect 24446 19294 24498 19346
rect 25230 19294 25282 19346
rect 26014 19294 26066 19346
rect 26910 19294 26962 19346
rect 28366 19294 28418 19346
rect 29486 19294 29538 19346
rect 31278 19294 31330 19346
rect 35310 19294 35362 19346
rect 38558 19294 38610 19346
rect 39118 19294 39170 19346
rect 41022 19294 41074 19346
rect 41470 19294 41522 19346
rect 43150 19294 43202 19346
rect 43710 19294 43762 19346
rect 44046 19294 44098 19346
rect 46174 19294 46226 19346
rect 47854 19294 47906 19346
rect 49982 19294 50034 19346
rect 1710 19182 1762 19234
rect 3390 19182 3442 19234
rect 3838 19182 3890 19234
rect 4174 19182 4226 19234
rect 5070 19182 5122 19234
rect 6078 19182 6130 19234
rect 7534 19182 7586 19234
rect 9886 19182 9938 19234
rect 13582 19182 13634 19234
rect 16046 19182 16098 19234
rect 17950 19182 18002 19234
rect 18174 19182 18226 19234
rect 18622 19182 18674 19234
rect 19966 19182 20018 19234
rect 21646 19182 21698 19234
rect 25678 19182 25730 19234
rect 28030 19182 28082 19234
rect 28590 19182 28642 19234
rect 29374 19182 29426 19234
rect 29710 19182 29762 19234
rect 31614 19182 31666 19234
rect 32286 19182 32338 19234
rect 32846 19182 32898 19234
rect 33294 19182 33346 19234
rect 33518 19182 33570 19234
rect 35758 19182 35810 19234
rect 37438 19182 37490 19234
rect 37886 19182 37938 19234
rect 38110 19182 38162 19234
rect 42142 19182 42194 19234
rect 43486 19182 43538 19234
rect 45166 19182 45218 19234
rect 47070 19182 47122 19234
rect 53678 19182 53730 19234
rect 53902 19182 53954 19234
rect 2382 19070 2434 19122
rect 2718 19070 2770 19122
rect 4510 19070 4562 19122
rect 5630 19070 5682 19122
rect 13694 19070 13746 19122
rect 14142 19070 14194 19122
rect 14478 19070 14530 19122
rect 14590 19070 14642 19122
rect 15710 19070 15762 19122
rect 17278 19070 17330 19122
rect 20750 19070 20802 19122
rect 26126 19070 26178 19122
rect 32398 19070 32450 19122
rect 36206 19070 36258 19122
rect 42702 19070 42754 19122
rect 53454 19070 53506 19122
rect 54574 19070 54626 19122
rect 2046 18958 2098 19010
rect 3614 18958 3666 19010
rect 4734 18958 4786 19010
rect 4958 18958 5010 19010
rect 10222 18958 10274 19010
rect 11118 18958 11170 19010
rect 13806 18958 13858 19010
rect 13918 18958 13970 19010
rect 15486 18958 15538 19010
rect 16158 18958 16210 19010
rect 16382 18958 16434 19010
rect 17502 18958 17554 19010
rect 18398 18958 18450 19010
rect 18958 18958 19010 19010
rect 19406 18958 19458 19010
rect 19742 18958 19794 19010
rect 20414 18958 20466 19010
rect 27246 18958 27298 19010
rect 29038 18958 29090 19010
rect 31838 18958 31890 19010
rect 32510 18958 32562 19010
rect 32958 18958 33010 19010
rect 33070 18958 33122 19010
rect 37102 18958 37154 19010
rect 37998 18958 38050 19010
rect 39566 18958 39618 19010
rect 40014 18958 40066 19010
rect 40462 18958 40514 19010
rect 43934 18958 43986 19010
rect 44158 18958 44210 19010
rect 45390 18958 45442 19010
rect 50430 18958 50482 19010
rect 53342 18958 53394 19010
rect 53566 18958 53618 19010
rect 54238 18958 54290 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 2718 18622 2770 18674
rect 3166 18622 3218 18674
rect 3614 18622 3666 18674
rect 5182 18622 5234 18674
rect 7870 18622 7922 18674
rect 8878 18622 8930 18674
rect 9998 18622 10050 18674
rect 15038 18622 15090 18674
rect 18958 18622 19010 18674
rect 19182 18622 19234 18674
rect 20862 18622 20914 18674
rect 21086 18622 21138 18674
rect 22094 18622 22146 18674
rect 22318 18622 22370 18674
rect 26798 18622 26850 18674
rect 36654 18622 36706 18674
rect 39902 18622 39954 18674
rect 42366 18622 42418 18674
rect 43038 18622 43090 18674
rect 43934 18622 43986 18674
rect 2046 18510 2098 18562
rect 5854 18510 5906 18562
rect 6078 18510 6130 18562
rect 8990 18510 9042 18562
rect 10334 18510 10386 18562
rect 21422 18510 21474 18562
rect 25790 18510 25842 18562
rect 28478 18510 28530 18562
rect 31614 18510 31666 18562
rect 32062 18510 32114 18562
rect 32286 18510 32338 18562
rect 36766 18510 36818 18562
rect 37886 18510 37938 18562
rect 38222 18510 38274 18562
rect 38334 18510 38386 18562
rect 44158 18510 44210 18562
rect 44270 18510 44322 18562
rect 44718 18510 44770 18562
rect 46062 18510 46114 18562
rect 1710 18398 1762 18450
rect 3838 18398 3890 18450
rect 4286 18398 4338 18450
rect 4398 18398 4450 18450
rect 6974 18398 7026 18450
rect 8094 18398 8146 18450
rect 8430 18398 8482 18450
rect 11342 18398 11394 18450
rect 11678 18398 11730 18450
rect 12462 18398 12514 18450
rect 14926 18398 14978 18450
rect 15822 18398 15874 18450
rect 16382 18398 16434 18450
rect 16494 18398 16546 18450
rect 17278 18398 17330 18450
rect 18062 18398 18114 18450
rect 18286 18398 18338 18450
rect 19630 18398 19682 18450
rect 21982 18398 22034 18450
rect 22206 18398 22258 18450
rect 22430 18398 22482 18450
rect 24222 18398 24274 18450
rect 24670 18398 24722 18450
rect 25230 18398 25282 18450
rect 25454 18398 25506 18450
rect 26350 18398 26402 18450
rect 26574 18398 26626 18450
rect 26686 18398 26738 18450
rect 27022 18398 27074 18450
rect 29374 18398 29426 18450
rect 29934 18398 29986 18450
rect 30942 18398 30994 18450
rect 31390 18398 31442 18450
rect 33070 18398 33122 18450
rect 33294 18398 33346 18450
rect 33630 18398 33682 18450
rect 36430 18398 36482 18450
rect 36878 18398 36930 18450
rect 37326 18398 37378 18450
rect 37550 18398 37602 18450
rect 38558 18398 38610 18450
rect 39230 18398 39282 18450
rect 39678 18398 39730 18450
rect 40350 18398 40402 18450
rect 42478 18398 42530 18450
rect 45390 18398 45442 18450
rect 48862 18398 48914 18450
rect 51998 18398 52050 18450
rect 55246 18398 55298 18450
rect 4062 18286 4114 18338
rect 5070 18286 5122 18338
rect 5742 18286 5794 18338
rect 6526 18286 6578 18338
rect 7422 18286 7474 18338
rect 7982 18286 8034 18338
rect 14590 18286 14642 18338
rect 18398 18286 18450 18338
rect 19070 18286 19122 18338
rect 23886 18286 23938 18338
rect 25342 18286 25394 18338
rect 27470 18286 27522 18338
rect 28030 18286 28082 18338
rect 29822 18286 29874 18338
rect 31950 18286 32002 18338
rect 33182 18286 33234 18338
rect 39790 18286 39842 18338
rect 43486 18286 43538 18338
rect 48190 18286 48242 18338
rect 52334 18286 52386 18338
rect 54462 18286 54514 18338
rect 5406 18174 5458 18226
rect 8878 18174 8930 18226
rect 15038 18174 15090 18226
rect 28030 18174 28082 18226
rect 28254 18174 28306 18226
rect 28926 18174 28978 18226
rect 42366 18174 42418 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 5518 17838 5570 17890
rect 6526 17838 6578 17890
rect 6862 17838 6914 17890
rect 33518 17838 33570 17890
rect 37438 17838 37490 17890
rect 42814 17838 42866 17890
rect 53566 17838 53618 17890
rect 4622 17726 4674 17778
rect 5070 17726 5122 17778
rect 5854 17726 5906 17778
rect 7646 17726 7698 17778
rect 11342 17726 11394 17778
rect 13694 17726 13746 17778
rect 15262 17726 15314 17778
rect 16494 17726 16546 17778
rect 17390 17726 17442 17778
rect 19518 17726 19570 17778
rect 20862 17726 20914 17778
rect 22094 17726 22146 17778
rect 24222 17726 24274 17778
rect 27022 17726 27074 17778
rect 32622 17726 32674 17778
rect 40350 17726 40402 17778
rect 42478 17726 42530 17778
rect 43598 17726 43650 17778
rect 44046 17726 44098 17778
rect 47630 17726 47682 17778
rect 49758 17726 49810 17778
rect 51214 17726 51266 17778
rect 51662 17726 51714 17778
rect 53454 17726 53506 17778
rect 1822 17614 1874 17666
rect 6190 17614 6242 17666
rect 8318 17614 8370 17666
rect 8878 17614 8930 17666
rect 9326 17614 9378 17666
rect 14030 17614 14082 17666
rect 14590 17614 14642 17666
rect 15934 17614 15986 17666
rect 20302 17614 20354 17666
rect 21422 17614 21474 17666
rect 25230 17614 25282 17666
rect 25566 17614 25618 17666
rect 25678 17614 25730 17666
rect 26126 17614 26178 17666
rect 26574 17614 26626 17666
rect 27582 17614 27634 17666
rect 28142 17614 28194 17666
rect 28366 17614 28418 17666
rect 29374 17614 29426 17666
rect 29822 17614 29874 17666
rect 30158 17614 30210 17666
rect 30270 17614 30322 17666
rect 31054 17614 31106 17666
rect 32398 17614 32450 17666
rect 33070 17614 33122 17666
rect 33294 17614 33346 17666
rect 37886 17614 37938 17666
rect 38222 17614 38274 17666
rect 38558 17614 38610 17666
rect 39230 17614 39282 17666
rect 39678 17614 39730 17666
rect 45614 17614 45666 17666
rect 46510 17614 46562 17666
rect 50766 17614 50818 17666
rect 2494 17502 2546 17554
rect 6974 17502 7026 17554
rect 7310 17502 7362 17554
rect 7534 17502 7586 17554
rect 7758 17502 7810 17554
rect 8094 17502 8146 17554
rect 10782 17502 10834 17554
rect 17054 17502 17106 17554
rect 27246 17502 27298 17554
rect 28590 17502 28642 17554
rect 29150 17502 29202 17554
rect 31726 17502 31778 17554
rect 37550 17502 37602 17554
rect 42926 17502 42978 17554
rect 43150 17502 43202 17554
rect 45278 17502 45330 17554
rect 45950 17502 46002 17554
rect 46174 17502 46226 17554
rect 51214 17502 51266 17554
rect 6862 17390 6914 17442
rect 9438 17390 9490 17442
rect 9886 17390 9938 17442
rect 10222 17390 10274 17442
rect 15598 17390 15650 17442
rect 16718 17390 16770 17442
rect 27470 17390 27522 17442
rect 28478 17390 28530 17442
rect 29262 17390 29314 17442
rect 30046 17390 30098 17442
rect 30494 17390 30546 17442
rect 31278 17390 31330 17442
rect 33966 17390 34018 17442
rect 34750 17390 34802 17442
rect 35086 17390 35138 17442
rect 36430 17390 36482 17442
rect 37438 17390 37490 17442
rect 37998 17390 38050 17442
rect 39006 17390 39058 17442
rect 39118 17390 39170 17442
rect 45166 17390 45218 17442
rect 45726 17390 45778 17442
rect 50878 17390 50930 17442
rect 51102 17390 51154 17442
rect 51774 17390 51826 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 1710 17054 1762 17106
rect 3166 17054 3218 17106
rect 3614 17054 3666 17106
rect 4286 17054 4338 17106
rect 11342 17054 11394 17106
rect 13358 17054 13410 17106
rect 19070 17054 19122 17106
rect 20078 17054 20130 17106
rect 20414 17054 20466 17106
rect 20750 17054 20802 17106
rect 25790 17054 25842 17106
rect 26686 17054 26738 17106
rect 26798 17054 26850 17106
rect 28254 17054 28306 17106
rect 37774 17054 37826 17106
rect 41694 17054 41746 17106
rect 42366 17054 42418 17106
rect 43486 17054 43538 17106
rect 46062 17054 46114 17106
rect 47070 17054 47122 17106
rect 47294 17054 47346 17106
rect 47966 17054 48018 17106
rect 2046 16942 2098 16994
rect 2718 16942 2770 16994
rect 4174 16942 4226 16994
rect 5630 16942 5682 16994
rect 9886 16942 9938 16994
rect 11678 16942 11730 16994
rect 13022 16942 13074 16994
rect 13134 16942 13186 16994
rect 15038 16942 15090 16994
rect 16270 16942 16322 16994
rect 18846 16942 18898 16994
rect 22878 16942 22930 16994
rect 24670 16942 24722 16994
rect 29486 16942 29538 16994
rect 30270 16942 30322 16994
rect 31054 16942 31106 16994
rect 39454 16942 39506 16994
rect 42142 16942 42194 16994
rect 42814 16942 42866 16994
rect 44046 16942 44098 16994
rect 44606 16942 44658 16994
rect 47742 16942 47794 16994
rect 48750 16942 48802 16994
rect 52222 16942 52274 16994
rect 2382 16830 2434 16882
rect 3278 16830 3330 16882
rect 3390 16830 3442 16882
rect 4062 16830 4114 16882
rect 5070 16830 5122 16882
rect 8654 16830 8706 16882
rect 10110 16830 10162 16882
rect 14366 16830 14418 16882
rect 14814 16830 14866 16882
rect 16158 16830 16210 16882
rect 18734 16830 18786 16882
rect 21198 16830 21250 16882
rect 24334 16830 24386 16882
rect 25566 16830 25618 16882
rect 26910 16830 26962 16882
rect 27246 16830 27298 16882
rect 28926 16830 28978 16882
rect 29374 16830 29426 16882
rect 34414 16830 34466 16882
rect 35198 16830 35250 16882
rect 42030 16830 42082 16882
rect 45166 16830 45218 16882
rect 45950 16830 46002 16882
rect 46734 16830 46786 16882
rect 47630 16830 47682 16882
rect 49422 16830 49474 16882
rect 53006 16830 53058 16882
rect 6638 16718 6690 16770
rect 14926 16718 14978 16770
rect 37326 16718 37378 16770
rect 42926 16718 42978 16770
rect 43262 16718 43314 16770
rect 44942 16718 44994 16770
rect 47182 16718 47234 16770
rect 49198 16718 49250 16770
rect 50094 16718 50146 16770
rect 16270 16606 16322 16658
rect 28590 16606 28642 16658
rect 42590 16606 42642 16658
rect 43598 16606 43650 16658
rect 46062 16606 46114 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 8766 16270 8818 16322
rect 9102 16270 9154 16322
rect 10782 16270 10834 16322
rect 17166 16270 17218 16322
rect 24670 16270 24722 16322
rect 25118 16270 25170 16322
rect 25790 16270 25842 16322
rect 26798 16270 26850 16322
rect 33070 16270 33122 16322
rect 43710 16270 43762 16322
rect 46510 16270 46562 16322
rect 48750 16270 48802 16322
rect 49086 16270 49138 16322
rect 4622 16158 4674 16210
rect 5070 16158 5122 16210
rect 9662 16158 9714 16210
rect 11118 16158 11170 16210
rect 12686 16158 12738 16210
rect 14702 16158 14754 16210
rect 15038 16158 15090 16210
rect 24334 16158 24386 16210
rect 25118 16158 25170 16210
rect 25678 16158 25730 16210
rect 27358 16158 27410 16210
rect 28366 16158 28418 16210
rect 35646 16158 35698 16210
rect 38222 16158 38274 16210
rect 39790 16158 39842 16210
rect 41918 16158 41970 16210
rect 45054 16158 45106 16210
rect 46734 16158 46786 16210
rect 47070 16158 47122 16210
rect 48414 16158 48466 16210
rect 49646 16158 49698 16210
rect 50094 16158 50146 16210
rect 1822 16046 1874 16098
rect 6750 16046 6802 16098
rect 6974 16046 7026 16098
rect 7870 16046 7922 16098
rect 8094 16046 8146 16098
rect 11790 16046 11842 16098
rect 12126 16046 12178 16098
rect 12350 16046 12402 16098
rect 14590 16046 14642 16098
rect 15262 16046 15314 16098
rect 16718 16046 16770 16098
rect 17614 16046 17666 16098
rect 17838 16046 17890 16098
rect 18062 16046 18114 16098
rect 21982 16046 22034 16098
rect 22206 16046 22258 16098
rect 22990 16046 23042 16098
rect 23662 16046 23714 16098
rect 26350 16046 26402 16098
rect 26574 16046 26626 16098
rect 31838 16046 31890 16098
rect 32062 16046 32114 16098
rect 32286 16046 32338 16098
rect 33182 16046 33234 16098
rect 34750 16046 34802 16098
rect 35534 16046 35586 16098
rect 35758 16046 35810 16098
rect 39118 16046 39170 16098
rect 42926 16046 42978 16098
rect 43262 16046 43314 16098
rect 45390 16046 45442 16098
rect 47182 16046 47234 16098
rect 47518 16046 47570 16098
rect 49198 16046 49250 16098
rect 50654 16046 50706 16098
rect 50766 16046 50818 16098
rect 2494 15934 2546 15986
rect 6190 15934 6242 15986
rect 6526 15934 6578 15986
rect 11454 15934 11506 15986
rect 13694 15934 13746 15986
rect 14030 15934 14082 15986
rect 15934 15934 15986 15986
rect 16830 15934 16882 15986
rect 22430 15934 22482 15986
rect 22766 15934 22818 15986
rect 24558 15934 24610 15986
rect 26126 15934 26178 15986
rect 27694 15934 27746 15986
rect 27806 15934 27858 15986
rect 32734 15934 32786 15986
rect 33070 15934 33122 15986
rect 33854 15934 33906 15986
rect 35198 15934 35250 15986
rect 36990 15934 37042 15986
rect 37550 15934 37602 15986
rect 37886 15934 37938 15986
rect 43374 15934 43426 15986
rect 43934 15934 43986 15986
rect 50990 15934 51042 15986
rect 51550 15934 51602 15986
rect 53454 15934 53506 15986
rect 5966 15822 6018 15874
rect 6078 15822 6130 15874
rect 7982 15822 8034 15874
rect 8318 15822 8370 15874
rect 8990 15822 9042 15874
rect 11006 15822 11058 15874
rect 11790 15822 11842 15874
rect 12574 15822 12626 15874
rect 17054 15822 17106 15874
rect 21870 15822 21922 15874
rect 22094 15822 22146 15874
rect 28030 15822 28082 15874
rect 34078 15822 34130 15874
rect 34190 15822 34242 15874
rect 34302 15822 34354 15874
rect 35982 15822 36034 15874
rect 37102 15822 37154 15874
rect 37326 15822 37378 15874
rect 37662 15822 37714 15874
rect 43822 15822 43874 15874
rect 45502 15822 45554 15874
rect 45726 15822 45778 15874
rect 46174 15822 46226 15874
rect 48526 15822 48578 15874
rect 49534 15822 49586 15874
rect 50878 15822 50930 15874
rect 51102 15822 51154 15874
rect 51662 15822 51714 15874
rect 52782 15822 52834 15874
rect 53118 15822 53170 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 2718 15486 2770 15538
rect 3166 15486 3218 15538
rect 3278 15486 3330 15538
rect 4734 15486 4786 15538
rect 4958 15486 5010 15538
rect 5518 15486 5570 15538
rect 8990 15486 9042 15538
rect 10446 15486 10498 15538
rect 16830 15486 16882 15538
rect 24446 15486 24498 15538
rect 32510 15486 32562 15538
rect 35982 15486 36034 15538
rect 38222 15486 38274 15538
rect 38334 15486 38386 15538
rect 39230 15486 39282 15538
rect 41246 15486 41298 15538
rect 42030 15486 42082 15538
rect 44158 15486 44210 15538
rect 44718 15486 44770 15538
rect 45614 15486 45666 15538
rect 45838 15486 45890 15538
rect 47966 15486 48018 15538
rect 1710 15374 1762 15426
rect 2046 15374 2098 15426
rect 2382 15374 2434 15426
rect 8094 15374 8146 15426
rect 8206 15374 8258 15426
rect 8654 15374 8706 15426
rect 13470 15374 13522 15426
rect 19294 15374 19346 15426
rect 19630 15374 19682 15426
rect 23662 15374 23714 15426
rect 23998 15374 24050 15426
rect 27582 15374 27634 15426
rect 28814 15374 28866 15426
rect 29038 15374 29090 15426
rect 32286 15374 32338 15426
rect 33070 15374 33122 15426
rect 38446 15374 38498 15426
rect 39006 15374 39058 15426
rect 42254 15374 42306 15426
rect 46958 15374 47010 15426
rect 47182 15374 47234 15426
rect 47742 15374 47794 15426
rect 48078 15374 48130 15426
rect 49422 15374 49474 15426
rect 49646 15374 49698 15426
rect 52558 15374 52610 15426
rect 3054 15262 3106 15314
rect 3726 15262 3778 15314
rect 3838 15262 3890 15314
rect 4062 15262 4114 15314
rect 4174 15262 4226 15314
rect 4510 15262 4562 15314
rect 5070 15262 5122 15314
rect 7086 15262 7138 15314
rect 7534 15262 7586 15314
rect 9438 15262 9490 15314
rect 9886 15262 9938 15314
rect 10110 15262 10162 15314
rect 10670 15262 10722 15314
rect 11342 15262 11394 15314
rect 11678 15262 11730 15314
rect 12798 15262 12850 15314
rect 13022 15262 13074 15314
rect 13134 15262 13186 15314
rect 13806 15262 13858 15314
rect 14030 15262 14082 15314
rect 14366 15262 14418 15314
rect 14702 15262 14754 15314
rect 14926 15262 14978 15314
rect 15150 15262 15202 15314
rect 16158 15262 16210 15314
rect 16606 15262 16658 15314
rect 17838 15262 17890 15314
rect 19070 15262 19122 15314
rect 20526 15262 20578 15314
rect 26910 15262 26962 15314
rect 27918 15262 27970 15314
rect 28478 15262 28530 15314
rect 31054 15262 31106 15314
rect 31838 15262 31890 15314
rect 33294 15262 33346 15314
rect 33518 15262 33570 15314
rect 34526 15262 34578 15314
rect 34974 15262 35026 15314
rect 35870 15262 35922 15314
rect 36206 15262 36258 15314
rect 36990 15262 37042 15314
rect 37326 15262 37378 15314
rect 38894 15262 38946 15314
rect 39342 15262 39394 15314
rect 42926 15262 42978 15314
rect 43150 15262 43202 15314
rect 43598 15262 43650 15314
rect 43822 15262 43874 15314
rect 44494 15262 44546 15314
rect 44606 15262 44658 15314
rect 45166 15262 45218 15314
rect 45390 15262 45442 15314
rect 46510 15262 46562 15314
rect 46622 15262 46674 15314
rect 47294 15262 47346 15314
rect 47518 15262 47570 15314
rect 49870 15262 49922 15314
rect 50094 15262 50146 15314
rect 53230 15262 53282 15314
rect 5966 15150 6018 15202
rect 6638 15150 6690 15202
rect 9998 15150 10050 15202
rect 11118 15150 11170 15202
rect 14254 15150 14306 15202
rect 15598 15150 15650 15202
rect 16718 15150 16770 15202
rect 17614 15150 17666 15202
rect 18510 15150 18562 15202
rect 19518 15150 19570 15202
rect 21198 15150 21250 15202
rect 23326 15150 23378 15202
rect 26798 15150 26850 15202
rect 29150 15150 29202 15202
rect 31166 15150 31218 15202
rect 32398 15150 32450 15202
rect 35422 15150 35474 15202
rect 37438 15150 37490 15202
rect 45502 15150 45554 15202
rect 49758 15150 49810 15202
rect 50430 15150 50482 15202
rect 8094 15038 8146 15090
rect 30606 15038 30658 15090
rect 33742 15038 33794 15090
rect 34190 15038 34242 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 4398 14702 4450 14754
rect 4958 14702 5010 14754
rect 6302 14702 6354 14754
rect 8430 14702 8482 14754
rect 9774 14702 9826 14754
rect 19070 14702 19122 14754
rect 21534 14702 21586 14754
rect 27694 14702 27746 14754
rect 28030 14702 28082 14754
rect 34302 14702 34354 14754
rect 45614 14702 45666 14754
rect 46846 14702 46898 14754
rect 47182 14702 47234 14754
rect 3166 14590 3218 14642
rect 3614 14590 3666 14642
rect 4622 14590 4674 14642
rect 5966 14590 6018 14642
rect 7534 14590 7586 14642
rect 10110 14590 10162 14642
rect 11790 14590 11842 14642
rect 13806 14590 13858 14642
rect 14926 14590 14978 14642
rect 16270 14590 16322 14642
rect 17502 14590 17554 14642
rect 21646 14590 21698 14642
rect 23214 14590 23266 14642
rect 25342 14590 25394 14642
rect 25902 14590 25954 14642
rect 31614 14590 31666 14642
rect 32622 14590 32674 14642
rect 33182 14590 33234 14642
rect 38670 14590 38722 14642
rect 40798 14590 40850 14642
rect 42030 14590 42082 14642
rect 42926 14590 42978 14642
rect 43822 14590 43874 14642
rect 45054 14590 45106 14642
rect 45278 14590 45330 14642
rect 48526 14590 48578 14642
rect 48862 14590 48914 14642
rect 1710 14478 1762 14530
rect 2494 14478 2546 14530
rect 4174 14478 4226 14530
rect 5070 14478 5122 14530
rect 6638 14478 6690 14530
rect 7310 14478 7362 14530
rect 7758 14478 7810 14530
rect 7982 14478 8034 14530
rect 9438 14478 9490 14530
rect 9774 14478 9826 14530
rect 11006 14478 11058 14530
rect 11902 14478 11954 14530
rect 13918 14478 13970 14530
rect 14814 14478 14866 14530
rect 16382 14478 16434 14530
rect 17950 14478 18002 14530
rect 18734 14478 18786 14530
rect 19742 14478 19794 14530
rect 22430 14478 22482 14530
rect 26350 14478 26402 14530
rect 26574 14478 26626 14530
rect 26686 14478 26738 14530
rect 26910 14478 26962 14530
rect 31166 14478 31218 14530
rect 33294 14478 33346 14530
rect 34750 14478 34802 14530
rect 34974 14478 35026 14530
rect 35198 14478 35250 14530
rect 35758 14478 35810 14530
rect 37214 14478 37266 14530
rect 37662 14478 37714 14530
rect 37886 14478 37938 14530
rect 41358 14478 41410 14530
rect 42254 14478 42306 14530
rect 43374 14478 43426 14530
rect 45614 14478 45666 14530
rect 51662 14478 51714 14530
rect 2046 14366 2098 14418
rect 2718 14366 2770 14418
rect 4062 14366 4114 14418
rect 6078 14366 6130 14418
rect 12574 14366 12626 14418
rect 13470 14366 13522 14418
rect 17054 14366 17106 14418
rect 18398 14366 18450 14418
rect 18958 14366 19010 14418
rect 19406 14366 19458 14418
rect 26014 14366 26066 14418
rect 26798 14366 26850 14418
rect 27806 14366 27858 14418
rect 30718 14366 30770 14418
rect 32846 14366 32898 14418
rect 35422 14366 35474 14418
rect 36206 14366 36258 14418
rect 41470 14366 41522 14418
rect 46622 14366 46674 14418
rect 50990 14366 51042 14418
rect 3838 14254 3890 14306
rect 6750 14254 6802 14306
rect 6862 14254 6914 14306
rect 11118 14254 11170 14306
rect 11342 14254 11394 14306
rect 15038 14254 15090 14306
rect 19518 14254 19570 14306
rect 22094 14254 22146 14306
rect 35870 14254 35922 14306
rect 35982 14254 36034 14306
rect 36990 14254 37042 14306
rect 37102 14254 37154 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 13022 13918 13074 13970
rect 18510 13918 18562 13970
rect 24670 13918 24722 13970
rect 25566 13918 25618 13970
rect 26014 13918 26066 13970
rect 28926 13918 28978 13970
rect 30942 13918 30994 13970
rect 33406 13918 33458 13970
rect 34974 13918 35026 13970
rect 37662 13918 37714 13970
rect 37774 13918 37826 13970
rect 37886 13918 37938 13970
rect 38782 13918 38834 13970
rect 39454 13918 39506 13970
rect 40014 13918 40066 13970
rect 43486 13918 43538 13970
rect 44830 13918 44882 13970
rect 45950 13918 46002 13970
rect 46174 13918 46226 13970
rect 47070 13918 47122 13970
rect 49422 13918 49474 13970
rect 49758 13918 49810 13970
rect 50878 13918 50930 13970
rect 5294 13806 5346 13858
rect 5518 13806 5570 13858
rect 7646 13806 7698 13858
rect 13134 13806 13186 13858
rect 18286 13806 18338 13858
rect 27134 13806 27186 13858
rect 27694 13806 27746 13858
rect 28366 13806 28418 13858
rect 29374 13806 29426 13858
rect 33294 13806 33346 13858
rect 39566 13806 39618 13858
rect 41134 13806 41186 13858
rect 41582 13806 41634 13858
rect 42702 13806 42754 13858
rect 46510 13806 46562 13858
rect 47294 13806 47346 13858
rect 47518 13806 47570 13858
rect 50094 13806 50146 13858
rect 50766 13806 50818 13858
rect 1822 13694 1874 13746
rect 4958 13694 5010 13746
rect 6974 13694 7026 13746
rect 7198 13694 7250 13746
rect 7870 13694 7922 13746
rect 8430 13694 8482 13746
rect 9998 13694 10050 13746
rect 13806 13694 13858 13746
rect 14254 13694 14306 13746
rect 22206 13694 22258 13746
rect 26014 13694 26066 13746
rect 26462 13694 26514 13746
rect 26798 13694 26850 13746
rect 27470 13694 27522 13746
rect 31166 13694 31218 13746
rect 31726 13694 31778 13746
rect 34078 13694 34130 13746
rect 34526 13694 34578 13746
rect 36206 13694 36258 13746
rect 36654 13694 36706 13746
rect 36766 13694 36818 13746
rect 37326 13694 37378 13746
rect 38334 13694 38386 13746
rect 38558 13694 38610 13746
rect 38894 13694 38946 13746
rect 42590 13694 42642 13746
rect 43486 13694 43538 13746
rect 44046 13694 44098 13746
rect 44270 13694 44322 13746
rect 44606 13694 44658 13746
rect 46846 13694 46898 13746
rect 50318 13694 50370 13746
rect 2494 13582 2546 13634
rect 4622 13582 4674 13634
rect 5070 13582 5122 13634
rect 6302 13582 6354 13634
rect 7982 13582 8034 13634
rect 9550 13582 9602 13634
rect 10334 13582 10386 13634
rect 14478 13582 14530 13634
rect 17390 13582 17442 13634
rect 17950 13582 18002 13634
rect 18398 13582 18450 13634
rect 19406 13582 19458 13634
rect 21534 13582 21586 13634
rect 22766 13582 22818 13634
rect 26686 13582 26738 13634
rect 28254 13582 28306 13634
rect 38110 13582 38162 13634
rect 47182 13582 47234 13634
rect 49086 13582 49138 13634
rect 8206 13470 8258 13522
rect 13022 13470 13074 13522
rect 17614 13470 17666 13522
rect 27806 13470 27858 13522
rect 28142 13470 28194 13522
rect 33406 13470 33458 13522
rect 34302 13470 34354 13522
rect 39454 13470 39506 13522
rect 41806 13470 41858 13522
rect 42142 13470 42194 13522
rect 44606 13470 44658 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 13470 13134 13522 13186
rect 25006 13134 25058 13186
rect 26238 13134 26290 13186
rect 27582 13134 27634 13186
rect 27806 13134 27858 13186
rect 41134 13134 41186 13186
rect 44270 13134 44322 13186
rect 3390 13022 3442 13074
rect 6638 13022 6690 13074
rect 7982 13022 8034 13074
rect 16830 13022 16882 13074
rect 20190 13022 20242 13074
rect 23886 13022 23938 13074
rect 26126 13022 26178 13074
rect 29934 13022 29986 13074
rect 37438 13022 37490 13074
rect 40686 13022 40738 13074
rect 41806 13022 41858 13074
rect 46958 13022 47010 13074
rect 1710 12910 1762 12962
rect 2382 12910 2434 12962
rect 3278 12910 3330 12962
rect 3838 12910 3890 12962
rect 4398 12910 4450 12962
rect 5742 12910 5794 12962
rect 6414 12910 6466 12962
rect 7758 12910 7810 12962
rect 10894 12910 10946 12962
rect 18846 12910 18898 12962
rect 19406 12910 19458 12962
rect 19630 12910 19682 12962
rect 20302 12910 20354 12962
rect 24334 12910 24386 12962
rect 25342 12910 25394 12962
rect 26686 12910 26738 12962
rect 26910 12910 26962 12962
rect 27022 12910 27074 12962
rect 27246 12910 27298 12962
rect 28142 12910 28194 12962
rect 28366 12910 28418 12962
rect 29150 12910 29202 12962
rect 29374 12910 29426 12962
rect 30942 12910 30994 12962
rect 31614 12910 31666 12962
rect 33854 12910 33906 12962
rect 38782 12910 38834 12962
rect 42142 12910 42194 12962
rect 42366 12910 42418 12962
rect 42590 12910 42642 12962
rect 43038 12910 43090 12962
rect 43374 12910 43426 12962
rect 2718 12798 2770 12850
rect 4286 12798 4338 12850
rect 4846 12798 4898 12850
rect 7086 12798 7138 12850
rect 8430 12798 8482 12850
rect 19182 12798 19234 12850
rect 24110 12798 24162 12850
rect 24670 12798 24722 12850
rect 25118 12798 25170 12850
rect 31390 12798 31442 12850
rect 31950 12798 32002 12850
rect 32062 12798 32114 12850
rect 33182 12798 33234 12850
rect 33406 12798 33458 12850
rect 41022 12798 41074 12850
rect 41134 12798 41186 12850
rect 44158 12798 44210 12850
rect 2046 12686 2098 12738
rect 3502 12686 3554 12738
rect 4062 12686 4114 12738
rect 10670 12686 10722 12738
rect 13582 12686 13634 12738
rect 13694 12686 13746 12738
rect 19070 12686 19122 12738
rect 20078 12686 20130 12738
rect 24222 12686 24274 12738
rect 26014 12686 26066 12738
rect 26798 12686 26850 12738
rect 28254 12686 28306 12738
rect 28478 12686 28530 12738
rect 31502 12686 31554 12738
rect 32286 12686 32338 12738
rect 33294 12686 33346 12738
rect 34302 12686 34354 12738
rect 38558 12686 38610 12738
rect 42366 12686 42418 12738
rect 43150 12686 43202 12738
rect 44046 12686 44098 12738
rect 47070 12686 47122 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 2046 12350 2098 12402
rect 2830 12350 2882 12402
rect 3390 12350 3442 12402
rect 4174 12350 4226 12402
rect 4510 12350 4562 12402
rect 5854 12350 5906 12402
rect 9774 12350 9826 12402
rect 13134 12350 13186 12402
rect 14702 12350 14754 12402
rect 17614 12350 17666 12402
rect 18622 12350 18674 12402
rect 19742 12350 19794 12402
rect 19966 12350 20018 12402
rect 26686 12350 26738 12402
rect 26798 12350 26850 12402
rect 26910 12350 26962 12402
rect 29822 12350 29874 12402
rect 30382 12350 30434 12402
rect 33182 12350 33234 12402
rect 33854 12350 33906 12402
rect 34750 12350 34802 12402
rect 38782 12350 38834 12402
rect 40350 12350 40402 12402
rect 4846 12238 4898 12290
rect 6414 12238 6466 12290
rect 6862 12238 6914 12290
rect 7086 12238 7138 12290
rect 8430 12238 8482 12290
rect 8766 12238 8818 12290
rect 9998 12238 10050 12290
rect 11790 12238 11842 12290
rect 12686 12238 12738 12290
rect 13918 12238 13970 12290
rect 14478 12238 14530 12290
rect 15822 12238 15874 12290
rect 16606 12238 16658 12290
rect 17950 12238 18002 12290
rect 19182 12238 19234 12290
rect 19294 12238 19346 12290
rect 19518 12238 19570 12290
rect 20638 12238 20690 12290
rect 20750 12238 20802 12290
rect 22542 12238 22594 12290
rect 26238 12238 26290 12290
rect 28814 12238 28866 12290
rect 29598 12238 29650 12290
rect 30718 12238 30770 12290
rect 32510 12238 32562 12290
rect 33294 12238 33346 12290
rect 33966 12238 34018 12290
rect 34974 12238 35026 12290
rect 35198 12238 35250 12290
rect 37102 12238 37154 12290
rect 37774 12238 37826 12290
rect 38670 12238 38722 12290
rect 39230 12238 39282 12290
rect 40910 12238 40962 12290
rect 42142 12238 42194 12290
rect 42366 12238 42418 12290
rect 43598 12238 43650 12290
rect 46174 12238 46226 12290
rect 1710 12126 1762 12178
rect 2494 12126 2546 12178
rect 3166 12126 3218 12178
rect 3838 12126 3890 12178
rect 5294 12126 5346 12178
rect 6078 12126 6130 12178
rect 8990 12126 9042 12178
rect 10334 12126 10386 12178
rect 12126 12126 12178 12178
rect 12238 12126 12290 12178
rect 12910 12126 12962 12178
rect 13246 12126 13298 12178
rect 13582 12126 13634 12178
rect 14142 12126 14194 12178
rect 15486 12126 15538 12178
rect 16382 12126 16434 12178
rect 17390 12126 17442 12178
rect 17726 12126 17778 12178
rect 18398 12126 18450 12178
rect 20414 12126 20466 12178
rect 21870 12126 21922 12178
rect 25342 12126 25394 12178
rect 25790 12126 25842 12178
rect 27358 12126 27410 12178
rect 27582 12126 27634 12178
rect 27918 12126 27970 12178
rect 29150 12126 29202 12178
rect 29486 12126 29538 12178
rect 30270 12126 30322 12178
rect 30494 12126 30546 12178
rect 31614 12126 31666 12178
rect 32958 12126 33010 12178
rect 33742 12126 33794 12178
rect 34414 12126 34466 12178
rect 34526 12126 34578 12178
rect 36206 12126 36258 12178
rect 36766 12126 36818 12178
rect 38222 12126 38274 12178
rect 38446 12126 38498 12178
rect 41470 12126 41522 12178
rect 42814 12126 42866 12178
rect 3278 12014 3330 12066
rect 8542 12014 8594 12066
rect 10110 12014 10162 12066
rect 11902 12014 11954 12066
rect 13694 12014 13746 12066
rect 14590 12014 14642 12066
rect 15598 12014 15650 12066
rect 19854 12014 19906 12066
rect 24670 12014 24722 12066
rect 29038 12014 29090 12066
rect 32062 12014 32114 12066
rect 39118 12014 39170 12066
rect 42478 12014 42530 12066
rect 45726 12014 45778 12066
rect 6078 11902 6130 11954
rect 6750 11902 6802 11954
rect 20750 11902 20802 11954
rect 37214 11902 37266 11954
rect 37886 11902 37938 11954
rect 39006 11902 39058 11954
rect 41022 11902 41074 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 9102 11566 9154 11618
rect 14814 11566 14866 11618
rect 27358 11566 27410 11618
rect 38222 11566 38274 11618
rect 41806 11566 41858 11618
rect 43038 11566 43090 11618
rect 2494 11454 2546 11506
rect 4622 11454 4674 11506
rect 5070 11454 5122 11506
rect 5742 11454 5794 11506
rect 9214 11454 9266 11506
rect 9998 11454 10050 11506
rect 11342 11454 11394 11506
rect 27134 11454 27186 11506
rect 28366 11454 28418 11506
rect 34302 11454 34354 11506
rect 35198 11454 35250 11506
rect 36094 11454 36146 11506
rect 41246 11454 41298 11506
rect 45838 11454 45890 11506
rect 49310 11454 49362 11506
rect 1822 11342 1874 11394
rect 6078 11342 6130 11394
rect 9438 11342 9490 11394
rect 11678 11342 11730 11394
rect 12238 11342 12290 11394
rect 12798 11342 12850 11394
rect 13582 11342 13634 11394
rect 13694 11342 13746 11394
rect 14030 11342 14082 11394
rect 14702 11342 14754 11394
rect 15038 11342 15090 11394
rect 15710 11342 15762 11394
rect 16942 11342 16994 11394
rect 20750 11342 20802 11394
rect 25342 11342 25394 11394
rect 25902 11342 25954 11394
rect 26014 11342 26066 11394
rect 26574 11342 26626 11394
rect 27470 11342 27522 11394
rect 30270 11342 30322 11394
rect 30942 11342 30994 11394
rect 31278 11342 31330 11394
rect 31838 11342 31890 11394
rect 32174 11342 32226 11394
rect 32846 11342 32898 11394
rect 33630 11342 33682 11394
rect 34078 11342 34130 11394
rect 34526 11342 34578 11394
rect 34638 11342 34690 11394
rect 35422 11342 35474 11394
rect 37102 11342 37154 11394
rect 37774 11342 37826 11394
rect 38222 11342 38274 11394
rect 38782 11342 38834 11394
rect 39118 11342 39170 11394
rect 39342 11342 39394 11394
rect 39790 11342 39842 11394
rect 40350 11342 40402 11394
rect 40798 11342 40850 11394
rect 41582 11342 41634 11394
rect 43374 11342 43426 11394
rect 47966 11342 48018 11394
rect 48750 11342 48802 11394
rect 5630 11230 5682 11282
rect 5966 11230 6018 11282
rect 15822 11230 15874 11282
rect 17054 11230 17106 11282
rect 19518 11230 19570 11282
rect 25566 11230 25618 11282
rect 29934 11230 29986 11282
rect 30046 11230 30098 11282
rect 30718 11230 30770 11282
rect 31502 11230 31554 11282
rect 37214 11230 37266 11282
rect 38894 11230 38946 11282
rect 39678 11230 39730 11282
rect 42142 11230 42194 11282
rect 42254 11230 42306 11282
rect 42366 11230 42418 11282
rect 42702 11230 42754 11282
rect 11790 11118 11842 11170
rect 11902 11118 11954 11170
rect 12014 11118 12066 11170
rect 12574 11118 12626 11170
rect 13806 11118 13858 11170
rect 13918 11118 13970 11170
rect 17166 11118 17218 11170
rect 24894 11118 24946 11170
rect 26126 11118 26178 11170
rect 30606 11118 30658 11170
rect 31390 11118 31442 11170
rect 32286 11118 32338 11170
rect 32398 11118 32450 11170
rect 33070 11118 33122 11170
rect 39902 11118 39954 11170
rect 42926 11118 42978 11170
rect 43486 11118 43538 11170
rect 44158 11118 44210 11170
rect 44942 11118 44994 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 2046 10782 2098 10834
rect 2718 10782 2770 10834
rect 3390 10782 3442 10834
rect 3950 10782 4002 10834
rect 4846 10782 4898 10834
rect 5518 10782 5570 10834
rect 7310 10782 7362 10834
rect 8654 10782 8706 10834
rect 13246 10782 13298 10834
rect 17950 10782 18002 10834
rect 26798 10782 26850 10834
rect 33742 10782 33794 10834
rect 34638 10782 34690 10834
rect 36206 10782 36258 10834
rect 37326 10782 37378 10834
rect 38558 10782 38610 10834
rect 39006 10782 39058 10834
rect 39566 10782 39618 10834
rect 42254 10782 42306 10834
rect 43598 10782 43650 10834
rect 1710 10670 1762 10722
rect 2382 10670 2434 10722
rect 4286 10670 4338 10722
rect 4398 10670 4450 10722
rect 5854 10670 5906 10722
rect 6750 10670 6802 10722
rect 9662 10670 9714 10722
rect 12126 10670 12178 10722
rect 13806 10670 13858 10722
rect 15374 10670 15426 10722
rect 16830 10670 16882 10722
rect 19966 10670 20018 10722
rect 27246 10670 27298 10722
rect 34526 10670 34578 10722
rect 36990 10670 37042 10722
rect 37102 10670 37154 10722
rect 37886 10670 37938 10722
rect 41470 10670 41522 10722
rect 42590 10670 42642 10722
rect 42814 10670 42866 10722
rect 43262 10670 43314 10722
rect 3054 10558 3106 10610
rect 5182 10558 5234 10610
rect 6190 10558 6242 10610
rect 6526 10558 6578 10610
rect 8430 10558 8482 10610
rect 8766 10558 8818 10610
rect 8990 10558 9042 10610
rect 9550 10558 9602 10610
rect 11566 10558 11618 10610
rect 14478 10558 14530 10610
rect 14814 10558 14866 10610
rect 16270 10558 16322 10610
rect 16606 10558 16658 10610
rect 18174 10558 18226 10610
rect 18510 10558 18562 10610
rect 19294 10558 19346 10610
rect 27582 10558 27634 10610
rect 33182 10558 33234 10610
rect 34862 10558 34914 10610
rect 35758 10558 35810 10610
rect 35982 10558 36034 10610
rect 36094 10558 36146 10610
rect 38222 10558 38274 10610
rect 39790 10558 39842 10610
rect 41246 10558 41298 10610
rect 44718 10558 44770 10610
rect 45166 10558 45218 10610
rect 6302 10446 6354 10498
rect 15038 10446 15090 10498
rect 16718 10446 16770 10498
rect 18062 10446 18114 10498
rect 22094 10446 22146 10498
rect 22542 10446 22594 10498
rect 23550 10446 23602 10498
rect 31278 10446 31330 10498
rect 33854 10446 33906 10498
rect 39118 10446 39170 10498
rect 42926 10446 42978 10498
rect 44046 10446 44098 10498
rect 4398 10334 4450 10386
rect 23438 10334 23490 10386
rect 30942 10334 30994 10386
rect 31278 10334 31330 10386
rect 35534 10334 35586 10386
rect 37662 10334 37714 10386
rect 38446 10334 38498 10386
rect 39454 10334 39506 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 7086 9998 7138 10050
rect 11902 9998 11954 10050
rect 14366 9998 14418 10050
rect 18510 9998 18562 10050
rect 35870 9998 35922 10050
rect 37550 9998 37602 10050
rect 4846 9886 4898 9938
rect 8542 9886 8594 9938
rect 10670 9886 10722 9938
rect 13582 9886 13634 9938
rect 16830 9886 16882 9938
rect 22990 9886 23042 9938
rect 25118 9886 25170 9938
rect 26686 9886 26738 9938
rect 29710 9886 29762 9938
rect 34190 9886 34242 9938
rect 34638 9886 34690 9938
rect 34862 9886 34914 9938
rect 36542 9886 36594 9938
rect 37214 9886 37266 9938
rect 38782 9886 38834 9938
rect 41246 9886 41298 9938
rect 2046 9774 2098 9826
rect 5518 9774 5570 9826
rect 5966 9774 6018 9826
rect 6190 9774 6242 9826
rect 7534 9774 7586 9826
rect 11342 9774 11394 9826
rect 11790 9774 11842 9826
rect 12350 9774 12402 9826
rect 12910 9774 12962 9826
rect 13358 9774 13410 9826
rect 13918 9774 13970 9826
rect 16270 9774 16322 9826
rect 17054 9774 17106 9826
rect 17726 9774 17778 9826
rect 18622 9774 18674 9826
rect 19070 9774 19122 9826
rect 19854 9774 19906 9826
rect 22206 9774 22258 9826
rect 27022 9774 27074 9826
rect 27246 9774 27298 9826
rect 27806 9774 27858 9826
rect 28030 9774 28082 9826
rect 32622 9774 32674 9826
rect 35422 9774 35474 9826
rect 39118 9774 39170 9826
rect 41134 9774 41186 9826
rect 43374 9774 43426 9826
rect 43486 9774 43538 9826
rect 43934 9774 43986 9826
rect 2718 9662 2770 9714
rect 6078 9662 6130 9714
rect 7758 9662 7810 9714
rect 12686 9662 12738 9714
rect 13806 9662 13858 9714
rect 14478 9662 14530 9714
rect 17502 9662 17554 9714
rect 18510 9662 18562 9714
rect 19406 9662 19458 9714
rect 28254 9662 28306 9714
rect 31838 9662 31890 9714
rect 35758 9662 35810 9714
rect 6750 9550 6802 9602
rect 12462 9550 12514 9602
rect 17614 9550 17666 9602
rect 21870 9550 21922 9602
rect 26686 9550 26738 9602
rect 26798 9550 26850 9602
rect 27694 9550 27746 9602
rect 27918 9550 27970 9602
rect 33070 9550 33122 9602
rect 37438 9606 37490 9658
rect 37550 9662 37602 9714
rect 39230 9662 39282 9714
rect 42814 9662 42866 9714
rect 43598 9550 43650 9602
rect 43710 9550 43762 9602
rect 44830 9550 44882 9602
rect 45166 9550 45218 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 2158 9214 2210 9266
rect 2494 9214 2546 9266
rect 3838 9214 3890 9266
rect 8430 9214 8482 9266
rect 9550 9214 9602 9266
rect 9774 9214 9826 9266
rect 10446 9214 10498 9266
rect 12574 9214 12626 9266
rect 16046 9214 16098 9266
rect 16270 9214 16322 9266
rect 22430 9214 22482 9266
rect 22654 9214 22706 9266
rect 22990 9214 23042 9266
rect 23662 9214 23714 9266
rect 23774 9214 23826 9266
rect 23886 9214 23938 9266
rect 24670 9214 24722 9266
rect 29150 9214 29202 9266
rect 33742 9214 33794 9266
rect 34526 9214 34578 9266
rect 34974 9214 35026 9266
rect 35086 9214 35138 9266
rect 35870 9214 35922 9266
rect 40014 9214 40066 9266
rect 40126 9214 40178 9266
rect 42366 9214 42418 9266
rect 46062 9214 46114 9266
rect 10782 9102 10834 9154
rect 19518 9102 19570 9154
rect 24110 9102 24162 9154
rect 28590 9102 28642 9154
rect 33966 9102 34018 9154
rect 35310 9102 35362 9154
rect 35534 9102 35586 9154
rect 39118 9102 39170 9154
rect 39790 9102 39842 9154
rect 40910 9102 40962 9154
rect 4622 8990 4674 9042
rect 5070 8990 5122 9042
rect 10222 8990 10274 9042
rect 12686 8990 12738 9042
rect 15934 8990 15986 9042
rect 20190 8990 20242 9042
rect 20750 8990 20802 9042
rect 23438 8990 23490 9042
rect 25230 8990 25282 9042
rect 29486 8990 29538 9042
rect 30270 8990 30322 9042
rect 36094 8990 36146 9042
rect 37214 8990 37266 9042
rect 37662 8990 37714 9042
rect 38222 8990 38274 9042
rect 39566 8990 39618 9042
rect 41022 8990 41074 9042
rect 41358 8990 41410 9042
rect 42702 8990 42754 9042
rect 5742 8878 5794 8930
rect 7870 8878 7922 8930
rect 8766 8878 8818 8930
rect 9662 8878 9714 8930
rect 17390 8878 17442 8930
rect 26014 8878 26066 8930
rect 28142 8878 28194 8930
rect 30046 8878 30098 8930
rect 30830 8878 30882 8930
rect 35086 8878 35138 8930
rect 39902 8878 39954 8930
rect 43486 8878 43538 8930
rect 45614 8878 45666 8930
rect 12574 8766 12626 8818
rect 28478 8766 28530 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 26126 8430 26178 8482
rect 43486 8430 43538 8482
rect 8094 8318 8146 8370
rect 10222 8318 10274 8370
rect 11230 8318 11282 8370
rect 15598 8318 15650 8370
rect 17726 8318 17778 8370
rect 26238 8318 26290 8370
rect 32174 8318 32226 8370
rect 34302 8318 34354 8370
rect 38334 8318 38386 8370
rect 39678 8318 39730 8370
rect 43598 8318 43650 8370
rect 6302 8206 6354 8258
rect 7310 8206 7362 8258
rect 10446 8206 10498 8258
rect 10782 8206 10834 8258
rect 12014 8206 12066 8258
rect 12238 8206 12290 8258
rect 12574 8206 12626 8258
rect 13470 8206 13522 8258
rect 13694 8206 13746 8258
rect 14030 8206 14082 8258
rect 14254 8206 14306 8258
rect 14590 8206 14642 8258
rect 18510 8206 18562 8258
rect 18958 8206 19010 8258
rect 31502 8206 31554 8258
rect 35422 8206 35474 8258
rect 35982 8206 36034 8258
rect 38894 8206 38946 8258
rect 42590 8206 42642 8258
rect 5966 8094 6018 8146
rect 10670 8094 10722 8146
rect 34750 8094 34802 8146
rect 38670 8094 38722 8146
rect 41806 8094 41858 8146
rect 42926 8094 42978 8146
rect 43038 8094 43090 8146
rect 12126 7982 12178 8034
rect 13582 7982 13634 8034
rect 14478 7982 14530 8034
rect 38222 7982 38274 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 8094 7646 8146 7698
rect 8990 7646 9042 7698
rect 27022 7646 27074 7698
rect 36430 7646 36482 7698
rect 40126 7646 40178 7698
rect 41134 7646 41186 7698
rect 41246 7646 41298 7698
rect 41358 7646 41410 7698
rect 41470 7646 41522 7698
rect 42814 7646 42866 7698
rect 10558 7534 10610 7586
rect 15150 7534 15202 7586
rect 28142 7534 28194 7586
rect 37550 7534 37602 7586
rect 41694 7534 41746 7586
rect 9774 7422 9826 7474
rect 15934 7422 15986 7474
rect 16382 7422 16434 7474
rect 27358 7422 27410 7474
rect 33182 7422 33234 7474
rect 36878 7422 36930 7474
rect 12686 7310 12738 7362
rect 13022 7310 13074 7362
rect 30270 7310 30322 7362
rect 33854 7310 33906 7362
rect 35982 7310 36034 7362
rect 39678 7310 39730 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 34638 6862 34690 6914
rect 35310 6750 35362 6802
rect 34862 6638 34914 6690
rect 35086 6638 35138 6690
rect 34750 6526 34802 6578
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 11454 6078 11506 6130
rect 12574 5966 12626 6018
rect 11790 5854 11842 5906
rect 14702 5742 14754 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 38558 4510 38610 4562
rect 38782 4286 38834 4338
rect 17614 4174 17666 4226
rect 18174 4174 18226 4226
rect 30942 4174 30994 4226
rect 31950 4174 32002 4226
rect 32622 4174 32674 4226
rect 33294 4174 33346 4226
rect 34190 4174 34242 4226
rect 34862 4174 34914 4226
rect 35758 4174 35810 4226
rect 36430 4174 36482 4226
rect 37102 4174 37154 4226
rect 37774 4174 37826 4226
rect 38334 4174 38386 4226
rect 39342 4174 39394 4226
rect 39790 4174 39842 4226
rect 40350 4174 40402 4226
rect 37774 4062 37826 4114
rect 38222 4062 38274 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 25006 3614 25058 3666
rect 33966 3614 34018 3666
rect 18622 3502 18674 3554
rect 29150 3502 29202 3554
rect 31166 3502 31218 3554
rect 32174 3502 32226 3554
rect 32846 3502 32898 3554
rect 33518 3502 33570 3554
rect 34414 3502 34466 3554
rect 36206 3502 36258 3554
rect 36878 3502 36930 3554
rect 37550 3502 37602 3554
rect 38222 3502 38274 3554
rect 39006 3502 39058 3554
rect 39790 3502 39842 3554
rect 40686 3502 40738 3554
rect 16494 3390 16546 3442
rect 17054 3390 17106 3442
rect 17390 3390 17442 3442
rect 17726 3390 17778 3442
rect 18062 3390 18114 3442
rect 18398 3390 18450 3442
rect 24110 3390 24162 3442
rect 24558 3390 24610 3442
rect 29822 3390 29874 3442
rect 30158 3390 30210 3442
rect 30494 3390 30546 3442
rect 30830 3390 30882 3442
rect 31502 3390 31554 3442
rect 32510 3390 32562 3442
rect 33182 3390 33234 3442
rect 34750 3390 34802 3442
rect 35086 3390 35138 3442
rect 35422 3390 35474 3442
rect 35982 3390 36034 3442
rect 36654 3390 36706 3442
rect 37326 3390 37378 3442
rect 37998 3390 38050 3442
rect 38670 3390 38722 3442
rect 40126 3390 40178 3442
rect 40462 3390 40514 3442
rect 29598 3278 29650 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 35646 2494 35698 2546
rect 36430 2494 36482 2546
rect 36878 2494 36930 2546
rect 36990 2382 37042 2434
rect 38222 2382 38274 2434
<< metal2 >>
rect 20160 59200 20272 60000
rect 23520 59200 23632 60000
rect 25536 59200 25648 60000
rect 27552 59200 27664 60000
rect 28896 59200 29008 60000
rect 29568 59200 29680 60000
rect 30240 59200 30352 60000
rect 30912 59200 31024 60000
rect 31584 59200 31696 60000
rect 32256 59200 32368 60000
rect 33600 59200 33712 60000
rect 36288 59200 36400 60000
rect 36960 59200 37072 60000
rect 37632 59200 37744 60000
rect 38304 59200 38416 60000
rect 19180 56642 19236 56654
rect 19180 56590 19182 56642
rect 19234 56590 19236 56642
rect 19180 56306 19236 56590
rect 20076 56644 20132 56654
rect 20188 56644 20244 59200
rect 23548 57428 23604 59200
rect 23548 57372 23716 57428
rect 20076 56642 20244 56644
rect 20076 56590 20078 56642
rect 20130 56590 20244 56642
rect 20076 56588 20244 56590
rect 20076 56578 20132 56588
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19180 56254 19182 56306
rect 19234 56254 19236 56306
rect 19180 56242 19236 56254
rect 20188 56084 20244 56094
rect 20188 55990 20244 56028
rect 20860 56084 20916 56094
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 14588 55410 14644 55422
rect 14588 55358 14590 55410
rect 14642 55358 14644 55410
rect 8764 55188 8820 55198
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 1932 50706 1988 50718
rect 1932 50654 1934 50706
rect 1986 50654 1988 50706
rect 1708 49810 1764 49822
rect 1708 49758 1710 49810
rect 1762 49758 1764 49810
rect 1708 49700 1764 49758
rect 1932 49812 1988 50654
rect 3836 50596 3892 50606
rect 3724 50594 3892 50596
rect 3724 50542 3838 50594
rect 3890 50542 3892 50594
rect 3724 50540 3892 50542
rect 2044 49924 2100 49934
rect 2044 49830 2100 49868
rect 1932 49746 1988 49756
rect 1708 49140 1764 49644
rect 2492 49700 2548 49710
rect 2492 49606 2548 49644
rect 1708 49074 1764 49084
rect 1708 48914 1764 48926
rect 1708 48862 1710 48914
rect 1762 48862 1764 48914
rect 1708 48468 1764 48862
rect 2044 48804 2100 48814
rect 2044 48802 2436 48804
rect 2044 48750 2046 48802
rect 2098 48750 2436 48802
rect 2044 48748 2436 48750
rect 2044 48738 2100 48748
rect 1708 48402 1764 48412
rect 2044 48356 2100 48366
rect 2044 48262 2100 48300
rect 1708 48242 1764 48254
rect 1708 48190 1710 48242
rect 1762 48190 1764 48242
rect 1708 47796 1764 48190
rect 1708 47730 1764 47740
rect 1708 47346 1764 47358
rect 1708 47294 1710 47346
rect 1762 47294 1764 47346
rect 1708 47124 1764 47294
rect 2044 47236 2100 47246
rect 2044 47142 2100 47180
rect 1708 47058 1764 47068
rect 2044 46788 2100 46798
rect 2380 46788 2436 48748
rect 2492 48802 2548 48814
rect 2492 48750 2494 48802
rect 2546 48750 2548 48802
rect 2492 48468 2548 48750
rect 2492 48402 2548 48412
rect 2492 48130 2548 48142
rect 2492 48078 2494 48130
rect 2546 48078 2548 48130
rect 2492 47796 2548 48078
rect 2492 47730 2548 47740
rect 2492 47234 2548 47246
rect 2492 47182 2494 47234
rect 2546 47182 2548 47234
rect 2492 47124 2548 47182
rect 2492 47058 2548 47068
rect 3612 47236 3668 47246
rect 2044 46786 2324 46788
rect 2044 46734 2046 46786
rect 2098 46734 2324 46786
rect 2044 46732 2324 46734
rect 2380 46732 2660 46788
rect 2044 46722 2100 46732
rect 1708 46674 1764 46686
rect 1708 46622 1710 46674
rect 1762 46622 1764 46674
rect 1708 46452 1764 46622
rect 1708 46386 1764 46396
rect 2268 46450 2324 46732
rect 2268 46398 2270 46450
rect 2322 46398 2324 46450
rect 2268 46386 2324 46398
rect 2492 46562 2548 46574
rect 2492 46510 2494 46562
rect 2546 46510 2548 46562
rect 2492 46004 2548 46510
rect 2268 45948 2548 46004
rect 1820 45892 1876 45902
rect 2268 45892 2324 45948
rect 1820 45890 2324 45892
rect 1820 45838 1822 45890
rect 1874 45838 2324 45890
rect 1820 45836 2324 45838
rect 1708 45106 1764 45118
rect 1708 45054 1710 45106
rect 1762 45054 1764 45106
rect 1708 44996 1764 45054
rect 1820 45108 1876 45836
rect 2380 45780 2436 45790
rect 2380 45686 2436 45724
rect 2044 45668 2100 45678
rect 2044 45666 2212 45668
rect 2044 45614 2046 45666
rect 2098 45614 2212 45666
rect 2044 45612 2212 45614
rect 2044 45602 2100 45612
rect 2044 45220 2100 45230
rect 2044 45126 2100 45164
rect 1820 45042 1876 45052
rect 1708 44436 1764 44940
rect 2156 44548 2212 45612
rect 2492 44996 2548 45006
rect 2492 44902 2548 44940
rect 2156 44482 2212 44492
rect 1708 44370 1764 44380
rect 1932 44434 1988 44446
rect 1932 44382 1934 44434
rect 1986 44382 1988 44434
rect 1932 43764 1988 44382
rect 1932 43698 1988 43708
rect 2044 43652 2100 43662
rect 2044 43558 2100 43596
rect 1708 43538 1764 43550
rect 1708 43486 1710 43538
rect 1762 43486 1764 43538
rect 1708 43092 1764 43486
rect 1708 43026 1764 43036
rect 2492 43426 2548 43438
rect 2492 43374 2494 43426
rect 2546 43374 2548 43426
rect 2492 43092 2548 43374
rect 2492 43026 2548 43036
rect 2156 42756 2212 42766
rect 1708 42642 1764 42654
rect 1708 42590 1710 42642
rect 1762 42590 1764 42642
rect 1708 42420 1764 42590
rect 2044 42644 2100 42654
rect 2044 42550 2100 42588
rect 1708 42354 1764 42364
rect 2044 42196 2100 42206
rect 2156 42196 2212 42700
rect 2492 42530 2548 42542
rect 2492 42478 2494 42530
rect 2546 42478 2548 42530
rect 2492 42420 2548 42478
rect 2492 42354 2548 42364
rect 2044 42194 2212 42196
rect 2044 42142 2046 42194
rect 2098 42142 2212 42194
rect 2044 42140 2212 42142
rect 2044 42130 2100 42140
rect 1708 41970 1764 41982
rect 1708 41918 1710 41970
rect 1762 41918 1764 41970
rect 1708 41748 1764 41918
rect 2604 41972 2660 46732
rect 2940 46562 2996 46574
rect 2940 46510 2942 46562
rect 2994 46510 2996 46562
rect 2940 46452 2996 46510
rect 2940 46386 2996 46396
rect 3052 46450 3108 46462
rect 3052 46398 3054 46450
rect 3106 46398 3108 46450
rect 2716 45666 2772 45678
rect 2716 45614 2718 45666
rect 2770 45614 2772 45666
rect 2716 43876 2772 45614
rect 2716 43810 2772 43820
rect 3052 43708 3108 46398
rect 3164 45780 3220 45790
rect 3164 45686 3220 45724
rect 3052 43652 3444 43708
rect 3388 42754 3444 43652
rect 3388 42702 3390 42754
rect 3442 42702 3444 42754
rect 3388 42690 3444 42702
rect 3612 41972 3668 47180
rect 3724 44100 3780 50540
rect 3836 50530 3892 50540
rect 3948 49924 4004 49934
rect 3724 44044 3892 44100
rect 3724 43876 3780 43886
rect 3724 42754 3780 43820
rect 3836 43428 3892 44044
rect 3836 43362 3892 43372
rect 3724 42702 3726 42754
rect 3778 42702 3780 42754
rect 3724 42690 3780 42702
rect 3948 42756 4004 49868
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 5964 48356 6020 48366
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 5292 44548 5348 44558
rect 4284 44322 4340 44334
rect 4284 44270 4286 44322
rect 4338 44270 4340 44322
rect 4284 43540 4340 44270
rect 4284 43474 4340 43484
rect 4844 43650 4900 43662
rect 4844 43598 4846 43650
rect 4898 43598 4900 43650
rect 4620 43316 4676 43326
rect 4060 43314 4676 43316
rect 4060 43262 4622 43314
rect 4674 43262 4676 43314
rect 4060 43260 4676 43262
rect 4060 42978 4116 43260
rect 4620 43250 4676 43260
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4060 42926 4062 42978
rect 4114 42926 4116 42978
rect 4060 42914 4116 42926
rect 3948 42700 4452 42756
rect 3948 42530 4004 42542
rect 3948 42478 3950 42530
rect 4002 42478 4004 42530
rect 3948 42194 4004 42478
rect 3948 42142 3950 42194
rect 4002 42142 4004 42194
rect 3948 42130 4004 42142
rect 4396 42082 4452 42700
rect 4844 42644 4900 43598
rect 5292 43650 5348 44492
rect 5292 43598 5294 43650
rect 5346 43598 5348 43650
rect 5292 43586 5348 43598
rect 5740 43428 5796 43438
rect 5740 43334 5796 43372
rect 4844 42578 4900 42588
rect 4956 43314 5012 43326
rect 4956 43262 4958 43314
rect 5010 43262 5012 43314
rect 4396 42030 4398 42082
rect 4450 42030 4452 42082
rect 4396 42018 4452 42030
rect 3836 41972 3892 41982
rect 3612 41970 3892 41972
rect 3612 41918 3838 41970
rect 3890 41918 3892 41970
rect 3612 41916 3892 41918
rect 2604 41906 2660 41916
rect 3836 41906 3892 41916
rect 4284 41972 4340 41982
rect 4284 41878 4340 41916
rect 4956 41972 5012 43262
rect 4956 41906 5012 41916
rect 5404 43314 5460 43326
rect 5404 43262 5406 43314
rect 5458 43262 5460 43314
rect 5404 41970 5460 43262
rect 5628 42756 5684 42766
rect 5404 41918 5406 41970
rect 5458 41918 5460 41970
rect 5404 41906 5460 41918
rect 5516 42754 5684 42756
rect 5516 42702 5630 42754
rect 5682 42702 5684 42754
rect 5516 42700 5684 42702
rect 1708 41682 1764 41692
rect 2492 41858 2548 41870
rect 2492 41806 2494 41858
rect 2546 41806 2548 41858
rect 2044 41412 2100 41422
rect 1820 41188 1876 41198
rect 1708 40402 1764 40414
rect 1708 40350 1710 40402
rect 1762 40350 1764 40402
rect 1708 40292 1764 40350
rect 1820 40404 1876 41132
rect 2044 41074 2100 41356
rect 2492 41188 2548 41806
rect 2492 41122 2548 41132
rect 2716 41860 2772 41870
rect 2044 41022 2046 41074
rect 2098 41022 2100 41074
rect 2044 41010 2100 41022
rect 2380 41076 2436 41086
rect 2380 40982 2436 41020
rect 2716 41074 2772 41804
rect 2940 41858 2996 41870
rect 2940 41806 2942 41858
rect 2994 41806 2996 41858
rect 2940 41748 2996 41806
rect 2940 41682 2996 41692
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 2716 41022 2718 41074
rect 2770 41022 2772 41074
rect 2716 41010 2772 41022
rect 3164 41076 3220 41086
rect 3164 40982 3220 41020
rect 1820 40338 1876 40348
rect 2044 40514 2100 40526
rect 5516 40516 5572 42700
rect 5628 42690 5684 42700
rect 5852 42756 5908 42766
rect 5852 42662 5908 42700
rect 5852 42196 5908 42206
rect 5852 42102 5908 42140
rect 5964 42082 6020 48300
rect 8428 47012 8484 47022
rect 8428 45892 8484 46956
rect 8204 45890 8484 45892
rect 8204 45838 8430 45890
rect 8482 45838 8484 45890
rect 8204 45836 8484 45838
rect 6748 45220 6804 45230
rect 6076 42868 6132 42878
rect 6076 42866 6692 42868
rect 6076 42814 6078 42866
rect 6130 42814 6692 42866
rect 6076 42812 6692 42814
rect 6076 42802 6132 42812
rect 6188 42642 6244 42654
rect 6188 42590 6190 42642
rect 6242 42590 6244 42642
rect 6188 42308 6244 42590
rect 6188 42252 6580 42308
rect 5964 42030 5966 42082
rect 6018 42030 6020 42082
rect 5964 42018 6020 42030
rect 6188 42082 6244 42094
rect 6188 42030 6190 42082
rect 6242 42030 6244 42082
rect 6188 41074 6244 42030
rect 6524 42082 6580 42252
rect 6524 42030 6526 42082
rect 6578 42030 6580 42082
rect 6524 42018 6580 42030
rect 6300 41972 6356 41982
rect 6300 41878 6356 41916
rect 6188 41022 6190 41074
rect 6242 41022 6244 41074
rect 6188 41010 6244 41022
rect 6300 40964 6356 40974
rect 6300 40962 6580 40964
rect 6300 40910 6302 40962
rect 6354 40910 6580 40962
rect 6300 40908 6580 40910
rect 6300 40898 6356 40908
rect 2044 40462 2046 40514
rect 2098 40462 2100 40514
rect 1708 39060 1764 40236
rect 2044 40180 2100 40462
rect 5180 40460 5572 40516
rect 2492 40402 2548 40414
rect 2492 40350 2494 40402
rect 2546 40350 2548 40402
rect 2492 40292 2548 40350
rect 4620 40404 4676 40414
rect 4620 40310 4676 40348
rect 2492 40226 2548 40236
rect 2044 40114 2100 40124
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 1932 39732 1988 39742
rect 1932 39638 1988 39676
rect 4284 39620 4340 39630
rect 4284 39526 4340 39564
rect 1708 38994 1764 39004
rect 2044 38948 2100 38958
rect 2044 38854 2100 38892
rect 4620 38948 4676 38958
rect 4620 38854 4676 38892
rect 1708 38834 1764 38846
rect 1708 38782 1710 38834
rect 1762 38782 1764 38834
rect 1708 38388 1764 38782
rect 4732 38836 4788 38846
rect 5180 38836 5236 40460
rect 5292 40290 5348 40302
rect 5292 40238 5294 40290
rect 5346 40238 5348 40290
rect 5292 39172 5348 40238
rect 6524 39732 6580 40908
rect 6076 39730 6580 39732
rect 6076 39678 6526 39730
rect 6578 39678 6580 39730
rect 6076 39676 6580 39678
rect 5292 39106 5348 39116
rect 5404 39564 6020 39620
rect 5180 38780 5348 38836
rect 4732 38742 4788 38780
rect 1708 38322 1764 38332
rect 2492 38722 2548 38734
rect 2492 38670 2494 38722
rect 2546 38670 2548 38722
rect 2492 38388 2548 38670
rect 5068 38722 5124 38734
rect 5068 38670 5070 38722
rect 5122 38670 5124 38722
rect 5068 38500 5124 38670
rect 5180 38612 5236 38622
rect 5180 38518 5236 38556
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 2492 38322 2548 38332
rect 1708 37938 1764 37950
rect 1708 37886 1710 37938
rect 1762 37886 1764 37938
rect 1708 37716 1764 37886
rect 2044 37940 2100 37950
rect 2044 37846 2100 37884
rect 1708 37650 1764 37660
rect 2492 37826 2548 37838
rect 2492 37774 2494 37826
rect 2546 37774 2548 37826
rect 2492 37716 2548 37774
rect 2492 37650 2548 37660
rect 2044 37492 2100 37502
rect 2044 37398 2100 37436
rect 5068 37492 5124 38444
rect 5068 37426 5124 37436
rect 1708 37266 1764 37278
rect 1708 37214 1710 37266
rect 1762 37214 1764 37266
rect 1708 37044 1764 37214
rect 1708 36978 1764 36988
rect 2492 37154 2548 37166
rect 2492 37102 2494 37154
rect 2546 37102 2548 37154
rect 1708 36484 1764 36494
rect 1708 36370 1764 36428
rect 2492 36484 2548 37102
rect 2940 37154 2996 37166
rect 2940 37102 2942 37154
rect 2994 37102 2996 37154
rect 2940 37044 2996 37102
rect 2940 36978 2996 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 2492 36418 2548 36428
rect 2716 36596 2772 36606
rect 1708 36318 1710 36370
rect 1762 36318 1764 36370
rect 1708 35700 1764 36318
rect 2380 36372 2436 36382
rect 2380 36278 2436 36316
rect 2716 36370 2772 36540
rect 2716 36318 2718 36370
rect 2770 36318 2772 36370
rect 2716 36306 2772 36318
rect 3164 36372 3220 36382
rect 3164 36278 3220 36316
rect 2044 36260 2100 36270
rect 2044 36166 2100 36204
rect 5292 36260 5348 38780
rect 5404 37940 5460 39564
rect 5964 39506 6020 39564
rect 6076 39618 6132 39676
rect 6524 39666 6580 39676
rect 6076 39566 6078 39618
rect 6130 39566 6132 39618
rect 6076 39554 6132 39566
rect 5964 39454 5966 39506
rect 6018 39454 6020 39506
rect 5964 39442 6020 39454
rect 5740 39396 5796 39406
rect 6412 39396 6468 39406
rect 5740 39394 5908 39396
rect 5740 39342 5742 39394
rect 5794 39342 5908 39394
rect 5740 39340 5908 39342
rect 5740 39330 5796 39340
rect 5740 38836 5796 38846
rect 5852 38836 5908 39340
rect 6076 39394 6468 39396
rect 6076 39342 6414 39394
rect 6466 39342 6468 39394
rect 6076 39340 6468 39342
rect 5964 38836 6020 38846
rect 5852 38780 5964 38836
rect 5740 38668 5796 38780
rect 5964 38742 6020 38780
rect 5404 37874 5460 37884
rect 5516 38610 5572 38622
rect 5516 38558 5518 38610
rect 5570 38558 5572 38610
rect 5292 36194 5348 36204
rect 5516 35812 5572 38558
rect 5628 38610 5684 38622
rect 5740 38612 5908 38668
rect 5628 38558 5630 38610
rect 5682 38558 5684 38610
rect 5628 38500 5684 38558
rect 5852 38610 6020 38612
rect 5852 38558 5854 38610
rect 5906 38558 6020 38610
rect 5852 38556 6020 38558
rect 5852 38546 5908 38556
rect 5628 38434 5684 38444
rect 5852 38276 5908 38286
rect 5852 37266 5908 38220
rect 5852 37214 5854 37266
rect 5906 37214 5908 37266
rect 5852 37202 5908 37214
rect 5964 38050 6020 38556
rect 6076 38276 6132 39340
rect 6412 39330 6468 39340
rect 6188 39172 6244 39182
rect 6244 39116 6468 39172
rect 6188 39106 6244 39116
rect 6412 38946 6468 39116
rect 6412 38894 6414 38946
rect 6466 38894 6468 38946
rect 6412 38882 6468 38894
rect 6188 38612 6244 38622
rect 6524 38612 6580 38622
rect 6244 38610 6580 38612
rect 6244 38558 6526 38610
rect 6578 38558 6580 38610
rect 6244 38556 6580 38558
rect 6188 38546 6244 38556
rect 6076 38210 6132 38220
rect 6188 38388 6244 38398
rect 6188 38274 6244 38332
rect 6188 38222 6190 38274
rect 6242 38222 6244 38274
rect 6188 38210 6244 38222
rect 5964 37998 5966 38050
rect 6018 37998 6020 38050
rect 5964 37266 6020 37998
rect 5964 37214 5966 37266
rect 6018 37214 6020 37266
rect 5964 37202 6020 37214
rect 6076 37940 6132 37950
rect 6076 37044 6132 37884
rect 6300 37828 6356 38556
rect 6524 38546 6580 38556
rect 6412 38050 6468 38062
rect 6412 37998 6414 38050
rect 6466 37998 6468 38050
rect 6412 37940 6468 37998
rect 6412 37874 6468 37884
rect 6524 37938 6580 37950
rect 6524 37886 6526 37938
rect 6578 37886 6580 37938
rect 6188 37772 6356 37828
rect 6188 37266 6244 37772
rect 6412 37604 6468 37614
rect 6300 37492 6356 37502
rect 6412 37492 6468 37548
rect 6300 37490 6468 37492
rect 6300 37438 6302 37490
rect 6354 37438 6468 37490
rect 6300 37436 6468 37438
rect 6300 37426 6356 37436
rect 6524 37380 6580 37886
rect 6524 37314 6580 37324
rect 6188 37214 6190 37266
rect 6242 37214 6244 37266
rect 6188 37202 6244 37214
rect 6412 37044 6468 37054
rect 6076 37042 6468 37044
rect 6076 36990 6414 37042
rect 6466 36990 6468 37042
rect 6076 36988 6468 36990
rect 6412 36978 6468 36988
rect 6636 36596 6692 42812
rect 6748 42754 6804 45164
rect 8204 44322 8260 45836
rect 8428 45798 8484 45836
rect 8204 44270 8206 44322
rect 8258 44270 8260 44322
rect 8204 44258 8260 44270
rect 8764 43708 8820 55132
rect 14588 54516 14644 55358
rect 20748 55410 20804 55422
rect 20748 55358 20750 55410
rect 20802 55358 20804 55410
rect 17500 55300 17556 55310
rect 17948 55300 18004 55310
rect 17500 55298 18004 55300
rect 17500 55246 17502 55298
rect 17554 55246 17950 55298
rect 18002 55246 18004 55298
rect 17500 55244 18004 55246
rect 17500 55234 17556 55244
rect 16716 55186 16772 55198
rect 16716 55134 16718 55186
rect 16770 55134 16772 55186
rect 16716 54738 16772 55134
rect 17724 54740 17780 54750
rect 16716 54686 16718 54738
rect 16770 54686 16772 54738
rect 16716 54674 16772 54686
rect 16828 54738 17780 54740
rect 16828 54686 17726 54738
rect 17778 54686 17780 54738
rect 16828 54684 17780 54686
rect 16828 54626 16884 54684
rect 17724 54674 17780 54684
rect 16828 54574 16830 54626
rect 16882 54574 16884 54626
rect 16828 54562 16884 54574
rect 14588 54450 14644 54460
rect 17052 54516 17108 54526
rect 15596 53844 15652 53854
rect 13804 53732 13860 53742
rect 13580 53730 13860 53732
rect 13580 53678 13806 53730
rect 13858 53678 13860 53730
rect 13580 53676 13860 53678
rect 13580 52164 13636 53676
rect 13804 53666 13860 53676
rect 14588 53620 14644 53630
rect 14588 53526 14644 53564
rect 15484 53620 15540 53630
rect 15484 53170 15540 53564
rect 15484 53118 15486 53170
rect 15538 53118 15540 53170
rect 15484 53106 15540 53118
rect 15596 53058 15652 53788
rect 16716 53844 16772 53854
rect 16716 53842 16884 53844
rect 16716 53790 16718 53842
rect 16770 53790 16884 53842
rect 16716 53788 16884 53790
rect 16716 53778 16772 53788
rect 16828 53508 16884 53788
rect 16828 53442 16884 53452
rect 17052 53618 17108 54460
rect 17500 54514 17556 54526
rect 17500 54462 17502 54514
rect 17554 54462 17556 54514
rect 17388 53844 17444 53854
rect 17388 53750 17444 53788
rect 17500 53732 17556 54462
rect 17612 54516 17668 54526
rect 17612 54422 17668 54460
rect 17836 54514 17892 54526
rect 17836 54462 17838 54514
rect 17890 54462 17892 54514
rect 17612 53732 17668 53742
rect 17500 53676 17612 53732
rect 17612 53638 17668 53676
rect 17052 53566 17054 53618
rect 17106 53566 17108 53618
rect 15596 53006 15598 53058
rect 15650 53006 15652 53058
rect 15596 52994 15652 53006
rect 16940 52836 16996 52846
rect 16380 52276 16436 52286
rect 13468 52162 13636 52164
rect 13468 52110 13582 52162
rect 13634 52110 13636 52162
rect 13468 52108 13636 52110
rect 12908 50484 12964 50494
rect 10108 49924 10164 49934
rect 10108 49026 10164 49868
rect 12236 49924 12292 49934
rect 12236 49810 12292 49868
rect 12908 49922 12964 50428
rect 12908 49870 12910 49922
rect 12962 49870 12964 49922
rect 12908 49858 12964 49870
rect 13468 49924 13524 52108
rect 13580 52098 13636 52108
rect 16044 52274 16436 52276
rect 16044 52222 16382 52274
rect 16434 52222 16436 52274
rect 16044 52220 16436 52222
rect 14252 52052 14308 52062
rect 14252 52050 14532 52052
rect 14252 51998 14254 52050
rect 14306 51998 14532 52050
rect 14252 51996 14532 51998
rect 14252 51986 14308 51996
rect 14476 51602 14532 51996
rect 14476 51550 14478 51602
rect 14530 51550 14532 51602
rect 14476 51538 14532 51550
rect 16044 51602 16100 52220
rect 16380 52210 16436 52220
rect 16828 52162 16884 52174
rect 16828 52110 16830 52162
rect 16882 52110 16884 52162
rect 16044 51550 16046 51602
rect 16098 51550 16100 51602
rect 15820 51380 15876 51390
rect 15708 51378 15876 51380
rect 15708 51326 15822 51378
rect 15874 51326 15876 51378
rect 15708 51324 15876 51326
rect 14588 51268 14644 51278
rect 14588 51174 14644 51212
rect 14700 50820 14756 50830
rect 13692 50708 13748 50718
rect 13692 50614 13748 50652
rect 13580 50484 13636 50494
rect 13580 50390 13636 50428
rect 13468 49858 13524 49868
rect 14028 49924 14084 49934
rect 12236 49758 12238 49810
rect 12290 49758 12292 49810
rect 12236 49746 12292 49758
rect 13356 49812 13412 49822
rect 11564 49700 11620 49710
rect 11564 49698 11732 49700
rect 11564 49646 11566 49698
rect 11618 49646 11732 49698
rect 11564 49644 11732 49646
rect 11564 49634 11620 49644
rect 11452 49588 11508 49598
rect 10780 49586 11508 49588
rect 10780 49534 11454 49586
rect 11506 49534 11508 49586
rect 10780 49532 11508 49534
rect 10780 49138 10836 49532
rect 11452 49522 11508 49532
rect 10780 49086 10782 49138
rect 10834 49086 10836 49138
rect 10780 49074 10836 49086
rect 10108 48974 10110 49026
rect 10162 48974 10164 49026
rect 10108 48692 10164 48974
rect 9660 48636 10164 48692
rect 9660 47458 9716 48636
rect 11676 48468 11732 49644
rect 12908 49138 12964 49150
rect 12908 49086 12910 49138
rect 12962 49086 12964 49138
rect 12236 48916 12292 48926
rect 12124 48468 12180 48478
rect 11676 48466 12180 48468
rect 11676 48414 12126 48466
rect 12178 48414 12180 48466
rect 11676 48412 12180 48414
rect 12124 48402 12180 48412
rect 12236 48466 12292 48860
rect 12236 48414 12238 48466
rect 12290 48414 12292 48466
rect 11788 48244 11844 48254
rect 9660 47406 9662 47458
rect 9714 47406 9716 47458
rect 9660 47012 9716 47406
rect 11564 48242 11844 48244
rect 11564 48190 11790 48242
rect 11842 48190 11844 48242
rect 11564 48188 11844 48190
rect 10332 47348 10388 47358
rect 10332 47346 10948 47348
rect 10332 47294 10334 47346
rect 10386 47294 10948 47346
rect 10332 47292 10948 47294
rect 10332 47282 10388 47292
rect 9660 46946 9716 46956
rect 10892 46898 10948 47292
rect 10892 46846 10894 46898
rect 10946 46846 10948 46898
rect 10892 46834 10948 46846
rect 11004 46788 11060 46798
rect 11004 46694 11060 46732
rect 11564 46674 11620 48188
rect 11788 48178 11844 48188
rect 12012 48244 12068 48254
rect 12012 48150 12068 48188
rect 12236 48020 12292 48414
rect 11900 47964 12292 48020
rect 12460 48242 12516 48254
rect 12460 48190 12462 48242
rect 12514 48190 12516 48242
rect 11900 46898 11956 47964
rect 11900 46846 11902 46898
rect 11954 46846 11956 46898
rect 11900 46834 11956 46846
rect 12460 47570 12516 48190
rect 12908 48244 12964 49086
rect 13356 48916 13412 49756
rect 13356 48468 13412 48860
rect 12908 48130 12964 48188
rect 12908 48078 12910 48130
rect 12962 48078 12964 48130
rect 12908 47796 12964 48078
rect 12908 47730 12964 47740
rect 13020 48466 13412 48468
rect 13020 48414 13358 48466
rect 13410 48414 13412 48466
rect 13020 48412 13412 48414
rect 12460 47518 12462 47570
rect 12514 47518 12516 47570
rect 11788 46788 11844 46798
rect 11788 46694 11844 46732
rect 11564 46622 11566 46674
rect 11618 46622 11620 46674
rect 9884 46564 9940 46574
rect 9884 46470 9940 46508
rect 9772 46452 9828 46462
rect 9100 46450 9828 46452
rect 9100 46398 9774 46450
rect 9826 46398 9828 46450
rect 9100 46396 9828 46398
rect 9100 46002 9156 46396
rect 9772 46386 9828 46396
rect 9100 45950 9102 46002
rect 9154 45950 9156 46002
rect 9100 45938 9156 45950
rect 11228 46004 11284 46014
rect 11228 45910 11284 45948
rect 11564 45892 11620 46622
rect 11340 45890 11620 45892
rect 11340 45838 11566 45890
rect 11618 45838 11620 45890
rect 11340 45836 11620 45838
rect 11340 45780 11396 45836
rect 11564 45826 11620 45836
rect 11676 46676 11732 46686
rect 10668 45724 11396 45780
rect 10668 45332 10724 45724
rect 10220 45330 10724 45332
rect 10220 45278 10670 45330
rect 10722 45278 10724 45330
rect 10220 45276 10724 45278
rect 9772 44996 9828 45006
rect 9772 44902 9828 44940
rect 9660 44884 9716 44894
rect 8876 44882 9716 44884
rect 8876 44830 9662 44882
rect 9714 44830 9716 44882
rect 8876 44828 9716 44830
rect 8876 44434 8932 44828
rect 9660 44818 9716 44828
rect 8876 44382 8878 44434
rect 8930 44382 8932 44434
rect 8876 44370 8932 44382
rect 10108 44660 10164 44670
rect 6748 42702 6750 42754
rect 6802 42702 6804 42754
rect 6748 42690 6804 42702
rect 6860 43652 6916 43662
rect 8764 43652 9716 43708
rect 6860 42642 6916 43596
rect 8092 43540 8148 43550
rect 7868 43426 7924 43438
rect 7868 43374 7870 43426
rect 7922 43374 7924 43426
rect 7868 42980 7924 43374
rect 7868 42914 7924 42924
rect 6860 42590 6862 42642
rect 6914 42590 6916 42642
rect 6860 42578 6916 42590
rect 7532 42644 7588 42654
rect 7532 42550 7588 42588
rect 8092 42642 8148 43484
rect 8652 43540 8708 43550
rect 8652 43446 8708 43484
rect 8204 43428 8260 43438
rect 8204 42868 8260 43372
rect 8876 42868 8932 42878
rect 8204 42866 8932 42868
rect 8204 42814 8878 42866
rect 8930 42814 8932 42866
rect 8204 42812 8932 42814
rect 8316 42754 8372 42812
rect 8876 42802 8932 42812
rect 8316 42702 8318 42754
rect 8370 42702 8372 42754
rect 8316 42690 8372 42702
rect 8092 42590 8094 42642
rect 8146 42590 8148 42642
rect 8092 42578 8148 42590
rect 8764 42644 8820 42654
rect 8764 42550 8820 42588
rect 7644 42530 7700 42542
rect 7644 42478 7646 42530
rect 7698 42478 7700 42530
rect 7084 42196 7140 42206
rect 7084 42082 7140 42140
rect 7084 42030 7086 42082
rect 7138 42030 7140 42082
rect 7084 42018 7140 42030
rect 7644 41186 7700 42478
rect 8204 42084 8260 42094
rect 8204 42082 8372 42084
rect 8204 42030 8206 42082
rect 8258 42030 8372 42082
rect 8204 42028 8372 42030
rect 8204 42018 8260 42028
rect 8092 41970 8148 41982
rect 8092 41918 8094 41970
rect 8146 41918 8148 41970
rect 8092 41412 8148 41918
rect 8092 41346 8148 41356
rect 8204 41746 8260 41758
rect 8204 41694 8206 41746
rect 8258 41694 8260 41746
rect 7644 41134 7646 41186
rect 7698 41134 7700 41186
rect 7644 41122 7700 41134
rect 8204 41186 8260 41694
rect 8204 41134 8206 41186
rect 8258 41134 8260 41186
rect 8204 41122 8260 41134
rect 8316 40516 8372 42028
rect 8652 41860 8708 41870
rect 8540 41858 8708 41860
rect 8540 41806 8654 41858
rect 8706 41806 8708 41858
rect 8540 41804 8708 41806
rect 8540 40628 8596 41804
rect 8652 41794 8708 41804
rect 8764 41748 8820 41758
rect 8764 41746 9268 41748
rect 8764 41694 8766 41746
rect 8818 41694 9268 41746
rect 8764 41692 9268 41694
rect 8764 41682 8820 41692
rect 8652 41076 8708 41086
rect 8652 41074 8820 41076
rect 8652 41022 8654 41074
rect 8706 41022 8820 41074
rect 8652 41020 8820 41022
rect 8652 41010 8708 41020
rect 8652 40628 8708 40638
rect 8540 40626 8708 40628
rect 8540 40574 8654 40626
rect 8706 40574 8708 40626
rect 8540 40572 8708 40574
rect 8652 40562 8708 40572
rect 7420 40460 7812 40516
rect 7420 40290 7476 40460
rect 7756 40404 7812 40460
rect 7980 40460 8316 40516
rect 7868 40404 7924 40414
rect 7756 40402 7924 40404
rect 7756 40350 7870 40402
rect 7922 40350 7924 40402
rect 7756 40348 7924 40350
rect 7868 40338 7924 40348
rect 7420 40238 7422 40290
rect 7474 40238 7476 40290
rect 7420 40226 7476 40238
rect 7644 40292 7700 40302
rect 7084 39730 7140 39742
rect 7084 39678 7086 39730
rect 7138 39678 7140 39730
rect 7084 39620 7140 39678
rect 7084 39554 7140 39564
rect 7644 39060 7700 40236
rect 7756 40180 7812 40190
rect 7980 40180 8036 40460
rect 8316 40450 8372 40460
rect 7756 40178 8036 40180
rect 7756 40126 7758 40178
rect 7810 40126 8036 40178
rect 7756 40124 8036 40126
rect 8316 40178 8372 40190
rect 8316 40126 8318 40178
rect 8370 40126 8372 40178
rect 7756 40114 7812 40124
rect 7644 39058 8036 39060
rect 7644 39006 7646 39058
rect 7698 39006 8036 39058
rect 7644 39004 8036 39006
rect 7644 38994 7700 39004
rect 6860 38836 6916 38846
rect 6860 38742 6916 38780
rect 6748 38724 6804 38734
rect 6748 38630 6804 38668
rect 7980 38052 8036 39004
rect 8092 38052 8148 38062
rect 7980 38050 8148 38052
rect 7980 37998 8094 38050
rect 8146 37998 8148 38050
rect 7980 37996 8148 37998
rect 7308 37938 7364 37950
rect 7308 37886 7310 37938
rect 7362 37886 7364 37938
rect 7308 37604 7364 37886
rect 7644 37940 7700 37950
rect 7644 37846 7700 37884
rect 7308 37538 7364 37548
rect 7532 37604 7588 37614
rect 6972 37380 7028 37390
rect 6972 37286 7028 37324
rect 7308 37378 7364 37390
rect 7308 37326 7310 37378
rect 7362 37326 7364 37378
rect 6636 36530 6692 36540
rect 7308 36596 7364 37326
rect 7308 36530 7364 36540
rect 5852 35812 5908 35822
rect 5516 35810 5908 35812
rect 5516 35758 5854 35810
rect 5906 35758 5908 35810
rect 5516 35756 5908 35758
rect 5852 35746 5908 35756
rect 1708 35634 1764 35644
rect 4284 35700 4340 35710
rect 4284 35606 4340 35644
rect 5180 35698 5236 35710
rect 5180 35646 5182 35698
rect 5234 35646 5236 35698
rect 5180 35588 5236 35646
rect 7532 35700 7588 37548
rect 7756 36484 7812 36494
rect 8092 36484 8148 37996
rect 7756 36482 8148 36484
rect 7756 36430 7758 36482
rect 7810 36430 8148 36482
rect 7756 36428 8148 36430
rect 7756 36418 7812 36428
rect 7532 35634 7588 35644
rect 7980 35812 8036 35822
rect 5068 35532 5180 35588
rect 1932 35474 1988 35486
rect 1932 35422 1934 35474
rect 1986 35422 1988 35474
rect 1932 35028 1988 35422
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 1932 34962 1988 34972
rect 1932 34132 1988 34142
rect 1820 34020 1876 34030
rect 1708 34018 1876 34020
rect 1708 33966 1822 34018
rect 1874 33966 1876 34018
rect 1708 33964 1876 33966
rect 1708 32340 1764 33964
rect 1820 33954 1876 33964
rect 1932 33346 1988 34076
rect 4284 34132 4340 34142
rect 4732 34132 4788 34142
rect 5068 34132 5124 35532
rect 5180 35522 5236 35532
rect 7980 35586 8036 35756
rect 7980 35534 7982 35586
rect 8034 35534 8036 35586
rect 7980 35522 8036 35534
rect 8092 35588 8148 36428
rect 8316 35812 8372 40126
rect 8540 40178 8596 40190
rect 8540 40126 8542 40178
rect 8594 40126 8596 40178
rect 8540 40068 8596 40126
rect 8764 40180 8820 41020
rect 8764 40114 8820 40124
rect 9100 40964 9156 40974
rect 8540 40002 8596 40012
rect 8988 40068 9044 40078
rect 8988 39058 9044 40012
rect 8988 39006 8990 39058
rect 9042 39006 9044 39058
rect 8988 38994 9044 39006
rect 9100 38836 9156 40908
rect 9212 39730 9268 41692
rect 9212 39678 9214 39730
rect 9266 39678 9268 39730
rect 9212 39666 9268 39678
rect 9548 40402 9604 40414
rect 9548 40350 9550 40402
rect 9602 40350 9604 40402
rect 9548 40292 9604 40350
rect 9548 39620 9604 40236
rect 9548 39554 9604 39564
rect 8988 38780 9156 38836
rect 8988 38668 9044 38780
rect 8988 38612 9268 38668
rect 8764 37940 8820 37950
rect 8764 37846 8820 37884
rect 8428 36596 8484 36606
rect 8428 36502 8484 36540
rect 8316 35746 8372 35756
rect 8428 35588 8484 35598
rect 8092 35532 8428 35588
rect 5852 34802 5908 34814
rect 5852 34750 5854 34802
rect 5906 34750 5908 34802
rect 5516 34692 5572 34702
rect 4284 34130 5068 34132
rect 4284 34078 4286 34130
rect 4338 34078 4734 34130
rect 4786 34078 5068 34130
rect 4284 34076 5068 34078
rect 4284 34066 4340 34076
rect 4732 34066 4788 34076
rect 5068 34038 5124 34076
rect 5180 34690 5572 34692
rect 5180 34638 5518 34690
rect 5570 34638 5572 34690
rect 5180 34636 5572 34638
rect 1932 33294 1934 33346
rect 1986 33294 1988 33346
rect 1820 32564 1876 32574
rect 1932 32564 1988 33294
rect 4284 33908 4340 33918
rect 2604 33236 2660 33246
rect 2604 33234 3108 33236
rect 2604 33182 2606 33234
rect 2658 33182 3108 33234
rect 2604 33180 3108 33182
rect 2604 33170 2660 33180
rect 1820 32562 1988 32564
rect 1820 32510 1822 32562
rect 1874 32510 1988 32562
rect 1820 32508 1988 32510
rect 1820 32498 1876 32508
rect 1708 31778 1764 32284
rect 2492 32450 2548 32462
rect 2492 32398 2494 32450
rect 2546 32398 2548 32450
rect 2492 31948 2548 32398
rect 2492 31892 2884 31948
rect 2828 31890 2884 31892
rect 2828 31838 2830 31890
rect 2882 31838 2884 31890
rect 2828 31826 2884 31838
rect 3052 31892 3108 33180
rect 3052 31826 3108 31836
rect 3388 31892 3444 31902
rect 1708 31726 1710 31778
rect 1762 31726 1764 31778
rect 1708 31714 1764 31726
rect 2940 31668 2996 31678
rect 2940 31574 2996 31612
rect 2044 31556 2100 31566
rect 2044 31462 2100 31500
rect 2716 31556 2772 31566
rect 3164 31556 3220 31566
rect 2716 31554 2884 31556
rect 2716 31502 2718 31554
rect 2770 31502 2884 31554
rect 2716 31500 2884 31502
rect 2716 31490 2772 31500
rect 1820 31220 1876 31230
rect 1820 30994 1876 31164
rect 2044 31108 2100 31118
rect 2044 31014 2100 31052
rect 2716 31106 2772 31118
rect 2716 31054 2718 31106
rect 2770 31054 2772 31106
rect 1820 30942 1822 30994
rect 1874 30942 1876 30994
rect 1820 30930 1876 30942
rect 2380 30996 2436 31006
rect 2380 30902 2436 30940
rect 2716 30772 2772 31054
rect 2716 30706 2772 30716
rect 1820 30210 1876 30222
rect 1820 30158 1822 30210
rect 1874 30158 1876 30210
rect 1708 29428 1764 29438
rect 1708 29334 1764 29372
rect 1820 28642 1876 30158
rect 2828 30212 2884 31500
rect 3164 31462 3220 31500
rect 3388 31444 3444 31836
rect 4060 31892 4116 31902
rect 3724 31780 3780 31790
rect 3612 31724 3724 31780
rect 3612 31666 3668 31724
rect 3724 31714 3780 31724
rect 3612 31614 3614 31666
rect 3666 31614 3668 31666
rect 3612 31602 3668 31614
rect 3836 31668 3892 31678
rect 3724 31554 3780 31566
rect 3724 31502 3726 31554
rect 3778 31502 3780 31554
rect 3724 31444 3780 31502
rect 3388 31388 3780 31444
rect 3388 31106 3444 31118
rect 3836 31108 3892 31612
rect 4060 31666 4116 31836
rect 4060 31614 4062 31666
rect 4114 31614 4116 31666
rect 4060 31602 4116 31614
rect 3388 31054 3390 31106
rect 3442 31054 3444 31106
rect 3052 30994 3108 31006
rect 3052 30942 3054 30994
rect 3106 30942 3108 30994
rect 3052 30884 3108 30942
rect 3052 30324 3108 30828
rect 3052 30258 3108 30268
rect 3164 30996 3220 31006
rect 2828 30146 2884 30156
rect 2492 30100 2548 30110
rect 2492 30006 2548 30044
rect 2044 29652 2100 29662
rect 2044 29558 2100 29596
rect 3164 29650 3220 30940
rect 3388 30436 3444 31054
rect 3388 30370 3444 30380
rect 3724 31052 3892 31108
rect 3164 29598 3166 29650
rect 3218 29598 3220 29650
rect 3164 29586 3220 29598
rect 3612 30100 3668 30110
rect 3612 29650 3668 30044
rect 3612 29598 3614 29650
rect 3666 29598 3668 29650
rect 3612 29586 3668 29598
rect 3724 29650 3780 31052
rect 4172 30996 4228 31006
rect 4284 30996 4340 33852
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4732 33460 4788 33470
rect 4732 33366 4788 33404
rect 4620 32676 4676 32686
rect 4620 32452 4676 32620
rect 4620 32450 4900 32452
rect 4620 32398 4622 32450
rect 4674 32398 4900 32450
rect 4620 32396 4900 32398
rect 4620 32386 4676 32396
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4620 31780 4676 31790
rect 4620 31686 4676 31724
rect 4844 31780 4900 32396
rect 5180 32004 5236 34636
rect 5516 34626 5572 34636
rect 5740 34690 5796 34702
rect 5740 34638 5742 34690
rect 5794 34638 5796 34690
rect 5628 34132 5684 34142
rect 5404 34020 5460 34030
rect 5404 34018 5572 34020
rect 5404 33966 5406 34018
rect 5458 33966 5572 34018
rect 5404 33964 5572 33966
rect 5404 33954 5460 33964
rect 5516 33570 5572 33964
rect 5516 33518 5518 33570
rect 5570 33518 5572 33570
rect 5516 33506 5572 33518
rect 5292 33460 5348 33470
rect 5292 32562 5348 33404
rect 5404 32676 5460 32686
rect 5404 32582 5460 32620
rect 5292 32510 5294 32562
rect 5346 32510 5348 32562
rect 5292 32004 5348 32510
rect 5404 32004 5460 32014
rect 5292 31948 5404 32004
rect 5180 31938 5236 31948
rect 5404 31938 5460 31948
rect 4844 31778 5012 31780
rect 4844 31726 4846 31778
rect 4898 31726 5012 31778
rect 4844 31724 5012 31726
rect 4844 31714 4900 31724
rect 4508 31668 4564 31678
rect 4508 31574 4564 31612
rect 4732 31556 4788 31566
rect 4732 31218 4788 31500
rect 4732 31166 4734 31218
rect 4786 31166 4788 31218
rect 4732 31154 4788 31166
rect 4956 31218 5012 31724
rect 5068 31666 5124 31678
rect 5068 31614 5070 31666
rect 5122 31614 5124 31666
rect 5068 31556 5124 31614
rect 5068 31490 5124 31500
rect 5516 31668 5572 31678
rect 4956 31166 4958 31218
rect 5010 31166 5012 31218
rect 4956 31154 5012 31166
rect 4172 30994 4340 30996
rect 4172 30942 4174 30994
rect 4226 30942 4340 30994
rect 4172 30940 4340 30942
rect 4508 31106 4564 31118
rect 4508 31054 4510 31106
rect 4562 31054 4564 31106
rect 4508 30996 4564 31054
rect 5068 30996 5124 31006
rect 4508 30994 5124 30996
rect 4508 30942 5070 30994
rect 5122 30942 5124 30994
rect 4508 30940 5124 30942
rect 3724 29598 3726 29650
rect 3778 29598 3780 29650
rect 2716 29540 2772 29550
rect 2716 29446 2772 29484
rect 2380 29426 2436 29438
rect 2380 29374 2382 29426
rect 2434 29374 2436 29426
rect 2380 29316 2436 29374
rect 2380 28980 2436 29260
rect 2380 28914 2436 28924
rect 3164 29428 3220 29438
rect 1820 28590 1822 28642
rect 1874 28590 1876 28642
rect 1708 28420 1764 28430
rect 1708 27970 1764 28364
rect 1708 27918 1710 27970
rect 1762 27918 1764 27970
rect 1708 27906 1764 27918
rect 1708 27412 1764 27422
rect 1708 27074 1764 27356
rect 1708 27022 1710 27074
rect 1762 27022 1764 27074
rect 1708 26964 1764 27022
rect 1708 26898 1764 26908
rect 1820 26290 1876 28590
rect 2492 28532 2548 28542
rect 2492 28438 2548 28476
rect 2716 28084 2772 28094
rect 2716 27990 2772 28028
rect 3164 28082 3220 29372
rect 3500 29426 3556 29438
rect 3500 29374 3502 29426
rect 3554 29374 3556 29426
rect 3500 28308 3556 29374
rect 3500 28242 3556 28252
rect 3612 28532 3668 28542
rect 3164 28030 3166 28082
rect 3218 28030 3220 28082
rect 3164 28018 3220 28030
rect 3612 28082 3668 28476
rect 3612 28030 3614 28082
rect 3666 28030 3668 28082
rect 3612 28018 3668 28030
rect 3724 28082 3780 29598
rect 3724 28030 3726 28082
rect 3778 28030 3780 28082
rect 2044 27970 2100 27982
rect 2044 27918 2046 27970
rect 2098 27918 2100 27970
rect 2044 27748 2100 27918
rect 3276 27972 3332 27982
rect 2492 27860 2548 27870
rect 2492 27858 2660 27860
rect 2492 27806 2494 27858
rect 2546 27806 2660 27858
rect 2492 27804 2660 27806
rect 2492 27794 2548 27804
rect 2044 27682 2100 27692
rect 2604 27636 2660 27804
rect 2044 27300 2100 27310
rect 2044 26962 2100 27244
rect 2044 26910 2046 26962
rect 2098 26910 2100 26962
rect 2044 26898 2100 26910
rect 2492 27074 2548 27086
rect 2492 27022 2494 27074
rect 2546 27022 2548 27074
rect 2492 26964 2548 27022
rect 1820 26238 1822 26290
rect 1874 26238 1876 26290
rect 1596 25844 1652 25854
rect 1596 17332 1652 25788
rect 1708 25620 1764 25630
rect 1708 25506 1764 25564
rect 1708 25454 1710 25506
rect 1762 25454 1764 25506
rect 1708 25442 1764 25454
rect 1820 25284 1876 26238
rect 1708 24948 1764 24958
rect 1708 24722 1764 24892
rect 1708 24670 1710 24722
rect 1762 24670 1764 24722
rect 1708 24052 1764 24670
rect 1708 23986 1764 23996
rect 1820 23938 1876 25228
rect 2044 26516 2100 26526
rect 2044 24946 2100 26460
rect 2492 26404 2548 26908
rect 2492 26338 2548 26348
rect 2492 26180 2548 26190
rect 2492 26086 2548 26124
rect 2268 25732 2324 25742
rect 2268 25618 2324 25676
rect 2268 25566 2270 25618
rect 2322 25566 2324 25618
rect 2268 25554 2324 25566
rect 2604 25620 2660 27580
rect 2716 27188 2772 27198
rect 2716 26962 2772 27132
rect 2716 26910 2718 26962
rect 2770 26910 2772 26962
rect 2716 26898 2772 26910
rect 3276 26962 3332 27916
rect 3724 27972 3780 28030
rect 3724 27906 3780 27916
rect 3836 30884 3892 30894
rect 4172 30884 4228 30940
rect 3836 30882 4228 30884
rect 3836 30830 3838 30882
rect 3890 30830 4228 30882
rect 3836 30828 4228 30830
rect 3500 27860 3556 27870
rect 3500 27858 3668 27860
rect 3500 27806 3502 27858
rect 3554 27806 3668 27858
rect 3500 27804 3668 27806
rect 3500 27794 3556 27804
rect 3276 26910 3278 26962
rect 3330 26910 3332 26962
rect 3276 26898 3332 26910
rect 3388 27412 3444 27422
rect 2604 25554 2660 25564
rect 3164 25506 3220 25518
rect 3388 25508 3444 27356
rect 3612 27188 3668 27804
rect 3724 27188 3780 27198
rect 3612 27132 3724 27188
rect 3724 27122 3780 27132
rect 3500 27074 3556 27086
rect 3500 27022 3502 27074
rect 3554 27022 3556 27074
rect 3500 26628 3556 27022
rect 3500 26562 3556 26572
rect 3836 26404 3892 30828
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4620 30324 4676 30334
rect 4508 30322 4676 30324
rect 4508 30270 4622 30322
rect 4674 30270 4676 30322
rect 4508 30268 4676 30270
rect 4508 30100 4564 30268
rect 4620 30258 4676 30268
rect 4284 29538 4340 29550
rect 4284 29486 4286 29538
rect 4338 29486 4340 29538
rect 4172 29428 4228 29438
rect 4284 29428 4340 29486
rect 4172 29426 4340 29428
rect 4172 29374 4174 29426
rect 4226 29374 4340 29426
rect 4172 29372 4340 29374
rect 4508 29538 4564 30044
rect 4508 29486 4510 29538
rect 4562 29486 4564 29538
rect 4172 29362 4228 29372
rect 4508 29204 4564 29486
rect 4620 29428 4676 29438
rect 4956 29428 5012 30940
rect 5068 30930 5124 30940
rect 5516 30210 5572 31612
rect 5628 31218 5684 34076
rect 5740 33460 5796 34638
rect 5852 33908 5908 34750
rect 7980 34356 8036 34366
rect 8092 34356 8148 35532
rect 8428 35494 8484 35532
rect 7644 34354 8148 34356
rect 7644 34302 7982 34354
rect 8034 34302 8148 34354
rect 7644 34300 8148 34302
rect 7532 34018 7588 34030
rect 7532 33966 7534 34018
rect 7586 33966 7588 34018
rect 5852 33842 5908 33852
rect 7196 33908 7252 33918
rect 5852 33572 5908 33582
rect 5852 33570 6244 33572
rect 5852 33518 5854 33570
rect 5906 33518 6244 33570
rect 5852 33516 6244 33518
rect 5852 33506 5908 33516
rect 5740 33394 5796 33404
rect 6188 33458 6244 33516
rect 7084 33460 7140 33470
rect 6188 33406 6190 33458
rect 6242 33406 6244 33458
rect 6188 33394 6244 33406
rect 6972 33404 7084 33460
rect 6636 33348 6692 33358
rect 6860 33348 6916 33358
rect 6636 33346 6916 33348
rect 6636 33294 6638 33346
rect 6690 33294 6862 33346
rect 6914 33294 6916 33346
rect 6636 33292 6916 33294
rect 6636 33282 6692 33292
rect 6860 33282 6916 33292
rect 5852 33124 5908 33134
rect 6076 33124 6132 33134
rect 5852 33030 5908 33068
rect 5964 33122 6132 33124
rect 5964 33070 6078 33122
rect 6130 33070 6132 33122
rect 5964 33068 6132 33070
rect 5628 31166 5630 31218
rect 5682 31166 5684 31218
rect 5628 31154 5684 31166
rect 5852 32450 5908 32462
rect 5852 32398 5854 32450
rect 5906 32398 5908 32450
rect 5516 30158 5518 30210
rect 5570 30158 5572 30210
rect 5516 30146 5572 30158
rect 5740 30212 5796 30222
rect 5740 30118 5796 30156
rect 5068 29988 5124 29998
rect 5068 29986 5236 29988
rect 5068 29934 5070 29986
rect 5122 29934 5236 29986
rect 5068 29932 5236 29934
rect 5068 29922 5124 29932
rect 4620 29426 5012 29428
rect 4620 29374 4622 29426
rect 4674 29374 5012 29426
rect 4620 29372 5012 29374
rect 4620 29362 4676 29372
rect 4508 29138 4564 29148
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4620 28756 4676 28766
rect 4620 28754 4788 28756
rect 4620 28702 4622 28754
rect 4674 28702 4788 28754
rect 4620 28700 4788 28702
rect 4620 28690 4676 28700
rect 3948 28532 4004 28542
rect 3948 27074 4004 28476
rect 4620 28308 4676 28318
rect 4620 28082 4676 28252
rect 4620 28030 4622 28082
rect 4674 28030 4676 28082
rect 4620 28018 4676 28030
rect 4172 27860 4228 27870
rect 4396 27860 4452 27870
rect 4172 27766 4228 27804
rect 4284 27858 4452 27860
rect 4284 27806 4398 27858
rect 4450 27806 4452 27858
rect 4284 27804 4452 27806
rect 4732 27860 4788 28700
rect 4844 28532 4900 29372
rect 5068 29316 5124 29326
rect 5068 29222 5124 29260
rect 5180 29316 5236 29932
rect 5516 29316 5572 29326
rect 5180 29314 5572 29316
rect 5180 29262 5518 29314
rect 5570 29262 5572 29314
rect 5180 29260 5572 29262
rect 4844 28466 4900 28476
rect 5068 28420 5124 28430
rect 5068 28326 5124 28364
rect 5068 27972 5124 27982
rect 5068 27878 5124 27916
rect 4844 27860 4900 27870
rect 4732 27858 4900 27860
rect 4732 27806 4846 27858
rect 4898 27806 4900 27858
rect 4732 27804 4900 27806
rect 3948 27022 3950 27074
rect 4002 27022 4004 27074
rect 3948 27010 4004 27022
rect 4284 27076 4340 27804
rect 4396 27794 4452 27804
rect 4844 27748 4900 27804
rect 4844 27682 4900 27692
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4508 27188 4564 27198
rect 4564 27132 4676 27188
rect 4508 27122 4564 27132
rect 4396 27076 4452 27086
rect 4284 27074 4452 27076
rect 4284 27022 4398 27074
rect 4450 27022 4452 27074
rect 4284 27020 4452 27022
rect 4396 26908 4452 27020
rect 4620 27074 4676 27132
rect 4620 27022 4622 27074
rect 4674 27022 4676 27074
rect 4620 27010 4676 27022
rect 4732 27074 4788 27086
rect 4732 27022 4734 27074
rect 4786 27022 4788 27074
rect 4060 26852 4116 26862
rect 4060 26758 4116 26796
rect 4284 26850 4340 26862
rect 4396 26852 4564 26908
rect 4284 26798 4286 26850
rect 4338 26798 4340 26850
rect 3164 25454 3166 25506
rect 3218 25454 3220 25506
rect 2716 25396 2772 25406
rect 2716 25302 2772 25340
rect 3164 25396 3220 25454
rect 3164 25330 3220 25340
rect 3276 25452 3444 25508
rect 3612 26348 3892 26404
rect 3948 26628 4004 26638
rect 3276 25060 3332 25452
rect 3388 25282 3444 25294
rect 3388 25230 3390 25282
rect 3442 25230 3444 25282
rect 3388 25172 3444 25230
rect 3500 25172 3556 25182
rect 3388 25116 3500 25172
rect 3500 25106 3556 25116
rect 3276 25004 3444 25060
rect 2044 24894 2046 24946
rect 2098 24894 2100 24946
rect 2044 24882 2100 24894
rect 2716 24948 2772 24958
rect 2716 24854 2772 24892
rect 2380 24724 2436 24734
rect 2380 24276 2436 24668
rect 2380 24210 2436 24220
rect 1820 23886 1822 23938
rect 1874 23886 1876 23938
rect 1708 23154 1764 23166
rect 1708 23102 1710 23154
rect 1762 23102 1764 23154
rect 1708 22932 1764 23102
rect 1708 22484 1764 22876
rect 1708 22418 1764 22428
rect 1820 22370 1876 23886
rect 2492 23826 2548 23838
rect 2492 23774 2494 23826
rect 2546 23774 2548 23826
rect 2492 23380 2548 23774
rect 2604 23380 2660 23390
rect 2492 23378 2660 23380
rect 2492 23326 2606 23378
rect 2658 23326 2660 23378
rect 2492 23324 2660 23326
rect 2604 23314 2660 23324
rect 2940 23156 2996 23166
rect 2940 23062 2996 23100
rect 3276 23154 3332 23166
rect 3276 23102 3278 23154
rect 3330 23102 3332 23154
rect 2268 23044 2324 23054
rect 2268 23042 2436 23044
rect 2268 22990 2270 23042
rect 2322 22990 2436 23042
rect 2268 22988 2436 22990
rect 2268 22978 2324 22988
rect 1820 22318 1822 22370
rect 1874 22318 1876 22370
rect 1708 22260 1764 22270
rect 1708 21812 1764 22204
rect 1708 21718 1764 21756
rect 1708 20916 1764 20926
rect 1708 20578 1764 20860
rect 1708 20526 1710 20578
rect 1762 20526 1764 20578
rect 1708 20244 1764 20526
rect 1708 20178 1764 20188
rect 1820 20018 1876 22318
rect 2268 21476 2324 21486
rect 2268 21382 2324 21420
rect 2380 21028 2436 22988
rect 2492 22258 2548 22270
rect 2492 22206 2494 22258
rect 2546 22206 2548 22258
rect 2492 21812 2548 22206
rect 2492 21746 2548 21756
rect 2940 22036 2996 22046
rect 2940 21810 2996 21980
rect 2940 21758 2942 21810
rect 2994 21758 2996 21810
rect 2940 21746 2996 21758
rect 2604 21588 2660 21598
rect 2604 21494 2660 21532
rect 3276 21364 3332 23102
rect 3388 21810 3444 25004
rect 3500 24948 3556 24958
rect 3612 24948 3668 26348
rect 3836 26180 3892 26190
rect 3724 26068 3780 26078
rect 3724 25506 3780 26012
rect 3836 25618 3892 26124
rect 3836 25566 3838 25618
rect 3890 25566 3892 25618
rect 3836 25554 3892 25566
rect 3724 25454 3726 25506
rect 3778 25454 3780 25506
rect 3724 25442 3780 25454
rect 3948 25508 4004 26572
rect 4060 26292 4116 26302
rect 4060 25732 4116 26236
rect 4060 25666 4116 25676
rect 3948 25452 4116 25508
rect 4060 25396 4116 25452
rect 4284 25506 4340 26798
rect 4508 26404 4564 26852
rect 4508 26338 4564 26348
rect 4732 26852 4788 27022
rect 5068 27076 5124 27086
rect 5068 26982 5124 27020
rect 4620 26180 4676 26190
rect 4732 26180 4788 26796
rect 4676 26124 4788 26180
rect 4844 26404 4900 26414
rect 4620 26086 4676 26124
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4844 25732 4900 26348
rect 5180 26292 5236 29260
rect 5516 29250 5572 29260
rect 5740 29204 5796 29214
rect 5628 28532 5684 28542
rect 5516 27972 5572 27982
rect 5404 27970 5572 27972
rect 5404 27918 5518 27970
rect 5570 27918 5572 27970
rect 5404 27916 5572 27918
rect 5292 27860 5348 27870
rect 5292 27766 5348 27804
rect 5404 27748 5460 27916
rect 5516 27906 5572 27916
rect 5628 27970 5684 28476
rect 5628 27918 5630 27970
rect 5682 27918 5684 27970
rect 5628 27906 5684 27918
rect 5740 27748 5796 29148
rect 5404 26908 5460 27692
rect 5628 27692 5796 27748
rect 5628 26908 5684 27692
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 4284 25442 4340 25454
rect 4620 25676 4900 25732
rect 4956 26236 5236 26292
rect 5292 26852 5460 26908
rect 5516 26852 5684 26908
rect 5740 26964 5796 26974
rect 5740 26870 5796 26908
rect 5852 26908 5908 32398
rect 5964 31892 6020 33068
rect 6076 33058 6132 33068
rect 6300 33124 6356 33134
rect 6300 32452 6356 33068
rect 6972 32900 7028 33404
rect 7084 33394 7140 33404
rect 7196 33346 7252 33852
rect 7196 33294 7198 33346
rect 7250 33294 7252 33346
rect 7196 33282 7252 33294
rect 6860 32844 7028 32900
rect 7084 33122 7140 33134
rect 7084 33070 7086 33122
rect 7138 33070 7140 33122
rect 6860 32674 6916 32844
rect 6860 32622 6862 32674
rect 6914 32622 6916 32674
rect 6860 32610 6916 32622
rect 6972 32676 7028 32686
rect 7084 32676 7140 33070
rect 7028 32620 7140 32676
rect 7532 32676 7588 33966
rect 7644 33346 7700 34300
rect 7980 34290 8036 34300
rect 8540 34242 8596 34254
rect 8540 34190 8542 34242
rect 8594 34190 8596 34242
rect 8316 34132 8372 34142
rect 7644 33294 7646 33346
rect 7698 33294 7700 33346
rect 7644 33282 7700 33294
rect 8092 34130 8372 34132
rect 8092 34078 8318 34130
rect 8370 34078 8372 34130
rect 8092 34076 8372 34078
rect 8092 32786 8148 34076
rect 8316 34066 8372 34076
rect 8540 33460 8596 34190
rect 8652 34130 8708 34142
rect 8652 34078 8654 34130
rect 8706 34078 8708 34130
rect 8652 33908 8708 34078
rect 8652 33842 8708 33852
rect 8540 33394 8596 33404
rect 8092 32734 8094 32786
rect 8146 32734 8148 32786
rect 8092 32722 8148 32734
rect 8316 33234 8372 33246
rect 8316 33182 8318 33234
rect 8370 33182 8372 33234
rect 8316 32788 8372 33182
rect 8428 32788 8484 32798
rect 8316 32786 8484 32788
rect 8316 32734 8430 32786
rect 8482 32734 8484 32786
rect 8316 32732 8484 32734
rect 8428 32722 8484 32732
rect 6972 32562 7028 32620
rect 7532 32610 7588 32620
rect 6972 32510 6974 32562
rect 7026 32510 7028 32562
rect 6972 32498 7028 32510
rect 8316 32562 8372 32574
rect 8316 32510 8318 32562
rect 8370 32510 8372 32562
rect 6300 32386 6356 32396
rect 7644 32452 7700 32462
rect 7644 32358 7700 32396
rect 8316 32452 8372 32510
rect 8540 32564 8596 32574
rect 8540 32470 8596 32508
rect 8316 32386 8372 32396
rect 9100 32450 9156 32462
rect 9100 32398 9102 32450
rect 9154 32398 9156 32450
rect 6188 32004 6244 32014
rect 6076 31892 6132 31902
rect 5964 31890 6132 31892
rect 5964 31838 6078 31890
rect 6130 31838 6132 31890
rect 5964 31836 6132 31838
rect 6076 31826 6132 31836
rect 6188 31778 6244 31948
rect 7644 32004 7700 32014
rect 7644 31890 7700 31948
rect 8876 31892 8932 31902
rect 7644 31838 7646 31890
rect 7698 31838 7700 31890
rect 7644 31826 7700 31838
rect 8764 31890 8932 31892
rect 8764 31838 8878 31890
rect 8930 31838 8932 31890
rect 8764 31836 8932 31838
rect 6188 31726 6190 31778
rect 6242 31726 6244 31778
rect 6188 31714 6244 31726
rect 6524 31780 6580 31790
rect 6524 31686 6580 31724
rect 8540 31778 8596 31790
rect 8540 31726 8542 31778
rect 8594 31726 8596 31778
rect 5964 31668 6020 31678
rect 5964 31574 6020 31612
rect 7756 31668 7812 31678
rect 8092 31668 8148 31678
rect 7756 31666 8148 31668
rect 7756 31614 7758 31666
rect 7810 31614 8094 31666
rect 8146 31614 8148 31666
rect 7756 31612 8148 31614
rect 7756 31602 7812 31612
rect 8092 31602 8148 31612
rect 7196 31556 7252 31566
rect 7532 31556 7588 31566
rect 7196 31554 7588 31556
rect 7196 31502 7198 31554
rect 7250 31502 7534 31554
rect 7586 31502 7588 31554
rect 7196 31500 7588 31502
rect 7196 31490 7252 31500
rect 7532 31444 7588 31500
rect 7532 31378 7588 31388
rect 8540 31332 8596 31726
rect 5964 31220 6020 31230
rect 5964 31126 6020 31164
rect 8428 31108 8484 31118
rect 8428 30994 8484 31052
rect 8428 30942 8430 30994
rect 8482 30942 8484 30994
rect 8428 30930 8484 30942
rect 6412 30884 6468 30894
rect 6412 30790 6468 30828
rect 8204 30882 8260 30894
rect 8204 30830 8206 30882
rect 8258 30830 8260 30882
rect 7980 30436 8036 30446
rect 6076 30210 6132 30222
rect 6076 30158 6078 30210
rect 6130 30158 6132 30210
rect 5964 30100 6020 30110
rect 5964 30006 6020 30044
rect 6076 29650 6132 30158
rect 7980 30210 8036 30380
rect 7980 30158 7982 30210
rect 8034 30158 8036 30210
rect 7980 30146 8036 30158
rect 8204 30212 8260 30830
rect 8540 30212 8596 31276
rect 8652 30212 8708 30222
rect 8540 30210 8708 30212
rect 8540 30158 8654 30210
rect 8706 30158 8708 30210
rect 8540 30156 8708 30158
rect 8204 30146 8260 30156
rect 8652 30100 8708 30156
rect 8652 30034 8708 30044
rect 7980 29988 8036 29998
rect 6076 29598 6078 29650
rect 6130 29598 6132 29650
rect 6076 29586 6132 29598
rect 6972 29652 7028 29662
rect 5964 29538 6020 29550
rect 5964 29486 5966 29538
rect 6018 29486 6020 29538
rect 5964 28980 6020 29486
rect 6972 29426 7028 29596
rect 7980 29650 8036 29932
rect 8316 29988 8372 29998
rect 8316 29986 8484 29988
rect 8316 29934 8318 29986
rect 8370 29934 8484 29986
rect 8316 29932 8484 29934
rect 8316 29922 8372 29932
rect 7980 29598 7982 29650
rect 8034 29598 8036 29650
rect 6972 29374 6974 29426
rect 7026 29374 7028 29426
rect 6188 29316 6244 29326
rect 6524 29316 6580 29326
rect 6188 29314 6580 29316
rect 6188 29262 6190 29314
rect 6242 29262 6526 29314
rect 6578 29262 6580 29314
rect 6188 29260 6580 29262
rect 6188 29250 6244 29260
rect 6524 29250 6580 29260
rect 5964 28924 6132 28980
rect 5964 28754 6020 28766
rect 5964 28702 5966 28754
rect 6018 28702 6020 28754
rect 5964 27972 6020 28702
rect 6076 28532 6132 28924
rect 6300 28644 6356 28654
rect 6636 28644 6692 28654
rect 6300 28642 6692 28644
rect 6300 28590 6302 28642
rect 6354 28590 6638 28642
rect 6690 28590 6692 28642
rect 6300 28588 6692 28590
rect 6300 28578 6356 28588
rect 6636 28578 6692 28588
rect 6972 28644 7028 29374
rect 7420 29428 7476 29438
rect 7756 29428 7812 29438
rect 7420 29426 7812 29428
rect 7420 29374 7422 29426
rect 7474 29374 7758 29426
rect 7810 29374 7812 29426
rect 7420 29372 7812 29374
rect 7420 29362 7476 29372
rect 7756 29362 7812 29372
rect 7868 29428 7924 29438
rect 7532 28756 7588 28766
rect 7756 28756 7812 28766
rect 7532 28754 7756 28756
rect 7532 28702 7534 28754
rect 7586 28702 7756 28754
rect 7532 28700 7756 28702
rect 7532 28690 7588 28700
rect 7756 28690 7812 28700
rect 6972 28578 7028 28588
rect 7308 28642 7364 28654
rect 7308 28590 7310 28642
rect 7362 28590 7364 28642
rect 6076 28530 6244 28532
rect 6076 28478 6078 28530
rect 6130 28478 6244 28530
rect 6076 28476 6244 28478
rect 6076 28466 6132 28476
rect 6188 27972 6244 28476
rect 6188 27916 6580 27972
rect 5964 27906 6020 27916
rect 6412 27186 6468 27198
rect 6412 27134 6414 27186
rect 6466 27134 6468 27186
rect 6188 27076 6244 27086
rect 6412 27076 6468 27134
rect 6244 27020 6468 27076
rect 6188 27010 6244 27020
rect 6524 26962 6580 27916
rect 7308 27748 7364 28590
rect 7420 28644 7476 28654
rect 7420 28420 7476 28588
rect 7420 28364 7700 28420
rect 7644 27858 7700 28364
rect 7644 27806 7646 27858
rect 7698 27806 7700 27858
rect 7644 27794 7700 27806
rect 7420 27748 7476 27758
rect 7308 27746 7476 27748
rect 7308 27694 7422 27746
rect 7474 27694 7476 27746
rect 7308 27692 7476 27694
rect 7420 27636 7476 27692
rect 7420 27570 7476 27580
rect 6524 26910 6526 26962
rect 6578 26910 6580 26962
rect 6524 26908 6580 26910
rect 6748 26962 6804 26974
rect 6748 26910 6750 26962
rect 6802 26910 6804 26962
rect 6748 26908 6804 26910
rect 7868 26962 7924 29372
rect 7980 28642 8036 29598
rect 8428 29652 8484 29932
rect 8540 29652 8596 29662
rect 8428 29596 8540 29652
rect 8540 29586 8596 29596
rect 8652 29652 8708 29662
rect 8764 29652 8820 31836
rect 8876 31826 8932 31836
rect 8988 31668 9044 31678
rect 8988 31106 9044 31612
rect 9100 31444 9156 32398
rect 9100 31378 9156 31388
rect 8988 31054 8990 31106
rect 9042 31054 9044 31106
rect 8988 31042 9044 31054
rect 9100 31108 9156 31118
rect 8876 30436 8932 30446
rect 8876 30342 8932 30380
rect 9100 30434 9156 31052
rect 9100 30382 9102 30434
rect 9154 30382 9156 30434
rect 9100 30370 9156 30382
rect 8652 29650 8820 29652
rect 8652 29598 8654 29650
rect 8706 29598 8820 29650
rect 8652 29596 8820 29598
rect 8876 29652 8932 29662
rect 8652 29586 8708 29596
rect 8876 29558 8932 29596
rect 8092 29428 8148 29438
rect 8092 29334 8148 29372
rect 8988 29428 9044 29438
rect 9044 29372 9156 29428
rect 8988 29334 9044 29372
rect 8092 28756 8148 28794
rect 8092 28690 8148 28700
rect 7980 28590 7982 28642
rect 8034 28590 8036 28642
rect 7980 28308 8036 28590
rect 8204 28644 8260 28654
rect 8204 28550 8260 28588
rect 8652 28642 8708 28654
rect 8652 28590 8654 28642
rect 8706 28590 8708 28642
rect 8652 28420 8708 28590
rect 9100 28530 9156 29372
rect 9100 28478 9102 28530
rect 9154 28478 9156 28530
rect 9100 28466 9156 28478
rect 8652 28354 8708 28364
rect 7980 28252 8484 28308
rect 8428 27970 8484 28252
rect 8428 27918 8430 27970
rect 8482 27918 8484 27970
rect 7980 27636 8036 27646
rect 7980 27542 8036 27580
rect 8428 27074 8484 27918
rect 8876 27860 8932 27870
rect 8428 27022 8430 27074
rect 8482 27022 8484 27074
rect 8428 27010 8484 27022
rect 8540 27636 8596 27646
rect 8652 27636 8708 27646
rect 8596 27634 8708 27636
rect 8596 27582 8654 27634
rect 8706 27582 8708 27634
rect 8596 27580 8708 27582
rect 7868 26910 7870 26962
rect 7922 26910 7924 26962
rect 5852 26852 6356 26908
rect 6524 26852 6692 26908
rect 6748 26852 7812 26908
rect 3500 24946 3612 24948
rect 3500 24894 3502 24946
rect 3554 24894 3612 24946
rect 3500 24892 3612 24894
rect 3500 24882 3556 24892
rect 3612 24854 3668 24892
rect 3948 25282 4004 25294
rect 3948 25230 3950 25282
rect 4002 25230 4004 25282
rect 3948 25172 4004 25230
rect 3836 24610 3892 24622
rect 3836 24558 3838 24610
rect 3890 24558 3892 24610
rect 3836 24498 3892 24558
rect 3836 24446 3838 24498
rect 3890 24446 3892 24498
rect 3836 24434 3892 24446
rect 3948 23940 4004 25116
rect 3836 23884 4004 23940
rect 4060 24498 4116 25340
rect 4172 24948 4228 24958
rect 4396 24948 4452 24958
rect 4228 24946 4452 24948
rect 4228 24894 4398 24946
rect 4450 24894 4452 24946
rect 4228 24892 4452 24894
rect 4172 24882 4228 24892
rect 4396 24882 4452 24892
rect 4620 24612 4676 25676
rect 4844 25284 4900 25294
rect 4956 25284 5012 26236
rect 5068 26066 5124 26078
rect 5068 26014 5070 26066
rect 5122 26014 5124 26066
rect 5068 25844 5124 26014
rect 5180 26068 5236 26078
rect 5292 26068 5348 26852
rect 5404 26180 5460 26190
rect 5404 26086 5460 26124
rect 5180 26066 5348 26068
rect 5180 26014 5182 26066
rect 5234 26014 5348 26066
rect 5180 26012 5348 26014
rect 5180 26002 5236 26012
rect 5516 25844 5572 26852
rect 5964 26404 6020 26414
rect 5964 26290 6020 26348
rect 5964 26238 5966 26290
rect 6018 26238 6020 26290
rect 5964 26226 6020 26238
rect 6188 26178 6244 26190
rect 6188 26126 6190 26178
rect 6242 26126 6244 26178
rect 5068 25788 5572 25844
rect 5628 26066 5684 26078
rect 5628 26014 5630 26066
rect 5682 26014 5684 26066
rect 5628 25620 5684 26014
rect 5740 26068 5796 26078
rect 6188 26068 6244 26126
rect 5740 26066 6132 26068
rect 5740 26014 5742 26066
rect 5794 26014 6132 26066
rect 5740 26012 6132 26014
rect 5740 26002 5796 26012
rect 5852 25732 5908 25742
rect 5628 25564 5796 25620
rect 4900 25228 5012 25284
rect 5628 25394 5684 25406
rect 5628 25342 5630 25394
rect 5682 25342 5684 25394
rect 4844 25190 4900 25228
rect 5516 25172 5572 25182
rect 5516 24946 5572 25116
rect 5516 24894 5518 24946
rect 5570 24894 5572 24946
rect 5516 24882 5572 24894
rect 4732 24836 4788 24846
rect 4788 24780 5012 24836
rect 4732 24742 4788 24780
rect 4620 24556 4900 24612
rect 4060 24446 4062 24498
rect 4114 24446 4116 24498
rect 3724 23828 3780 23838
rect 3724 23378 3780 23772
rect 3724 23326 3726 23378
rect 3778 23326 3780 23378
rect 3724 23314 3780 23326
rect 3612 23154 3668 23166
rect 3612 23102 3614 23154
rect 3666 23102 3668 23154
rect 3612 23044 3668 23102
rect 3612 22978 3668 22988
rect 3836 22036 3892 23884
rect 3948 23716 4004 23726
rect 3948 23154 4004 23660
rect 3948 23102 3950 23154
rect 4002 23102 4004 23154
rect 3948 23090 4004 23102
rect 3388 21758 3390 21810
rect 3442 21758 3444 21810
rect 3388 21746 3444 21758
rect 3612 21980 4004 22036
rect 3276 21298 3332 21308
rect 2380 20962 2436 20972
rect 2268 20916 2324 20926
rect 2268 20822 2324 20860
rect 2716 20802 2772 20814
rect 2716 20750 2718 20802
rect 2770 20750 2772 20802
rect 2492 20580 2548 20590
rect 2492 20130 2548 20524
rect 2716 20356 2772 20750
rect 2940 20804 2996 20814
rect 2940 20690 2996 20748
rect 3612 20802 3668 21980
rect 3836 21812 3892 21822
rect 3836 21718 3892 21756
rect 3948 21810 4004 21980
rect 3948 21758 3950 21810
rect 4002 21758 4004 21810
rect 3948 21746 4004 21758
rect 3724 21586 3780 21598
rect 4060 21588 4116 24446
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4620 24050 4676 24062
rect 4620 23998 4622 24050
rect 4674 23998 4676 24050
rect 3724 21534 3726 21586
rect 3778 21534 3780 21586
rect 3724 21252 3780 21534
rect 3724 21186 3780 21196
rect 3948 21532 4116 21588
rect 4284 23266 4340 23278
rect 4284 23214 4286 23266
rect 4338 23214 4340 23266
rect 3612 20750 3614 20802
rect 3666 20750 3668 20802
rect 3612 20738 3668 20750
rect 2940 20638 2942 20690
rect 2994 20638 2996 20690
rect 2940 20626 2996 20638
rect 2492 20078 2494 20130
rect 2546 20078 2548 20130
rect 2492 20066 2548 20078
rect 2604 20244 2660 20254
rect 1820 19966 1822 20018
rect 1874 19966 1876 20018
rect 1708 19572 1764 19582
rect 1708 19234 1764 19516
rect 1708 19182 1710 19234
rect 1762 19182 1764 19234
rect 1708 19170 1764 19182
rect 1708 18450 1764 18462
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1708 18228 1764 18398
rect 1708 17780 1764 18172
rect 1708 17714 1764 17724
rect 1820 17666 1876 19966
rect 2380 19122 2436 19134
rect 2380 19070 2382 19122
rect 2434 19070 2436 19122
rect 2044 19012 2100 19022
rect 2044 18918 2100 18956
rect 2380 18900 2436 19070
rect 2380 18834 2436 18844
rect 2604 18676 2660 20188
rect 2716 19460 2772 20300
rect 3388 20578 3444 20590
rect 3388 20526 3390 20578
rect 3442 20526 3444 20578
rect 3388 19908 3444 20526
rect 3500 20580 3556 20590
rect 3500 20486 3556 20524
rect 3948 20244 4004 21532
rect 4284 21364 4340 23214
rect 4620 23044 4676 23998
rect 4844 23716 4900 24556
rect 4844 23650 4900 23660
rect 4620 22978 4676 22988
rect 4844 23380 4900 23390
rect 4844 23154 4900 23324
rect 4844 23102 4846 23154
rect 4898 23102 4900 23154
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4844 22596 4900 23102
rect 4620 22540 4900 22596
rect 4620 22482 4676 22540
rect 4620 22430 4622 22482
rect 4674 22430 4676 22482
rect 4620 22418 4676 22430
rect 4732 21810 4788 22540
rect 4732 21758 4734 21810
rect 4786 21758 4788 21810
rect 4732 21746 4788 21758
rect 4508 21698 4564 21710
rect 4508 21646 4510 21698
rect 4562 21646 4564 21698
rect 4396 21588 4452 21598
rect 4508 21588 4564 21646
rect 4844 21700 4900 21710
rect 4956 21700 5012 24780
rect 5292 24722 5348 24734
rect 5292 24670 5294 24722
rect 5346 24670 5348 24722
rect 5068 24052 5124 24062
rect 5068 23958 5124 23996
rect 5292 23828 5348 24670
rect 5404 24612 5460 24622
rect 5404 24518 5460 24556
rect 5628 24276 5684 25342
rect 5740 25172 5796 25564
rect 5852 25506 5908 25676
rect 5852 25454 5854 25506
rect 5906 25454 5908 25506
rect 5852 25442 5908 25454
rect 6076 25506 6132 26012
rect 6188 26002 6244 26012
rect 6188 25732 6244 25742
rect 6188 25638 6244 25676
rect 6076 25454 6078 25506
rect 6130 25454 6132 25506
rect 6076 25442 6132 25454
rect 6300 25506 6356 26852
rect 6636 26628 6692 26852
rect 6636 26572 7140 26628
rect 7084 26514 7140 26572
rect 7084 26462 7086 26514
rect 7138 26462 7140 26514
rect 6300 25454 6302 25506
rect 6354 25454 6356 25506
rect 6300 25442 6356 25454
rect 6412 26290 6468 26302
rect 6412 26238 6414 26290
rect 6466 26238 6468 26290
rect 5964 25284 6020 25294
rect 6020 25228 6132 25284
rect 5964 25218 6020 25228
rect 5852 25172 5908 25182
rect 5740 25116 5852 25172
rect 5852 25106 5908 25116
rect 5740 24834 5796 24846
rect 5740 24782 5742 24834
rect 5794 24782 5796 24834
rect 5740 24500 5796 24782
rect 5740 24434 5796 24444
rect 5292 23762 5348 23772
rect 5516 24220 5684 24276
rect 5516 23380 5572 24220
rect 6076 24052 6132 25228
rect 6412 25172 6468 26238
rect 6636 26290 6692 26302
rect 6636 26238 6638 26290
rect 6690 26238 6692 26290
rect 6636 26180 6692 26238
rect 6972 26180 7028 26190
rect 6636 26178 7028 26180
rect 6636 26126 6974 26178
rect 7026 26126 7028 26178
rect 6636 26124 7028 26126
rect 6972 26114 7028 26124
rect 7084 25956 7140 26462
rect 7756 26516 7812 26852
rect 7868 26740 7924 26910
rect 7980 26964 8036 27002
rect 7980 26898 8036 26908
rect 8540 26962 8596 27580
rect 8652 27570 8708 27580
rect 8540 26910 8542 26962
rect 8594 26910 8596 26962
rect 8540 26898 8596 26910
rect 8876 26908 8932 27804
rect 8204 26850 8260 26862
rect 8204 26798 8206 26850
rect 8258 26798 8260 26850
rect 7868 26684 8148 26740
rect 7756 26460 8036 26516
rect 7980 26402 8036 26460
rect 7980 26350 7982 26402
rect 8034 26350 8036 26402
rect 7980 26338 8036 26350
rect 7308 26180 7364 26190
rect 7308 26086 7364 26124
rect 6748 25900 7140 25956
rect 6748 25394 6804 25900
rect 7980 25620 8036 25630
rect 7980 25526 8036 25564
rect 6972 25508 7028 25518
rect 7644 25508 7700 25518
rect 6748 25342 6750 25394
rect 6802 25342 6804 25394
rect 6748 25330 6804 25342
rect 6860 25506 7700 25508
rect 6860 25454 6974 25506
rect 7026 25454 7646 25506
rect 7698 25454 7700 25506
rect 6860 25452 7700 25454
rect 6412 25060 6468 25116
rect 6412 25004 6692 25060
rect 6188 24836 6244 24846
rect 6188 24742 6244 24780
rect 6300 24836 6356 24846
rect 6300 24834 6468 24836
rect 6300 24782 6302 24834
rect 6354 24782 6468 24834
rect 6300 24780 6468 24782
rect 6300 24770 6356 24780
rect 6300 24500 6356 24510
rect 6300 24406 6356 24444
rect 5852 23996 6356 24052
rect 5740 23938 5796 23950
rect 5740 23886 5742 23938
rect 5794 23886 5796 23938
rect 5740 23828 5796 23886
rect 5740 23762 5796 23772
rect 5740 23604 5796 23614
rect 5628 23380 5684 23390
rect 5516 23378 5684 23380
rect 5516 23326 5630 23378
rect 5682 23326 5684 23378
rect 5516 23324 5684 23326
rect 5628 23314 5684 23324
rect 5740 23266 5796 23548
rect 5740 23214 5742 23266
rect 5794 23214 5796 23266
rect 5740 23202 5796 23214
rect 5292 23154 5348 23166
rect 5292 23102 5294 23154
rect 5346 23102 5348 23154
rect 5292 23044 5348 23102
rect 5292 22978 5348 22988
rect 5068 22484 5124 22494
rect 5740 22484 5796 22494
rect 5852 22484 5908 23996
rect 6300 23938 6356 23996
rect 6300 23886 6302 23938
rect 6354 23886 6356 23938
rect 6300 23874 6356 23886
rect 5964 23716 6020 23726
rect 5964 23622 6020 23660
rect 6300 23604 6356 23614
rect 6412 23604 6468 24780
rect 6636 24052 6692 25004
rect 6636 23986 6692 23996
rect 6356 23548 6468 23604
rect 6636 23828 6692 23838
rect 6300 23538 6356 23548
rect 6636 23268 6692 23772
rect 6524 23212 6692 23268
rect 6300 23156 6356 23166
rect 6300 23062 6356 23100
rect 5068 22482 5908 22484
rect 5068 22430 5070 22482
rect 5122 22430 5742 22482
rect 5794 22430 5908 22482
rect 5068 22428 5908 22430
rect 5068 22418 5124 22428
rect 5740 22418 5796 22428
rect 4844 21698 5012 21700
rect 4844 21646 4846 21698
rect 4898 21646 5012 21698
rect 4844 21644 5012 21646
rect 4844 21634 4900 21644
rect 4396 21586 4564 21588
rect 4396 21534 4398 21586
rect 4450 21534 4564 21586
rect 4396 21532 4564 21534
rect 4396 21522 4452 21532
rect 4284 21308 4900 21364
rect 4172 21252 4228 21262
rect 4228 21196 4340 21252
rect 4172 21186 4228 21196
rect 4284 20916 4340 21196
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4844 21028 4900 21308
rect 4956 21140 5012 21644
rect 5740 21700 5796 21710
rect 5740 21606 5796 21644
rect 5292 21588 5348 21598
rect 5292 21494 5348 21532
rect 4956 21084 5236 21140
rect 4620 20972 5012 21028
rect 4396 20916 4452 20926
rect 4284 20914 4452 20916
rect 4284 20862 4398 20914
rect 4450 20862 4452 20914
rect 4284 20860 4452 20862
rect 4396 20850 4452 20860
rect 4060 20802 4116 20814
rect 4060 20750 4062 20802
rect 4114 20750 4116 20802
rect 4060 20356 4116 20750
rect 4172 20804 4228 20814
rect 4172 20710 4228 20748
rect 4620 20802 4676 20972
rect 4620 20750 4622 20802
rect 4674 20750 4676 20802
rect 4620 20738 4676 20750
rect 4844 20804 4900 20814
rect 4844 20710 4900 20748
rect 4060 20300 4900 20356
rect 3948 20188 4228 20244
rect 3388 19852 4116 19908
rect 3388 19460 3444 19470
rect 2716 19404 2996 19460
rect 2716 19124 2772 19134
rect 2716 19030 2772 19068
rect 2716 18676 2772 18686
rect 2604 18674 2772 18676
rect 2604 18622 2718 18674
rect 2770 18622 2772 18674
rect 2604 18620 2772 18622
rect 2716 18610 2772 18620
rect 2044 18562 2100 18574
rect 2044 18510 2046 18562
rect 2098 18510 2100 18562
rect 2044 17892 2100 18510
rect 2044 17826 2100 17836
rect 1820 17614 1822 17666
rect 1874 17614 1876 17666
rect 1820 17602 1876 17614
rect 2940 17668 2996 19404
rect 3388 19236 3444 19404
rect 4060 19346 4116 19852
rect 4172 19796 4228 20188
rect 4844 20242 4900 20300
rect 4844 20190 4846 20242
rect 4898 20190 4900 20242
rect 4844 20178 4900 20190
rect 4956 20132 5012 20972
rect 5068 20132 5124 20142
rect 4956 20130 5124 20132
rect 4956 20078 5070 20130
rect 5122 20078 5124 20130
rect 4956 20076 5124 20078
rect 4620 19908 4676 19918
rect 4956 19908 5012 20076
rect 5068 20066 5124 20076
rect 5180 20130 5236 21084
rect 5852 20244 5908 22428
rect 6188 22484 6244 22494
rect 6188 22390 6244 22428
rect 6412 21698 6468 21710
rect 6412 21646 6414 21698
rect 6466 21646 6468 21698
rect 6300 21364 6356 21374
rect 6300 21270 6356 21308
rect 5964 20914 6020 20926
rect 5964 20862 5966 20914
rect 6018 20862 6020 20914
rect 5964 20804 6020 20862
rect 5964 20738 6020 20748
rect 6188 20692 6244 20702
rect 6188 20690 6356 20692
rect 6188 20638 6190 20690
rect 6242 20638 6356 20690
rect 6188 20636 6356 20638
rect 6188 20626 6244 20636
rect 5964 20578 6020 20590
rect 5964 20526 5966 20578
rect 6018 20526 6020 20578
rect 5964 20356 6020 20526
rect 6300 20356 6356 20636
rect 5964 20300 6244 20356
rect 5852 20188 6132 20244
rect 5180 20078 5182 20130
rect 5234 20078 5236 20130
rect 4620 19906 5012 19908
rect 4620 19854 4622 19906
rect 4674 19854 5012 19906
rect 4620 19852 5012 19854
rect 4620 19842 4676 19852
rect 4172 19730 4228 19740
rect 4844 19684 4900 19694
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4060 19294 4062 19346
rect 4114 19294 4116 19346
rect 4060 19282 4116 19294
rect 3836 19236 3892 19246
rect 3388 19234 3556 19236
rect 3388 19182 3390 19234
rect 3442 19182 3556 19234
rect 3388 19180 3556 19182
rect 3388 19170 3444 19180
rect 3164 18900 3220 18910
rect 3164 18674 3220 18844
rect 3164 18622 3166 18674
rect 3218 18622 3220 18674
rect 3164 18610 3220 18622
rect 3500 18676 3556 19180
rect 3612 19012 3668 19022
rect 3836 19012 3892 19180
rect 3612 19010 3892 19012
rect 3612 18958 3614 19010
rect 3666 18958 3892 19010
rect 3612 18956 3892 18958
rect 3612 18946 3668 18956
rect 3612 18676 3668 18686
rect 3500 18674 3668 18676
rect 3500 18622 3614 18674
rect 3666 18622 3668 18674
rect 3500 18620 3668 18622
rect 2940 17602 2996 17612
rect 1596 17266 1652 17276
rect 1708 17556 1764 17566
rect 1708 17108 1764 17500
rect 2492 17554 2548 17566
rect 2492 17502 2494 17554
rect 2546 17502 2548 17554
rect 1708 17106 1988 17108
rect 1708 17054 1710 17106
rect 1762 17054 1988 17106
rect 1708 17052 1988 17054
rect 1708 17042 1764 17052
rect 1708 16212 1764 16222
rect 1708 15652 1764 16156
rect 1708 15426 1764 15596
rect 1708 15374 1710 15426
rect 1762 15374 1764 15426
rect 1708 15362 1764 15374
rect 1820 16098 1876 16110
rect 1820 16046 1822 16098
rect 1874 16046 1876 16098
rect 1708 15092 1764 15102
rect 1708 14530 1764 15036
rect 1708 14478 1710 14530
rect 1762 14478 1764 14530
rect 1708 14466 1764 14478
rect 1820 13746 1876 16046
rect 1932 15148 1988 17052
rect 2044 16994 2100 17006
rect 2044 16942 2046 16994
rect 2098 16942 2100 16994
rect 2044 16660 2100 16942
rect 2380 16884 2436 16894
rect 2380 16790 2436 16828
rect 2492 16772 2548 17502
rect 3164 17108 3220 17118
rect 3164 17014 3220 17052
rect 2492 16706 2548 16716
rect 2716 16994 2772 17006
rect 2716 16942 2718 16994
rect 2770 16942 2772 16994
rect 2044 16594 2100 16604
rect 2716 16324 2772 16942
rect 3276 16882 3332 16894
rect 3276 16830 3278 16882
rect 3330 16830 3332 16882
rect 3276 16772 3332 16830
rect 3276 16706 3332 16716
rect 3388 16882 3444 16894
rect 3388 16830 3390 16882
rect 3442 16830 3444 16882
rect 3388 16548 3444 16830
rect 2716 16258 2772 16268
rect 3276 16492 3444 16548
rect 2492 15988 2548 15998
rect 2492 15986 3220 15988
rect 2492 15934 2494 15986
rect 2546 15934 3220 15986
rect 2492 15932 3220 15934
rect 2492 15922 2548 15932
rect 2380 15540 2436 15550
rect 2044 15428 2100 15438
rect 2044 15334 2100 15372
rect 2380 15426 2436 15484
rect 2716 15540 2772 15550
rect 2716 15446 2772 15484
rect 3164 15538 3220 15932
rect 3164 15486 3166 15538
rect 3218 15486 3220 15538
rect 3164 15474 3220 15486
rect 3276 15538 3332 16492
rect 3276 15486 3278 15538
rect 3330 15486 3332 15538
rect 2380 15374 2382 15426
rect 2434 15374 2436 15426
rect 2380 15362 2436 15374
rect 3052 15316 3108 15326
rect 3052 15222 3108 15260
rect 1932 15092 2884 15148
rect 2044 14756 2100 14766
rect 2044 14418 2100 14700
rect 2716 14644 2772 14654
rect 2828 14644 2884 15092
rect 3164 14644 3220 14654
rect 2828 14642 3220 14644
rect 2828 14590 3166 14642
rect 3218 14590 3220 14642
rect 2828 14588 3220 14590
rect 2492 14532 2548 14542
rect 2492 14438 2548 14476
rect 2044 14366 2046 14418
rect 2098 14366 2100 14418
rect 2044 14354 2100 14366
rect 2716 14418 2772 14588
rect 3164 14578 3220 14588
rect 2716 14366 2718 14418
rect 2770 14366 2772 14418
rect 2716 14354 2772 14366
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1708 13412 1764 13422
rect 1708 12962 1764 13356
rect 1708 12910 1710 12962
rect 1762 12910 1764 12962
rect 1708 12628 1764 12910
rect 1708 12562 1764 12572
rect 1708 12180 1764 12190
rect 1708 12086 1764 12124
rect 1708 11508 1764 11518
rect 1708 10724 1764 11452
rect 1708 10630 1764 10668
rect 1820 11394 1876 13694
rect 2716 13748 2772 13758
rect 3276 13748 3332 15486
rect 3276 13692 3444 13748
rect 2492 13634 2548 13646
rect 2492 13582 2494 13634
rect 2546 13582 2548 13634
rect 2492 13076 2548 13582
rect 2492 13010 2548 13020
rect 2380 12964 2436 12974
rect 2380 12870 2436 12908
rect 2716 12850 2772 13692
rect 3276 13524 3332 13534
rect 3276 12962 3332 13468
rect 3388 13300 3444 13692
rect 3500 13412 3556 18620
rect 3612 18610 3668 18620
rect 3612 18452 3668 18462
rect 3612 17106 3668 18396
rect 3612 17054 3614 17106
rect 3666 17054 3668 17106
rect 3612 17042 3668 17054
rect 3836 18450 3892 18956
rect 4172 19234 4228 19246
rect 4172 19182 4174 19234
rect 4226 19182 4228 19234
rect 3836 18398 3838 18450
rect 3890 18398 3892 18450
rect 3724 15764 3780 15774
rect 3612 15428 3668 15438
rect 3612 14642 3668 15372
rect 3724 15314 3780 15708
rect 3724 15262 3726 15314
rect 3778 15262 3780 15314
rect 3724 15250 3780 15262
rect 3836 15314 3892 18398
rect 3948 18452 4004 18462
rect 3948 16884 4004 18396
rect 4060 18338 4116 18350
rect 4060 18286 4062 18338
rect 4114 18286 4116 18338
rect 4060 17108 4116 18286
rect 4060 17042 4116 17052
rect 4172 17668 4228 19182
rect 4508 19122 4564 19134
rect 4508 19070 4510 19122
rect 4562 19070 4564 19122
rect 4284 18452 4340 18462
rect 4284 18358 4340 18396
rect 4396 18450 4452 18462
rect 4396 18398 4398 18450
rect 4450 18398 4452 18450
rect 4396 18340 4452 18398
rect 4508 18452 4564 19070
rect 4732 19012 4788 19022
rect 4620 19010 4788 19012
rect 4620 18958 4734 19010
rect 4786 18958 4788 19010
rect 4620 18956 4788 18958
rect 4620 18564 4676 18956
rect 4732 18946 4788 18956
rect 4620 18498 4676 18508
rect 4844 18564 4900 19628
rect 5068 19236 5124 19246
rect 5180 19236 5236 20078
rect 6076 20130 6132 20188
rect 6076 20078 6078 20130
rect 6130 20078 6132 20130
rect 5628 19908 5684 19918
rect 5628 19814 5684 19852
rect 5068 19234 5236 19236
rect 5068 19182 5070 19234
rect 5122 19182 5236 19234
rect 5068 19180 5236 19182
rect 5516 19794 5572 19806
rect 5516 19742 5518 19794
rect 5570 19742 5572 19794
rect 5068 19170 5124 19180
rect 4844 18498 4900 18508
rect 4956 19010 5012 19022
rect 4956 18958 4958 19010
rect 5010 18958 5012 19010
rect 4508 18386 4564 18396
rect 4396 18274 4452 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4620 17780 4676 17790
rect 4956 17780 5012 18958
rect 5180 18676 5236 18686
rect 5516 18676 5572 19742
rect 6076 19460 6132 20078
rect 6188 20132 6244 20300
rect 6300 20290 6356 20300
rect 6412 20132 6468 21646
rect 6188 20130 6468 20132
rect 6188 20078 6414 20130
rect 6466 20078 6468 20130
rect 6188 20076 6468 20078
rect 6188 19794 6244 20076
rect 6412 20066 6468 20076
rect 6188 19742 6190 19794
rect 6242 19742 6244 19794
rect 6188 19730 6244 19742
rect 6524 19572 6580 23212
rect 6636 23044 6692 23054
rect 6636 22950 6692 22988
rect 6636 22260 6692 22270
rect 6636 21698 6692 22204
rect 6636 21646 6638 21698
rect 6690 21646 6692 21698
rect 6636 21634 6692 21646
rect 6748 20244 6804 20254
rect 6860 20244 6916 25452
rect 6972 25442 7028 25452
rect 7644 25442 7700 25452
rect 7756 25508 7812 25518
rect 7756 24946 7812 25452
rect 7756 24894 7758 24946
rect 7810 24894 7812 24946
rect 7756 24882 7812 24894
rect 7308 24724 7364 24734
rect 7308 24630 7364 24668
rect 6972 24610 7028 24622
rect 6972 24558 6974 24610
rect 7026 24558 7028 24610
rect 6972 23716 7028 24558
rect 7084 24612 7140 24622
rect 7084 24050 7140 24556
rect 7084 23998 7086 24050
rect 7138 23998 7140 24050
rect 7084 23986 7140 23998
rect 6972 23650 7028 23660
rect 7420 23268 7476 23278
rect 8092 23268 8148 26684
rect 8204 26290 8260 26798
rect 8652 26852 8932 26908
rect 8988 27636 9044 27646
rect 8988 26964 9044 27580
rect 8988 26898 9044 26908
rect 8204 26238 8206 26290
rect 8258 26238 8260 26290
rect 8204 26226 8260 26238
rect 8428 26292 8484 26302
rect 8652 26292 8708 26852
rect 8484 26236 8708 26292
rect 8428 26198 8484 26236
rect 9212 25508 9268 38612
rect 9548 35698 9604 35710
rect 9548 35646 9550 35698
rect 9602 35646 9604 35698
rect 9548 35588 9604 35646
rect 9548 35522 9604 35532
rect 9548 32562 9604 32574
rect 9548 32510 9550 32562
rect 9602 32510 9604 32562
rect 9548 32004 9604 32510
rect 9548 31938 9604 31948
rect 9436 31890 9492 31902
rect 9436 31838 9438 31890
rect 9490 31838 9492 31890
rect 9436 31780 9492 31838
rect 9436 31714 9492 31724
rect 9660 31780 9716 43652
rect 9996 43538 10052 43550
rect 9996 43486 9998 43538
rect 10050 43486 10052 43538
rect 9996 42868 10052 43486
rect 9996 42802 10052 42812
rect 9996 39620 10052 39630
rect 9996 39060 10052 39564
rect 9996 38994 10052 39004
rect 10108 32788 10164 44604
rect 10220 43762 10276 45276
rect 10668 45266 10724 45276
rect 10780 45556 10836 45566
rect 10780 45106 10836 45500
rect 11676 45556 11732 46620
rect 12012 46674 12068 46686
rect 12012 46622 12014 46674
rect 12066 46622 12068 46674
rect 11788 46564 11844 46574
rect 11788 46002 11844 46508
rect 11788 45950 11790 46002
rect 11842 45950 11844 46002
rect 11788 45938 11844 45950
rect 12012 45892 12068 46622
rect 12460 46676 12516 47518
rect 12908 47572 12964 47582
rect 13020 47572 13076 48412
rect 13356 48402 13412 48412
rect 13468 48804 13524 48814
rect 13916 48804 13972 48814
rect 12908 47570 13076 47572
rect 12908 47518 12910 47570
rect 12962 47518 13076 47570
rect 12908 47516 13076 47518
rect 13132 47796 13188 47806
rect 12908 47506 12964 47516
rect 12460 46610 12516 46620
rect 12684 46562 12740 46574
rect 12684 46510 12686 46562
rect 12738 46510 12740 46562
rect 12684 46004 12740 46510
rect 13132 46116 13188 47740
rect 11900 45836 12068 45892
rect 12124 45948 12740 46004
rect 13020 46004 13076 46014
rect 13132 46004 13188 46060
rect 13020 46002 13188 46004
rect 13020 45950 13022 46002
rect 13074 45950 13188 46002
rect 13020 45948 13188 45950
rect 13244 47012 13300 47022
rect 13244 46674 13300 46956
rect 13244 46622 13246 46674
rect 13298 46622 13300 46674
rect 11788 45780 11844 45790
rect 11900 45780 11956 45836
rect 11844 45724 11956 45780
rect 11788 45686 11844 45724
rect 11676 45490 11732 45500
rect 12012 45668 12068 45678
rect 12124 45668 12180 45948
rect 13020 45938 13076 45948
rect 12012 45666 12180 45668
rect 12012 45614 12014 45666
rect 12066 45614 12180 45666
rect 12012 45612 12180 45614
rect 12236 45778 12292 45790
rect 12236 45726 12238 45778
rect 12290 45726 12292 45778
rect 12236 45668 12292 45726
rect 11228 45220 11284 45230
rect 11228 45126 11284 45164
rect 10780 45054 10782 45106
rect 10834 45054 10836 45106
rect 10780 44436 10836 45054
rect 11004 45108 11060 45118
rect 11004 45106 11172 45108
rect 11004 45054 11006 45106
rect 11058 45054 11172 45106
rect 11004 45052 11172 45054
rect 11004 45042 11060 45052
rect 10892 44996 10948 45006
rect 10892 44902 10948 44940
rect 11004 44436 11060 44446
rect 10780 44434 11060 44436
rect 10780 44382 11006 44434
rect 11058 44382 11060 44434
rect 10780 44380 11060 44382
rect 11004 44370 11060 44380
rect 11116 44100 11172 45052
rect 11452 44100 11508 44110
rect 11116 44044 11452 44100
rect 11452 44006 11508 44044
rect 12012 44100 12068 45612
rect 12236 45602 12292 45612
rect 12572 45780 12628 45790
rect 12236 45444 12292 45454
rect 12124 45332 12180 45342
rect 12124 45106 12180 45276
rect 12124 45054 12126 45106
rect 12178 45054 12180 45106
rect 12124 45042 12180 45054
rect 12012 44034 12068 44044
rect 10220 43710 10222 43762
rect 10274 43710 10276 43762
rect 10220 43698 10276 43710
rect 12012 43652 12068 43662
rect 10556 43540 10612 43550
rect 10556 43446 10612 43484
rect 11340 43428 11396 43438
rect 11340 43334 11396 43372
rect 11228 42980 11284 42990
rect 11228 42886 11284 42924
rect 12012 42978 12068 43596
rect 12236 43540 12292 45388
rect 12236 43474 12292 43484
rect 12460 44322 12516 44334
rect 12460 44270 12462 44322
rect 12514 44270 12516 44322
rect 12460 43204 12516 44270
rect 12572 44322 12628 45724
rect 13244 45444 13300 46622
rect 13244 44994 13300 45388
rect 13244 44942 13246 44994
rect 13298 44942 13300 44994
rect 13244 44930 13300 44942
rect 12572 44270 12574 44322
rect 12626 44270 12628 44322
rect 12572 44258 12628 44270
rect 13020 44324 13076 44334
rect 13020 44230 13076 44268
rect 12460 43138 12516 43148
rect 12796 44098 12852 44110
rect 12796 44046 12798 44098
rect 12850 44046 12852 44098
rect 12012 42926 12014 42978
rect 12066 42926 12068 42978
rect 10444 42868 10500 42878
rect 10444 42774 10500 42812
rect 11004 42868 11060 42878
rect 10332 42082 10388 42094
rect 10332 42030 10334 42082
rect 10386 42030 10388 42082
rect 10332 40514 10388 42030
rect 10556 41972 10612 41982
rect 10332 40462 10334 40514
rect 10386 40462 10388 40514
rect 10332 40450 10388 40462
rect 10444 41970 10612 41972
rect 10444 41918 10558 41970
rect 10610 41918 10612 41970
rect 10444 41916 10612 41918
rect 10332 39844 10388 39854
rect 10444 39844 10500 41916
rect 10556 41906 10612 41916
rect 10892 41188 10948 41198
rect 10892 41094 10948 41132
rect 10332 39842 10500 39844
rect 10332 39790 10334 39842
rect 10386 39790 10500 39842
rect 10332 39788 10500 39790
rect 10668 40516 10724 40526
rect 10668 39842 10724 40460
rect 10668 39790 10670 39842
rect 10722 39790 10724 39842
rect 10332 39778 10388 39788
rect 10668 39778 10724 39790
rect 10892 39732 10948 39742
rect 10892 39638 10948 39676
rect 10220 39060 10276 39070
rect 10220 38966 10276 39004
rect 10892 38162 10948 38174
rect 10892 38110 10894 38162
rect 10946 38110 10948 38162
rect 10892 38052 10948 38110
rect 10892 37986 10948 37996
rect 11004 36820 11060 42812
rect 11340 42756 11396 42766
rect 11340 42642 11396 42700
rect 12012 42756 12068 42926
rect 12796 42980 12852 44046
rect 12796 42914 12852 42924
rect 13132 44100 13188 44110
rect 12012 42690 12068 42700
rect 11340 42590 11342 42642
rect 11394 42590 11396 42642
rect 11340 42578 11396 42590
rect 11564 42644 11620 42654
rect 11900 42644 11956 42654
rect 11564 42550 11620 42588
rect 11788 42642 11956 42644
rect 11788 42590 11902 42642
rect 11954 42590 11956 42642
rect 11788 42588 11956 42590
rect 11452 42082 11508 42094
rect 11452 42030 11454 42082
rect 11506 42030 11508 42082
rect 11116 41970 11172 41982
rect 11116 41918 11118 41970
rect 11170 41918 11172 41970
rect 11116 41860 11172 41918
rect 11116 41794 11172 41804
rect 11452 41972 11508 42030
rect 11788 41972 11844 42588
rect 11900 42578 11956 42588
rect 12572 42644 12628 42654
rect 12124 42196 12180 42206
rect 11452 41916 11844 41972
rect 11900 42194 12180 42196
rect 11900 42142 12126 42194
rect 12178 42142 12180 42194
rect 11900 42140 12180 42142
rect 11452 40516 11508 41916
rect 11452 40450 11508 40460
rect 11116 39732 11172 39742
rect 11116 39060 11172 39676
rect 11564 39732 11620 39742
rect 11564 39638 11620 39676
rect 11900 39620 11956 42140
rect 12124 42130 12180 42140
rect 12572 42084 12628 42588
rect 12572 41990 12628 42028
rect 12684 42084 12740 42094
rect 12684 42082 12852 42084
rect 12684 42030 12686 42082
rect 12738 42030 12852 42082
rect 12684 42028 12852 42030
rect 12684 42018 12740 42028
rect 12012 41970 12068 41982
rect 12012 41918 12014 41970
rect 12066 41918 12068 41970
rect 12012 40516 12068 41918
rect 12348 41972 12404 41982
rect 12348 41878 12404 41916
rect 12796 41860 12852 42028
rect 12908 41972 12964 41982
rect 12908 41970 13076 41972
rect 12908 41918 12910 41970
rect 12962 41918 13076 41970
rect 12908 41916 13076 41918
rect 12908 41906 12964 41916
rect 12796 41794 12852 41804
rect 12684 41300 12740 41310
rect 12684 41298 12964 41300
rect 12684 41246 12686 41298
rect 12738 41246 12964 41298
rect 12684 41244 12964 41246
rect 12684 41234 12740 41244
rect 12908 40628 12964 41244
rect 12908 40562 12964 40572
rect 12796 40516 12852 40526
rect 12012 40514 12852 40516
rect 12012 40462 12798 40514
rect 12850 40462 12852 40514
rect 12012 40460 12852 40462
rect 12012 39844 12068 40460
rect 12796 40450 12852 40460
rect 12460 40292 12516 40302
rect 12908 40292 12964 40302
rect 12460 40290 12964 40292
rect 12460 40238 12462 40290
rect 12514 40238 12910 40290
rect 12962 40238 12964 40290
rect 12460 40236 12964 40238
rect 12460 40226 12516 40236
rect 12908 40226 12964 40236
rect 12124 39844 12180 39854
rect 12012 39842 12180 39844
rect 12012 39790 12126 39842
rect 12178 39790 12180 39842
rect 12012 39788 12180 39790
rect 12124 39778 12180 39788
rect 11900 39526 11956 39564
rect 12908 39620 12964 39630
rect 12908 39526 12964 39564
rect 11116 38966 11172 39004
rect 12460 39394 12516 39406
rect 12460 39342 12462 39394
rect 12514 39342 12516 39394
rect 12460 39060 12516 39342
rect 11564 38052 11620 38062
rect 11340 37940 11396 37950
rect 11228 37378 11284 37390
rect 11228 37326 11230 37378
rect 11282 37326 11284 37378
rect 11228 36820 11284 37326
rect 10220 36764 11284 36820
rect 10220 34130 10276 36764
rect 11340 36708 11396 37884
rect 11564 37938 11620 37996
rect 12012 38052 12068 38062
rect 12012 37958 12068 37996
rect 12236 38050 12292 38062
rect 12236 37998 12238 38050
rect 12290 37998 12292 38050
rect 11564 37886 11566 37938
rect 11618 37886 11620 37938
rect 11564 37874 11620 37886
rect 12236 37940 12292 37998
rect 12236 37874 12292 37884
rect 11452 37826 11508 37838
rect 11452 37774 11454 37826
rect 11506 37774 11508 37826
rect 11452 37492 11508 37774
rect 11452 37426 11508 37436
rect 12460 37378 12516 39004
rect 13020 39058 13076 41916
rect 13020 39006 13022 39058
rect 13074 39006 13076 39058
rect 12684 38946 12740 38958
rect 12684 38894 12686 38946
rect 12738 38894 12740 38946
rect 12572 38388 12628 38398
rect 12572 38274 12628 38332
rect 12572 38222 12574 38274
rect 12626 38222 12628 38274
rect 12572 38210 12628 38222
rect 12460 37326 12462 37378
rect 12514 37326 12516 37378
rect 11116 36652 11396 36708
rect 11564 37266 11620 37278
rect 11564 37214 11566 37266
rect 11618 37214 11620 37266
rect 10556 36594 10612 36606
rect 10556 36542 10558 36594
rect 10610 36542 10612 36594
rect 10556 36484 10612 36542
rect 11116 36484 11172 36652
rect 10556 36428 11172 36484
rect 11564 36484 11620 37214
rect 12236 37042 12292 37054
rect 12236 36990 12238 37042
rect 12290 36990 12292 37042
rect 11788 36484 11844 36494
rect 11564 36428 11788 36484
rect 11004 36258 11060 36270
rect 11004 36206 11006 36258
rect 11058 36206 11060 36258
rect 10332 35588 10388 35598
rect 11004 35588 11060 36206
rect 10332 35586 10724 35588
rect 10332 35534 10334 35586
rect 10386 35534 10724 35586
rect 10332 35532 10724 35534
rect 10332 35522 10388 35532
rect 10668 35140 10724 35532
rect 11004 35522 11060 35532
rect 11004 35364 11060 35374
rect 10892 35140 10948 35150
rect 10668 35138 10948 35140
rect 10668 35086 10894 35138
rect 10946 35086 10948 35138
rect 10668 35084 10948 35086
rect 10892 35074 10948 35084
rect 11004 35026 11060 35308
rect 11004 34974 11006 35026
rect 11058 34974 11060 35026
rect 11004 34962 11060 34974
rect 11004 34356 11060 34366
rect 10892 34300 11004 34356
rect 10220 34078 10222 34130
rect 10274 34078 10276 34130
rect 10220 34020 10276 34078
rect 10220 33954 10276 33964
rect 10556 34242 10612 34254
rect 10556 34190 10558 34242
rect 10610 34190 10612 34242
rect 10556 33908 10612 34190
rect 10556 33842 10612 33852
rect 10444 33460 10500 33470
rect 10892 33460 10948 34300
rect 11004 34290 11060 34300
rect 11004 34020 11060 34030
rect 11004 33926 11060 33964
rect 10444 33366 10500 33404
rect 10556 33458 10948 33460
rect 10556 33406 10894 33458
rect 10946 33406 10948 33458
rect 10556 33404 10948 33406
rect 10108 32732 10500 32788
rect 9772 32676 9828 32686
rect 9772 32582 9828 32620
rect 9996 32564 10052 32574
rect 9996 32470 10052 32508
rect 10220 32562 10276 32574
rect 10220 32510 10222 32562
rect 10274 32510 10276 32562
rect 10220 31892 10276 32510
rect 10220 31826 10276 31836
rect 9660 31714 9716 31724
rect 9772 31666 9828 31678
rect 9772 31614 9774 31666
rect 9826 31614 9828 31666
rect 9548 31554 9604 31566
rect 9548 31502 9550 31554
rect 9602 31502 9604 31554
rect 9548 31444 9604 31502
rect 9548 31378 9604 31388
rect 9548 31108 9604 31118
rect 9772 31108 9828 31614
rect 10108 31668 10164 31678
rect 10108 31574 10164 31612
rect 10332 31668 10388 31678
rect 10332 31574 10388 31612
rect 10220 31556 10276 31566
rect 10220 31462 10276 31500
rect 10444 31332 10500 32732
rect 10556 32562 10612 33404
rect 10892 33394 10948 33404
rect 11116 33236 11172 36428
rect 11788 36390 11844 36428
rect 12236 36258 12292 36990
rect 12236 36206 12238 36258
rect 12290 36206 12292 36258
rect 12012 35812 12068 35822
rect 11564 33908 11620 33918
rect 10556 32510 10558 32562
rect 10610 32510 10612 32562
rect 10556 32498 10612 32510
rect 10892 33180 11172 33236
rect 11452 33460 11508 33470
rect 9548 31106 9828 31108
rect 9548 31054 9550 31106
rect 9602 31054 9828 31106
rect 9548 31052 9828 31054
rect 10332 31276 10500 31332
rect 10668 31668 10724 31678
rect 9548 31042 9604 31052
rect 9996 30994 10052 31006
rect 9996 30942 9998 30994
rect 10050 30942 10052 30994
rect 9884 30882 9940 30894
rect 9884 30830 9886 30882
rect 9938 30830 9940 30882
rect 9324 30772 9380 30782
rect 9324 30434 9380 30716
rect 9324 30382 9326 30434
rect 9378 30382 9380 30434
rect 9324 30370 9380 30382
rect 9548 30324 9604 30334
rect 9436 28644 9492 28654
rect 9548 28644 9604 30268
rect 9660 30100 9716 30110
rect 9660 29764 9716 30044
rect 9772 29988 9828 29998
rect 9772 29894 9828 29932
rect 9660 29708 9828 29764
rect 9660 29538 9716 29550
rect 9660 29486 9662 29538
rect 9714 29486 9716 29538
rect 9660 28756 9716 29486
rect 9772 29428 9828 29708
rect 9884 29652 9940 30830
rect 9996 30772 10052 30942
rect 9996 30706 10052 30716
rect 10220 30324 10276 30334
rect 10220 30230 10276 30268
rect 9996 29652 10052 29662
rect 9884 29650 10052 29652
rect 9884 29598 9998 29650
rect 10050 29598 10052 29650
rect 9884 29596 10052 29598
rect 9996 29586 10052 29596
rect 10108 29652 10164 29662
rect 10108 29558 10164 29596
rect 9884 29428 9940 29438
rect 9772 29426 9940 29428
rect 9772 29374 9886 29426
rect 9938 29374 9940 29426
rect 9772 29372 9940 29374
rect 9884 29362 9940 29372
rect 9660 28700 10052 28756
rect 9436 28642 9940 28644
rect 9436 28590 9438 28642
rect 9490 28590 9940 28642
rect 9436 28588 9940 28590
rect 9436 28578 9492 28588
rect 9548 27858 9604 27870
rect 9548 27806 9550 27858
rect 9602 27806 9604 27858
rect 9548 27636 9604 27806
rect 9772 27860 9828 27870
rect 9772 27766 9828 27804
rect 9548 27570 9604 27580
rect 9660 27746 9716 27758
rect 9660 27694 9662 27746
rect 9714 27694 9716 27746
rect 9212 25442 9268 25452
rect 9436 26850 9492 26862
rect 9436 26798 9438 26850
rect 9490 26798 9492 26850
rect 9212 24050 9268 24062
rect 9212 23998 9214 24050
rect 9266 23998 9268 24050
rect 9212 23604 9268 23998
rect 9212 23538 9268 23548
rect 9436 23492 9492 26798
rect 9660 26290 9716 27694
rect 9660 26238 9662 26290
rect 9714 26238 9716 26290
rect 9660 26226 9716 26238
rect 9548 26180 9604 26190
rect 9548 26086 9604 26124
rect 9884 25396 9940 28588
rect 9996 28420 10052 28700
rect 9996 27860 10052 28364
rect 10220 27860 10276 27870
rect 9996 27858 10276 27860
rect 9996 27806 10222 27858
rect 10274 27806 10276 27858
rect 9996 27804 10276 27806
rect 10220 27412 10276 27804
rect 10220 27346 10276 27356
rect 10332 26908 10388 31276
rect 10556 30212 10612 30222
rect 10556 30118 10612 30156
rect 10444 30100 10500 30110
rect 10444 30006 10500 30044
rect 10668 29314 10724 31612
rect 10780 30996 10836 31006
rect 10780 30434 10836 30940
rect 10780 30382 10782 30434
rect 10834 30382 10836 30434
rect 10780 29652 10836 30382
rect 10780 29586 10836 29596
rect 10668 29262 10670 29314
rect 10722 29262 10724 29314
rect 10444 27860 10500 27870
rect 10444 27074 10500 27804
rect 10444 27022 10446 27074
rect 10498 27022 10500 27074
rect 10444 27010 10500 27022
rect 10668 26908 10724 29262
rect 10892 28308 10948 33180
rect 11228 32450 11284 32462
rect 11228 32398 11230 32450
rect 11282 32398 11284 32450
rect 11228 31890 11284 32398
rect 11228 31838 11230 31890
rect 11282 31838 11284 31890
rect 11228 31826 11284 31838
rect 11340 31668 11396 31678
rect 11340 31574 11396 31612
rect 11116 31556 11172 31566
rect 11116 31462 11172 31500
rect 11340 30996 11396 31006
rect 11452 30996 11508 33404
rect 11564 33346 11620 33852
rect 11564 33294 11566 33346
rect 11618 33294 11620 33346
rect 11564 33282 11620 33294
rect 11676 33124 11732 33134
rect 11900 33124 11956 33134
rect 11676 33030 11732 33068
rect 11788 33122 11956 33124
rect 11788 33070 11902 33122
rect 11954 33070 11956 33122
rect 11788 33068 11956 33070
rect 11788 32340 11844 33068
rect 11900 33058 11956 33068
rect 11676 32284 11844 32340
rect 11564 31892 11620 31902
rect 11564 31556 11620 31836
rect 11676 31778 11732 32284
rect 12012 32228 12068 35756
rect 12236 35252 12292 36206
rect 12460 36036 12516 37326
rect 12684 37380 12740 38894
rect 13020 38052 13076 39006
rect 13020 37986 13076 37996
rect 12572 37156 12628 37166
rect 12572 37062 12628 37100
rect 12684 36482 12740 37324
rect 12908 37156 12964 37166
rect 13132 37156 13188 44044
rect 13468 43708 13524 48748
rect 13804 48802 13972 48804
rect 13804 48750 13918 48802
rect 13970 48750 13972 48802
rect 13804 48748 13972 48750
rect 13580 46116 13636 46126
rect 13580 46022 13636 46060
rect 13692 45890 13748 45902
rect 13692 45838 13694 45890
rect 13746 45838 13748 45890
rect 13692 45556 13748 45838
rect 13692 45490 13748 45500
rect 13580 44212 13636 44222
rect 13580 44118 13636 44156
rect 13468 43652 13748 43708
rect 13468 43426 13524 43438
rect 13468 43374 13470 43426
rect 13522 43374 13524 43426
rect 13468 43204 13524 43374
rect 13468 43138 13524 43148
rect 13580 43428 13636 43438
rect 13468 42980 13524 42990
rect 13468 42886 13524 42924
rect 13580 42866 13636 43372
rect 13580 42814 13582 42866
rect 13634 42814 13636 42866
rect 13580 42802 13636 42814
rect 13692 42756 13748 43652
rect 13692 42690 13748 42700
rect 13692 42532 13748 42542
rect 13356 42476 13692 42532
rect 13244 41076 13300 41086
rect 13244 38948 13300 41020
rect 13356 40626 13412 42476
rect 13692 42438 13748 42476
rect 13804 42308 13860 48748
rect 13916 48738 13972 48748
rect 14028 48242 14084 49868
rect 14700 49026 14756 50764
rect 15372 50596 15428 50606
rect 15708 50596 15764 51324
rect 15820 51314 15876 51324
rect 15820 50708 15876 50718
rect 15820 50614 15876 50652
rect 16044 50596 16100 51550
rect 16268 52052 16324 52062
rect 16268 51378 16324 51996
rect 16492 52052 16548 52062
rect 16492 51490 16548 51996
rect 16492 51438 16494 51490
rect 16546 51438 16548 51490
rect 16492 51426 16548 51438
rect 16268 51326 16270 51378
rect 16322 51326 16324 51378
rect 16156 51268 16212 51278
rect 16156 51174 16212 51212
rect 16156 50596 16212 50606
rect 15372 50594 15708 50596
rect 15372 50542 15374 50594
rect 15426 50542 15708 50594
rect 15372 50540 15708 50542
rect 15372 50530 15428 50540
rect 15708 50502 15764 50540
rect 15932 50594 16212 50596
rect 15932 50542 16158 50594
rect 16210 50542 16212 50594
rect 15932 50540 16212 50542
rect 14924 50482 14980 50494
rect 14924 50430 14926 50482
rect 14978 50430 14980 50482
rect 14924 49924 14980 50430
rect 15820 50482 15876 50494
rect 15820 50430 15822 50482
rect 15874 50430 15876 50482
rect 14924 49868 15316 49924
rect 15260 49812 15316 49868
rect 15708 49922 15764 49934
rect 15708 49870 15710 49922
rect 15762 49870 15764 49922
rect 15372 49812 15428 49822
rect 15260 49810 15428 49812
rect 15260 49758 15374 49810
rect 15426 49758 15428 49810
rect 15260 49756 15428 49758
rect 15036 49698 15092 49710
rect 15036 49646 15038 49698
rect 15090 49646 15092 49698
rect 15036 49588 15092 49646
rect 15036 49522 15092 49532
rect 14700 48974 14702 49026
rect 14754 48974 14756 49026
rect 14700 48962 14756 48974
rect 14812 49026 14868 49038
rect 14812 48974 14814 49026
rect 14866 48974 14868 49026
rect 14028 48190 14030 48242
rect 14082 48190 14084 48242
rect 14028 47012 14084 48190
rect 14700 48132 14756 48142
rect 14700 48038 14756 48076
rect 14028 46946 14084 46956
rect 13916 46564 13972 46574
rect 13916 46562 14644 46564
rect 13916 46510 13918 46562
rect 13970 46510 14644 46562
rect 13916 46508 14644 46510
rect 13916 46498 13972 46508
rect 14588 46114 14644 46508
rect 14588 46062 14590 46114
rect 14642 46062 14644 46114
rect 14588 46050 14644 46062
rect 14140 46004 14196 46014
rect 14700 46004 14756 46014
rect 14140 46002 14532 46004
rect 14140 45950 14142 46002
rect 14194 45950 14532 46002
rect 14140 45948 14532 45950
rect 14140 45938 14196 45948
rect 13916 45890 13972 45902
rect 13916 45838 13918 45890
rect 13970 45838 13972 45890
rect 13916 45780 13972 45838
rect 13916 45714 13972 45724
rect 14252 45780 14308 45790
rect 14252 45778 14420 45780
rect 14252 45726 14254 45778
rect 14306 45726 14420 45778
rect 14252 45724 14420 45726
rect 14252 45714 14308 45724
rect 14252 45556 14308 45566
rect 14140 45332 14196 45342
rect 13916 44772 13972 44782
rect 13916 44324 13972 44716
rect 13916 44230 13972 44268
rect 14140 44212 14196 45276
rect 14252 44322 14308 45500
rect 14364 45106 14420 45724
rect 14364 45054 14366 45106
rect 14418 45054 14420 45106
rect 14364 45042 14420 45054
rect 14476 45668 14532 45948
rect 14700 45910 14756 45948
rect 14476 44884 14532 45612
rect 14700 45108 14756 45118
rect 14700 45014 14756 45052
rect 14812 44994 14868 48974
rect 15148 49028 15204 49066
rect 15148 48962 15204 48972
rect 15036 48916 15092 48926
rect 14812 44942 14814 44994
rect 14866 44942 14868 44994
rect 14812 44930 14868 44942
rect 14924 45218 14980 45230
rect 14924 45166 14926 45218
rect 14978 45166 14980 45218
rect 14252 44270 14254 44322
rect 14306 44270 14308 44322
rect 14252 44258 14308 44270
rect 14364 44828 14532 44884
rect 14028 44098 14084 44110
rect 14028 44046 14030 44098
rect 14082 44046 14084 44098
rect 13916 43540 13972 43550
rect 13916 43446 13972 43484
rect 14028 42980 14084 44046
rect 14028 42914 14084 42924
rect 13692 42252 13860 42308
rect 13580 42084 13636 42094
rect 13468 41972 13524 41982
rect 13468 41076 13524 41916
rect 13580 41410 13636 42028
rect 13580 41358 13582 41410
rect 13634 41358 13636 41410
rect 13580 41346 13636 41358
rect 13692 41186 13748 42252
rect 13692 41134 13694 41186
rect 13746 41134 13748 41186
rect 13580 41076 13636 41086
rect 13468 41074 13636 41076
rect 13468 41022 13582 41074
rect 13634 41022 13636 41074
rect 13468 41020 13636 41022
rect 13580 41010 13636 41020
rect 13692 41076 13748 41134
rect 13692 41010 13748 41020
rect 13804 42082 13860 42094
rect 13804 42030 13806 42082
rect 13858 42030 13860 42082
rect 13804 41972 13860 42030
rect 13804 40964 13860 41916
rect 14140 41860 14196 44156
rect 14364 43204 14420 44828
rect 14924 44660 14980 45166
rect 14924 44594 14980 44604
rect 15036 44436 15092 48860
rect 15148 48804 15204 48814
rect 15260 48804 15316 49756
rect 15372 49746 15428 49756
rect 15708 49812 15764 49870
rect 15708 49746 15764 49756
rect 15820 49588 15876 50430
rect 15932 49812 15988 50540
rect 16156 50530 16212 50540
rect 16268 50428 16324 51326
rect 16828 50708 16884 52110
rect 16716 50652 16884 50708
rect 16044 50372 16324 50428
rect 16380 50596 16436 50606
rect 16716 50596 16772 50652
rect 16940 50596 16996 52780
rect 17052 51716 17108 53566
rect 17388 53620 17444 53630
rect 17276 53508 17332 53518
rect 17388 53508 17444 53564
rect 17836 53620 17892 54462
rect 17948 54516 18004 55244
rect 18620 55188 18676 55198
rect 18508 55186 18676 55188
rect 18508 55134 18622 55186
rect 18674 55134 18676 55186
rect 18508 55132 18676 55134
rect 18508 54738 18564 55132
rect 18620 55122 18676 55132
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 18508 54686 18510 54738
rect 18562 54686 18564 54738
rect 18508 54674 18564 54686
rect 17948 54450 18004 54460
rect 18060 54516 18116 54526
rect 18956 54516 19012 54526
rect 18060 54514 18228 54516
rect 18060 54462 18062 54514
rect 18114 54462 18228 54514
rect 18060 54460 18228 54462
rect 18060 54450 18116 54460
rect 17836 53554 17892 53564
rect 18172 53620 18228 54460
rect 18396 54404 18452 54414
rect 18396 54310 18452 54348
rect 18956 53844 19012 54460
rect 18956 53778 19012 53788
rect 19628 54402 19684 54414
rect 19628 54350 19630 54402
rect 19682 54350 19684 54402
rect 18396 53732 18452 53742
rect 18228 53564 18340 53620
rect 18172 53554 18228 53564
rect 17276 53506 17444 53508
rect 17276 53454 17278 53506
rect 17330 53454 17444 53506
rect 17276 53452 17444 53454
rect 17276 53442 17332 53452
rect 17388 53058 17444 53452
rect 17388 53006 17390 53058
rect 17442 53006 17444 53058
rect 17388 52164 17444 53006
rect 17500 53508 17556 53518
rect 17500 52164 17556 53452
rect 18060 53506 18116 53518
rect 18060 53454 18062 53506
rect 18114 53454 18116 53506
rect 17724 53060 17780 53070
rect 17724 52388 17780 53004
rect 18060 52836 18116 53454
rect 18172 53060 18228 53098
rect 18172 52994 18228 53004
rect 18172 52836 18228 52846
rect 18060 52780 18172 52836
rect 18172 52770 18228 52780
rect 17724 52322 17780 52332
rect 18060 52388 18116 52398
rect 17836 52164 17892 52202
rect 17500 52108 17836 52164
rect 17388 52098 17444 52108
rect 17836 52098 17892 52108
rect 17948 52162 18004 52174
rect 17948 52110 17950 52162
rect 18002 52110 18004 52162
rect 17836 51940 17892 51950
rect 17500 51938 17892 51940
rect 17500 51886 17838 51938
rect 17890 51886 17892 51938
rect 17500 51884 17892 51886
rect 17500 51716 17556 51884
rect 17836 51874 17892 51884
rect 17052 51650 17108 51660
rect 17164 51660 17556 51716
rect 17948 51716 18004 52110
rect 17052 50820 17108 50830
rect 17052 50706 17108 50764
rect 17052 50654 17054 50706
rect 17106 50654 17108 50706
rect 17052 50642 17108 50654
rect 16436 50540 16772 50596
rect 16828 50540 16996 50596
rect 17164 50594 17220 51660
rect 17948 51650 18004 51660
rect 17612 51604 17668 51614
rect 17164 50542 17166 50594
rect 17218 50542 17220 50594
rect 16380 50428 16436 50540
rect 16380 50372 16660 50428
rect 16044 50370 16100 50372
rect 16044 50318 16046 50370
rect 16098 50318 16100 50370
rect 16044 50306 16100 50318
rect 15932 49746 15988 49756
rect 16492 50036 16548 50046
rect 16492 49810 16548 49980
rect 16492 49758 16494 49810
rect 16546 49758 16548 49810
rect 15820 49522 15876 49532
rect 16156 49700 16212 49710
rect 16492 49700 16548 49758
rect 16156 49698 16548 49700
rect 16156 49646 16158 49698
rect 16210 49646 16548 49698
rect 16156 49644 16548 49646
rect 15820 49028 15876 49038
rect 15820 48934 15876 48972
rect 16156 48916 16212 49644
rect 16604 49588 16660 50372
rect 16156 48850 16212 48860
rect 16268 49532 16660 49588
rect 16828 49922 16884 50540
rect 17164 50530 17220 50542
rect 17500 51548 17612 51604
rect 17500 50594 17556 51548
rect 17612 51538 17668 51548
rect 17500 50542 17502 50594
rect 17554 50542 17556 50594
rect 17500 50530 17556 50542
rect 17612 51378 17668 51390
rect 17612 51326 17614 51378
rect 17666 51326 17668 51378
rect 16828 49870 16830 49922
rect 16882 49870 16884 49922
rect 15204 48748 15316 48804
rect 15148 48738 15204 48748
rect 15260 46900 15316 46910
rect 15148 46004 15204 46014
rect 15148 45910 15204 45948
rect 15260 45890 15316 46844
rect 16044 46900 16100 46910
rect 16044 46562 16100 46844
rect 16044 46510 16046 46562
rect 16098 46510 16100 46562
rect 16044 46498 16100 46510
rect 15260 45838 15262 45890
rect 15314 45838 15316 45890
rect 15260 45826 15316 45838
rect 15708 45892 15764 45902
rect 15708 45798 15764 45836
rect 15148 45666 15204 45678
rect 15148 45614 15150 45666
rect 15202 45614 15204 45666
rect 15148 44548 15204 45614
rect 15484 45666 15540 45678
rect 15484 45614 15486 45666
rect 15538 45614 15540 45666
rect 15372 45220 15428 45230
rect 15260 45108 15316 45118
rect 15260 45014 15316 45052
rect 15148 44482 15204 44492
rect 15372 44994 15428 45164
rect 15372 44942 15374 44994
rect 15426 44942 15428 44994
rect 14700 44380 15092 44436
rect 14476 44210 14532 44222
rect 14476 44158 14478 44210
rect 14530 44158 14532 44210
rect 14476 43652 14532 44158
rect 14700 43708 14756 44380
rect 14476 43586 14532 43596
rect 14588 43652 14756 43708
rect 14924 44212 14980 44222
rect 15260 44212 15316 44222
rect 14924 44210 15316 44212
rect 14924 44158 14926 44210
rect 14978 44158 15262 44210
rect 15314 44158 15316 44210
rect 14924 44156 15316 44158
rect 14924 43708 14980 44156
rect 15260 44146 15316 44156
rect 14924 43652 15092 43708
rect 14364 43148 14532 43204
rect 14364 42980 14420 42990
rect 14364 42886 14420 42924
rect 14476 42756 14532 43148
rect 14364 42700 14532 42756
rect 14252 41860 14308 41870
rect 14140 41858 14308 41860
rect 14140 41806 14254 41858
rect 14306 41806 14308 41858
rect 14140 41804 14308 41806
rect 14028 41300 14084 41310
rect 14028 41186 14084 41244
rect 14028 41134 14030 41186
rect 14082 41134 14084 41186
rect 14028 41122 14084 41134
rect 14252 41188 14308 41804
rect 14252 41122 14308 41132
rect 14364 41186 14420 42700
rect 14588 42644 14644 43652
rect 14700 43426 14756 43438
rect 14700 43374 14702 43426
rect 14754 43374 14756 43426
rect 14700 42978 14756 43374
rect 14700 42926 14702 42978
rect 14754 42926 14756 42978
rect 14700 42914 14756 42926
rect 14364 41134 14366 41186
rect 14418 41134 14420 41186
rect 14364 41122 14420 41134
rect 14476 42588 14644 42644
rect 14700 42754 14756 42766
rect 14700 42702 14702 42754
rect 14754 42702 14756 42754
rect 13804 40898 13860 40908
rect 14140 40962 14196 40974
rect 14140 40910 14142 40962
rect 14194 40910 14196 40962
rect 14140 40740 14196 40910
rect 13356 40574 13358 40626
rect 13410 40574 13412 40626
rect 13356 40562 13412 40574
rect 13580 40684 14196 40740
rect 13580 40514 13636 40684
rect 13580 40462 13582 40514
rect 13634 40462 13636 40514
rect 13580 40450 13636 40462
rect 14028 40516 14084 40526
rect 14028 40404 14084 40460
rect 13692 40402 14196 40404
rect 13692 40350 14030 40402
rect 14082 40350 14196 40402
rect 13692 40348 14196 40350
rect 13468 40292 13524 40302
rect 13468 40198 13524 40236
rect 13580 39620 13636 39630
rect 13692 39620 13748 40348
rect 14028 40338 14084 40348
rect 13636 39564 13748 39620
rect 13580 39526 13636 39564
rect 13580 39060 13636 39070
rect 13580 38966 13636 39004
rect 14140 39058 14196 40348
rect 14252 40292 14308 40302
rect 14252 39730 14308 40236
rect 14252 39678 14254 39730
rect 14306 39678 14308 39730
rect 14252 39666 14308 39678
rect 14140 39006 14142 39058
rect 14194 39006 14196 39058
rect 13356 38948 13412 38958
rect 13244 38946 13412 38948
rect 13244 38894 13358 38946
rect 13410 38894 13412 38946
rect 13244 38892 13412 38894
rect 13356 38882 13412 38892
rect 13692 38612 13748 38622
rect 13916 38612 13972 38622
rect 13692 38610 13972 38612
rect 13692 38558 13694 38610
rect 13746 38558 13918 38610
rect 13970 38558 13972 38610
rect 13692 38556 13972 38558
rect 13692 38546 13748 38556
rect 13916 38546 13972 38556
rect 14140 38164 14196 39006
rect 14140 38098 14196 38108
rect 14252 38610 14308 38622
rect 14252 38558 14254 38610
rect 14306 38558 14308 38610
rect 13804 38052 13860 38062
rect 14252 38052 14308 38558
rect 14364 38052 14420 38062
rect 14252 38050 14420 38052
rect 14252 37998 14366 38050
rect 14418 37998 14420 38050
rect 14252 37996 14420 37998
rect 13804 37958 13860 37996
rect 14364 37986 14420 37996
rect 14028 37938 14084 37950
rect 14028 37886 14030 37938
rect 14082 37886 14084 37938
rect 12684 36430 12686 36482
rect 12738 36430 12740 36482
rect 12460 35980 12628 36036
rect 12460 35812 12516 35822
rect 12460 35586 12516 35756
rect 12460 35534 12462 35586
rect 12514 35534 12516 35586
rect 12460 35522 12516 35534
rect 12572 35476 12628 35980
rect 12572 35410 12628 35420
rect 12684 35252 12740 36430
rect 12796 37154 13188 37156
rect 12796 37102 12910 37154
rect 12962 37102 13188 37154
rect 12796 37100 13188 37102
rect 13356 37268 13412 37278
rect 13804 37268 13860 37278
rect 13356 37266 13860 37268
rect 13356 37214 13358 37266
rect 13410 37214 13806 37266
rect 13858 37214 13860 37266
rect 13356 37212 13860 37214
rect 13356 37156 13412 37212
rect 13804 37202 13860 37212
rect 12796 36148 12852 37100
rect 12908 37090 12964 37100
rect 13356 37090 13412 37100
rect 13356 36484 13412 36494
rect 12908 36372 12964 36382
rect 13356 36372 13412 36428
rect 13804 36484 13860 36494
rect 13804 36390 13860 36428
rect 12908 36370 13412 36372
rect 12908 36318 12910 36370
rect 12962 36318 13412 36370
rect 12908 36316 13412 36318
rect 12908 36306 12964 36316
rect 12796 36092 13076 36148
rect 12236 35196 12740 35252
rect 12908 35588 12964 35598
rect 12236 34356 12292 34366
rect 12236 34262 12292 34300
rect 12572 33908 12628 35196
rect 12684 34356 12740 34366
rect 12908 34356 12964 35532
rect 12740 34300 12964 34356
rect 12684 34130 12740 34300
rect 12684 34078 12686 34130
rect 12738 34078 12740 34130
rect 12684 34066 12740 34078
rect 12572 33852 12740 33908
rect 11676 31726 11678 31778
rect 11730 31726 11732 31778
rect 11676 31714 11732 31726
rect 11788 32172 12068 32228
rect 12348 33346 12404 33358
rect 12348 33294 12350 33346
rect 12402 33294 12404 33346
rect 12348 32452 12404 33294
rect 11564 31500 11732 31556
rect 11340 30994 11508 30996
rect 11340 30942 11342 30994
rect 11394 30942 11508 30994
rect 11340 30940 11508 30942
rect 11340 30930 11396 30940
rect 11116 30882 11172 30894
rect 11116 30830 11118 30882
rect 11170 30830 11172 30882
rect 11004 30772 11060 30782
rect 11004 30434 11060 30716
rect 11116 30660 11172 30830
rect 11564 30770 11620 30782
rect 11564 30718 11566 30770
rect 11618 30718 11620 30770
rect 11564 30660 11620 30718
rect 11116 30604 11620 30660
rect 11004 30382 11006 30434
rect 11058 30382 11060 30434
rect 11004 30370 11060 30382
rect 11564 30436 11620 30604
rect 11564 30370 11620 30380
rect 11676 30098 11732 31500
rect 11676 30046 11678 30098
rect 11730 30046 11732 30098
rect 11676 30034 11732 30046
rect 11004 28308 11060 28318
rect 10892 28252 11004 28308
rect 11004 28242 11060 28252
rect 11564 28308 11620 28318
rect 11564 27970 11620 28252
rect 11564 27918 11566 27970
rect 11618 27918 11620 27970
rect 11564 27906 11620 27918
rect 11788 27860 11844 32172
rect 12124 31668 12180 31678
rect 12124 31554 12180 31612
rect 12124 31502 12126 31554
rect 12178 31502 12180 31554
rect 12124 31444 12180 31502
rect 12348 31444 12404 32396
rect 12684 31668 12740 33852
rect 12796 31892 12852 34300
rect 12908 33348 12964 33358
rect 12908 33254 12964 33292
rect 12908 31892 12964 31902
rect 12796 31890 12964 31892
rect 12796 31838 12910 31890
rect 12962 31838 12964 31890
rect 12796 31836 12964 31838
rect 12908 31826 12964 31836
rect 12684 31612 12964 31668
rect 12124 31388 12404 31444
rect 11900 30996 11956 31006
rect 12236 30996 12292 31006
rect 11900 30994 12292 30996
rect 11900 30942 11902 30994
rect 11954 30942 12238 30994
rect 12290 30942 12292 30994
rect 11900 30940 12292 30942
rect 11900 30930 11956 30940
rect 12236 30930 12292 30940
rect 12012 29988 12068 29998
rect 12012 29894 12068 29932
rect 12236 29426 12292 29438
rect 12236 29374 12238 29426
rect 12290 29374 12292 29426
rect 11788 27766 11844 27804
rect 11900 29316 11956 29326
rect 12236 29316 12292 29374
rect 11900 29314 12292 29316
rect 11900 29262 11902 29314
rect 11954 29262 12292 29314
rect 11900 29260 12292 29262
rect 11788 27412 11844 27422
rect 11004 26962 11060 26974
rect 11004 26910 11006 26962
rect 11058 26910 11060 26962
rect 10332 26852 10612 26908
rect 10668 26852 10948 26908
rect 9996 26516 10052 26526
rect 9996 26290 10052 26460
rect 9996 26238 9998 26290
rect 10050 26238 10052 26290
rect 9996 26226 10052 26238
rect 10444 26068 10500 26078
rect 10332 26012 10444 26068
rect 10332 25506 10388 26012
rect 10444 26002 10500 26012
rect 10332 25454 10334 25506
rect 10386 25454 10388 25506
rect 10332 25442 10388 25454
rect 9996 25396 10052 25406
rect 9772 25394 10052 25396
rect 9772 25342 9998 25394
rect 10050 25342 10052 25394
rect 9772 25340 10052 25342
rect 9660 25172 9716 25182
rect 9660 24946 9716 25116
rect 9660 24894 9662 24946
rect 9714 24894 9716 24946
rect 9660 24882 9716 24894
rect 9548 24052 9604 24062
rect 9548 23958 9604 23996
rect 9436 23426 9492 23436
rect 8764 23380 8820 23390
rect 8764 23286 8820 23324
rect 7420 23174 7476 23212
rect 7644 23212 8148 23268
rect 9660 23268 9716 23278
rect 7308 23154 7364 23166
rect 7308 23102 7310 23154
rect 7362 23102 7364 23154
rect 7308 22484 7364 23102
rect 7532 22484 7588 22494
rect 7308 22482 7588 22484
rect 7308 22430 7534 22482
rect 7586 22430 7588 22482
rect 7308 22428 7588 22430
rect 7532 22372 7588 22428
rect 7532 22306 7588 22316
rect 7308 21924 7364 21934
rect 7308 20916 7364 21868
rect 6972 20578 7028 20590
rect 6972 20526 6974 20578
rect 7026 20526 7028 20578
rect 6972 20244 7028 20526
rect 7308 20580 7364 20860
rect 7420 20804 7476 20814
rect 7420 20710 7476 20748
rect 7308 20514 7364 20524
rect 7532 20578 7588 20590
rect 7532 20526 7534 20578
rect 7586 20526 7588 20578
rect 7532 20356 7588 20526
rect 7532 20290 7588 20300
rect 6804 20188 7028 20244
rect 6748 20130 6804 20188
rect 6748 20078 6750 20130
rect 6802 20078 6804 20130
rect 6748 20066 6804 20078
rect 7308 20130 7364 20142
rect 7308 20078 7310 20130
rect 7362 20078 7364 20130
rect 7084 20020 7140 20030
rect 6412 19516 6580 19572
rect 6860 20018 7140 20020
rect 6860 19966 7086 20018
rect 7138 19966 7140 20018
rect 6860 19964 7140 19966
rect 6412 19460 6468 19516
rect 6860 19460 6916 19964
rect 7084 19954 7140 19964
rect 6076 19404 6244 19460
rect 6188 19348 6244 19404
rect 6412 19394 6468 19404
rect 6524 19404 6916 19460
rect 6972 19796 7028 19806
rect 6076 19234 6132 19246
rect 6076 19182 6078 19234
rect 6130 19182 6132 19234
rect 5628 19124 5684 19134
rect 6076 19124 6132 19182
rect 5628 19122 6020 19124
rect 5628 19070 5630 19122
rect 5682 19070 6020 19122
rect 5628 19068 6020 19070
rect 5628 19058 5684 19068
rect 5964 18900 6020 19068
rect 6076 19058 6132 19068
rect 5964 18844 6132 18900
rect 5180 18674 5908 18676
rect 5180 18622 5182 18674
rect 5234 18622 5908 18674
rect 5180 18620 5908 18622
rect 5180 18610 5236 18620
rect 5852 18562 5908 18620
rect 5852 18510 5854 18562
rect 5906 18510 5908 18562
rect 5852 18498 5908 18510
rect 6076 18562 6132 18844
rect 6076 18510 6078 18562
rect 6130 18510 6132 18562
rect 6076 18498 6132 18510
rect 5740 18452 5796 18462
rect 5068 18340 5124 18350
rect 5068 18246 5124 18284
rect 5740 18338 5796 18396
rect 6188 18340 6244 19292
rect 6524 19346 6580 19404
rect 6524 19294 6526 19346
rect 6578 19294 6580 19346
rect 6524 19282 6580 19294
rect 6972 18450 7028 19740
rect 7308 19460 7364 20078
rect 7420 20132 7476 20142
rect 7644 20132 7700 23212
rect 9660 23174 9716 23212
rect 8876 23156 8932 23166
rect 8876 23062 8932 23100
rect 9548 23154 9604 23166
rect 9548 23102 9550 23154
rect 9602 23102 9604 23154
rect 8428 23042 8484 23054
rect 8428 22990 8430 23042
rect 8482 22990 8484 23042
rect 8428 22932 8484 22990
rect 8988 22932 9044 22942
rect 8428 22930 9044 22932
rect 8428 22878 8990 22930
rect 9042 22878 9044 22930
rect 8428 22876 9044 22878
rect 7980 22370 8036 22382
rect 7980 22318 7982 22370
rect 8034 22318 8036 22370
rect 7868 22260 7924 22270
rect 7868 22166 7924 22204
rect 7980 21476 8036 22318
rect 8316 22370 8372 22382
rect 8316 22318 8318 22370
rect 8370 22318 8372 22370
rect 8316 21924 8372 22318
rect 8316 21858 8372 21868
rect 8316 21588 8372 21598
rect 8204 21586 8372 21588
rect 8204 21534 8318 21586
rect 8370 21534 8372 21586
rect 8204 21532 8372 21534
rect 7756 21420 8036 21476
rect 8092 21476 8148 21486
rect 7756 20802 7812 21420
rect 7756 20750 7758 20802
rect 7810 20750 7812 20802
rect 7756 20738 7812 20750
rect 7980 21028 8036 21038
rect 7980 20802 8036 20972
rect 7980 20750 7982 20802
rect 8034 20750 8036 20802
rect 7980 20738 8036 20750
rect 8092 20804 8148 21420
rect 8204 21028 8260 21532
rect 8316 21522 8372 21532
rect 8428 21028 8484 22876
rect 8988 22866 9044 22876
rect 9212 22148 9268 22158
rect 8652 22146 9268 22148
rect 8652 22094 9214 22146
rect 9266 22094 9268 22146
rect 8652 22092 9268 22094
rect 8204 20962 8260 20972
rect 8316 20972 8484 21028
rect 8540 21588 8596 21598
rect 8540 21026 8596 21532
rect 8540 20974 8542 21026
rect 8594 20974 8596 21026
rect 8204 20804 8260 20814
rect 8092 20802 8260 20804
rect 8092 20750 8206 20802
rect 8258 20750 8260 20802
rect 8092 20748 8260 20750
rect 8204 20738 8260 20748
rect 8316 20580 8372 20972
rect 8540 20962 8596 20974
rect 8428 20804 8484 20814
rect 8652 20804 8708 22092
rect 9212 22082 9268 22092
rect 9324 22146 9380 22158
rect 9324 22094 9326 22146
rect 9378 22094 9380 22146
rect 9324 21924 9380 22094
rect 9436 22146 9492 22158
rect 9436 22094 9438 22146
rect 9490 22094 9492 22146
rect 9436 22036 9492 22094
rect 9436 21970 9492 21980
rect 8876 21868 9380 21924
rect 8876 21586 8932 21868
rect 9548 21812 9604 23102
rect 8988 21756 9604 21812
rect 9660 22146 9716 22158
rect 9660 22094 9662 22146
rect 9714 22094 9716 22146
rect 8988 21698 9044 21756
rect 8988 21646 8990 21698
rect 9042 21646 9044 21698
rect 8988 21634 9044 21646
rect 8876 21534 8878 21586
rect 8930 21534 8932 21586
rect 8876 21522 8932 21534
rect 9436 21588 9492 21598
rect 9436 21494 9492 21532
rect 9436 21364 9492 21374
rect 8876 21028 8932 21038
rect 8932 20972 9044 21028
rect 8876 20962 8932 20972
rect 8428 20802 8596 20804
rect 8428 20750 8430 20802
rect 8482 20750 8596 20802
rect 8428 20748 8596 20750
rect 8428 20738 8484 20748
rect 8540 20580 8596 20748
rect 8316 20524 8484 20580
rect 7420 20130 7700 20132
rect 7420 20078 7422 20130
rect 7474 20078 7700 20130
rect 7420 20076 7700 20078
rect 7420 20066 7476 20076
rect 7756 20018 7812 20030
rect 7756 19966 7758 20018
rect 7810 19966 7812 20018
rect 7420 19908 7476 19918
rect 7756 19908 7812 19966
rect 7980 20020 8036 20030
rect 7980 20018 8260 20020
rect 7980 19966 7982 20018
rect 8034 19966 8260 20018
rect 7980 19964 8260 19966
rect 7980 19954 8036 19964
rect 7476 19852 7812 19908
rect 7420 19842 7476 19852
rect 8092 19794 8148 19806
rect 8092 19742 8094 19794
rect 8146 19742 8148 19794
rect 7308 19404 7924 19460
rect 7532 19234 7588 19246
rect 7532 19182 7534 19234
rect 7586 19182 7588 19234
rect 7532 19012 7588 19182
rect 7532 18946 7588 18956
rect 7868 18674 7924 19404
rect 7868 18622 7870 18674
rect 7922 18622 7924 18674
rect 6972 18398 6974 18450
rect 7026 18398 7028 18450
rect 5740 18286 5742 18338
rect 5794 18286 5796 18338
rect 5740 18274 5796 18286
rect 5852 18284 6244 18340
rect 6524 18338 6580 18350
rect 6524 18286 6526 18338
rect 6578 18286 6580 18338
rect 5404 18226 5460 18238
rect 5404 18174 5406 18226
rect 5458 18174 5460 18226
rect 5404 18116 5460 18174
rect 5404 18060 5572 18116
rect 5516 17890 5572 18060
rect 5516 17838 5518 17890
rect 5570 17838 5572 17890
rect 5516 17826 5572 17838
rect 4620 17778 5012 17780
rect 4620 17726 4622 17778
rect 4674 17726 5012 17778
rect 4620 17724 5012 17726
rect 5068 17780 5124 17790
rect 4620 17668 4676 17724
rect 5068 17686 5124 17724
rect 5852 17778 5908 18284
rect 6524 17890 6580 18286
rect 6972 18228 7028 18398
rect 6972 18162 7028 18172
rect 7308 18564 7364 18574
rect 7308 18116 7364 18508
rect 7868 18452 7924 18622
rect 7868 18386 7924 18396
rect 8092 19124 8148 19742
rect 8092 18450 8148 19068
rect 8092 18398 8094 18450
rect 8146 18398 8148 18450
rect 8092 18386 8148 18398
rect 7420 18340 7476 18350
rect 7420 18338 7812 18340
rect 7420 18286 7422 18338
rect 7474 18286 7812 18338
rect 7420 18284 7812 18286
rect 7420 18274 7476 18284
rect 7756 18228 7812 18284
rect 7980 18338 8036 18350
rect 7980 18286 7982 18338
rect 8034 18286 8036 18338
rect 7980 18228 8036 18286
rect 7756 18172 8036 18228
rect 7308 18060 7476 18116
rect 6860 17892 6916 17902
rect 6524 17838 6526 17890
rect 6578 17838 6580 17890
rect 6524 17826 6580 17838
rect 6748 17890 6916 17892
rect 6748 17838 6862 17890
rect 6914 17838 6916 17890
rect 6748 17836 6916 17838
rect 5852 17726 5854 17778
rect 5906 17726 5908 17778
rect 5852 17714 5908 17726
rect 4172 17612 4676 17668
rect 6188 17668 6244 17678
rect 4172 16994 4228 17612
rect 6188 17574 6244 17612
rect 4284 17108 4340 17118
rect 4284 17014 4340 17052
rect 4172 16942 4174 16994
rect 4226 16942 4228 16994
rect 4172 16930 4228 16942
rect 5628 16994 5684 17006
rect 5628 16942 5630 16994
rect 5682 16942 5684 16994
rect 4060 16884 4116 16894
rect 3948 16882 4116 16884
rect 3948 16830 4062 16882
rect 4114 16830 4116 16882
rect 3948 16828 4116 16830
rect 4060 16212 4116 16828
rect 5068 16882 5124 16894
rect 5068 16830 5070 16882
rect 5122 16830 5124 16882
rect 4284 16772 4340 16782
rect 4060 16146 4116 16156
rect 4172 16716 4284 16772
rect 3836 15262 3838 15314
rect 3890 15262 3892 15314
rect 3836 15250 3892 15262
rect 4060 15316 4116 15326
rect 4060 15222 4116 15260
rect 4172 15314 4228 16716
rect 4284 16706 4340 16716
rect 5068 16772 5124 16830
rect 5068 16706 5124 16716
rect 5180 16884 5236 16894
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4620 16212 4676 16222
rect 5068 16212 5124 16222
rect 5180 16212 5236 16828
rect 4676 16156 5012 16212
rect 4620 16118 4676 16156
rect 4732 15764 4788 15774
rect 4732 15538 4788 15708
rect 4732 15486 4734 15538
rect 4786 15486 4788 15538
rect 4732 15474 4788 15486
rect 4844 15652 4900 15662
rect 4172 15262 4174 15314
rect 4226 15262 4228 15314
rect 4172 14980 4228 15262
rect 4508 15316 4564 15326
rect 4508 15222 4564 15260
rect 3612 14590 3614 14642
rect 3666 14590 3668 14642
rect 3612 14578 3668 14590
rect 4060 14924 4228 14980
rect 4476 14924 4740 14934
rect 4060 14418 4116 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4396 14754 4452 14766
rect 4396 14702 4398 14754
rect 4450 14702 4452 14754
rect 4172 14532 4228 14542
rect 4396 14532 4452 14702
rect 4620 14644 4676 14654
rect 4844 14644 4900 15596
rect 4956 15538 5012 16156
rect 5068 16210 5236 16212
rect 5068 16158 5070 16210
rect 5122 16158 5236 16210
rect 5068 16156 5236 16158
rect 5516 16772 5572 16782
rect 5068 16146 5124 16156
rect 4956 15486 4958 15538
rect 5010 15486 5012 15538
rect 4956 15474 5012 15486
rect 5516 15538 5572 16716
rect 5516 15486 5518 15538
rect 5570 15486 5572 15538
rect 5068 15314 5124 15326
rect 5068 15262 5070 15314
rect 5122 15262 5124 15314
rect 5068 15148 5124 15262
rect 5516 15148 5572 15486
rect 4620 14642 4900 14644
rect 4620 14590 4622 14642
rect 4674 14590 4900 14642
rect 4620 14588 4900 14590
rect 4956 15092 5124 15148
rect 5180 15092 5572 15148
rect 4956 14754 5012 15092
rect 4956 14702 4958 14754
rect 5010 14702 5012 14754
rect 4620 14578 4676 14588
rect 4172 14530 4452 14532
rect 4172 14478 4174 14530
rect 4226 14478 4452 14530
rect 4172 14476 4452 14478
rect 4172 14466 4228 14476
rect 4060 14366 4062 14418
rect 4114 14366 4116 14418
rect 3836 14306 3892 14318
rect 3836 14254 3838 14306
rect 3890 14254 3892 14306
rect 3500 13356 3668 13412
rect 3388 13244 3556 13300
rect 3388 13076 3444 13086
rect 3388 12982 3444 13020
rect 3276 12910 3278 12962
rect 3330 12910 3332 12962
rect 3276 12898 3332 12910
rect 2716 12798 2718 12850
rect 2770 12798 2772 12850
rect 2716 12786 2772 12798
rect 2044 12740 2100 12750
rect 2044 12646 2100 12684
rect 3500 12738 3556 13244
rect 3500 12686 3502 12738
rect 3554 12686 3556 12738
rect 2044 12516 2100 12526
rect 2044 12402 2100 12460
rect 2044 12350 2046 12402
rect 2098 12350 2100 12402
rect 2044 12338 2100 12350
rect 2828 12404 2884 12414
rect 3388 12404 3444 12414
rect 3500 12404 3556 12686
rect 2828 12402 3556 12404
rect 2828 12350 2830 12402
rect 2882 12350 3390 12402
rect 3442 12350 3556 12402
rect 2828 12348 3556 12350
rect 3612 12404 3668 13356
rect 3836 12962 3892 14254
rect 4060 14308 4116 14366
rect 4060 14252 4676 14308
rect 4620 13634 4676 14252
rect 4956 13972 5012 14702
rect 5068 14532 5124 14542
rect 5068 14438 5124 14476
rect 4620 13582 4622 13634
rect 4674 13582 4676 13634
rect 4620 13570 4676 13582
rect 4844 13916 5012 13972
rect 3836 12910 3838 12962
rect 3890 12910 3892 12962
rect 3836 12898 3892 12910
rect 4284 13412 4340 13422
rect 4284 12850 4340 13356
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4844 13188 4900 13916
rect 4396 13132 4900 13188
rect 4956 13746 5012 13758
rect 4956 13694 4958 13746
rect 5010 13694 5012 13746
rect 4396 12962 4452 13132
rect 4396 12910 4398 12962
rect 4450 12910 4452 12962
rect 4396 12898 4452 12910
rect 4284 12798 4286 12850
rect 4338 12798 4340 12850
rect 4060 12740 4116 12750
rect 2828 12338 2884 12348
rect 3388 12310 3444 12348
rect 3612 12338 3668 12348
rect 3836 12738 4116 12740
rect 3836 12686 4062 12738
rect 4114 12686 4116 12738
rect 3836 12684 4116 12686
rect 2492 12178 2548 12190
rect 2492 12126 2494 12178
rect 2546 12126 2548 12178
rect 2492 11732 2548 12126
rect 3164 12178 3220 12190
rect 3164 12126 3166 12178
rect 3218 12126 3220 12178
rect 2492 11666 2548 11676
rect 2604 12068 2660 12078
rect 1820 11342 1822 11394
rect 1874 11342 1876 11394
rect 1820 9828 1876 11342
rect 2044 11620 2100 11630
rect 2044 10834 2100 11564
rect 2492 11508 2548 11518
rect 2604 11508 2660 12012
rect 2492 11506 2660 11508
rect 2492 11454 2494 11506
rect 2546 11454 2660 11506
rect 2492 11452 2660 11454
rect 3164 11508 3220 12126
rect 3836 12178 3892 12684
rect 4060 12674 4116 12684
rect 4172 12628 4228 12638
rect 4172 12402 4228 12572
rect 4172 12350 4174 12402
rect 4226 12350 4228 12402
rect 4172 12338 4228 12350
rect 3836 12126 3838 12178
rect 3890 12126 3892 12178
rect 3836 12114 3892 12126
rect 3276 12068 3332 12078
rect 3276 11974 3332 12012
rect 2492 11442 2548 11452
rect 3164 11442 3220 11452
rect 3388 11956 3444 11966
rect 2716 11396 2772 11406
rect 2044 10782 2046 10834
rect 2098 10782 2100 10834
rect 2044 10770 2100 10782
rect 2380 10836 2436 10846
rect 2380 10724 2436 10780
rect 2716 10834 2772 11340
rect 2716 10782 2718 10834
rect 2770 10782 2772 10834
rect 2716 10770 2772 10782
rect 3388 10834 3444 11900
rect 3388 10782 3390 10834
rect 3442 10782 3444 10834
rect 3388 10770 3444 10782
rect 3948 11732 4004 11742
rect 3948 10836 4004 11676
rect 4284 11620 4340 12798
rect 4508 12404 4564 12414
rect 4508 12310 4564 12348
rect 4732 12068 4788 13132
rect 4956 13076 5012 13694
rect 5068 13636 5124 13646
rect 5068 13542 5124 13580
rect 4956 13010 5012 13020
rect 4844 12852 4900 12862
rect 5180 12852 5236 15092
rect 5628 14756 5684 16942
rect 6636 16772 6692 16782
rect 6636 16678 6692 16716
rect 6748 16098 6804 17836
rect 6860 17826 6916 17836
rect 7308 17780 7364 17790
rect 6972 17554 7028 17566
rect 6972 17502 6974 17554
rect 7026 17502 7028 17554
rect 6860 17442 6916 17454
rect 6860 17390 6862 17442
rect 6914 17390 6916 17442
rect 6860 17332 6916 17390
rect 6860 17266 6916 17276
rect 6972 16548 7028 17502
rect 7308 17554 7364 17724
rect 7308 17502 7310 17554
rect 7362 17502 7364 17554
rect 7308 17490 7364 17502
rect 6972 16482 7028 16492
rect 6748 16046 6750 16098
rect 6802 16046 6804 16098
rect 6748 16034 6804 16046
rect 6972 16324 7028 16334
rect 6972 16098 7028 16268
rect 6972 16046 6974 16098
rect 7026 16046 7028 16098
rect 6972 16034 7028 16046
rect 6188 15988 6244 15998
rect 6524 15988 6580 15998
rect 6188 15986 6580 15988
rect 6188 15934 6190 15986
rect 6242 15934 6526 15986
rect 6578 15934 6580 15986
rect 6188 15932 6580 15934
rect 6188 15922 6244 15932
rect 6524 15922 6580 15932
rect 5964 15874 6020 15886
rect 5964 15822 5966 15874
rect 6018 15822 6020 15874
rect 5964 15540 6020 15822
rect 5964 15474 6020 15484
rect 6076 15874 6132 15886
rect 6076 15822 6078 15874
rect 6130 15822 6132 15874
rect 6076 15316 6132 15822
rect 7084 15876 7140 15886
rect 6076 15250 6132 15260
rect 6188 15540 6244 15550
rect 5964 15202 6020 15214
rect 5964 15150 5966 15202
rect 6018 15150 6020 15202
rect 5964 15092 6020 15150
rect 6188 15148 6244 15484
rect 6748 15316 6804 15326
rect 6636 15202 6692 15214
rect 6636 15150 6638 15202
rect 6690 15150 6692 15202
rect 6636 15148 6692 15150
rect 5964 15026 6020 15036
rect 6076 15092 6244 15148
rect 6300 15092 6692 15148
rect 5292 14700 5684 14756
rect 5292 13858 5348 14700
rect 5964 14644 6020 14654
rect 5292 13806 5294 13858
rect 5346 13806 5348 13858
rect 5292 13524 5348 13806
rect 5516 14642 6020 14644
rect 5516 14590 5966 14642
rect 6018 14590 6020 14642
rect 5516 14588 6020 14590
rect 5516 13858 5572 14588
rect 5964 14578 6020 14588
rect 5516 13806 5518 13858
rect 5570 13806 5572 13858
rect 5516 13794 5572 13806
rect 6076 14418 6132 15092
rect 6300 14754 6356 15092
rect 6748 14980 6804 15260
rect 7084 15314 7140 15820
rect 7084 15262 7086 15314
rect 7138 15262 7140 15314
rect 7084 15204 7140 15262
rect 7084 15138 7140 15148
rect 6300 14702 6302 14754
rect 6354 14702 6356 14754
rect 6300 14690 6356 14702
rect 6636 14924 6804 14980
rect 6972 15092 7028 15102
rect 6636 14530 6692 14924
rect 6636 14478 6638 14530
rect 6690 14478 6692 14530
rect 6636 14466 6692 14478
rect 6076 14366 6078 14418
rect 6130 14366 6132 14418
rect 5292 13458 5348 13468
rect 5740 12964 5796 12974
rect 5740 12870 5796 12908
rect 4844 12850 5236 12852
rect 4844 12798 4846 12850
rect 4898 12798 5236 12850
rect 4844 12796 5236 12798
rect 4844 12786 4900 12796
rect 4844 12292 4900 12302
rect 4900 12236 5012 12292
rect 4844 12198 4900 12236
rect 4732 12012 4900 12068
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4284 11564 4676 11620
rect 4620 11506 4676 11564
rect 4620 11454 4622 11506
rect 4674 11454 4676 11506
rect 4620 11442 4676 11454
rect 4844 10948 4900 12012
rect 4956 11284 5012 12236
rect 4956 11218 5012 11228
rect 5068 11506 5124 12796
rect 5852 12404 5908 12414
rect 5852 12310 5908 12348
rect 6076 12292 6132 14366
rect 6748 14308 6804 14318
rect 6636 14306 6804 14308
rect 6636 14254 6750 14306
rect 6802 14254 6804 14306
rect 6636 14252 6804 14254
rect 6300 13634 6356 13646
rect 6300 13582 6302 13634
rect 6354 13582 6356 13634
rect 6300 12292 6356 13582
rect 6636 13074 6692 14252
rect 6748 14242 6804 14252
rect 6860 14306 6916 14318
rect 6860 14254 6862 14306
rect 6914 14254 6916 14306
rect 6860 13748 6916 14254
rect 6972 13972 7028 15036
rect 7420 15092 7476 18060
rect 7644 17780 7700 17790
rect 7644 17778 7924 17780
rect 7644 17726 7646 17778
rect 7698 17726 7924 17778
rect 7644 17724 7924 17726
rect 7644 17714 7700 17724
rect 7532 17556 7588 17566
rect 7532 17462 7588 17500
rect 7756 17556 7812 17566
rect 7756 17462 7812 17500
rect 7868 17332 7924 17724
rect 8092 17556 8148 17566
rect 8204 17556 8260 19964
rect 8428 19796 8484 20524
rect 8540 20514 8596 20524
rect 8652 20130 8708 20748
rect 8876 20802 8932 20814
rect 8876 20750 8878 20802
rect 8930 20750 8932 20802
rect 8876 20692 8932 20750
rect 8876 20626 8932 20636
rect 8988 20690 9044 20972
rect 8988 20638 8990 20690
rect 9042 20638 9044 20690
rect 8988 20626 9044 20638
rect 8652 20078 8654 20130
rect 8706 20078 8708 20130
rect 8652 20066 8708 20078
rect 8876 20132 8932 20142
rect 8876 20038 8932 20076
rect 8988 20020 9044 20030
rect 8988 20018 9268 20020
rect 8988 19966 8990 20018
rect 9042 19966 9268 20018
rect 8988 19964 9268 19966
rect 8988 19954 9044 19964
rect 9212 19908 9268 19964
rect 8428 19740 9156 19796
rect 8428 19348 8484 19358
rect 8484 19292 8596 19348
rect 8428 19254 8484 19292
rect 8316 19236 8372 19246
rect 8316 17780 8372 19180
rect 8316 17666 8372 17724
rect 8316 17614 8318 17666
rect 8370 17614 8372 17666
rect 8316 17602 8372 17614
rect 8428 18450 8484 18462
rect 8428 18398 8430 18450
rect 8482 18398 8484 18450
rect 8148 17500 8260 17556
rect 8092 17462 8148 17500
rect 7868 16098 7924 17276
rect 8204 16548 8260 16558
rect 7868 16046 7870 16098
rect 7922 16046 7924 16098
rect 7868 16034 7924 16046
rect 8092 16324 8148 16334
rect 8092 16098 8148 16268
rect 8092 16046 8094 16098
rect 8146 16046 8148 16098
rect 8092 16034 8148 16046
rect 7980 15874 8036 15886
rect 7980 15822 7982 15874
rect 8034 15822 8036 15874
rect 7532 15316 7588 15326
rect 7980 15316 8036 15822
rect 7532 15314 8036 15316
rect 7532 15262 7534 15314
rect 7586 15262 8036 15314
rect 7532 15260 8036 15262
rect 8092 15426 8148 15438
rect 8092 15374 8094 15426
rect 8146 15374 8148 15426
rect 8092 15316 8148 15374
rect 8204 15426 8260 16492
rect 8204 15374 8206 15426
rect 8258 15374 8260 15426
rect 8204 15362 8260 15374
rect 8316 15876 8372 15886
rect 8428 15876 8484 18398
rect 8540 18452 8596 19292
rect 8540 18386 8596 18396
rect 8652 19012 8708 19022
rect 8652 16882 8708 18956
rect 8988 18788 9044 18798
rect 8876 18676 8932 18686
rect 8876 18582 8932 18620
rect 8988 18562 9044 18732
rect 8988 18510 8990 18562
rect 9042 18510 9044 18562
rect 8988 18498 9044 18510
rect 8764 18340 8820 18350
rect 8820 18284 8932 18340
rect 8764 18274 8820 18284
rect 8876 18226 8932 18284
rect 9100 18228 9156 19740
rect 9212 18676 9268 19852
rect 9436 19796 9492 21308
rect 9660 20356 9716 22094
rect 9772 22148 9828 25340
rect 9996 25330 10052 25340
rect 10108 25172 10164 25182
rect 10108 24946 10164 25116
rect 10108 24894 10110 24946
rect 10162 24894 10164 24946
rect 10108 24882 10164 24894
rect 10556 24724 10612 26852
rect 10556 24658 10612 24668
rect 9884 23716 9940 23726
rect 9884 23380 9940 23660
rect 9884 23314 9940 23324
rect 9884 23154 9940 23166
rect 9884 23102 9886 23154
rect 9938 23102 9940 23154
rect 9884 22596 9940 23102
rect 9996 23156 10052 23166
rect 9996 23062 10052 23100
rect 10556 23042 10612 23054
rect 10556 22990 10558 23042
rect 10610 22990 10612 23042
rect 10556 22932 10612 22990
rect 9884 22540 10052 22596
rect 9996 22484 10052 22540
rect 9996 22418 10052 22428
rect 10556 22484 10612 22876
rect 10556 22418 10612 22428
rect 9772 22092 10052 22148
rect 9660 20290 9716 20300
rect 9772 21810 9828 21822
rect 9772 21758 9774 21810
rect 9826 21758 9828 21810
rect 9548 20020 9604 20030
rect 9548 19926 9604 19964
rect 9772 20018 9828 21758
rect 9772 19966 9774 20018
rect 9826 19966 9828 20018
rect 9772 19954 9828 19966
rect 9884 21586 9940 21598
rect 9884 21534 9886 21586
rect 9938 21534 9940 21586
rect 9884 20020 9940 21534
rect 9884 19954 9940 19964
rect 9436 19740 9604 19796
rect 9212 18610 9268 18620
rect 9324 18788 9380 18798
rect 8876 18174 8878 18226
rect 8930 18174 8932 18226
rect 8876 18162 8932 18174
rect 8988 18172 9156 18228
rect 8876 18004 8932 18014
rect 8876 17668 8932 17948
rect 8876 17574 8932 17612
rect 8988 17444 9044 18172
rect 9324 18004 9380 18732
rect 9324 17938 9380 17948
rect 9324 17668 9380 17678
rect 8652 16830 8654 16882
rect 8706 16830 8708 16882
rect 8652 16818 8708 16830
rect 8876 17388 9044 17444
rect 9100 17666 9380 17668
rect 9100 17614 9326 17666
rect 9378 17614 9380 17666
rect 9100 17612 9380 17614
rect 8764 16324 8820 16334
rect 8764 16230 8820 16268
rect 8316 15874 8484 15876
rect 8316 15822 8318 15874
rect 8370 15822 8484 15874
rect 8316 15820 8484 15822
rect 8316 15652 8372 15820
rect 7532 15250 7588 15260
rect 8092 15250 8148 15260
rect 7420 15026 7476 15036
rect 8092 15090 8148 15102
rect 8092 15038 8094 15090
rect 8146 15038 8148 15090
rect 7532 14700 7924 14756
rect 7532 14642 7588 14700
rect 7532 14590 7534 14642
rect 7586 14590 7588 14642
rect 7532 14578 7588 14590
rect 7308 14530 7364 14542
rect 7308 14478 7310 14530
rect 7362 14478 7364 14530
rect 7308 14420 7364 14478
rect 7756 14532 7812 14542
rect 7756 14438 7812 14476
rect 7308 14354 7364 14364
rect 7756 14196 7812 14206
rect 7196 14084 7252 14094
rect 6972 13916 7140 13972
rect 6972 13748 7028 13758
rect 6860 13746 7028 13748
rect 6860 13694 6974 13746
rect 7026 13694 7028 13746
rect 6860 13692 7028 13694
rect 6636 13022 6638 13074
rect 6690 13022 6692 13074
rect 6636 13010 6692 13022
rect 6972 13412 7028 13692
rect 6412 12962 6468 12974
rect 6412 12910 6414 12962
rect 6466 12910 6468 12962
rect 6412 12516 6468 12910
rect 6412 12450 6468 12460
rect 6412 12292 6468 12302
rect 6300 12290 6468 12292
rect 6300 12238 6414 12290
rect 6466 12238 6468 12290
rect 6300 12236 6468 12238
rect 5292 12180 5348 12190
rect 5292 12086 5348 12124
rect 6076 12178 6132 12236
rect 6412 12226 6468 12236
rect 6860 12292 6916 12302
rect 6860 12198 6916 12236
rect 6076 12126 6078 12178
rect 6130 12126 6132 12178
rect 6076 12114 6132 12126
rect 6076 11954 6132 11966
rect 6076 11902 6078 11954
rect 6130 11902 6132 11954
rect 5068 11454 5070 11506
rect 5122 11454 5124 11506
rect 3948 10742 4004 10780
rect 4284 10892 4900 10948
rect 2156 10722 2436 10724
rect 2156 10670 2382 10722
rect 2434 10670 2436 10722
rect 2156 10668 2436 10670
rect 2044 9828 2100 9838
rect 1820 9772 2044 9828
rect 2044 9734 2100 9772
rect 2156 9266 2212 10668
rect 2380 10658 2436 10668
rect 2492 10724 2548 10734
rect 2156 9214 2158 9266
rect 2210 9214 2212 9266
rect 2156 9202 2212 9214
rect 2492 9266 2548 10668
rect 4284 10722 4340 10892
rect 4844 10834 4900 10892
rect 4844 10782 4846 10834
rect 4898 10782 4900 10834
rect 4844 10770 4900 10782
rect 4284 10670 4286 10722
rect 4338 10670 4340 10722
rect 4284 10658 4340 10670
rect 4396 10724 4452 10734
rect 4396 10630 4452 10668
rect 4956 10724 5012 10734
rect 3052 10610 3108 10622
rect 3052 10558 3054 10610
rect 3106 10558 3108 10610
rect 3052 10164 3108 10558
rect 4396 10388 4452 10398
rect 4284 10386 4452 10388
rect 4284 10334 4398 10386
rect 4450 10334 4452 10386
rect 4284 10332 4452 10334
rect 3052 10098 3108 10108
rect 3836 10164 3892 10174
rect 2716 9716 2772 9726
rect 2716 9622 2772 9660
rect 2492 9214 2494 9266
rect 2546 9214 2548 9266
rect 2492 9202 2548 9214
rect 3836 9266 3892 10108
rect 4284 9940 4340 10332
rect 4396 10322 4452 10332
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4284 9874 4340 9884
rect 4844 9940 4900 9950
rect 4956 9940 5012 10668
rect 4844 9938 5012 9940
rect 4844 9886 4846 9938
rect 4898 9886 5012 9938
rect 4844 9884 5012 9886
rect 4844 9874 4900 9884
rect 3836 9214 3838 9266
rect 3890 9214 3892 9266
rect 3836 9202 3892 9214
rect 5068 9828 5124 11454
rect 5740 11508 5796 11518
rect 5740 11414 5796 11452
rect 6076 11394 6132 11902
rect 6076 11342 6078 11394
rect 6130 11342 6132 11394
rect 6076 11330 6132 11342
rect 6748 11954 6804 11966
rect 6748 11902 6750 11954
rect 6802 11902 6804 11954
rect 5628 11284 5684 11294
rect 5516 10836 5572 10846
rect 5516 10742 5572 10780
rect 5180 10610 5236 10622
rect 5180 10558 5182 10610
rect 5234 10558 5236 10610
rect 5180 10388 5236 10558
rect 5628 10500 5684 11228
rect 5964 11282 6020 11294
rect 5964 11230 5966 11282
rect 6018 11230 6020 11282
rect 5628 10434 5684 10444
rect 5852 10722 5908 10734
rect 5852 10670 5854 10722
rect 5906 10670 5908 10722
rect 5180 10322 5236 10332
rect 4620 9044 4676 9054
rect 5068 9044 5124 9772
rect 5516 9940 5572 9950
rect 5516 9826 5572 9884
rect 5516 9774 5518 9826
rect 5570 9774 5572 9826
rect 5516 9762 5572 9774
rect 5852 9828 5908 10670
rect 5964 10724 6020 11230
rect 5964 10658 6020 10668
rect 6748 10722 6804 11902
rect 6860 11956 6916 11966
rect 6972 11956 7028 13356
rect 7084 13076 7140 13916
rect 7196 13746 7252 14028
rect 7644 13860 7700 13870
rect 7644 13766 7700 13804
rect 7196 13694 7198 13746
rect 7250 13694 7252 13746
rect 7196 13682 7252 13694
rect 7084 13020 7364 13076
rect 7084 12850 7140 12862
rect 7084 12798 7086 12850
rect 7138 12798 7140 12850
rect 7084 12290 7140 12798
rect 7084 12238 7086 12290
rect 7138 12238 7140 12290
rect 7084 12226 7140 12238
rect 6916 11900 7028 11956
rect 6860 11890 6916 11900
rect 7308 10836 7364 13020
rect 7756 12964 7812 14140
rect 7644 12962 7812 12964
rect 7644 12910 7758 12962
rect 7810 12910 7812 12962
rect 7644 12908 7812 12910
rect 7644 11620 7700 12908
rect 7756 12898 7812 12908
rect 7868 13746 7924 14700
rect 7980 14530 8036 14542
rect 7980 14478 7982 14530
rect 8034 14478 8036 14530
rect 7980 14308 8036 14478
rect 7980 14242 8036 14252
rect 7980 14084 8036 14094
rect 8092 14084 8148 15038
rect 8036 14028 8148 14084
rect 8204 14532 8260 14542
rect 7980 14018 8036 14028
rect 7868 13694 7870 13746
rect 7922 13694 7924 13746
rect 7756 12516 7812 12526
rect 7868 12516 7924 13694
rect 7980 13634 8036 13646
rect 7980 13582 7982 13634
rect 8034 13582 8036 13634
rect 7980 13074 8036 13582
rect 8204 13522 8260 14476
rect 8316 14420 8372 15596
rect 8652 15426 8708 15438
rect 8652 15374 8654 15426
rect 8706 15374 8708 15426
rect 8652 15316 8708 15374
rect 8428 15204 8484 15214
rect 8652 15148 8708 15260
rect 8428 14754 8484 15148
rect 8428 14702 8430 14754
rect 8482 14702 8484 14754
rect 8428 14690 8484 14702
rect 8540 15092 8708 15148
rect 8316 14354 8372 14364
rect 8428 13748 8484 13758
rect 8540 13748 8596 15092
rect 8428 13746 8596 13748
rect 8428 13694 8430 13746
rect 8482 13694 8596 13746
rect 8428 13692 8596 13694
rect 8428 13682 8484 13692
rect 8204 13470 8206 13522
rect 8258 13470 8260 13522
rect 8092 13412 8148 13422
rect 8204 13412 8260 13470
rect 8148 13356 8260 13412
rect 8092 13346 8148 13356
rect 8876 13188 8932 17388
rect 9100 16322 9156 17612
rect 9324 17602 9380 17612
rect 9436 17444 9492 17454
rect 9100 16270 9102 16322
rect 9154 16270 9156 16322
rect 9100 16258 9156 16270
rect 9324 17442 9492 17444
rect 9324 17390 9438 17442
rect 9490 17390 9492 17442
rect 9324 17388 9492 17390
rect 8988 15876 9044 15886
rect 8988 15782 9044 15820
rect 8988 15540 9044 15550
rect 9324 15540 9380 17388
rect 9436 17378 9492 17388
rect 8988 15538 9380 15540
rect 8988 15486 8990 15538
rect 9042 15486 9380 15538
rect 8988 15484 9380 15486
rect 8988 15474 9044 15484
rect 9324 15148 9380 15484
rect 9436 15652 9492 15662
rect 9436 15314 9492 15596
rect 9436 15262 9438 15314
rect 9490 15262 9492 15314
rect 9436 15250 9492 15262
rect 9324 15092 9492 15148
rect 9436 14530 9492 15092
rect 9436 14478 9438 14530
rect 9490 14478 9492 14530
rect 9436 14466 9492 14478
rect 9548 13860 9604 19740
rect 9884 19236 9940 19246
rect 9884 19142 9940 19180
rect 9660 19012 9716 19022
rect 9660 16210 9716 18956
rect 9996 18674 10052 22092
rect 10108 21588 10164 21598
rect 10108 21586 10276 21588
rect 10108 21534 10110 21586
rect 10162 21534 10276 21586
rect 10108 21532 10276 21534
rect 10108 21522 10164 21532
rect 10108 20692 10164 20702
rect 10108 20018 10164 20636
rect 10108 19966 10110 20018
rect 10162 19966 10164 20018
rect 10108 19954 10164 19966
rect 10220 19796 10276 21532
rect 10780 21586 10836 21598
rect 10780 21534 10782 21586
rect 10834 21534 10836 21586
rect 10780 21476 10836 21534
rect 10892 21588 10948 26852
rect 11004 26516 11060 26910
rect 11004 26450 11060 26460
rect 11676 26068 11732 26078
rect 11564 26012 11676 26068
rect 11116 25172 11172 25182
rect 11116 24948 11172 25116
rect 11116 24946 11508 24948
rect 11116 24894 11118 24946
rect 11170 24894 11508 24946
rect 11116 24892 11508 24894
rect 11116 24882 11172 24892
rect 11452 24722 11508 24892
rect 11452 24670 11454 24722
rect 11506 24670 11508 24722
rect 11452 24658 11508 24670
rect 11564 23492 11620 26012
rect 11676 25974 11732 26012
rect 11564 23426 11620 23436
rect 11676 23826 11732 23838
rect 11676 23774 11678 23826
rect 11730 23774 11732 23826
rect 11676 23266 11732 23774
rect 11788 23380 11844 27356
rect 11900 25172 11956 29260
rect 12348 28196 12404 31388
rect 12572 31556 12628 31566
rect 12572 31218 12628 31500
rect 12572 31166 12574 31218
rect 12626 31166 12628 31218
rect 12572 31154 12628 31166
rect 12460 30996 12516 31006
rect 12460 30902 12516 30940
rect 12796 30994 12852 31006
rect 12796 30942 12798 30994
rect 12850 30942 12852 30994
rect 12796 30884 12852 30942
rect 12796 30818 12852 30828
rect 12572 29988 12628 29998
rect 12572 29894 12628 29932
rect 12460 28644 12516 28654
rect 12460 28642 12628 28644
rect 12460 28590 12462 28642
rect 12514 28590 12628 28642
rect 12460 28588 12628 28590
rect 12460 28578 12516 28588
rect 12572 28420 12628 28588
rect 12796 28532 12852 28542
rect 12796 28438 12852 28476
rect 12572 28354 12628 28364
rect 12684 28418 12740 28430
rect 12684 28366 12686 28418
rect 12738 28366 12740 28418
rect 12684 28308 12740 28366
rect 12684 28242 12740 28252
rect 12348 28140 12628 28196
rect 12572 28084 12628 28140
rect 12572 28028 12740 28084
rect 12460 27858 12516 27870
rect 12460 27806 12462 27858
rect 12514 27806 12516 27858
rect 12124 27636 12180 27646
rect 12012 27634 12180 27636
rect 12012 27582 12126 27634
rect 12178 27582 12180 27634
rect 12012 27580 12180 27582
rect 12012 27188 12068 27580
rect 12124 27570 12180 27580
rect 12460 27412 12516 27806
rect 12460 27346 12516 27356
rect 12012 27132 12628 27188
rect 12012 26290 12068 27132
rect 12572 27074 12628 27132
rect 12572 27022 12574 27074
rect 12626 27022 12628 27074
rect 12572 27010 12628 27022
rect 12124 26964 12180 26974
rect 12684 26908 12740 28028
rect 12796 27972 12852 27982
rect 12796 27878 12852 27916
rect 12908 27860 12964 31612
rect 13020 30324 13076 36092
rect 13356 35924 13412 36316
rect 13468 36260 13524 36270
rect 13468 36258 13636 36260
rect 13468 36206 13470 36258
rect 13522 36206 13636 36258
rect 13468 36204 13636 36206
rect 13468 36194 13524 36204
rect 13468 35924 13524 35934
rect 13356 35922 13524 35924
rect 13356 35870 13470 35922
rect 13522 35870 13524 35922
rect 13356 35868 13524 35870
rect 13468 35858 13524 35868
rect 13356 34692 13412 34702
rect 13356 34242 13412 34636
rect 13356 34190 13358 34242
rect 13410 34190 13412 34242
rect 13356 34178 13412 34190
rect 13580 33348 13636 36204
rect 13580 33282 13636 33292
rect 13692 35476 13748 35486
rect 13468 33124 13524 33134
rect 13468 33030 13524 33068
rect 13356 32450 13412 32462
rect 13356 32398 13358 32450
rect 13410 32398 13412 32450
rect 13356 32116 13412 32398
rect 13356 32050 13412 32060
rect 13692 31668 13748 35420
rect 14028 35028 14084 37886
rect 14252 37828 14308 37838
rect 14252 37734 14308 37772
rect 14364 37268 14420 37278
rect 14364 37174 14420 37212
rect 14476 36484 14532 42588
rect 14700 42532 14756 42702
rect 14700 42466 14756 42476
rect 14812 42756 14868 42766
rect 14588 41076 14644 41086
rect 14588 40982 14644 41020
rect 14700 40964 14756 40974
rect 14700 40514 14756 40908
rect 14700 40462 14702 40514
rect 14754 40462 14756 40514
rect 14700 40450 14756 40462
rect 14812 38668 14868 42700
rect 15036 41972 15092 43652
rect 15148 42532 15204 42542
rect 15148 42438 15204 42476
rect 15036 41906 15092 41916
rect 14924 41858 14980 41870
rect 14924 41806 14926 41858
rect 14978 41806 14980 41858
rect 14924 41300 14980 41806
rect 14924 41074 14980 41244
rect 15036 41188 15092 41198
rect 15036 41094 15092 41132
rect 15148 41188 15204 41198
rect 15372 41188 15428 44942
rect 15484 44772 15540 45614
rect 16268 45332 16324 49532
rect 16828 49140 16884 49870
rect 16940 50370 16996 50382
rect 16940 50318 16942 50370
rect 16994 50318 16996 50370
rect 16940 49924 16996 50318
rect 17388 49924 17444 49934
rect 16940 49922 17444 49924
rect 16940 49870 17390 49922
rect 17442 49870 17444 49922
rect 16940 49868 17444 49870
rect 17388 49858 17444 49868
rect 17500 49812 17556 49822
rect 17500 49718 17556 49756
rect 17052 49700 17108 49710
rect 16828 49084 16996 49140
rect 16828 48914 16884 48926
rect 16828 48862 16830 48914
rect 16882 48862 16884 48914
rect 16716 48804 16772 48814
rect 16492 48356 16548 48366
rect 16380 48132 16436 48142
rect 16380 47682 16436 48076
rect 16380 47630 16382 47682
rect 16434 47630 16436 47682
rect 16380 47618 16436 47630
rect 16492 47348 16548 48300
rect 16716 47682 16772 48748
rect 16716 47630 16718 47682
rect 16770 47630 16772 47682
rect 16716 47618 16772 47630
rect 16828 48130 16884 48862
rect 16828 48078 16830 48130
rect 16882 48078 16884 48130
rect 16492 47346 16660 47348
rect 16492 47294 16494 47346
rect 16546 47294 16660 47346
rect 16492 47292 16660 47294
rect 16492 47282 16548 47292
rect 16380 46676 16436 46686
rect 16380 46582 16436 46620
rect 16268 45276 16548 45332
rect 16268 45108 16324 45118
rect 15932 45106 16324 45108
rect 15932 45054 16270 45106
rect 16322 45054 16324 45106
rect 15932 45052 16324 45054
rect 15484 44706 15540 44716
rect 15820 44994 15876 45006
rect 15820 44942 15822 44994
rect 15874 44942 15876 44994
rect 15820 44660 15876 44942
rect 15820 44594 15876 44604
rect 15484 44548 15540 44558
rect 15484 44210 15540 44492
rect 15596 44434 15652 44446
rect 15596 44382 15598 44434
rect 15650 44382 15652 44434
rect 15596 44324 15652 44382
rect 15596 44258 15652 44268
rect 15484 44158 15486 44210
rect 15538 44158 15540 44210
rect 15484 43764 15540 44158
rect 15932 44100 15988 45052
rect 16268 45042 16324 45052
rect 16380 44324 16436 44334
rect 16268 44212 16324 44222
rect 16380 44212 16436 44268
rect 16268 44210 16436 44212
rect 16268 44158 16270 44210
rect 16322 44158 16436 44210
rect 16268 44156 16436 44158
rect 16268 44146 16324 44156
rect 15484 43698 15540 43708
rect 15596 44098 15988 44100
rect 15596 44046 15934 44098
rect 15986 44046 15988 44098
rect 15596 44044 15988 44046
rect 15484 42756 15540 42766
rect 15596 42756 15652 44044
rect 15932 44034 15988 44044
rect 15484 42754 15652 42756
rect 15484 42702 15486 42754
rect 15538 42702 15652 42754
rect 15484 42700 15652 42702
rect 15484 42690 15540 42700
rect 15148 41186 15428 41188
rect 15148 41134 15150 41186
rect 15202 41134 15428 41186
rect 15148 41132 15428 41134
rect 14924 41022 14926 41074
rect 14978 41022 14980 41074
rect 14924 40628 14980 41022
rect 14924 40562 14980 40572
rect 14700 38612 14868 38668
rect 14700 37268 14756 38612
rect 14812 38164 14868 38174
rect 14812 38070 14868 38108
rect 14812 37380 14868 37390
rect 14812 37286 14868 37324
rect 14700 37202 14756 37212
rect 14476 36418 14532 36428
rect 15148 36260 15204 41132
rect 15484 41074 15540 41086
rect 15484 41022 15486 41074
rect 15538 41022 15540 41074
rect 15484 40292 15540 41022
rect 15484 40226 15540 40236
rect 15596 39058 15652 42700
rect 16044 42532 16100 42542
rect 15820 41188 15876 41198
rect 15820 41094 15876 41132
rect 16044 41074 16100 42476
rect 16044 41022 16046 41074
rect 16098 41022 16100 41074
rect 16044 41010 16100 41022
rect 16380 41076 16436 41086
rect 15932 40964 15988 40974
rect 15932 40870 15988 40908
rect 16380 40404 16436 41020
rect 16380 39730 16436 40348
rect 16380 39678 16382 39730
rect 16434 39678 16436 39730
rect 16380 39666 16436 39678
rect 16492 39508 16548 45276
rect 16604 45330 16660 47292
rect 16716 46788 16772 46798
rect 16716 46694 16772 46732
rect 16828 45668 16884 48078
rect 16940 46452 16996 49084
rect 17052 49026 17108 49644
rect 17388 49700 17444 49710
rect 17052 48974 17054 49026
rect 17106 48974 17108 49026
rect 17052 48962 17108 48974
rect 17276 49588 17332 49598
rect 17164 48804 17220 48814
rect 17164 48710 17220 48748
rect 17164 47460 17220 47470
rect 17164 47366 17220 47404
rect 17276 46564 17332 49532
rect 17388 49026 17444 49644
rect 17388 48974 17390 49026
rect 17442 48974 17444 49026
rect 17388 46786 17444 48974
rect 17612 48916 17668 51326
rect 17836 50594 17892 50606
rect 17836 50542 17838 50594
rect 17890 50542 17892 50594
rect 17836 50036 17892 50542
rect 18060 50482 18116 52332
rect 18172 52388 18228 52398
rect 18284 52388 18340 53564
rect 18396 53618 18452 53676
rect 18844 53732 18900 53742
rect 18844 53638 18900 53676
rect 19292 53730 19348 53742
rect 19292 53678 19294 53730
rect 19346 53678 19348 53730
rect 18396 53566 18398 53618
rect 18450 53566 18452 53618
rect 18396 53554 18452 53566
rect 18956 53620 19012 53630
rect 18172 52386 18340 52388
rect 18172 52334 18174 52386
rect 18226 52334 18340 52386
rect 18172 52332 18340 52334
rect 18396 53396 18452 53406
rect 18396 52386 18452 53340
rect 18956 53172 19012 53564
rect 19180 53620 19236 53630
rect 19180 53526 19236 53564
rect 19068 53506 19124 53518
rect 19068 53454 19070 53506
rect 19122 53454 19124 53506
rect 19068 53172 19124 53454
rect 19292 53396 19348 53678
rect 19292 53330 19348 53340
rect 19068 53116 19572 53172
rect 18956 53106 19012 53116
rect 19516 52948 19572 53116
rect 19628 53170 19684 54350
rect 19852 54404 19908 54414
rect 19852 53842 19908 54348
rect 20748 54180 20804 55358
rect 19852 53790 19854 53842
rect 19906 53790 19908 53842
rect 19852 53778 19908 53790
rect 20300 54124 20804 54180
rect 19740 53732 19796 53742
rect 19740 53638 19796 53676
rect 19964 53732 20020 53742
rect 19964 53508 20020 53676
rect 20300 53732 20356 54124
rect 20860 54068 20916 56028
rect 22988 55858 23044 55870
rect 22988 55806 22990 55858
rect 23042 55806 23044 55858
rect 22988 55300 23044 55806
rect 22988 55234 23044 55244
rect 23548 55298 23604 55310
rect 23548 55246 23550 55298
rect 23602 55246 23604 55298
rect 23324 54740 23380 54750
rect 20300 53666 20356 53676
rect 20524 54012 20916 54068
rect 21756 54402 21812 54414
rect 21756 54350 21758 54402
rect 21810 54350 21812 54402
rect 20188 53620 20244 53630
rect 20188 53526 20244 53564
rect 20412 53618 20468 53630
rect 20412 53566 20414 53618
rect 20466 53566 20468 53618
rect 19964 53442 20020 53452
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19628 53118 19630 53170
rect 19682 53118 19684 53170
rect 19628 53106 19684 53118
rect 19740 52948 19796 52958
rect 19516 52946 19796 52948
rect 19516 52894 19742 52946
rect 19794 52894 19796 52946
rect 19516 52892 19796 52894
rect 19740 52882 19796 52892
rect 18620 52836 18676 52846
rect 18620 52742 18676 52780
rect 20412 52612 20468 53566
rect 20412 52546 20468 52556
rect 18396 52334 18398 52386
rect 18450 52334 18452 52386
rect 18172 52322 18228 52332
rect 18396 52322 18452 52334
rect 18956 52276 19012 52286
rect 18508 52274 19012 52276
rect 18508 52222 18958 52274
rect 19010 52222 19012 52274
rect 18508 52220 19012 52222
rect 18172 52164 18228 52174
rect 18228 52108 18340 52164
rect 18172 52098 18228 52108
rect 18060 50430 18062 50482
rect 18114 50430 18116 50482
rect 18060 50418 18116 50430
rect 17836 49970 17892 49980
rect 17948 49810 18004 49822
rect 17948 49758 17950 49810
rect 18002 49758 18004 49810
rect 17724 49588 17780 49598
rect 17724 49494 17780 49532
rect 17500 48860 17668 48916
rect 17500 47460 17556 48860
rect 17836 48356 17892 48366
rect 17836 48262 17892 48300
rect 17836 48130 17892 48142
rect 17836 48078 17838 48130
rect 17890 48078 17892 48130
rect 17612 48020 17668 48030
rect 17612 48018 17780 48020
rect 17612 47966 17614 48018
rect 17666 47966 17780 48018
rect 17612 47964 17780 47966
rect 17612 47954 17668 47964
rect 17612 47460 17668 47470
rect 17500 47404 17612 47460
rect 17612 47394 17668 47404
rect 17612 46900 17668 46910
rect 17724 46900 17780 47964
rect 17836 47570 17892 48078
rect 17836 47518 17838 47570
rect 17890 47518 17892 47570
rect 17836 47506 17892 47518
rect 17612 46898 17780 46900
rect 17612 46846 17614 46898
rect 17666 46846 17780 46898
rect 17612 46844 17780 46846
rect 17948 46900 18004 49758
rect 17612 46834 17668 46844
rect 17948 46834 18004 46844
rect 18060 48356 18116 48366
rect 17388 46734 17390 46786
rect 17442 46734 17444 46786
rect 17388 46722 17444 46734
rect 17612 46674 17668 46686
rect 17612 46622 17614 46674
rect 17666 46622 17668 46674
rect 17612 46564 17668 46622
rect 17948 46676 18004 46686
rect 17948 46582 18004 46620
rect 17276 46508 17668 46564
rect 16940 46396 17444 46452
rect 16828 45602 16884 45612
rect 16604 45278 16606 45330
rect 16658 45278 16660 45330
rect 16604 45266 16660 45278
rect 17276 44772 17332 44782
rect 17276 44098 17332 44716
rect 17276 44046 17278 44098
rect 17330 44046 17332 44098
rect 16828 43426 16884 43438
rect 16828 43374 16830 43426
rect 16882 43374 16884 43426
rect 16828 43316 16884 43374
rect 16828 43250 16884 43260
rect 17276 42868 17332 44046
rect 17388 44100 17444 46396
rect 17612 45892 17668 46508
rect 17612 45826 17668 45836
rect 17948 46116 18004 46126
rect 17500 45108 17556 45118
rect 17500 45014 17556 45052
rect 17612 44324 17668 44334
rect 17612 44322 17780 44324
rect 17612 44270 17614 44322
rect 17666 44270 17780 44322
rect 17612 44268 17780 44270
rect 17612 44258 17668 44268
rect 17724 44100 17780 44268
rect 17948 44100 18004 46060
rect 18060 45778 18116 48300
rect 18284 46116 18340 52108
rect 18508 51940 18564 52220
rect 18956 52210 19012 52220
rect 19180 52164 19236 52174
rect 19740 52164 19796 52174
rect 19180 52070 19236 52108
rect 19628 52108 19740 52164
rect 18844 52052 18900 52062
rect 18396 51884 18564 51940
rect 18620 52050 18900 52052
rect 18620 51998 18846 52050
rect 18898 51998 18900 52050
rect 18620 51996 18900 51998
rect 18396 51490 18452 51884
rect 18396 51438 18398 51490
rect 18450 51438 18452 51490
rect 18396 51426 18452 51438
rect 18620 50706 18676 51996
rect 18844 51986 18900 51996
rect 18620 50654 18622 50706
rect 18674 50654 18676 50706
rect 18620 50642 18676 50654
rect 18732 51828 18788 51838
rect 18732 50594 18788 51772
rect 19516 51716 19572 51726
rect 19404 51268 19460 51278
rect 18732 50542 18734 50594
rect 18786 50542 18788 50594
rect 18732 50530 18788 50542
rect 19068 50596 19124 50606
rect 19068 50502 19124 50540
rect 18508 50482 18564 50494
rect 18508 50430 18510 50482
rect 18562 50430 18564 50482
rect 18396 50036 18452 50046
rect 18396 49942 18452 49980
rect 18508 49812 18564 50430
rect 18508 49746 18564 49756
rect 19404 50370 19460 51212
rect 19404 50318 19406 50370
rect 19458 50318 19460 50370
rect 19068 49700 19124 49710
rect 19404 49700 19460 50318
rect 19516 50036 19572 51660
rect 19628 50484 19684 52108
rect 19740 52098 19796 52108
rect 20412 52164 20468 52174
rect 20412 52070 20468 52108
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 20524 51492 20580 54012
rect 21756 53956 21812 54350
rect 21756 53900 22148 53956
rect 20748 53844 20804 53854
rect 20748 52948 20804 53788
rect 21980 53732 22036 53742
rect 22092 53732 22148 53900
rect 22652 53732 22708 53742
rect 22092 53676 22260 53732
rect 21644 53506 21700 53518
rect 21644 53454 21646 53506
rect 21698 53454 21700 53506
rect 21644 53396 21700 53454
rect 20748 52946 20916 52948
rect 20748 52894 20750 52946
rect 20802 52894 20916 52946
rect 20748 52892 20916 52894
rect 20748 52882 20804 52892
rect 20636 52276 20692 52286
rect 20636 52182 20692 52220
rect 20748 52164 20804 52174
rect 20748 52070 20804 52108
rect 20524 51436 20804 51492
rect 20524 51266 20580 51278
rect 20524 51214 20526 51266
rect 20578 51214 20580 51266
rect 20188 50596 20244 50606
rect 20524 50596 20580 51214
rect 20244 50540 20580 50596
rect 19740 50484 19796 50494
rect 19628 50482 19796 50484
rect 19628 50430 19742 50482
rect 19794 50430 19796 50482
rect 19628 50428 19796 50430
rect 19740 50372 19796 50428
rect 19740 50306 19796 50316
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19516 49980 19796 50036
rect 19516 49812 19572 49822
rect 19516 49718 19572 49756
rect 19740 49810 19796 49980
rect 19740 49758 19742 49810
rect 19794 49758 19796 49810
rect 19740 49746 19796 49758
rect 20076 49810 20132 49822
rect 20076 49758 20078 49810
rect 20130 49758 20132 49810
rect 19068 49698 19460 49700
rect 19068 49646 19070 49698
rect 19122 49646 19460 49698
rect 19068 49644 19460 49646
rect 19628 49700 19684 49710
rect 18284 46050 18340 46060
rect 18620 46900 18676 46910
rect 18060 45726 18062 45778
rect 18114 45726 18116 45778
rect 18060 45714 18116 45726
rect 18284 45780 18340 45790
rect 18284 45778 18564 45780
rect 18284 45726 18286 45778
rect 18338 45726 18564 45778
rect 18284 45724 18564 45726
rect 18284 45714 18340 45724
rect 18172 45666 18228 45678
rect 18172 45614 18174 45666
rect 18226 45614 18228 45666
rect 18172 45218 18228 45614
rect 18172 45166 18174 45218
rect 18226 45166 18228 45218
rect 18172 45154 18228 45166
rect 18508 44434 18564 45724
rect 18508 44382 18510 44434
rect 18562 44382 18564 44434
rect 18508 44370 18564 44382
rect 18620 44322 18676 46844
rect 18620 44270 18622 44322
rect 18674 44270 18676 44322
rect 18620 44258 18676 44270
rect 18396 44212 18452 44222
rect 18396 44118 18452 44156
rect 18956 44210 19012 44222
rect 18956 44158 18958 44210
rect 19010 44158 19012 44210
rect 18060 44100 18116 44110
rect 17388 44044 17668 44100
rect 17724 44098 18116 44100
rect 17724 44046 18062 44098
rect 18114 44046 18116 44098
rect 17724 44044 18116 44046
rect 17500 43652 17556 43662
rect 17500 43558 17556 43596
rect 17276 42812 17556 42868
rect 17388 41970 17444 41982
rect 17388 41918 17390 41970
rect 17442 41918 17444 41970
rect 16940 41860 16996 41870
rect 17388 41860 17444 41918
rect 16940 41858 17444 41860
rect 16940 41806 16942 41858
rect 16994 41806 17444 41858
rect 16940 41804 17444 41806
rect 16604 40964 16660 40974
rect 16604 40870 16660 40908
rect 16940 40516 16996 41804
rect 16940 40450 16996 40460
rect 16828 40292 16884 40302
rect 16828 39620 16884 40236
rect 16828 39554 16884 39564
rect 15596 39006 15598 39058
rect 15650 39006 15652 39058
rect 15260 38052 15316 38062
rect 15260 38050 15428 38052
rect 15260 37998 15262 38050
rect 15314 37998 15428 38050
rect 15260 37996 15428 37998
rect 15260 37986 15316 37996
rect 15372 37490 15428 37996
rect 15484 37940 15540 37950
rect 15484 37846 15540 37884
rect 15372 37438 15374 37490
rect 15426 37438 15428 37490
rect 15372 37426 15428 37438
rect 15596 37380 15652 39006
rect 16380 39452 16548 39508
rect 15932 38948 15988 38958
rect 16044 38948 16100 38958
rect 15932 38946 16044 38948
rect 15932 38894 15934 38946
rect 15986 38894 16044 38946
rect 15932 38892 16044 38894
rect 15932 38882 15988 38892
rect 15820 38052 15876 38062
rect 15820 37958 15876 37996
rect 15932 37380 15988 37390
rect 15596 37378 15988 37380
rect 15596 37326 15934 37378
rect 15986 37326 15988 37378
rect 15596 37324 15988 37326
rect 15932 37314 15988 37324
rect 15708 37044 15764 37054
rect 15708 36950 15764 36988
rect 16044 36708 16100 38892
rect 15036 36204 15204 36260
rect 15596 36652 16100 36708
rect 16156 37268 16212 37278
rect 14588 35924 14644 35934
rect 14364 35812 14420 35822
rect 14140 35700 14196 35710
rect 14140 35606 14196 35644
rect 14364 35698 14420 35756
rect 14364 35646 14366 35698
rect 14418 35646 14420 35698
rect 14364 35634 14420 35646
rect 14588 35698 14644 35868
rect 15036 35812 15092 36204
rect 15596 35924 15652 36652
rect 16044 36260 16100 36270
rect 16156 36260 16212 37212
rect 16100 36204 16212 36260
rect 16380 36370 16436 39452
rect 16604 37940 16660 37950
rect 16604 37846 16660 37884
rect 16492 37378 16548 37390
rect 16492 37326 16494 37378
rect 16546 37326 16548 37378
rect 16492 37044 16548 37326
rect 17500 37380 17556 42812
rect 17612 38668 17668 44044
rect 17836 43538 17892 43550
rect 17836 43486 17838 43538
rect 17890 43486 17892 43538
rect 17836 43316 17892 43486
rect 17724 43204 17780 43214
rect 17724 38948 17780 43148
rect 17836 42980 17892 43260
rect 17948 42980 18004 42990
rect 17836 42978 18004 42980
rect 17836 42926 17950 42978
rect 18002 42926 18004 42978
rect 17836 42924 18004 42926
rect 17948 42914 18004 42924
rect 17836 42644 17892 42654
rect 18060 42644 18116 44044
rect 18956 43652 19012 44158
rect 18956 43586 19012 43596
rect 19068 43204 19124 49644
rect 19628 49606 19684 49644
rect 20076 48916 20132 49758
rect 20076 48850 20132 48860
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19516 48244 19572 48254
rect 19516 47460 19572 48188
rect 20188 47684 20244 50540
rect 20748 50428 20804 51436
rect 20860 50596 20916 52892
rect 21420 52834 21476 52846
rect 21420 52782 21422 52834
rect 21474 52782 21476 52834
rect 21420 52276 21476 52782
rect 21644 52836 21700 53340
rect 21980 52836 22036 53676
rect 22092 53508 22148 53518
rect 22092 53060 22148 53452
rect 22092 52994 22148 53004
rect 22204 53172 22260 53676
rect 22652 53618 22708 53676
rect 23212 53730 23268 53742
rect 23212 53678 23214 53730
rect 23266 53678 23268 53730
rect 22652 53566 22654 53618
rect 22706 53566 22708 53618
rect 22652 53554 22708 53566
rect 22988 53620 23044 53630
rect 22316 53506 22372 53518
rect 22316 53454 22318 53506
rect 22370 53454 22372 53506
rect 22316 53396 22372 53454
rect 22316 53330 22372 53340
rect 22988 53506 23044 53564
rect 22988 53454 22990 53506
rect 23042 53454 23044 53506
rect 21980 52780 22148 52836
rect 21644 52770 21700 52780
rect 21420 52210 21476 52220
rect 21868 52500 21924 52510
rect 21868 52050 21924 52444
rect 21980 52164 22036 52174
rect 21980 52070 22036 52108
rect 22092 52162 22148 52780
rect 22092 52110 22094 52162
rect 22146 52110 22148 52162
rect 22092 52098 22148 52110
rect 21868 51998 21870 52050
rect 21922 51998 21924 52050
rect 21868 51378 21924 51998
rect 21868 51326 21870 51378
rect 21922 51326 21924 51378
rect 21868 51314 21924 51326
rect 22204 51378 22260 53116
rect 22988 53060 23044 53454
rect 23212 53508 23268 53678
rect 23212 53442 23268 53452
rect 22988 52994 23044 53004
rect 22428 52164 22484 52174
rect 22428 52070 22484 52108
rect 23324 51604 23380 54684
rect 23548 53732 23604 55246
rect 23660 54738 23716 57372
rect 23996 56642 24052 56654
rect 23996 56590 23998 56642
rect 24050 56590 24052 56642
rect 23996 56082 24052 56590
rect 23996 56030 23998 56082
rect 24050 56030 24052 56082
rect 23996 56018 24052 56030
rect 25004 56642 25060 56654
rect 25004 56590 25006 56642
rect 25058 56590 25060 56642
rect 24668 55970 24724 55982
rect 24668 55918 24670 55970
rect 24722 55918 24724 55970
rect 24556 55860 24612 55870
rect 24220 55858 24612 55860
rect 24220 55806 24558 55858
rect 24610 55806 24612 55858
rect 24220 55804 24612 55806
rect 24220 55410 24276 55804
rect 24556 55794 24612 55804
rect 24668 55468 24724 55918
rect 24220 55358 24222 55410
rect 24274 55358 24276 55410
rect 24220 55346 24276 55358
rect 24332 55412 24724 55468
rect 23660 54686 23662 54738
rect 23714 54686 23716 54738
rect 23660 54674 23716 54686
rect 23772 53732 23828 53742
rect 23548 53730 23828 53732
rect 23548 53678 23774 53730
rect 23826 53678 23828 53730
rect 23548 53676 23828 53678
rect 23548 52834 23604 52846
rect 23548 52782 23550 52834
rect 23602 52782 23604 52834
rect 23548 52164 23604 52782
rect 23548 52098 23604 52108
rect 23324 51538 23380 51548
rect 23660 51492 23716 51502
rect 23660 51398 23716 51436
rect 22204 51326 22206 51378
rect 22258 51326 22260 51378
rect 22204 51314 22260 51326
rect 22540 51378 22596 51390
rect 22540 51326 22542 51378
rect 22594 51326 22596 51378
rect 22092 51266 22148 51278
rect 22092 51214 22094 51266
rect 22146 51214 22148 51266
rect 22092 50708 22148 51214
rect 21980 50652 22148 50708
rect 21420 50596 21476 50606
rect 20860 50594 21476 50596
rect 20860 50542 21422 50594
rect 21474 50542 21476 50594
rect 20860 50540 21476 50542
rect 21420 50484 21476 50540
rect 21420 50428 21924 50484
rect 20636 50372 20692 50382
rect 20748 50372 20916 50428
rect 20636 50036 20692 50316
rect 20636 49942 20692 49980
rect 20412 49700 20468 49710
rect 20412 49606 20468 49644
rect 20524 49698 20580 49710
rect 20524 49646 20526 49698
rect 20578 49646 20580 49698
rect 20300 48356 20356 48366
rect 20524 48356 20580 49646
rect 20300 48354 20580 48356
rect 20300 48302 20302 48354
rect 20354 48302 20580 48354
rect 20300 48300 20580 48302
rect 20300 48290 20356 48300
rect 20188 47628 20580 47684
rect 19964 47572 20020 47582
rect 19964 47570 20356 47572
rect 19964 47518 19966 47570
rect 20018 47518 20356 47570
rect 19964 47516 20356 47518
rect 19964 47506 20020 47516
rect 19516 47394 19572 47404
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20188 46900 20244 47516
rect 20300 47458 20356 47516
rect 20300 47406 20302 47458
rect 20354 47406 20356 47458
rect 20300 47394 20356 47406
rect 20076 46844 20244 46900
rect 19852 46674 19908 46686
rect 19852 46622 19854 46674
rect 19906 46622 19908 46674
rect 19628 46116 19684 46126
rect 19628 46002 19684 46060
rect 19628 45950 19630 46002
rect 19682 45950 19684 46002
rect 19628 45938 19684 45950
rect 19852 46004 19908 46622
rect 20076 46674 20132 46844
rect 20076 46622 20078 46674
rect 20130 46622 20132 46674
rect 20076 46610 20132 46622
rect 20188 46676 20244 46686
rect 19852 45938 19908 45948
rect 20188 46114 20244 46620
rect 20524 46676 20580 47628
rect 20524 46582 20580 46620
rect 20636 47234 20692 47246
rect 20636 47182 20638 47234
rect 20690 47182 20692 47234
rect 20636 46564 20692 47182
rect 20636 46498 20692 46508
rect 20188 46062 20190 46114
rect 20242 46062 20244 46114
rect 19964 45890 20020 45902
rect 19964 45838 19966 45890
rect 20018 45838 20020 45890
rect 19964 45668 20020 45838
rect 19964 45602 20020 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19404 44212 19460 44222
rect 19404 44118 19460 44156
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19964 43764 20020 43774
rect 19068 43138 19124 43148
rect 19628 43650 19684 43662
rect 19628 43598 19630 43650
rect 19682 43598 19684 43650
rect 19628 43316 19684 43598
rect 19852 43652 19908 43662
rect 19852 43558 19908 43596
rect 19964 43650 20020 43708
rect 19964 43598 19966 43650
rect 20018 43598 20020 43650
rect 19964 43586 20020 43598
rect 20076 43652 20132 43662
rect 20188 43652 20244 46062
rect 20300 46450 20356 46462
rect 20300 46398 20302 46450
rect 20354 46398 20356 46450
rect 20300 45668 20356 46398
rect 20524 46004 20580 46014
rect 20412 45892 20468 45902
rect 20412 45798 20468 45836
rect 20524 45892 20580 45948
rect 20748 46004 20804 46014
rect 20748 45910 20804 45948
rect 20524 45890 20692 45892
rect 20524 45838 20526 45890
rect 20578 45838 20692 45890
rect 20524 45836 20692 45838
rect 20524 45826 20580 45836
rect 20300 45602 20356 45612
rect 20636 45332 20692 45836
rect 20300 45330 20692 45332
rect 20300 45278 20638 45330
rect 20690 45278 20692 45330
rect 20300 45276 20692 45278
rect 20300 44994 20356 45276
rect 20636 45266 20692 45276
rect 20300 44942 20302 44994
rect 20354 44942 20356 44994
rect 20300 44930 20356 44942
rect 20748 45108 20804 45118
rect 20748 44434 20804 45052
rect 20748 44382 20750 44434
rect 20802 44382 20804 44434
rect 20748 44370 20804 44382
rect 20860 44212 20916 50372
rect 21756 50260 21812 50270
rect 21644 50204 21756 50260
rect 21308 49812 21364 49822
rect 21308 47346 21364 49756
rect 21644 49698 21700 50204
rect 21756 50194 21812 50204
rect 21756 50036 21812 50046
rect 21756 49942 21812 49980
rect 21644 49646 21646 49698
rect 21698 49646 21700 49698
rect 21644 49634 21700 49646
rect 21308 47294 21310 47346
rect 21362 47294 21364 47346
rect 21308 47282 21364 47294
rect 21868 48244 21924 50428
rect 21980 49922 22036 50652
rect 22092 50484 22148 50494
rect 22092 50390 22148 50428
rect 22540 50428 22596 51326
rect 23436 51378 23492 51390
rect 23436 51326 23438 51378
rect 23490 51326 23492 51378
rect 22988 51268 23044 51278
rect 22988 51174 23044 51212
rect 23436 51268 23492 51326
rect 23436 51202 23492 51212
rect 23772 50596 23828 53676
rect 24108 53620 24164 53630
rect 24108 53170 24164 53564
rect 24108 53118 24110 53170
rect 24162 53118 24164 53170
rect 24108 53106 24164 53118
rect 24332 53170 24388 55412
rect 24668 54516 24724 54526
rect 24668 54514 24836 54516
rect 24668 54462 24670 54514
rect 24722 54462 24836 54514
rect 24668 54460 24836 54462
rect 24668 54450 24724 54460
rect 24444 53620 24500 53630
rect 24444 53618 24612 53620
rect 24444 53566 24446 53618
rect 24498 53566 24612 53618
rect 24444 53564 24612 53566
rect 24444 53554 24500 53564
rect 24332 53118 24334 53170
rect 24386 53118 24388 53170
rect 24332 53106 24388 53118
rect 24444 53060 24500 53070
rect 24444 52966 24500 53004
rect 24220 52946 24276 52958
rect 24220 52894 24222 52946
rect 24274 52894 24276 52946
rect 24220 52612 24276 52894
rect 24220 52546 24276 52556
rect 24220 52388 24276 52398
rect 24220 52274 24276 52332
rect 24556 52386 24612 53564
rect 24668 52946 24724 52958
rect 24668 52894 24670 52946
rect 24722 52894 24724 52946
rect 24668 52724 24724 52894
rect 24668 52658 24724 52668
rect 24556 52334 24558 52386
rect 24610 52334 24612 52386
rect 24556 52322 24612 52334
rect 24220 52222 24222 52274
rect 24274 52222 24276 52274
rect 24220 52210 24276 52222
rect 24668 52276 24724 52286
rect 24668 52182 24724 52220
rect 23772 50530 23828 50540
rect 24220 50706 24276 50718
rect 24220 50654 24222 50706
rect 24274 50654 24276 50706
rect 24220 50428 24276 50654
rect 22540 50372 23268 50428
rect 23212 50036 23268 50372
rect 23548 50372 24276 50428
rect 24556 50596 24612 50606
rect 23212 50034 23380 50036
rect 23212 49982 23214 50034
rect 23266 49982 23380 50034
rect 23212 49980 23380 49982
rect 23212 49970 23268 49980
rect 21980 49870 21982 49922
rect 22034 49870 22036 49922
rect 21980 49858 22036 49870
rect 22764 49026 22820 49038
rect 22764 48974 22766 49026
rect 22818 48974 22820 49026
rect 21644 47234 21700 47246
rect 21644 47182 21646 47234
rect 21698 47182 21700 47234
rect 21084 46900 21140 46910
rect 21084 46786 21140 46844
rect 21084 46734 21086 46786
rect 21138 46734 21140 46786
rect 21084 46722 21140 46734
rect 21420 45666 21476 45678
rect 21420 45614 21422 45666
rect 21474 45614 21476 45666
rect 21420 45556 21476 45614
rect 21420 45332 21476 45500
rect 21644 45444 21700 47182
rect 21868 46562 21924 48188
rect 22204 48916 22260 48926
rect 21868 46510 21870 46562
rect 21922 46510 21924 46562
rect 21868 46498 21924 46510
rect 22092 46676 22148 46686
rect 21868 45892 21924 45902
rect 21868 45798 21924 45836
rect 22092 45890 22148 46620
rect 22092 45838 22094 45890
rect 22146 45838 22148 45890
rect 22092 45826 22148 45838
rect 21644 45378 21700 45388
rect 21868 45668 21924 45678
rect 21420 45330 21588 45332
rect 21420 45278 21422 45330
rect 21474 45278 21588 45330
rect 21420 45276 21588 45278
rect 21420 45266 21476 45276
rect 20636 44156 20916 44212
rect 20972 45218 21028 45230
rect 20972 45166 20974 45218
rect 21026 45166 21028 45218
rect 20412 44100 20468 44110
rect 20076 43650 20244 43652
rect 20076 43598 20078 43650
rect 20130 43598 20244 43650
rect 20076 43596 20244 43598
rect 20076 43586 20132 43596
rect 20188 43540 20244 43596
rect 20188 43474 20244 43484
rect 20300 44098 20468 44100
rect 20300 44046 20414 44098
rect 20466 44046 20468 44098
rect 20300 44044 20468 44046
rect 20300 43316 20356 44044
rect 20412 44034 20468 44044
rect 20524 43652 20580 43662
rect 19628 43260 20356 43316
rect 20412 43596 20524 43652
rect 18172 42980 18228 42990
rect 18172 42886 18228 42924
rect 18284 42868 18340 42878
rect 18284 42774 18340 42812
rect 17836 42550 17892 42588
rect 17948 42588 18116 42644
rect 19068 42642 19124 42654
rect 19068 42590 19070 42642
rect 19122 42590 19124 42642
rect 17724 38882 17780 38892
rect 17612 38612 17892 38668
rect 17500 37324 17668 37380
rect 16492 36978 16548 36988
rect 16940 37156 16996 37166
rect 16716 36484 16772 36494
rect 16716 36390 16772 36428
rect 16380 36318 16382 36370
rect 16434 36318 16436 36370
rect 16044 36166 16100 36204
rect 15596 35830 15652 35868
rect 15036 35746 15092 35756
rect 14588 35646 14590 35698
rect 14642 35646 14644 35698
rect 14252 35586 14308 35598
rect 14252 35534 14254 35586
rect 14306 35534 14308 35586
rect 14252 35364 14308 35534
rect 14252 35298 14308 35308
rect 14028 34972 14532 35028
rect 14252 34802 14308 34814
rect 14252 34750 14254 34802
rect 14306 34750 14308 34802
rect 14140 34692 14196 34702
rect 14140 34598 14196 34636
rect 14252 33460 14308 34750
rect 14252 33394 14308 33404
rect 14028 33348 14084 33358
rect 14084 33292 14196 33348
rect 14028 33282 14084 33292
rect 14140 33236 14196 33292
rect 14252 33236 14308 33246
rect 14140 33234 14308 33236
rect 14140 33182 14254 33234
rect 14306 33182 14308 33234
rect 14140 33180 14308 33182
rect 13804 33122 13860 33134
rect 13804 33070 13806 33122
rect 13858 33070 13860 33122
rect 13804 32116 13860 33070
rect 14252 33012 14308 33180
rect 14252 32946 14308 32956
rect 14364 33124 14420 33134
rect 14364 32786 14420 33068
rect 14476 32900 14532 34972
rect 14476 32834 14532 32844
rect 14364 32734 14366 32786
rect 14418 32734 14420 32786
rect 14364 32722 14420 32734
rect 14588 32788 14644 35646
rect 15148 35588 15204 35598
rect 16156 35588 16212 35598
rect 15204 35532 15316 35588
rect 15148 35494 15204 35532
rect 15148 34914 15204 34926
rect 15148 34862 15150 34914
rect 15202 34862 15204 34914
rect 14700 34692 14756 34702
rect 15148 34692 15204 34862
rect 14700 34690 15204 34692
rect 14700 34638 14702 34690
rect 14754 34638 15204 34690
rect 14700 34636 15204 34638
rect 14700 34626 14756 34636
rect 15148 34356 15204 34636
rect 15148 34290 15204 34300
rect 14924 33234 14980 33246
rect 14924 33182 14926 33234
rect 14978 33182 14980 33234
rect 14924 33124 14980 33182
rect 15148 33124 15204 33134
rect 14980 33068 15092 33124
rect 14924 33058 14980 33068
rect 14588 32722 14644 32732
rect 14700 32564 14756 32574
rect 14364 32562 14756 32564
rect 14364 32510 14702 32562
rect 14754 32510 14756 32562
rect 14364 32508 14756 32510
rect 13916 32450 13972 32462
rect 13916 32398 13918 32450
rect 13970 32398 13972 32450
rect 13916 32340 13972 32398
rect 13916 32274 13972 32284
rect 14140 32340 14196 32350
rect 14140 32246 14196 32284
rect 14364 32340 14420 32508
rect 14700 32498 14756 32508
rect 15036 32562 15092 33068
rect 15148 33030 15204 33068
rect 15036 32510 15038 32562
rect 15090 32510 15092 32562
rect 15036 32498 15092 32510
rect 15148 32900 15204 32910
rect 14924 32450 14980 32462
rect 14924 32398 14926 32450
rect 14978 32398 14980 32450
rect 13804 32050 13860 32060
rect 14140 32116 14196 32126
rect 14140 31778 14196 32060
rect 14140 31726 14142 31778
rect 14194 31726 14196 31778
rect 14140 31714 14196 31726
rect 14364 31780 14420 32284
rect 14476 32340 14532 32350
rect 14476 32338 14868 32340
rect 14476 32286 14478 32338
rect 14530 32286 14868 32338
rect 14476 32284 14868 32286
rect 14476 32274 14532 32284
rect 14588 31780 14644 31790
rect 14364 31778 14644 31780
rect 14364 31726 14590 31778
rect 14642 31726 14644 31778
rect 14364 31724 14644 31726
rect 13692 31612 14084 31668
rect 14028 31556 14084 31612
rect 14028 31500 14308 31556
rect 13916 31444 13972 31454
rect 13244 30884 13300 30894
rect 13244 30790 13300 30828
rect 13020 30258 13076 30268
rect 13804 30100 13860 30110
rect 13804 30006 13860 30044
rect 13468 29988 13524 29998
rect 13020 29986 13524 29988
rect 13020 29934 13470 29986
rect 13522 29934 13524 29986
rect 13020 29932 13524 29934
rect 13020 29538 13076 29932
rect 13468 29922 13524 29932
rect 13020 29486 13022 29538
rect 13074 29486 13076 29538
rect 13020 29474 13076 29486
rect 13916 28754 13972 31388
rect 13916 28702 13918 28754
rect 13970 28702 13972 28754
rect 13916 28690 13972 28702
rect 13356 28644 13412 28654
rect 13020 28642 13412 28644
rect 13020 28590 13358 28642
rect 13410 28590 13412 28642
rect 13020 28588 13412 28590
rect 13020 28082 13076 28588
rect 13356 28578 13412 28588
rect 13020 28030 13022 28082
rect 13074 28030 13076 28082
rect 13020 28018 13076 28030
rect 13580 28532 13636 28542
rect 13580 28082 13636 28476
rect 13804 28418 13860 28430
rect 13804 28366 13806 28418
rect 13858 28366 13860 28418
rect 13804 28196 13860 28366
rect 14028 28420 14084 28430
rect 14028 28326 14084 28364
rect 13804 28140 14196 28196
rect 13580 28030 13582 28082
rect 13634 28030 13636 28082
rect 13580 28018 13636 28030
rect 13244 27970 13300 27982
rect 13804 27972 13860 27982
rect 13244 27918 13246 27970
rect 13298 27918 13300 27970
rect 13132 27860 13188 27870
rect 13244 27860 13300 27918
rect 13692 27970 13860 27972
rect 13692 27918 13806 27970
rect 13858 27918 13860 27970
rect 13692 27916 13860 27918
rect 12908 27804 13076 27860
rect 12124 26852 12292 26908
rect 12012 26238 12014 26290
rect 12066 26238 12068 26290
rect 12012 26226 12068 26238
rect 12236 26290 12292 26852
rect 12236 26238 12238 26290
rect 12290 26238 12292 26290
rect 12236 26226 12292 26238
rect 12460 26852 12740 26908
rect 12908 27076 12964 27086
rect 12908 26962 12964 27020
rect 12908 26910 12910 26962
rect 12962 26910 12964 26962
rect 12908 26898 12964 26910
rect 11956 25116 12404 25172
rect 11900 25106 11956 25116
rect 12236 24612 12292 24622
rect 12236 24518 12292 24556
rect 12348 23938 12404 25116
rect 12460 24388 12516 26852
rect 12460 24322 12516 24332
rect 12908 24052 12964 24062
rect 12908 23958 12964 23996
rect 12348 23886 12350 23938
rect 12402 23886 12404 23938
rect 12348 23874 12404 23886
rect 12796 23714 12852 23726
rect 12796 23662 12798 23714
rect 12850 23662 12852 23714
rect 12572 23604 12628 23614
rect 11788 23314 11844 23324
rect 12012 23380 12068 23390
rect 11676 23214 11678 23266
rect 11730 23214 11732 23266
rect 11676 23202 11732 23214
rect 11900 23268 11956 23278
rect 12012 23268 12068 23324
rect 12348 23268 12404 23278
rect 11900 23266 12068 23268
rect 11900 23214 11902 23266
rect 11954 23214 12068 23266
rect 11900 23212 12068 23214
rect 12124 23266 12404 23268
rect 12124 23214 12350 23266
rect 12402 23214 12404 23266
rect 12124 23212 12404 23214
rect 11900 23202 11956 23212
rect 11340 23154 11396 23166
rect 11564 23156 11620 23166
rect 11340 23102 11342 23154
rect 11394 23102 11396 23154
rect 11340 22484 11396 23102
rect 11452 23154 11620 23156
rect 11452 23102 11566 23154
rect 11618 23102 11620 23154
rect 11452 23100 11620 23102
rect 11452 22594 11508 23100
rect 11564 23090 11620 23100
rect 11788 23154 11844 23166
rect 11788 23102 11790 23154
rect 11842 23102 11844 23154
rect 11788 23044 11844 23102
rect 11900 23044 11956 23054
rect 11788 22988 11900 23044
rect 11900 22978 11956 22988
rect 11564 22820 11620 22830
rect 11620 22764 11732 22820
rect 11564 22754 11620 22764
rect 11452 22542 11454 22594
rect 11506 22542 11508 22594
rect 11452 22530 11508 22542
rect 11564 22596 11620 22606
rect 11340 22418 11396 22428
rect 11340 22258 11396 22270
rect 11340 22206 11342 22258
rect 11394 22206 11396 22258
rect 11340 21700 11396 22206
rect 11452 22148 11508 22158
rect 11564 22148 11620 22540
rect 11452 22146 11620 22148
rect 11452 22094 11454 22146
rect 11506 22094 11620 22146
rect 11452 22092 11620 22094
rect 11452 22082 11508 22092
rect 11452 21700 11508 21710
rect 11340 21698 11508 21700
rect 11340 21646 11454 21698
rect 11506 21646 11508 21698
rect 11340 21644 11508 21646
rect 11452 21634 11508 21644
rect 10892 21532 11172 21588
rect 10836 21420 10948 21476
rect 10780 21410 10836 21420
rect 10892 20804 10948 21420
rect 10668 20802 10948 20804
rect 10668 20750 10894 20802
rect 10946 20750 10948 20802
rect 10668 20748 10948 20750
rect 10220 19730 10276 19740
rect 10332 20578 10388 20590
rect 10332 20526 10334 20578
rect 10386 20526 10388 20578
rect 9996 18622 9998 18674
rect 10050 18622 10052 18674
rect 9884 17444 9940 17454
rect 9660 16158 9662 16210
rect 9714 16158 9716 16210
rect 9660 16146 9716 16158
rect 9772 17442 9940 17444
rect 9772 17390 9886 17442
rect 9938 17390 9940 17442
rect 9772 17388 9940 17390
rect 9772 15988 9828 17388
rect 9884 17378 9940 17388
rect 9884 16994 9940 17006
rect 9884 16942 9886 16994
rect 9938 16942 9940 16994
rect 9884 16548 9940 16942
rect 9996 16884 10052 18622
rect 10220 19010 10276 19022
rect 10220 18958 10222 19010
rect 10274 18958 10276 19010
rect 10220 18676 10276 18958
rect 10332 18788 10388 20526
rect 10556 20132 10612 20142
rect 10556 19458 10612 20076
rect 10556 19406 10558 19458
rect 10610 19406 10612 19458
rect 10556 19394 10612 19406
rect 10668 19346 10724 20748
rect 10892 20738 10948 20748
rect 10668 19294 10670 19346
rect 10722 19294 10724 19346
rect 10668 19282 10724 19294
rect 11004 20018 11060 20030
rect 11004 19966 11006 20018
rect 11058 19966 11060 20018
rect 10332 18722 10388 18732
rect 10220 18610 10276 18620
rect 11004 18676 11060 19966
rect 11116 20020 11172 21532
rect 11228 21586 11284 21598
rect 11228 21534 11230 21586
rect 11282 21534 11284 21586
rect 11228 20242 11284 21534
rect 11228 20190 11230 20242
rect 11282 20190 11284 20242
rect 11228 20178 11284 20190
rect 11116 19964 11284 20020
rect 11116 19012 11172 19022
rect 11116 18918 11172 18956
rect 11004 18610 11060 18620
rect 10332 18562 10388 18574
rect 10332 18510 10334 18562
rect 10386 18510 10388 18562
rect 10332 18228 10388 18510
rect 10332 18162 10388 18172
rect 11228 17780 11284 19964
rect 11340 19796 11396 19806
rect 11452 19796 11508 19806
rect 11340 19794 11452 19796
rect 11340 19742 11342 19794
rect 11394 19742 11452 19794
rect 11340 19740 11452 19742
rect 11340 19730 11396 19740
rect 11340 18452 11396 18462
rect 11340 18358 11396 18396
rect 11340 17780 11396 17790
rect 11228 17778 11396 17780
rect 11228 17726 11342 17778
rect 11394 17726 11396 17778
rect 11228 17724 11396 17726
rect 10780 17556 10836 17566
rect 10668 17554 10948 17556
rect 10668 17502 10782 17554
rect 10834 17502 10948 17554
rect 10668 17500 10948 17502
rect 10220 17442 10276 17454
rect 10220 17390 10222 17442
rect 10274 17390 10276 17442
rect 10220 17108 10276 17390
rect 10220 17042 10276 17052
rect 10108 16884 10164 16894
rect 9996 16882 10164 16884
rect 9996 16830 10110 16882
rect 10162 16830 10164 16882
rect 9996 16828 10164 16830
rect 10108 16818 10164 16828
rect 9884 16482 9940 16492
rect 9660 15932 9828 15988
rect 9660 15652 9716 15932
rect 9884 15652 9940 15662
rect 9660 15586 9716 15596
rect 9772 15596 9884 15652
rect 9772 14754 9828 15596
rect 9884 15586 9940 15596
rect 10444 15540 10500 15550
rect 10444 15446 10500 15484
rect 9884 15316 9940 15326
rect 9884 15222 9940 15260
rect 10108 15314 10164 15326
rect 10108 15262 10110 15314
rect 10162 15262 10164 15314
rect 9772 14702 9774 14754
rect 9826 14702 9828 14754
rect 9772 14690 9828 14702
rect 9996 15202 10052 15214
rect 9996 15150 9998 15202
rect 10050 15150 10052 15202
rect 7980 13022 7982 13074
rect 8034 13022 8036 13074
rect 7980 13010 8036 13022
rect 8652 13132 8932 13188
rect 9436 13804 9604 13860
rect 9772 14530 9828 14542
rect 9772 14478 9774 14530
rect 9826 14478 9828 14530
rect 7812 12460 7924 12516
rect 8428 12850 8484 12862
rect 8428 12798 8430 12850
rect 8482 12798 8484 12850
rect 7756 12450 7812 12460
rect 8428 12290 8484 12798
rect 8428 12238 8430 12290
rect 8482 12238 8484 12290
rect 8428 12226 8484 12238
rect 7644 11554 7700 11564
rect 8540 12066 8596 12078
rect 8540 12014 8542 12066
rect 8594 12014 8596 12066
rect 7868 10836 7924 10846
rect 7308 10742 7364 10780
rect 7756 10780 7868 10836
rect 6748 10670 6750 10722
rect 6802 10670 6804 10722
rect 6748 10658 6804 10670
rect 6188 10610 6244 10622
rect 6188 10558 6190 10610
rect 6242 10558 6244 10610
rect 6188 10500 6244 10558
rect 6524 10612 6580 10622
rect 6524 10518 6580 10556
rect 7084 10612 7140 10622
rect 6188 10434 6244 10444
rect 6300 10498 6356 10510
rect 6300 10446 6302 10498
rect 6354 10446 6356 10498
rect 5964 9828 6020 9838
rect 5852 9826 6020 9828
rect 5852 9774 5966 9826
rect 6018 9774 6020 9826
rect 5852 9772 6020 9774
rect 5964 9268 6020 9772
rect 6188 9828 6244 9838
rect 6300 9828 6356 10446
rect 7084 10050 7140 10556
rect 7084 9998 7086 10050
rect 7138 9998 7140 10050
rect 7084 9986 7140 9998
rect 6188 9826 6356 9828
rect 6188 9774 6190 9826
rect 6242 9774 6356 9826
rect 6188 9772 6356 9774
rect 7532 9826 7588 9838
rect 7532 9774 7534 9826
rect 7586 9774 7588 9826
rect 6188 9762 6244 9772
rect 6076 9716 6132 9726
rect 6076 9622 6132 9660
rect 6748 9604 6804 9614
rect 5964 9202 6020 9212
rect 6300 9602 6804 9604
rect 6300 9550 6750 9602
rect 6802 9550 6804 9602
rect 6300 9548 6804 9550
rect 4620 9042 5124 9044
rect 4620 8990 4622 9042
rect 4674 8990 5070 9042
rect 5122 8990 5124 9042
rect 4620 8988 5124 8990
rect 4620 8978 4676 8988
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 5068 8484 5124 8988
rect 5740 8932 5796 8942
rect 5740 8930 6020 8932
rect 5740 8878 5742 8930
rect 5794 8878 6020 8930
rect 5740 8876 6020 8878
rect 5740 8866 5796 8876
rect 5068 8418 5124 8428
rect 5964 8146 6020 8876
rect 6300 8258 6356 9548
rect 6748 9538 6804 9548
rect 7532 9380 7588 9774
rect 7756 9714 7812 10780
rect 7868 10770 7924 10780
rect 8540 10836 8596 12014
rect 8652 11956 8708 13132
rect 9436 13076 9492 13804
rect 9772 13748 9828 14478
rect 9996 14420 10052 15150
rect 10108 15204 10164 15262
rect 10668 15316 10724 17500
rect 10780 17490 10836 17500
rect 10892 17444 10948 17500
rect 10892 17378 10948 17388
rect 11340 17332 11396 17724
rect 11340 17266 11396 17276
rect 11340 17108 11396 17118
rect 11340 17014 11396 17052
rect 11452 16884 11508 19740
rect 11004 16828 11508 16884
rect 10780 16324 10836 16334
rect 11004 16324 11060 16828
rect 10780 16322 11060 16324
rect 10780 16270 10782 16322
rect 10834 16270 11060 16322
rect 10780 16268 11060 16270
rect 10780 16258 10836 16268
rect 11116 16210 11172 16222
rect 11116 16158 11118 16210
rect 11170 16158 11172 16210
rect 11116 15988 11172 16158
rect 11452 15988 11508 15998
rect 11116 15986 11508 15988
rect 11116 15934 11454 15986
rect 11506 15934 11508 15986
rect 11116 15932 11508 15934
rect 11004 15874 11060 15886
rect 11004 15822 11006 15874
rect 11058 15822 11060 15874
rect 11004 15652 11060 15822
rect 11004 15586 11060 15596
rect 10668 15314 10948 15316
rect 10668 15262 10670 15314
rect 10722 15262 10948 15314
rect 10668 15260 10948 15262
rect 10668 15250 10724 15260
rect 10108 14642 10164 15148
rect 10108 14590 10110 14642
rect 10162 14590 10164 14642
rect 10108 14578 10164 14590
rect 10444 14532 10500 14542
rect 9996 14364 10164 14420
rect 9996 13748 10052 13758
rect 9772 13692 9996 13748
rect 9996 13654 10052 13692
rect 9548 13636 9604 13646
rect 10108 13636 10164 14364
rect 10332 13636 10388 13646
rect 9548 13634 9940 13636
rect 9548 13582 9550 13634
rect 9602 13582 9940 13634
rect 9548 13580 9940 13582
rect 10108 13634 10388 13636
rect 10108 13582 10334 13634
rect 10386 13582 10388 13634
rect 10108 13580 10388 13582
rect 9548 13570 9604 13580
rect 8764 13020 9828 13076
rect 8764 12290 8820 13020
rect 9772 12402 9828 13020
rect 9772 12350 9774 12402
rect 9826 12350 9828 12402
rect 9772 12338 9828 12350
rect 8764 12238 8766 12290
rect 8818 12238 8820 12290
rect 8764 12226 8820 12238
rect 9884 12292 9940 13580
rect 10332 13570 10388 13580
rect 10444 12740 10500 14476
rect 10892 12962 10948 15260
rect 11340 15314 11396 15932
rect 11452 15922 11508 15932
rect 11564 15764 11620 22092
rect 11676 20242 11732 22764
rect 12124 22708 12180 23212
rect 12348 23202 12404 23212
rect 12572 23044 12628 23548
rect 11676 20190 11678 20242
rect 11730 20190 11732 20242
rect 11676 18676 11732 20190
rect 11676 18610 11732 18620
rect 11900 22652 12180 22708
rect 12236 22988 12628 23044
rect 12684 23154 12740 23166
rect 12684 23102 12686 23154
rect 12738 23102 12740 23154
rect 12684 23044 12740 23102
rect 12796 23156 12852 23662
rect 13020 23548 13076 27804
rect 13188 27804 13300 27860
rect 13356 27860 13412 27870
rect 13692 27860 13748 27916
rect 13804 27906 13860 27916
rect 13916 27972 13972 27982
rect 13356 27858 13748 27860
rect 13356 27806 13358 27858
rect 13410 27806 13748 27858
rect 13356 27804 13748 27806
rect 13132 27794 13188 27804
rect 13356 27794 13412 27804
rect 13692 27188 13748 27804
rect 13916 27300 13972 27916
rect 13692 27122 13748 27132
rect 13804 27244 13972 27300
rect 13244 27076 13300 27086
rect 13244 26402 13300 27020
rect 13804 27074 13860 27244
rect 13804 27022 13806 27074
rect 13858 27022 13860 27074
rect 13804 26908 13860 27022
rect 14028 27188 14084 27198
rect 14028 27074 14084 27132
rect 14140 27186 14196 28140
rect 14252 28082 14308 31500
rect 14588 31220 14644 31724
rect 14700 31668 14756 31678
rect 14812 31668 14868 32284
rect 14924 31892 14980 32398
rect 15148 32002 15204 32844
rect 15260 32228 15316 35532
rect 16156 35586 16324 35588
rect 16156 35534 16158 35586
rect 16210 35534 16324 35586
rect 16156 35532 16324 35534
rect 16156 35522 16212 35532
rect 16044 35476 16100 35486
rect 15820 35474 16100 35476
rect 15820 35422 16046 35474
rect 16098 35422 16100 35474
rect 15820 35420 16100 35422
rect 15820 35026 15876 35420
rect 16044 35410 16100 35420
rect 15820 34974 15822 35026
rect 15874 34974 15876 35026
rect 15820 34962 15876 34974
rect 16268 34354 16324 35532
rect 16380 35308 16436 36318
rect 16380 35252 16548 35308
rect 16268 34302 16270 34354
rect 16322 34302 16324 34354
rect 16268 34290 16324 34302
rect 16492 34356 16548 35252
rect 16492 34354 16660 34356
rect 16492 34302 16494 34354
rect 16546 34302 16660 34354
rect 16492 34300 16660 34302
rect 16492 34290 16548 34300
rect 16156 34244 16212 34254
rect 15932 34132 15988 34142
rect 15484 34130 15988 34132
rect 15484 34078 15934 34130
rect 15986 34078 15988 34130
rect 15484 34076 15988 34078
rect 15484 34020 15540 34076
rect 15372 34018 15540 34020
rect 15372 33966 15486 34018
rect 15538 33966 15540 34018
rect 15372 33964 15540 33966
rect 15372 33346 15428 33964
rect 15484 33954 15540 33964
rect 15484 33460 15540 33470
rect 15484 33366 15540 33404
rect 15932 33458 15988 34076
rect 15932 33406 15934 33458
rect 15986 33406 15988 33458
rect 15932 33394 15988 33406
rect 15372 33294 15374 33346
rect 15426 33294 15428 33346
rect 15372 33282 15428 33294
rect 15484 33236 15540 33246
rect 15484 33142 15540 33180
rect 16044 33124 16100 33134
rect 15820 33122 16100 33124
rect 15820 33070 16046 33122
rect 16098 33070 16100 33122
rect 15820 33068 16100 33070
rect 15820 32786 15876 33068
rect 15820 32734 15822 32786
rect 15874 32734 15876 32786
rect 15820 32722 15876 32734
rect 15708 32676 15764 32686
rect 15484 32674 15764 32676
rect 15484 32622 15710 32674
rect 15762 32622 15764 32674
rect 15484 32620 15764 32622
rect 15372 32564 15428 32574
rect 15372 32470 15428 32508
rect 15484 32452 15540 32620
rect 15708 32610 15764 32620
rect 15932 32564 15988 32574
rect 15484 32396 15764 32452
rect 15260 32172 15540 32228
rect 15148 31950 15150 32002
rect 15202 31950 15204 32002
rect 15148 31938 15204 31950
rect 14924 31826 14980 31836
rect 14924 31668 14980 31678
rect 14812 31612 14924 31668
rect 14700 31574 14756 31612
rect 14924 31602 14980 31612
rect 15036 31666 15092 31678
rect 15036 31614 15038 31666
rect 15090 31614 15092 31666
rect 14924 31220 14980 31230
rect 14588 31218 14980 31220
rect 14588 31166 14926 31218
rect 14978 31166 14980 31218
rect 14588 31164 14980 31166
rect 14924 31154 14980 31164
rect 14252 28030 14254 28082
rect 14306 28030 14308 28082
rect 14252 28018 14308 28030
rect 14364 30884 14420 30894
rect 14364 27636 14420 30828
rect 14700 29764 14756 29774
rect 14756 29708 14868 29764
rect 14700 29698 14756 29708
rect 14140 27134 14142 27186
rect 14194 27134 14196 27186
rect 14140 27122 14196 27134
rect 14252 27580 14420 27636
rect 14588 27970 14644 27982
rect 14588 27918 14590 27970
rect 14642 27918 14644 27970
rect 14028 27022 14030 27074
rect 14082 27022 14084 27074
rect 14028 27010 14084 27022
rect 14252 26908 14308 27580
rect 14588 27412 14644 27918
rect 14588 27346 14644 27356
rect 14364 27074 14420 27086
rect 14364 27022 14366 27074
rect 14418 27022 14420 27074
rect 14364 26964 14420 27022
rect 14700 27076 14756 27086
rect 14588 26964 14644 26974
rect 14364 26962 14644 26964
rect 14364 26910 14590 26962
rect 14642 26910 14644 26962
rect 14364 26908 14644 26910
rect 13356 26852 13972 26908
rect 13356 26514 13412 26852
rect 13916 26740 13972 26852
rect 14140 26852 14308 26908
rect 14028 26740 14084 26750
rect 13916 26684 14028 26740
rect 14028 26674 14084 26684
rect 13356 26462 13358 26514
rect 13410 26462 13412 26514
rect 13356 26450 13412 26462
rect 13244 26350 13246 26402
rect 13298 26350 13300 26402
rect 13244 26338 13300 26350
rect 13580 26290 13636 26302
rect 13580 26238 13582 26290
rect 13634 26238 13636 26290
rect 13468 25284 13524 25294
rect 13132 24388 13188 24398
rect 13188 24332 13300 24388
rect 13132 24322 13188 24332
rect 12796 23090 12852 23100
rect 12908 23492 13076 23548
rect 11900 22370 11956 22652
rect 12012 22484 12068 22494
rect 12012 22390 12068 22428
rect 11900 22318 11902 22370
rect 11954 22318 11956 22370
rect 11676 18452 11732 18462
rect 11676 18358 11732 18396
rect 11676 16994 11732 17006
rect 11676 16942 11678 16994
rect 11730 16942 11732 16994
rect 11676 16324 11732 16942
rect 11676 16258 11732 16268
rect 11788 16100 11844 16138
rect 11340 15262 11342 15314
rect 11394 15262 11396 15314
rect 11340 15250 11396 15262
rect 11452 15708 11620 15764
rect 11676 16044 11788 16100
rect 11116 15202 11172 15214
rect 11116 15150 11118 15202
rect 11170 15150 11172 15202
rect 11116 15148 11172 15150
rect 11452 15148 11508 15708
rect 11004 15092 11172 15148
rect 11228 15092 11508 15148
rect 11676 15314 11732 16044
rect 11788 16034 11844 16044
rect 11676 15262 11678 15314
rect 11730 15262 11732 15314
rect 11004 14530 11060 15092
rect 11004 14478 11006 14530
rect 11058 14478 11060 14530
rect 11004 14466 11060 14478
rect 11116 14308 11172 14318
rect 11228 14308 11284 15092
rect 11676 14756 11732 15262
rect 11676 14690 11732 14700
rect 11788 15874 11844 15886
rect 11788 15822 11790 15874
rect 11842 15822 11844 15874
rect 11788 14642 11844 15822
rect 11900 15148 11956 22318
rect 12236 22370 12292 22988
rect 12684 22978 12740 22988
rect 12236 22318 12238 22370
rect 12290 22318 12292 22370
rect 12236 22306 12292 22318
rect 12348 22370 12404 22382
rect 12348 22318 12350 22370
rect 12402 22318 12404 22370
rect 12348 21924 12404 22318
rect 12908 22148 12964 23492
rect 13132 23044 13188 23054
rect 13132 22950 13188 22988
rect 12236 21868 12348 21924
rect 12012 20690 12068 20702
rect 12012 20638 12014 20690
rect 12066 20638 12068 20690
rect 12012 20580 12068 20638
rect 12012 20514 12068 20524
rect 12012 20132 12068 20142
rect 12012 19236 12068 20076
rect 12012 19170 12068 19180
rect 12124 16212 12180 16222
rect 12124 16098 12180 16156
rect 12124 16046 12126 16098
rect 12178 16046 12180 16098
rect 12124 16034 12180 16046
rect 11900 15092 12068 15148
rect 11788 14590 11790 14642
rect 11842 14590 11844 14642
rect 11788 14578 11844 14590
rect 11900 14644 11956 14654
rect 11900 14530 11956 14588
rect 11900 14478 11902 14530
rect 11954 14478 11956 14530
rect 11900 14466 11956 14478
rect 11116 14306 11284 14308
rect 11116 14254 11118 14306
rect 11170 14254 11284 14306
rect 11116 14252 11284 14254
rect 11340 14308 11396 14318
rect 12012 14308 12068 15092
rect 11340 14306 11620 14308
rect 11340 14254 11342 14306
rect 11394 14254 11620 14306
rect 11340 14252 11620 14254
rect 11116 13972 11172 14252
rect 11340 14242 11396 14252
rect 11116 13906 11172 13916
rect 10892 12910 10894 12962
rect 10946 12910 10948 12962
rect 10892 12898 10948 12910
rect 11452 13748 11508 13758
rect 10444 12674 10500 12684
rect 10668 12740 10724 12750
rect 9996 12292 10052 12302
rect 9884 12290 10052 12292
rect 9884 12238 9998 12290
rect 10050 12238 10052 12290
rect 9884 12236 10052 12238
rect 9996 12226 10052 12236
rect 8988 12180 9044 12190
rect 10332 12180 10388 12190
rect 10668 12180 10724 12684
rect 8988 12178 9268 12180
rect 8988 12126 8990 12178
rect 9042 12126 9268 12178
rect 8988 12124 9268 12126
rect 8988 12114 9044 12124
rect 8652 11890 8708 11900
rect 9100 11956 9156 11966
rect 8988 11844 9044 11854
rect 8540 10770 8596 10780
rect 8652 10836 8708 10846
rect 8652 10834 8932 10836
rect 8652 10782 8654 10834
rect 8706 10782 8932 10834
rect 8652 10780 8932 10782
rect 8652 10770 8708 10780
rect 7756 9662 7758 9714
rect 7810 9662 7812 9714
rect 7756 9650 7812 9662
rect 7868 10612 7924 10622
rect 7532 9314 7588 9324
rect 7868 8930 7924 10556
rect 8428 10610 8484 10622
rect 8428 10558 8430 10610
rect 8482 10558 8484 10610
rect 8428 10500 8484 10558
rect 8428 10434 8484 10444
rect 8764 10610 8820 10622
rect 8764 10558 8766 10610
rect 8818 10558 8820 10610
rect 8540 9940 8596 9950
rect 8764 9940 8820 10558
rect 8540 9938 8820 9940
rect 8540 9886 8542 9938
rect 8594 9886 8820 9938
rect 8540 9884 8820 9886
rect 8540 9874 8596 9884
rect 8764 9828 8820 9884
rect 8876 9828 8932 10780
rect 8988 10610 9044 11788
rect 9100 11618 9156 11900
rect 9100 11566 9102 11618
rect 9154 11566 9156 11618
rect 9100 11554 9156 11566
rect 9212 11506 9268 12124
rect 10332 12178 10724 12180
rect 10332 12126 10334 12178
rect 10386 12126 10724 12178
rect 10332 12124 10724 12126
rect 10332 12114 10388 12124
rect 9212 11454 9214 11506
rect 9266 11454 9268 11506
rect 9212 11442 9268 11454
rect 9996 12068 10052 12078
rect 9996 11506 10052 12012
rect 10108 12066 10164 12078
rect 10108 12014 10110 12066
rect 10162 12014 10164 12066
rect 10108 11844 10164 12014
rect 10108 11778 10164 11788
rect 9996 11454 9998 11506
rect 10050 11454 10052 11506
rect 9996 11442 10052 11454
rect 11340 11508 11396 11518
rect 11340 11414 11396 11452
rect 9436 11396 9492 11406
rect 11452 11396 11508 13692
rect 9436 11394 9604 11396
rect 9436 11342 9438 11394
rect 9490 11342 9604 11394
rect 9436 11340 9604 11342
rect 9436 11330 9492 11340
rect 9548 10836 9604 11340
rect 11452 11330 11508 11340
rect 10668 11172 10724 11182
rect 11564 11172 11620 14252
rect 11788 14252 12068 14308
rect 11788 12290 11844 14252
rect 11788 12238 11790 12290
rect 11842 12238 11844 12290
rect 11788 12180 11844 12238
rect 12236 12292 12292 21868
rect 12348 21858 12404 21868
rect 12460 22146 12964 22148
rect 12460 22094 12910 22146
rect 12962 22094 12964 22146
rect 12460 22092 12964 22094
rect 12348 21588 12404 21598
rect 12460 21588 12516 22092
rect 12908 22082 12964 22092
rect 13020 21924 13076 21934
rect 12348 21586 12516 21588
rect 12348 21534 12350 21586
rect 12402 21534 12516 21586
rect 12348 21532 12516 21534
rect 12684 21812 12740 21822
rect 12684 21698 12740 21756
rect 13020 21810 13076 21868
rect 13020 21758 13022 21810
rect 13074 21758 13076 21810
rect 13020 21746 13076 21758
rect 12684 21646 12686 21698
rect 12738 21646 12740 21698
rect 12348 18228 12404 21532
rect 12460 20130 12516 20142
rect 12460 20078 12462 20130
rect 12514 20078 12516 20130
rect 12460 18788 12516 20078
rect 12684 20018 12740 21646
rect 13244 21476 13300 24332
rect 13468 23826 13524 25228
rect 13468 23774 13470 23826
rect 13522 23774 13524 23826
rect 13468 22596 13524 23774
rect 13468 22530 13524 22540
rect 13468 22372 13524 22382
rect 13468 22146 13524 22316
rect 13468 22094 13470 22146
rect 13522 22094 13524 22146
rect 13468 21924 13524 22094
rect 13468 21858 13524 21868
rect 13356 21812 13412 21822
rect 13356 21718 13412 21756
rect 12684 19966 12686 20018
rect 12738 19966 12740 20018
rect 12684 19954 12740 19966
rect 12908 21420 13300 21476
rect 12908 19348 12964 21420
rect 13244 20130 13300 20142
rect 13580 20132 13636 26238
rect 13916 25732 13972 25742
rect 13916 25638 13972 25676
rect 14140 25508 14196 26852
rect 14476 26516 14532 26908
rect 14588 26898 14644 26908
rect 14700 26962 14756 27020
rect 14700 26910 14702 26962
rect 14754 26910 14756 26962
rect 14700 26898 14756 26910
rect 14476 26450 14532 26460
rect 14588 26740 14644 26750
rect 14588 26514 14644 26684
rect 14812 26516 14868 29708
rect 14588 26462 14590 26514
rect 14642 26462 14644 26514
rect 14588 26450 14644 26462
rect 14700 26514 14868 26516
rect 14700 26462 14814 26514
rect 14866 26462 14868 26514
rect 14700 26460 14868 26462
rect 14252 26292 14308 26302
rect 14252 25730 14308 26236
rect 14364 26292 14420 26302
rect 14700 26292 14756 26460
rect 14812 26450 14868 26460
rect 14924 26850 14980 26862
rect 14924 26798 14926 26850
rect 14978 26798 14980 26850
rect 14924 26404 14980 26798
rect 15036 26628 15092 31614
rect 15260 31668 15316 31678
rect 15260 31574 15316 31612
rect 15148 30884 15204 30894
rect 15148 29314 15204 30828
rect 15148 29262 15150 29314
rect 15202 29262 15204 29314
rect 15148 29250 15204 29262
rect 15372 30324 15428 30334
rect 15260 27074 15316 27086
rect 15260 27022 15262 27074
rect 15314 27022 15316 27074
rect 15260 26908 15316 27022
rect 15036 26562 15092 26572
rect 15148 26852 15316 26908
rect 15036 26404 15092 26414
rect 14924 26402 15092 26404
rect 14924 26350 15038 26402
rect 15090 26350 15092 26402
rect 14924 26348 15092 26350
rect 15036 26338 15092 26348
rect 14364 26290 14756 26292
rect 14364 26238 14366 26290
rect 14418 26238 14756 26290
rect 14364 26236 14756 26238
rect 14364 26226 14420 26236
rect 14252 25678 14254 25730
rect 14306 25678 14308 25730
rect 14252 25666 14308 25678
rect 14476 26068 14532 26078
rect 14028 25452 14196 25508
rect 13692 24724 13748 24734
rect 13692 23826 13748 24668
rect 13916 24388 13972 24398
rect 13804 24332 13916 24388
rect 13804 24162 13860 24332
rect 13916 24322 13972 24332
rect 13804 24110 13806 24162
rect 13858 24110 13860 24162
rect 13804 24098 13860 24110
rect 13692 23774 13694 23826
rect 13746 23774 13748 23826
rect 13692 23762 13748 23774
rect 13804 23380 13860 23390
rect 13804 22146 13860 23324
rect 13804 22094 13806 22146
rect 13858 22094 13860 22146
rect 13692 21812 13748 21822
rect 13692 21476 13748 21756
rect 13692 21410 13748 21420
rect 13244 20078 13246 20130
rect 13298 20078 13300 20130
rect 13244 19796 13300 20078
rect 13244 19730 13300 19740
rect 13468 20130 13636 20132
rect 13468 20078 13582 20130
rect 13634 20078 13636 20130
rect 13468 20076 13636 20078
rect 12908 19254 12964 19292
rect 12460 18722 12516 18732
rect 12460 18564 12516 18574
rect 12460 18450 12516 18508
rect 12460 18398 12462 18450
rect 12514 18398 12516 18450
rect 12460 18386 12516 18398
rect 12348 18172 12516 18228
rect 12348 16100 12404 16110
rect 12348 16006 12404 16044
rect 12460 12964 12516 18172
rect 13020 18116 13076 18126
rect 13020 16994 13076 18060
rect 13356 17780 13412 17790
rect 13356 17106 13412 17724
rect 13356 17054 13358 17106
rect 13410 17054 13412 17106
rect 13356 17042 13412 17054
rect 13020 16942 13022 16994
rect 13074 16942 13076 16994
rect 13020 16930 13076 16942
rect 13132 16996 13188 17006
rect 13132 16902 13188 16940
rect 12684 16212 12740 16222
rect 12684 16210 12852 16212
rect 12684 16158 12686 16210
rect 12738 16158 12852 16210
rect 12684 16156 12852 16158
rect 12684 16146 12740 16156
rect 12796 15988 12852 16156
rect 12572 15874 12628 15886
rect 12572 15822 12574 15874
rect 12626 15822 12628 15874
rect 12572 14644 12628 15822
rect 12796 15314 12852 15932
rect 13132 15652 13188 15662
rect 12796 15262 12798 15314
rect 12850 15262 12852 15314
rect 12796 15250 12852 15262
rect 13020 15316 13076 15326
rect 13020 15222 13076 15260
rect 13132 15314 13188 15596
rect 13468 15426 13524 20076
rect 13580 20066 13636 20076
rect 13580 19348 13636 19358
rect 13580 19234 13636 19292
rect 13580 19182 13582 19234
rect 13634 19182 13636 19234
rect 13580 19170 13636 19182
rect 13804 19236 13860 22094
rect 14028 20132 14084 25452
rect 14028 20066 14084 20076
rect 14140 25282 14196 25294
rect 14140 25230 14142 25282
rect 14194 25230 14196 25282
rect 14140 19908 14196 25230
rect 14364 24724 14420 24734
rect 14364 24612 14420 24668
rect 14252 24610 14420 24612
rect 14252 24558 14366 24610
rect 14418 24558 14420 24610
rect 14252 24556 14420 24558
rect 14252 24050 14308 24556
rect 14364 24546 14420 24556
rect 14252 23998 14254 24050
rect 14306 23998 14308 24050
rect 14252 23986 14308 23998
rect 14476 22370 14532 26012
rect 14924 26066 14980 26078
rect 14924 26014 14926 26066
rect 14978 26014 14980 26066
rect 14700 25284 14756 25294
rect 14700 25190 14756 25228
rect 14924 25172 14980 26014
rect 15036 25620 15092 25630
rect 15036 25506 15092 25564
rect 15036 25454 15038 25506
rect 15090 25454 15092 25506
rect 15036 25442 15092 25454
rect 14924 25106 14980 25116
rect 15148 25284 15204 26852
rect 14924 24834 14980 24846
rect 14924 24782 14926 24834
rect 14978 24782 14980 24834
rect 14812 24612 14868 24622
rect 14812 24518 14868 24556
rect 14700 24498 14756 24510
rect 14700 24446 14702 24498
rect 14754 24446 14756 24498
rect 14700 24388 14756 24446
rect 14700 24322 14756 24332
rect 14924 24164 14980 24782
rect 14812 24108 14980 24164
rect 14812 23380 14868 24108
rect 15148 24052 15204 25228
rect 15036 23996 15204 24052
rect 14924 23940 14980 23950
rect 15036 23940 15092 23996
rect 14924 23938 15092 23940
rect 14924 23886 14926 23938
rect 14978 23886 15092 23938
rect 14924 23884 15092 23886
rect 14924 23874 14980 23884
rect 14812 23314 14868 23324
rect 14476 22318 14478 22370
rect 14530 22318 14532 22370
rect 14476 22306 14532 22318
rect 14812 22258 14868 22270
rect 14812 22206 14814 22258
rect 14866 22206 14868 22258
rect 14252 22146 14308 22158
rect 14252 22094 14254 22146
rect 14306 22094 14308 22146
rect 14252 21924 14308 22094
rect 14252 21858 14308 21868
rect 14700 22148 14756 22158
rect 14700 21812 14756 22092
rect 14364 21756 14756 21812
rect 14252 21588 14308 21598
rect 14252 21494 14308 21532
rect 14364 20802 14420 21756
rect 14588 21586 14644 21598
rect 14588 21534 14590 21586
rect 14642 21534 14644 21586
rect 14588 21476 14644 21534
rect 14588 21410 14644 21420
rect 14364 20750 14366 20802
rect 14418 20750 14420 20802
rect 14364 20738 14420 20750
rect 14476 20914 14532 20926
rect 14476 20862 14478 20914
rect 14530 20862 14532 20914
rect 14476 20242 14532 20862
rect 14476 20190 14478 20242
rect 14530 20190 14532 20242
rect 14476 20178 14532 20190
rect 14700 20020 14756 20030
rect 14812 20020 14868 22206
rect 15036 21812 15092 23884
rect 15260 22260 15316 22270
rect 15260 22166 15316 22204
rect 15148 22148 15204 22158
rect 15148 22054 15204 22092
rect 15036 21756 15316 21812
rect 14924 21588 14980 21598
rect 14924 20914 14980 21532
rect 15148 21476 15204 21486
rect 15148 21382 15204 21420
rect 14924 20862 14926 20914
rect 14978 20862 14980 20914
rect 14924 20850 14980 20862
rect 15260 20802 15316 21756
rect 15260 20750 15262 20802
rect 15314 20750 15316 20802
rect 15260 20738 15316 20750
rect 15372 20356 15428 30268
rect 15484 26908 15540 32172
rect 15596 31778 15652 31790
rect 15596 31726 15598 31778
rect 15650 31726 15652 31778
rect 15596 31668 15652 31726
rect 15596 31602 15652 31612
rect 15708 31332 15764 32396
rect 15820 32340 15876 32350
rect 15932 32340 15988 32508
rect 15820 32338 15988 32340
rect 15820 32286 15822 32338
rect 15874 32286 15988 32338
rect 15820 32284 15988 32286
rect 15820 32274 15876 32284
rect 15820 31892 15876 31902
rect 15820 31798 15876 31836
rect 15596 30884 15652 30894
rect 15708 30884 15764 31276
rect 15652 30828 15764 30884
rect 15596 30790 15652 30828
rect 15932 30324 15988 32284
rect 16044 30994 16100 33068
rect 16156 33124 16212 34188
rect 16380 34132 16436 34142
rect 16380 34038 16436 34076
rect 16604 33460 16660 34300
rect 16156 33058 16212 33068
rect 16492 33458 16660 33460
rect 16492 33406 16606 33458
rect 16658 33406 16660 33458
rect 16492 33404 16660 33406
rect 16492 33236 16548 33404
rect 16604 33394 16660 33404
rect 16492 32786 16548 33180
rect 16492 32734 16494 32786
rect 16546 32734 16548 32786
rect 16492 32722 16548 32734
rect 16828 33124 16884 33134
rect 16828 32786 16884 33068
rect 16828 32734 16830 32786
rect 16882 32734 16884 32786
rect 16828 32452 16884 32734
rect 16828 32386 16884 32396
rect 16268 31780 16324 31790
rect 16268 31778 16548 31780
rect 16268 31726 16270 31778
rect 16322 31726 16548 31778
rect 16268 31724 16548 31726
rect 16268 31714 16324 31724
rect 16044 30942 16046 30994
rect 16098 30942 16100 30994
rect 16044 30930 16100 30942
rect 16380 31556 16436 31566
rect 16380 30996 16436 31500
rect 16380 30930 16436 30940
rect 16492 31106 16548 31724
rect 16604 31668 16660 31678
rect 16828 31668 16884 31678
rect 16604 31666 16884 31668
rect 16604 31614 16606 31666
rect 16658 31614 16830 31666
rect 16882 31614 16884 31666
rect 16604 31612 16884 31614
rect 16604 31602 16660 31612
rect 16828 31602 16884 31612
rect 16940 31444 16996 37100
rect 17500 37154 17556 37166
rect 17500 37102 17502 37154
rect 17554 37102 17556 37154
rect 17500 37044 17556 37102
rect 17500 36978 17556 36988
rect 17164 36708 17220 36718
rect 17164 36482 17220 36652
rect 17164 36430 17166 36482
rect 17218 36430 17220 36482
rect 17164 36260 17220 36430
rect 17388 36372 17444 36382
rect 17388 36278 17444 36316
rect 17164 36194 17220 36204
rect 17052 34356 17108 34366
rect 17052 33348 17108 34300
rect 17612 34356 17668 37324
rect 17836 36594 17892 38612
rect 17836 36542 17838 36594
rect 17890 36542 17892 36594
rect 17836 36484 17892 36542
rect 17836 36418 17892 36428
rect 17948 36372 18004 42588
rect 18732 42532 18788 42542
rect 18172 42530 18788 42532
rect 18172 42478 18734 42530
rect 18786 42478 18788 42530
rect 18172 42476 18788 42478
rect 18172 41970 18228 42476
rect 18732 42466 18788 42476
rect 18172 41918 18174 41970
rect 18226 41918 18228 41970
rect 18172 41906 18228 41918
rect 19068 41972 19124 42590
rect 19404 42644 19460 42654
rect 19404 42550 19460 42588
rect 19068 41906 19124 41916
rect 19516 42530 19572 42542
rect 19516 42478 19518 42530
rect 19570 42478 19572 42530
rect 19180 41188 19236 41198
rect 19516 41188 19572 42478
rect 19180 41186 19572 41188
rect 19180 41134 19182 41186
rect 19234 41134 19518 41186
rect 19570 41134 19572 41186
rect 19180 41132 19572 41134
rect 19180 41122 19236 41132
rect 19516 41122 19572 41132
rect 19628 41524 19684 43260
rect 20076 43092 20132 43102
rect 20076 42868 20132 43036
rect 20076 42866 20356 42868
rect 20076 42814 20078 42866
rect 20130 42814 20356 42866
rect 20076 42812 20356 42814
rect 20076 42802 20132 42812
rect 20300 42644 20356 42812
rect 20412 42756 20468 43596
rect 20524 43586 20580 43596
rect 20524 43426 20580 43438
rect 20524 43374 20526 43426
rect 20578 43374 20580 43426
rect 20524 42978 20580 43374
rect 20524 42926 20526 42978
rect 20578 42926 20580 42978
rect 20524 42914 20580 42926
rect 20412 42700 20580 42756
rect 20300 42588 20468 42644
rect 20412 42586 20468 42588
rect 20412 42534 20414 42586
rect 20466 42534 20468 42586
rect 20524 42642 20580 42700
rect 20524 42590 20526 42642
rect 20578 42590 20580 42642
rect 20524 42578 20580 42590
rect 20412 42522 20468 42534
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 20300 41860 20356 41870
rect 20636 41860 20692 44156
rect 20972 43652 21028 45166
rect 21420 44322 21476 44334
rect 21420 44270 21422 44322
rect 21474 44270 21476 44322
rect 21420 43764 21476 44270
rect 21420 43698 21476 43708
rect 21028 43596 21140 43652
rect 20972 43586 21028 43596
rect 20748 43540 20804 43550
rect 20748 43446 20804 43484
rect 20748 41972 20804 41982
rect 20748 41878 20804 41916
rect 21084 41970 21140 43596
rect 21420 43426 21476 43438
rect 21420 43374 21422 43426
rect 21474 43374 21476 43426
rect 21308 42532 21364 42542
rect 21308 42084 21364 42476
rect 21084 41918 21086 41970
rect 21138 41918 21140 41970
rect 21084 41906 21140 41918
rect 21196 42082 21364 42084
rect 21196 42030 21310 42082
rect 21362 42030 21364 42082
rect 21196 42028 21364 42030
rect 20300 41858 20692 41860
rect 20300 41806 20302 41858
rect 20354 41806 20692 41858
rect 20300 41804 20692 41806
rect 20300 41794 20356 41804
rect 19628 41074 19684 41468
rect 20188 41524 20244 41534
rect 20188 41298 20244 41468
rect 20188 41246 20190 41298
rect 20242 41246 20244 41298
rect 20188 41234 20244 41246
rect 19628 41022 19630 41074
rect 19682 41022 19684 41074
rect 19628 41010 19684 41022
rect 19852 41076 19908 41086
rect 19852 40982 19908 41020
rect 18396 40964 18452 40974
rect 18732 40964 18788 40974
rect 18956 40964 19012 40974
rect 18396 40962 18788 40964
rect 18396 40910 18398 40962
rect 18450 40910 18734 40962
rect 18786 40910 18788 40962
rect 18396 40908 18788 40910
rect 18396 40898 18452 40908
rect 18732 40516 18788 40908
rect 18732 40450 18788 40460
rect 18844 40962 19012 40964
rect 18844 40910 18958 40962
rect 19010 40910 19012 40962
rect 18844 40908 19012 40910
rect 18844 40404 18900 40908
rect 18956 40898 19012 40908
rect 19068 40962 19124 40974
rect 19068 40910 19070 40962
rect 19122 40910 19124 40962
rect 19068 40404 19124 40910
rect 19836 40796 20100 40806
rect 18844 40310 18900 40348
rect 18956 40348 19124 40404
rect 19404 40740 19460 40750
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19404 40402 19460 40684
rect 19404 40350 19406 40402
rect 19458 40350 19460 40402
rect 18396 39620 18452 39630
rect 18396 39526 18452 39564
rect 18956 39618 19012 40348
rect 19404 40338 19460 40350
rect 21196 40404 21252 42028
rect 21308 42018 21364 42028
rect 21420 42084 21476 43374
rect 21420 42018 21476 42028
rect 21420 41300 21476 41310
rect 21196 40310 21252 40348
rect 21308 40628 21364 40638
rect 18956 39566 18958 39618
rect 19010 39566 19012 39618
rect 18956 39554 19012 39566
rect 19516 40290 19572 40302
rect 19516 40238 19518 40290
rect 19570 40238 19572 40290
rect 19068 39508 19124 39518
rect 19068 39414 19124 39452
rect 19516 38668 19572 40238
rect 21308 39620 21364 40572
rect 21420 40626 21476 41244
rect 21420 40574 21422 40626
rect 21474 40574 21476 40626
rect 21420 40562 21476 40574
rect 20972 39618 21364 39620
rect 20972 39566 21310 39618
rect 21362 39566 21364 39618
rect 20972 39564 21364 39566
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19404 38612 19572 38668
rect 20860 38834 20916 38846
rect 20860 38782 20862 38834
rect 20914 38782 20916 38834
rect 18732 38500 18788 38510
rect 18732 38162 18788 38444
rect 18732 38110 18734 38162
rect 18786 38110 18788 38162
rect 18732 38098 18788 38110
rect 18060 37604 18116 37614
rect 18060 37154 18116 37548
rect 18060 37102 18062 37154
rect 18114 37102 18116 37154
rect 18060 37090 18116 37102
rect 17948 36306 18004 36316
rect 18508 36484 18564 36494
rect 18508 35924 18564 36428
rect 19404 36148 19460 38612
rect 19964 38052 20020 38062
rect 19964 37958 20020 37996
rect 20188 37938 20244 37950
rect 20188 37886 20190 37938
rect 20242 37886 20244 37938
rect 19628 37826 19684 37838
rect 19628 37774 19630 37826
rect 19682 37774 19684 37826
rect 19516 36596 19572 36606
rect 19516 36482 19572 36540
rect 19516 36430 19518 36482
rect 19570 36430 19572 36482
rect 19516 36418 19572 36430
rect 19628 36484 19684 37774
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37380 20244 37886
rect 20860 37940 20916 38782
rect 20860 37846 20916 37884
rect 20188 37314 20244 37324
rect 20524 37268 20580 37278
rect 20300 37212 20524 37268
rect 20188 37156 20244 37166
rect 20076 37154 20244 37156
rect 20076 37102 20190 37154
rect 20242 37102 20244 37154
rect 20076 37100 20244 37102
rect 20076 36594 20132 37100
rect 20188 37090 20244 37100
rect 20076 36542 20078 36594
rect 20130 36542 20132 36594
rect 20076 36530 20132 36542
rect 19964 36484 20020 36494
rect 19628 36482 20020 36484
rect 19628 36430 19966 36482
rect 20018 36430 20020 36482
rect 19628 36428 20020 36430
rect 19964 36418 20020 36428
rect 20188 36484 20244 36494
rect 20300 36484 20356 37212
rect 20524 37202 20580 37212
rect 20972 37268 21028 39564
rect 21308 39554 21364 39564
rect 21420 38946 21476 38958
rect 21420 38894 21422 38946
rect 21474 38894 21476 38946
rect 21196 38834 21252 38846
rect 21196 38782 21198 38834
rect 21250 38782 21252 38834
rect 21196 38668 21252 38782
rect 21196 38612 21364 38668
rect 21196 38052 21252 38062
rect 21196 37604 21252 37996
rect 21308 37828 21364 38612
rect 21420 38612 21476 38894
rect 21420 38546 21476 38556
rect 21308 37734 21364 37772
rect 21532 37716 21588 45276
rect 21756 45218 21812 45230
rect 21756 45166 21758 45218
rect 21810 45166 21812 45218
rect 21756 44884 21812 45166
rect 21756 44818 21812 44828
rect 21868 44322 21924 45612
rect 22092 45332 22148 45342
rect 22092 45106 22148 45276
rect 22092 45054 22094 45106
rect 22146 45054 22148 45106
rect 22092 45042 22148 45054
rect 21868 44270 21870 44322
rect 21922 44270 21924 44322
rect 21868 44258 21924 44270
rect 22204 43652 22260 48860
rect 22540 48916 22596 48926
rect 22540 48822 22596 48860
rect 22428 48130 22484 48142
rect 22428 48078 22430 48130
rect 22482 48078 22484 48130
rect 22428 48020 22484 48078
rect 22764 48020 22820 48974
rect 22428 47964 22820 48020
rect 22764 47346 22820 47964
rect 22764 47294 22766 47346
rect 22818 47294 22820 47346
rect 22764 47282 22820 47294
rect 23324 47124 23380 49980
rect 23436 49812 23492 49822
rect 23548 49812 23604 50372
rect 23436 49810 23604 49812
rect 23436 49758 23438 49810
rect 23490 49758 23604 49810
rect 23436 49756 23604 49758
rect 23436 49746 23492 49756
rect 23548 48804 23604 49756
rect 23548 48738 23604 48748
rect 24108 49028 24164 49038
rect 24556 49028 24612 50540
rect 24668 49924 24724 49934
rect 24668 49830 24724 49868
rect 24108 49026 24612 49028
rect 24108 48974 24110 49026
rect 24162 48974 24612 49026
rect 24108 48972 24612 48974
rect 24108 48244 24164 48972
rect 24108 48178 24164 48188
rect 24332 48804 24388 48814
rect 24332 47458 24388 48748
rect 24668 48130 24724 48142
rect 24668 48078 24670 48130
rect 24722 48078 24724 48130
rect 24668 47796 24724 48078
rect 24668 47730 24724 47740
rect 24332 47406 24334 47458
rect 24386 47406 24388 47458
rect 24332 47394 24388 47406
rect 23324 47068 23604 47124
rect 23212 45890 23268 45902
rect 23212 45838 23214 45890
rect 23266 45838 23268 45890
rect 22764 45780 22820 45790
rect 22764 45686 22820 45724
rect 22764 45444 22820 45454
rect 22316 44210 22372 44222
rect 22316 44158 22318 44210
rect 22370 44158 22372 44210
rect 22316 43876 22372 44158
rect 22652 44212 22708 44222
rect 22652 44118 22708 44156
rect 22764 44212 22820 45388
rect 23212 45108 23268 45838
rect 23212 44994 23268 45052
rect 23212 44942 23214 44994
rect 23266 44942 23268 44994
rect 23212 44930 23268 44942
rect 23548 44996 23604 47068
rect 23660 46674 23716 46686
rect 23660 46622 23662 46674
rect 23714 46622 23716 46674
rect 23660 46564 23716 46622
rect 24444 46564 24500 46574
rect 23660 46562 24500 46564
rect 23660 46510 24446 46562
rect 24498 46510 24500 46562
rect 23660 46508 24500 46510
rect 23660 45332 23716 46508
rect 24444 46498 24500 46508
rect 23884 46004 23940 46014
rect 23884 45910 23940 45948
rect 24332 45780 24388 45790
rect 23660 45266 23716 45276
rect 23772 45556 23828 45566
rect 23548 44930 23604 44940
rect 23660 44436 23716 44446
rect 23772 44436 23828 45500
rect 23660 44434 23828 44436
rect 23660 44382 23662 44434
rect 23714 44382 23828 44434
rect 23660 44380 23828 44382
rect 23884 44996 23940 45006
rect 23660 44370 23716 44380
rect 23100 44322 23156 44334
rect 23100 44270 23102 44322
rect 23154 44270 23156 44322
rect 23100 44212 23156 44270
rect 22764 44156 23156 44212
rect 23548 44210 23604 44222
rect 23548 44158 23550 44210
rect 23602 44158 23604 44210
rect 22316 43810 22372 43820
rect 22316 43652 22372 43662
rect 22204 43650 22708 43652
rect 22204 43598 22318 43650
rect 22370 43598 22708 43650
rect 22204 43596 22708 43598
rect 22316 43586 22372 43596
rect 22540 43316 22596 43326
rect 22540 42754 22596 43260
rect 22540 42702 22542 42754
rect 22594 42702 22596 42754
rect 21868 42532 21924 42542
rect 21644 42530 21924 42532
rect 21644 42478 21870 42530
rect 21922 42478 21924 42530
rect 21644 42476 21924 42478
rect 21644 42082 21700 42476
rect 21868 42466 21924 42476
rect 22316 42532 22372 42542
rect 22316 42438 22372 42476
rect 21644 42030 21646 42082
rect 21698 42030 21700 42082
rect 21644 41860 21700 42030
rect 22540 41970 22596 42702
rect 22652 42756 22708 43596
rect 22764 43204 22820 44156
rect 23548 44100 23604 44158
rect 23212 44044 23604 44100
rect 23772 44212 23828 44222
rect 23884 44212 23940 44940
rect 24332 44546 24388 45724
rect 24780 45220 24836 54460
rect 24892 48914 24948 48926
rect 24892 48862 24894 48914
rect 24946 48862 24948 48914
rect 24892 48020 24948 48862
rect 24892 47954 24948 47964
rect 24892 47460 24948 47470
rect 24892 47366 24948 47404
rect 24332 44494 24334 44546
rect 24386 44494 24388 44546
rect 24332 44482 24388 44494
rect 24444 45164 24836 45220
rect 24220 44436 24276 44446
rect 24220 44322 24276 44380
rect 24220 44270 24222 44322
rect 24274 44270 24276 44322
rect 24220 44258 24276 44270
rect 23772 44210 23940 44212
rect 23772 44158 23774 44210
rect 23826 44158 23940 44210
rect 23772 44156 23940 44158
rect 23212 43652 23268 44044
rect 23772 43876 23828 44156
rect 23548 43820 23828 43876
rect 23436 43652 23492 43662
rect 23548 43652 23604 43820
rect 22876 43650 23380 43652
rect 22876 43598 23214 43650
rect 23266 43598 23380 43650
rect 22876 43596 23380 43598
rect 22876 43426 22932 43596
rect 23212 43586 23268 43596
rect 22876 43374 22878 43426
rect 22930 43374 22932 43426
rect 22876 43362 22932 43374
rect 22764 43148 22932 43204
rect 22764 42756 22820 42766
rect 22652 42700 22764 42756
rect 22764 42662 22820 42700
rect 22540 41918 22542 41970
rect 22594 41918 22596 41970
rect 22540 41906 22596 41918
rect 21644 41804 21924 41860
rect 21644 40962 21700 40974
rect 21644 40910 21646 40962
rect 21698 40910 21700 40962
rect 21644 40404 21700 40910
rect 21868 40852 21924 41804
rect 22764 41858 22820 41870
rect 22764 41806 22766 41858
rect 22818 41806 22820 41858
rect 22092 41300 22148 41310
rect 22092 41206 22148 41244
rect 22428 41188 22484 41198
rect 22428 41094 22484 41132
rect 22540 41188 22596 41198
rect 22764 41188 22820 41806
rect 22540 41186 22820 41188
rect 22540 41134 22542 41186
rect 22594 41134 22820 41186
rect 22540 41132 22820 41134
rect 22540 41122 22596 41132
rect 21868 40786 21924 40796
rect 22652 40962 22708 40974
rect 22652 40910 22654 40962
rect 22706 40910 22708 40962
rect 22204 40628 22260 40638
rect 22092 40572 22204 40628
rect 22092 40516 22148 40572
rect 22204 40562 22260 40572
rect 21644 40338 21700 40348
rect 21868 40460 22148 40516
rect 22540 40516 22596 40526
rect 21868 40402 21924 40460
rect 22540 40422 22596 40460
rect 21868 40350 21870 40402
rect 21922 40350 21924 40402
rect 21868 40338 21924 40350
rect 22652 40180 22708 40910
rect 22764 40964 22820 40974
rect 22764 40870 22820 40908
rect 22092 40124 22708 40180
rect 22764 40740 22820 40750
rect 22092 39730 22148 40124
rect 22092 39678 22094 39730
rect 22146 39678 22148 39730
rect 22092 39666 22148 39678
rect 21980 39284 22036 39294
rect 21868 38834 21924 38846
rect 21868 38782 21870 38834
rect 21922 38782 21924 38834
rect 21868 38668 21924 38782
rect 21756 38612 21924 38668
rect 21756 37940 21812 38556
rect 21756 37874 21812 37884
rect 21868 38050 21924 38062
rect 21868 37998 21870 38050
rect 21922 37998 21924 38050
rect 21868 37716 21924 37998
rect 21532 37660 21924 37716
rect 21196 37548 21364 37604
rect 20972 37266 21252 37268
rect 20972 37214 20974 37266
rect 21026 37214 21252 37266
rect 20972 37212 21252 37214
rect 20972 37202 21028 37212
rect 21196 36932 21252 37212
rect 21308 37266 21364 37548
rect 21308 37214 21310 37266
rect 21362 37214 21364 37266
rect 21308 37156 21364 37214
rect 21420 37268 21476 37278
rect 21420 37174 21476 37212
rect 21308 37090 21364 37100
rect 21196 36876 21476 36932
rect 20636 36596 20692 36606
rect 20636 36502 20692 36540
rect 21420 36594 21476 36876
rect 21420 36542 21422 36594
rect 21474 36542 21476 36594
rect 21420 36530 21476 36542
rect 20188 36482 20356 36484
rect 20188 36430 20190 36482
rect 20242 36430 20356 36482
rect 20188 36428 20356 36430
rect 20188 36418 20244 36428
rect 19740 36260 19796 36270
rect 19628 36258 19796 36260
rect 19628 36206 19742 36258
rect 19794 36206 19796 36258
rect 19628 36204 19796 36206
rect 19628 36148 19684 36204
rect 19740 36194 19796 36204
rect 19404 36092 19684 36148
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 18732 35924 18788 35934
rect 18508 35922 18788 35924
rect 18508 35870 18510 35922
rect 18562 35870 18734 35922
rect 18786 35870 18788 35922
rect 18508 35868 18788 35870
rect 18508 35858 18564 35868
rect 18732 35858 18788 35868
rect 19068 35810 19124 35822
rect 19068 35758 19070 35810
rect 19122 35758 19124 35810
rect 17612 34290 17668 34300
rect 17948 35026 18004 35038
rect 17948 34974 17950 35026
rect 18002 34974 18004 35026
rect 17948 34132 18004 34974
rect 18396 34356 18452 34366
rect 18396 34262 18452 34300
rect 18284 34132 18340 34142
rect 18004 34130 18340 34132
rect 18004 34078 18286 34130
rect 18338 34078 18340 34130
rect 18004 34076 18340 34078
rect 17948 34038 18004 34076
rect 17724 34020 17780 34030
rect 17724 33926 17780 33964
rect 17836 33908 17892 33918
rect 17836 33906 18228 33908
rect 17836 33854 17838 33906
rect 17890 33854 18228 33906
rect 17836 33852 18228 33854
rect 17836 33842 17892 33852
rect 18172 33458 18228 33852
rect 18284 33684 18340 34076
rect 18620 34130 18676 34142
rect 18620 34078 18622 34130
rect 18674 34078 18676 34130
rect 18508 34020 18564 34030
rect 18508 33926 18564 33964
rect 18284 33618 18340 33628
rect 18508 33796 18564 33806
rect 18172 33406 18174 33458
rect 18226 33406 18228 33458
rect 18172 33394 18228 33406
rect 17388 33348 17444 33358
rect 17052 33346 17444 33348
rect 17052 33294 17054 33346
rect 17106 33294 17390 33346
rect 17442 33294 17444 33346
rect 17052 33292 17444 33294
rect 17052 33282 17108 33292
rect 17388 33282 17444 33292
rect 17612 33124 17668 33134
rect 17276 33012 17332 33022
rect 16940 31378 16996 31388
rect 17052 31666 17108 31678
rect 17052 31614 17054 31666
rect 17106 31614 17108 31666
rect 17052 31220 17108 31614
rect 17164 31668 17220 31678
rect 17164 31554 17220 31612
rect 17164 31502 17166 31554
rect 17218 31502 17220 31554
rect 17164 31490 17220 31502
rect 17164 31220 17220 31230
rect 17052 31164 17164 31220
rect 17164 31154 17220 31164
rect 16492 31054 16494 31106
rect 16546 31054 16548 31106
rect 16492 30548 16548 31054
rect 17276 30996 17332 32956
rect 17388 31668 17444 31678
rect 17388 31574 17444 31612
rect 16492 30482 16548 30492
rect 16828 30940 17332 30996
rect 16156 30324 16212 30334
rect 15932 30322 16212 30324
rect 15932 30270 16158 30322
rect 16210 30270 16212 30322
rect 15932 30268 16212 30270
rect 16156 30258 16212 30268
rect 16268 30100 16324 30110
rect 16604 30100 16660 30110
rect 16268 30098 16660 30100
rect 16268 30046 16270 30098
rect 16322 30046 16606 30098
rect 16658 30046 16660 30098
rect 16268 30044 16660 30046
rect 16268 30034 16324 30044
rect 16604 30034 16660 30044
rect 15932 27412 15988 27422
rect 15484 26852 15876 26908
rect 15484 26178 15540 26190
rect 15484 26126 15486 26178
rect 15538 26126 15540 26178
rect 15484 25620 15540 26126
rect 15820 25620 15876 26852
rect 15932 26514 15988 27356
rect 16044 26962 16100 26974
rect 16044 26910 16046 26962
rect 16098 26910 16100 26962
rect 16044 26908 16100 26910
rect 16828 26908 16884 30940
rect 17500 30884 17556 30894
rect 17052 30882 17556 30884
rect 17052 30830 17502 30882
rect 17554 30830 17556 30882
rect 17052 30828 17556 30830
rect 17052 30322 17108 30828
rect 17500 30818 17556 30828
rect 17612 30660 17668 33068
rect 17724 31554 17780 31566
rect 17724 31502 17726 31554
rect 17778 31502 17780 31554
rect 17724 31332 17780 31502
rect 18060 31554 18116 31566
rect 18060 31502 18062 31554
rect 18114 31502 18116 31554
rect 18060 31444 18116 31502
rect 18508 31444 18564 33740
rect 18620 32788 18676 34078
rect 18844 34132 18900 34142
rect 19068 34132 19124 35758
rect 21308 34692 21364 34702
rect 20188 34690 21364 34692
rect 20188 34638 21310 34690
rect 21362 34638 21364 34690
rect 20188 34636 21364 34638
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20188 34242 20244 34636
rect 21308 34626 21364 34636
rect 21532 34468 21588 37660
rect 21644 37380 21700 37390
rect 21644 37268 21700 37324
rect 21868 37268 21924 37278
rect 21644 37266 21812 37268
rect 21644 37214 21646 37266
rect 21698 37214 21812 37266
rect 21644 37212 21812 37214
rect 21644 37202 21700 37212
rect 21644 34804 21700 34814
rect 21644 34710 21700 34748
rect 20188 34190 20190 34242
rect 20242 34190 20244 34242
rect 20188 34178 20244 34190
rect 20636 34412 21588 34468
rect 18844 34130 19124 34132
rect 18844 34078 18846 34130
rect 18898 34078 19124 34130
rect 18844 34076 19124 34078
rect 19516 34130 19572 34142
rect 19516 34078 19518 34130
rect 19570 34078 19572 34130
rect 18844 33572 18900 34076
rect 18844 33506 18900 33516
rect 19068 33684 19124 33694
rect 18620 32722 18676 32732
rect 18060 31388 18564 31444
rect 17724 31266 17780 31276
rect 17724 30996 17780 31006
rect 17724 30902 17780 30940
rect 17500 30604 17668 30660
rect 18396 30882 18452 30894
rect 18396 30830 18398 30882
rect 18450 30830 18452 30882
rect 17052 30270 17054 30322
rect 17106 30270 17108 30322
rect 17052 30258 17108 30270
rect 17164 30548 17220 30558
rect 16940 30212 16996 30222
rect 16940 30118 16996 30156
rect 17164 30210 17220 30492
rect 17388 30436 17444 30446
rect 17164 30158 17166 30210
rect 17218 30158 17220 30210
rect 17164 30146 17220 30158
rect 17276 30380 17388 30436
rect 17276 26908 17332 30380
rect 17388 30370 17444 30380
rect 17500 30212 17556 30604
rect 18060 30548 18116 30558
rect 17388 30156 17556 30212
rect 17836 30212 17892 30222
rect 17388 27970 17444 30156
rect 17836 30118 17892 30156
rect 18060 30210 18116 30492
rect 18060 30158 18062 30210
rect 18114 30158 18116 30210
rect 18060 30146 18116 30158
rect 18396 30212 18452 30830
rect 18508 30772 18564 31388
rect 18620 31666 18676 31678
rect 18620 31614 18622 31666
rect 18674 31614 18676 31666
rect 18620 30996 18676 31614
rect 18732 31668 18788 31678
rect 18732 31106 18788 31612
rect 18956 31666 19012 31678
rect 18956 31614 18958 31666
rect 19010 31614 19012 31666
rect 18956 31332 19012 31614
rect 19068 31556 19124 33628
rect 19516 33348 19572 34078
rect 20300 33460 20356 33470
rect 20300 33366 20356 33404
rect 19516 33282 19572 33292
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19740 32788 19796 32798
rect 19740 32562 19796 32732
rect 19740 32510 19742 32562
rect 19794 32510 19796 32562
rect 19740 32498 19796 32510
rect 19740 32338 19796 32350
rect 19740 32286 19742 32338
rect 19794 32286 19796 32338
rect 19740 32228 19796 32286
rect 19628 32172 19796 32228
rect 20076 32338 20132 32350
rect 20076 32286 20078 32338
rect 20130 32286 20132 32338
rect 19628 32116 19684 32172
rect 19180 32060 19684 32116
rect 19180 31778 19236 32060
rect 19180 31726 19182 31778
rect 19234 31726 19236 31778
rect 19180 31714 19236 31726
rect 19516 31892 19908 31948
rect 19516 31556 19572 31892
rect 19068 31500 19572 31556
rect 18956 31276 19460 31332
rect 18844 31220 18900 31230
rect 18900 31164 19236 31220
rect 18844 31126 18900 31164
rect 18732 31054 18734 31106
rect 18786 31054 18788 31106
rect 18732 31042 18788 31054
rect 18620 30930 18676 30940
rect 19068 30996 19124 31006
rect 18844 30772 18900 30782
rect 18508 30716 18676 30772
rect 18396 30156 18564 30212
rect 17724 30100 17780 30110
rect 17612 29988 17668 29998
rect 17612 29894 17668 29932
rect 17500 29652 17556 29662
rect 17724 29652 17780 30044
rect 17500 29650 17780 29652
rect 17500 29598 17502 29650
rect 17554 29598 17780 29650
rect 17500 29596 17780 29598
rect 17948 29986 18004 29998
rect 17948 29934 17950 29986
rect 18002 29934 18004 29986
rect 17500 29586 17556 29596
rect 17836 29204 17892 29214
rect 17836 29110 17892 29148
rect 17948 28868 18004 29934
rect 18396 29986 18452 29998
rect 18396 29934 18398 29986
rect 18450 29934 18452 29986
rect 18060 29540 18116 29550
rect 18060 29538 18228 29540
rect 18060 29486 18062 29538
rect 18114 29486 18228 29538
rect 18060 29484 18228 29486
rect 18060 29474 18116 29484
rect 18060 28868 18116 28878
rect 17948 28866 18116 28868
rect 17948 28814 18062 28866
rect 18114 28814 18116 28866
rect 17948 28812 18116 28814
rect 18060 28802 18116 28812
rect 18172 28644 18228 29484
rect 18396 29428 18452 29934
rect 18284 29372 18452 29428
rect 18284 28754 18340 29372
rect 18508 29316 18564 30156
rect 18620 29538 18676 30716
rect 18844 30770 19012 30772
rect 18844 30718 18846 30770
rect 18898 30718 19012 30770
rect 18844 30716 19012 30718
rect 18844 30706 18900 30716
rect 18732 30548 18788 30558
rect 18732 30434 18788 30492
rect 18732 30382 18734 30434
rect 18786 30382 18788 30434
rect 18732 30370 18788 30382
rect 18956 30322 19012 30716
rect 18956 30270 18958 30322
rect 19010 30270 19012 30322
rect 18956 30212 19012 30270
rect 18956 30146 19012 30156
rect 18620 29486 18622 29538
rect 18674 29486 18676 29538
rect 18620 29474 18676 29486
rect 18284 28702 18286 28754
rect 18338 28702 18340 28754
rect 18284 28690 18340 28702
rect 18396 29260 18564 29316
rect 19068 29314 19124 30940
rect 19180 30772 19236 31164
rect 19404 31218 19460 31276
rect 19404 31166 19406 31218
rect 19458 31166 19460 31218
rect 19404 30772 19460 31166
rect 19516 31106 19572 31500
rect 19516 31054 19518 31106
rect 19570 31054 19572 31106
rect 19516 31042 19572 31054
rect 19628 31778 19684 31790
rect 19628 31726 19630 31778
rect 19682 31726 19684 31778
rect 19628 30996 19684 31726
rect 19852 31778 19908 31892
rect 19852 31726 19854 31778
rect 19906 31726 19908 31778
rect 19852 31714 19908 31726
rect 20076 31556 20132 32286
rect 20524 31668 20580 31678
rect 20524 31574 20580 31612
rect 20076 31500 20244 31556
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19964 31220 20020 31230
rect 20188 31220 20244 31500
rect 19964 31218 20244 31220
rect 19964 31166 19966 31218
rect 20018 31166 20244 31218
rect 19964 31164 20244 31166
rect 20300 31220 20356 31230
rect 19964 31154 20020 31164
rect 20300 31126 20356 31164
rect 19628 30930 19684 30940
rect 19852 30996 19908 31006
rect 19852 30902 19908 30940
rect 20076 30994 20132 31006
rect 20076 30942 20078 30994
rect 20130 30942 20132 30994
rect 20076 30772 20132 30942
rect 19404 30716 20132 30772
rect 19180 30706 19236 30716
rect 19068 29262 19070 29314
rect 19122 29262 19124 29314
rect 17388 27918 17390 27970
rect 17442 27918 17444 27970
rect 17388 27906 17444 27918
rect 17500 28588 18228 28644
rect 16044 26852 16436 26908
rect 16828 26852 16996 26908
rect 17276 26852 17444 26908
rect 15932 26462 15934 26514
rect 15986 26462 15988 26514
rect 15932 26450 15988 26462
rect 16380 26514 16436 26852
rect 16380 26462 16382 26514
rect 16434 26462 16436 26514
rect 16380 26450 16436 26462
rect 16716 26292 16772 26302
rect 16716 26198 16772 26236
rect 16044 25620 16100 25630
rect 15820 25618 16660 25620
rect 15820 25566 16046 25618
rect 16098 25566 16660 25618
rect 15820 25564 16660 25566
rect 15484 25526 15540 25564
rect 16044 25554 16100 25564
rect 15596 25172 15652 25182
rect 15596 24834 15652 25116
rect 15596 24782 15598 24834
rect 15650 24782 15652 24834
rect 15596 24770 15652 24782
rect 15708 24836 15764 24846
rect 16268 24836 16324 24846
rect 15708 24834 16324 24836
rect 15708 24782 15710 24834
rect 15762 24782 16270 24834
rect 16322 24782 16324 24834
rect 15708 24780 16324 24782
rect 15708 24770 15764 24780
rect 16268 24770 16324 24780
rect 16492 24834 16548 24846
rect 16492 24782 16494 24834
rect 16546 24782 16548 24834
rect 15708 24498 15764 24510
rect 15708 24446 15710 24498
rect 15762 24446 15764 24498
rect 15596 24052 15652 24062
rect 15708 24052 15764 24446
rect 15596 24050 15764 24052
rect 15596 23998 15598 24050
rect 15650 23998 15764 24050
rect 15596 23996 15764 23998
rect 16492 24052 16548 24782
rect 15596 23986 15652 23996
rect 16492 23986 16548 23996
rect 16604 24836 16660 25564
rect 16492 23268 16548 23278
rect 15932 22260 15988 22270
rect 15596 22258 15988 22260
rect 15596 22206 15934 22258
rect 15986 22206 15988 22258
rect 15596 22204 15988 22206
rect 15596 21810 15652 22204
rect 15932 22194 15988 22204
rect 16268 22148 16324 22158
rect 15596 21758 15598 21810
rect 15650 21758 15652 21810
rect 15596 21746 15652 21758
rect 16044 22146 16324 22148
rect 16044 22094 16270 22146
rect 16322 22094 16324 22146
rect 16044 22092 16324 22094
rect 15932 21364 15988 21374
rect 15932 21270 15988 21308
rect 16044 20914 16100 22092
rect 16268 22082 16324 22092
rect 16044 20862 16046 20914
rect 16098 20862 16100 20914
rect 16044 20850 16100 20862
rect 16156 21924 16212 21934
rect 16156 21698 16212 21868
rect 16156 21646 16158 21698
rect 16210 21646 16212 21698
rect 16156 20356 16212 21646
rect 16492 20580 16548 23212
rect 16604 21812 16660 24780
rect 16828 23380 16884 23390
rect 16828 23286 16884 23324
rect 16604 21252 16660 21756
rect 16716 21700 16772 21710
rect 16716 21606 16772 21644
rect 16604 21186 16660 21196
rect 15372 20300 15652 20356
rect 14700 20018 14812 20020
rect 14700 19966 14702 20018
rect 14754 19966 14812 20018
rect 14700 19964 14812 19966
rect 14700 19954 14756 19964
rect 14812 19926 14868 19964
rect 15036 20132 15092 20142
rect 14140 19852 14308 19908
rect 14252 19236 14308 19852
rect 14364 19796 14420 19806
rect 14364 19702 14420 19740
rect 13804 19180 14084 19236
rect 14252 19180 14420 19236
rect 13692 19124 13748 19134
rect 13692 19030 13748 19068
rect 13804 19010 13860 19022
rect 13804 18958 13806 19010
rect 13858 18958 13860 19010
rect 13804 18564 13860 18958
rect 13804 18498 13860 18508
rect 13916 19010 13972 19022
rect 13916 18958 13918 19010
rect 13970 18958 13972 19010
rect 13916 18228 13972 18958
rect 13916 18162 13972 18172
rect 14028 18004 14084 19180
rect 14140 19124 14196 19134
rect 14140 19122 14308 19124
rect 14140 19070 14142 19122
rect 14194 19070 14308 19122
rect 14140 19068 14308 19070
rect 14140 19058 14196 19068
rect 13468 15374 13470 15426
rect 13522 15374 13524 15426
rect 13468 15362 13524 15374
rect 13580 17948 14084 18004
rect 13132 15262 13134 15314
rect 13186 15262 13188 15314
rect 13132 15250 13188 15262
rect 12572 14578 12628 14588
rect 12572 14418 12628 14430
rect 13468 14420 13524 14430
rect 12572 14366 12574 14418
rect 12626 14366 12628 14418
rect 12572 13188 12628 14366
rect 13132 14418 13524 14420
rect 13132 14366 13470 14418
rect 13522 14366 13524 14418
rect 13132 14364 13524 14366
rect 13020 13972 13076 13982
rect 13020 13878 13076 13916
rect 13132 13858 13188 14364
rect 13468 14354 13524 14364
rect 13132 13806 13134 13858
rect 13186 13806 13188 13858
rect 13132 13794 13188 13806
rect 12572 13122 12628 13132
rect 13020 13522 13076 13534
rect 13020 13470 13022 13522
rect 13074 13470 13076 13522
rect 12460 12908 12852 12964
rect 12684 12292 12740 12302
rect 12236 12290 12740 12292
rect 12236 12238 12686 12290
rect 12738 12238 12740 12290
rect 12236 12236 12740 12238
rect 11788 12114 11844 12124
rect 12124 12178 12180 12190
rect 12124 12126 12126 12178
rect 12178 12126 12180 12178
rect 11900 12066 11956 12078
rect 11900 12014 11902 12066
rect 11954 12014 11956 12066
rect 11900 11844 11956 12014
rect 11676 11788 11956 11844
rect 11676 11394 11732 11788
rect 11676 11342 11678 11394
rect 11730 11342 11732 11394
rect 11676 11330 11732 11342
rect 11788 11172 11844 11182
rect 11564 11170 11844 11172
rect 11564 11118 11790 11170
rect 11842 11118 11844 11170
rect 11564 11116 11844 11118
rect 9548 10770 9604 10780
rect 10220 10836 10276 10846
rect 9660 10724 9716 10734
rect 9660 10630 9716 10668
rect 8988 10558 8990 10610
rect 9042 10558 9044 10610
rect 8988 10546 9044 10558
rect 9548 10612 9604 10622
rect 9548 10518 9604 10556
rect 8876 9772 9604 9828
rect 8764 9762 8820 9772
rect 8428 9380 8484 9390
rect 8428 9266 8484 9324
rect 8428 9214 8430 9266
rect 8482 9214 8484 9266
rect 8428 9202 8484 9214
rect 9548 9266 9604 9772
rect 10220 9604 10276 10780
rect 10108 9548 10276 9604
rect 10444 10388 10500 10398
rect 9548 9214 9550 9266
rect 9602 9214 9604 9266
rect 9548 9202 9604 9214
rect 9772 9268 9828 9278
rect 9828 9212 9940 9268
rect 9772 9174 9828 9212
rect 7868 8878 7870 8930
rect 7922 8878 7924 8930
rect 7868 8866 7924 8878
rect 8092 8932 8148 8942
rect 6300 8206 6302 8258
rect 6354 8206 6356 8258
rect 6300 8194 6356 8206
rect 7308 8372 7364 8382
rect 7308 8258 7364 8316
rect 7308 8206 7310 8258
rect 7362 8206 7364 8258
rect 7308 8194 7364 8206
rect 7980 8372 8036 8382
rect 5964 8094 5966 8146
rect 6018 8094 6020 8146
rect 5964 8082 6020 8094
rect 7980 7700 8036 8316
rect 8092 8370 8148 8876
rect 8092 8318 8094 8370
rect 8146 8318 8148 8370
rect 8092 8306 8148 8318
rect 8764 8930 8820 8942
rect 8764 8878 8766 8930
rect 8818 8878 8820 8930
rect 8764 8372 8820 8878
rect 9660 8932 9716 8942
rect 9660 8838 9716 8876
rect 9772 8484 9828 8494
rect 8820 8316 9044 8372
rect 8764 8306 8820 8316
rect 8092 7700 8148 7710
rect 7980 7698 8148 7700
rect 7980 7646 8094 7698
rect 8146 7646 8148 7698
rect 7980 7644 8148 7646
rect 8092 7634 8148 7644
rect 8988 7700 9044 8316
rect 8988 7606 9044 7644
rect 9772 7700 9828 8428
rect 9884 8260 9940 9212
rect 10108 8372 10164 9548
rect 10444 9266 10500 10332
rect 10668 9938 10724 11116
rect 11788 11106 11844 11116
rect 11900 11172 11956 11182
rect 11900 11078 11956 11116
rect 12012 11170 12068 11182
rect 12012 11118 12014 11170
rect 12066 11118 12068 11170
rect 11564 10836 11620 10846
rect 11564 10610 11620 10780
rect 11564 10558 11566 10610
rect 11618 10558 11620 10610
rect 11564 10546 11620 10558
rect 11900 10052 11956 10062
rect 12012 10052 12068 11118
rect 12124 10948 12180 12126
rect 12236 12178 12292 12236
rect 12236 12126 12238 12178
rect 12290 12126 12292 12178
rect 12236 12114 12292 12126
rect 12348 11844 12404 11854
rect 12236 11396 12292 11406
rect 12236 11302 12292 11340
rect 12124 10882 12180 10892
rect 11900 10050 12068 10052
rect 11900 9998 11902 10050
rect 11954 9998 12068 10050
rect 11900 9996 12068 9998
rect 12124 10722 12180 10734
rect 12124 10670 12126 10722
rect 12178 10670 12180 10722
rect 11900 9986 11956 9996
rect 10668 9886 10670 9938
rect 10722 9886 10724 9938
rect 10668 9874 10724 9886
rect 11340 9828 11396 9838
rect 10444 9214 10446 9266
rect 10498 9214 10500 9266
rect 10444 9202 10500 9214
rect 11228 9826 11396 9828
rect 11228 9774 11342 9826
rect 11394 9774 11396 9826
rect 11228 9772 11396 9774
rect 10780 9154 10836 9166
rect 10780 9102 10782 9154
rect 10834 9102 10836 9154
rect 10220 9044 10276 9054
rect 10220 9042 10388 9044
rect 10220 8990 10222 9042
rect 10274 8990 10388 9042
rect 10220 8988 10388 8990
rect 10220 8978 10276 8988
rect 10220 8372 10276 8382
rect 10108 8370 10276 8372
rect 10108 8318 10222 8370
rect 10274 8318 10276 8370
rect 10108 8316 10276 8318
rect 9884 8194 9940 8204
rect 10220 8148 10276 8316
rect 10332 8260 10388 8988
rect 10780 8372 10836 9102
rect 10444 8260 10500 8270
rect 10332 8258 10500 8260
rect 10332 8206 10446 8258
rect 10498 8206 10500 8258
rect 10332 8204 10500 8206
rect 10444 8194 10500 8204
rect 10780 8258 10836 8316
rect 11228 8484 11284 9772
rect 11340 9762 11396 9772
rect 11788 9828 11844 9838
rect 12124 9828 12180 10670
rect 11844 9772 12180 9828
rect 12348 9826 12404 11788
rect 12572 11172 12628 11182
rect 12460 11170 12628 11172
rect 12460 11118 12574 11170
rect 12626 11118 12628 11170
rect 12460 11116 12628 11118
rect 12460 11060 12516 11116
rect 12572 11106 12628 11116
rect 12460 10388 12516 11004
rect 12460 10322 12516 10332
rect 12572 10948 12628 10958
rect 12348 9774 12350 9826
rect 12402 9774 12404 9826
rect 11788 9734 11844 9772
rect 12348 9762 12404 9774
rect 12460 9602 12516 9614
rect 12460 9550 12462 9602
rect 12514 9550 12516 9602
rect 12460 8820 12516 9550
rect 12572 9268 12628 10892
rect 12684 10724 12740 12236
rect 12796 11508 12852 12908
rect 13020 12292 13076 13470
rect 13580 13300 13636 17948
rect 13692 17780 13748 17790
rect 13692 17686 13748 17724
rect 14028 17666 14084 17678
rect 14028 17614 14030 17666
rect 14082 17614 14084 17666
rect 13916 17556 13972 17566
rect 13692 15988 13748 15998
rect 13692 15894 13748 15932
rect 13916 15764 13972 17500
rect 14028 16660 14084 17614
rect 14028 16594 14084 16604
rect 13580 13234 13636 13244
rect 13692 15708 13972 15764
rect 14028 15986 14084 15998
rect 14028 15934 14030 15986
rect 14082 15934 14084 15986
rect 13468 13188 13524 13198
rect 13468 13094 13524 13132
rect 13692 12964 13748 15708
rect 14028 15652 14084 15934
rect 14252 15764 14308 19068
rect 14364 17108 14420 19180
rect 14476 19124 14532 19134
rect 14476 19030 14532 19068
rect 14588 19122 14644 19134
rect 14588 19070 14590 19122
rect 14642 19070 14644 19122
rect 14588 18340 14644 19070
rect 15036 18676 15092 20076
rect 15372 20020 15428 20030
rect 15372 19458 15428 19964
rect 15372 19406 15374 19458
rect 15426 19406 15428 19458
rect 15372 19394 15428 19406
rect 15036 18582 15092 18620
rect 15484 19010 15540 19022
rect 15484 18958 15486 19010
rect 15538 18958 15540 19010
rect 15484 18900 15540 18958
rect 15484 18564 15540 18844
rect 15596 18788 15652 20300
rect 16156 20290 16212 20300
rect 16268 20524 16548 20580
rect 16044 19236 16100 19274
rect 16044 19170 16100 19180
rect 15708 19124 15764 19134
rect 15708 19030 15764 19068
rect 15596 18722 15652 18732
rect 16156 19010 16212 19022
rect 16156 18958 16158 19010
rect 16210 18958 16212 19010
rect 16156 18900 16212 18958
rect 15484 18498 15540 18508
rect 15820 18564 15876 18574
rect 14476 18338 14644 18340
rect 14476 18286 14590 18338
rect 14642 18286 14644 18338
rect 14476 18284 14644 18286
rect 14476 17556 14532 18284
rect 14588 18274 14644 18284
rect 14924 18450 14980 18462
rect 14924 18398 14926 18450
rect 14978 18398 14980 18450
rect 14588 17668 14644 17678
rect 14924 17668 14980 18398
rect 15260 18452 15316 18462
rect 15036 18228 15092 18238
rect 15036 18134 15092 18172
rect 15260 17778 15316 18396
rect 15820 18450 15876 18508
rect 15820 18398 15822 18450
rect 15874 18398 15876 18450
rect 15820 18386 15876 18398
rect 15932 18452 15988 18462
rect 15260 17726 15262 17778
rect 15314 17726 15316 17778
rect 15260 17714 15316 17726
rect 14588 17666 14980 17668
rect 14588 17614 14590 17666
rect 14642 17614 14980 17666
rect 14588 17612 14980 17614
rect 15932 17666 15988 18396
rect 16156 18004 16212 18844
rect 16156 17938 16212 17948
rect 15932 17614 15934 17666
rect 15986 17614 15988 17666
rect 14588 17602 14644 17612
rect 15932 17602 15988 17614
rect 16268 17556 16324 20524
rect 16492 19124 16548 19134
rect 16380 19010 16436 19022
rect 16380 18958 16382 19010
rect 16434 18958 16436 19010
rect 16380 18450 16436 18958
rect 16380 18398 16382 18450
rect 16434 18398 16436 18450
rect 16380 18386 16436 18398
rect 16492 18450 16548 19068
rect 16492 18398 16494 18450
rect 16546 18398 16548 18450
rect 16492 18386 16548 18398
rect 16604 18676 16660 18686
rect 16492 17780 16548 17790
rect 16604 17780 16660 18620
rect 16940 18564 16996 26852
rect 17388 24724 17444 26852
rect 17500 26516 17556 28588
rect 18396 28532 18452 29260
rect 19068 29250 19124 29262
rect 19292 30100 19348 30110
rect 18620 29204 18676 29214
rect 18508 28756 18564 28766
rect 18508 28642 18564 28700
rect 18620 28754 18676 29148
rect 18620 28702 18622 28754
rect 18674 28702 18676 28754
rect 18620 28690 18676 28702
rect 19292 28756 19348 30044
rect 19516 29988 19572 29998
rect 19516 29894 19572 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19292 28662 19348 28700
rect 18508 28590 18510 28642
rect 18562 28590 18564 28642
rect 18508 28578 18564 28590
rect 18060 28476 18452 28532
rect 18732 28532 18788 28542
rect 18732 28530 19236 28532
rect 18732 28478 18734 28530
rect 18786 28478 19236 28530
rect 18732 28476 19236 28478
rect 17836 28418 17892 28430
rect 17836 28366 17838 28418
rect 17890 28366 17892 28418
rect 17836 27860 17892 28366
rect 18060 28082 18116 28476
rect 18732 28466 18788 28476
rect 18060 28030 18062 28082
rect 18114 28030 18116 28082
rect 18060 28018 18116 28030
rect 19068 28084 19124 28094
rect 17836 27794 17892 27804
rect 18284 27860 18340 27870
rect 17500 26450 17556 26460
rect 17612 27748 17668 27758
rect 17500 26292 17556 26302
rect 17612 26292 17668 27692
rect 17724 27746 17780 27758
rect 17724 27694 17726 27746
rect 17778 27694 17780 27746
rect 17724 27188 17780 27694
rect 18172 27748 18228 27758
rect 18172 27654 18228 27692
rect 18284 27524 18340 27804
rect 18284 27458 18340 27468
rect 18620 27858 18676 27870
rect 18620 27806 18622 27858
rect 18674 27806 18676 27858
rect 18620 27298 18676 27806
rect 18620 27246 18622 27298
rect 18674 27246 18676 27298
rect 18620 27234 18676 27246
rect 18172 27188 18228 27198
rect 17724 27186 18228 27188
rect 17724 27134 18174 27186
rect 18226 27134 18228 27186
rect 17724 27132 18228 27134
rect 18060 26516 18116 26526
rect 18060 26402 18116 26460
rect 18060 26350 18062 26402
rect 18114 26350 18116 26402
rect 18060 26338 18116 26350
rect 18172 26404 18228 27132
rect 18732 27188 18788 27198
rect 18732 26850 18788 27132
rect 18732 26798 18734 26850
rect 18786 26798 18788 26850
rect 18508 26740 18564 26750
rect 18396 26404 18452 26414
rect 18172 26402 18452 26404
rect 18172 26350 18398 26402
rect 18450 26350 18452 26402
rect 18172 26348 18452 26350
rect 18396 26338 18452 26348
rect 17836 26292 17892 26302
rect 17612 26290 17892 26292
rect 17612 26238 17838 26290
rect 17890 26238 17892 26290
rect 17612 26236 17892 26238
rect 17500 26198 17556 26236
rect 17836 26226 17892 26236
rect 18396 25620 18452 25630
rect 18508 25620 18564 26684
rect 18732 26516 18788 26798
rect 18956 27188 19012 27198
rect 18956 27074 19012 27132
rect 18956 27022 18958 27074
rect 19010 27022 19012 27074
rect 18956 26740 19012 27022
rect 19068 26908 19124 28028
rect 19180 27970 19236 28476
rect 19852 28420 19908 28430
rect 19180 27918 19182 27970
rect 19234 27918 19236 27970
rect 19180 27906 19236 27918
rect 19628 28418 20244 28420
rect 19628 28366 19854 28418
rect 19906 28366 20244 28418
rect 19628 28364 20244 28366
rect 19628 28084 19684 28364
rect 19852 28354 19908 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19628 27858 19684 28028
rect 19628 27806 19630 27858
rect 19682 27806 19684 27858
rect 19628 27794 19684 27806
rect 20076 27748 20132 27758
rect 20076 27654 20132 27692
rect 19740 27300 19796 27310
rect 19292 27298 19796 27300
rect 19292 27246 19742 27298
rect 19794 27246 19796 27298
rect 19292 27244 19796 27246
rect 19292 27074 19348 27244
rect 19740 27234 19796 27244
rect 19852 27300 19908 27310
rect 19292 27022 19294 27074
rect 19346 27022 19348 27074
rect 19292 27010 19348 27022
rect 19628 27076 19684 27086
rect 19628 26962 19684 27020
rect 19628 26910 19630 26962
rect 19682 26910 19684 26962
rect 19068 26852 19236 26908
rect 18956 26674 19012 26684
rect 19068 26516 19124 26526
rect 18732 26514 19124 26516
rect 18732 26462 19070 26514
rect 19122 26462 19124 26514
rect 18732 26460 19124 26462
rect 19068 26450 19124 26460
rect 18452 25564 18564 25620
rect 19068 25620 19124 25630
rect 19180 25620 19236 26852
rect 19068 25618 19236 25620
rect 19068 25566 19070 25618
rect 19122 25566 19236 25618
rect 19068 25564 19236 25566
rect 19292 26290 19348 26302
rect 19292 26238 19294 26290
rect 19346 26238 19348 26290
rect 18396 25526 18452 25564
rect 19068 25554 19124 25564
rect 17612 25508 17668 25518
rect 17500 24724 17556 24734
rect 17388 24722 17556 24724
rect 17388 24670 17502 24722
rect 17554 24670 17556 24722
rect 17388 24668 17556 24670
rect 17500 24658 17556 24668
rect 17388 23380 17444 23390
rect 17388 23286 17444 23324
rect 17612 23154 17668 25452
rect 19292 25508 19348 26238
rect 19516 25732 19572 25742
rect 19628 25732 19684 26910
rect 19852 27074 19908 27244
rect 20188 27298 20244 28364
rect 20188 27246 20190 27298
rect 20242 27246 20244 27298
rect 20188 27234 20244 27246
rect 20300 28418 20356 28430
rect 20300 28366 20302 28418
rect 20354 28366 20356 28418
rect 19852 27022 19854 27074
rect 19906 27022 19908 27074
rect 19852 26908 19908 27022
rect 20188 26964 20244 26974
rect 20300 26964 20356 28366
rect 20412 27076 20468 27086
rect 20412 26982 20468 27020
rect 20244 26908 20356 26964
rect 19852 26852 20244 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19964 26516 20020 26526
rect 20188 26516 20244 26852
rect 19964 26514 20244 26516
rect 19964 26462 19966 26514
rect 20018 26462 20244 26514
rect 19964 26460 20244 26462
rect 19964 26450 20020 26460
rect 20636 26178 20692 34412
rect 20972 34244 21028 34254
rect 20860 32788 20916 32798
rect 20860 32694 20916 32732
rect 20972 26908 21028 34188
rect 21756 33796 21812 37212
rect 21868 37174 21924 37212
rect 21756 33730 21812 33740
rect 21084 33460 21140 33470
rect 21084 32562 21140 33404
rect 21868 33460 21924 33470
rect 21868 33346 21924 33404
rect 21868 33294 21870 33346
rect 21922 33294 21924 33346
rect 21868 33282 21924 33294
rect 21084 32510 21086 32562
rect 21138 32510 21140 32562
rect 21084 32498 21140 32510
rect 21532 31444 21588 31454
rect 21532 31218 21588 31388
rect 21532 31166 21534 31218
rect 21586 31166 21588 31218
rect 21532 30436 21588 31166
rect 21868 30996 21924 31006
rect 21868 30902 21924 30940
rect 21980 30772 22036 39228
rect 22428 38948 22484 38958
rect 22428 38834 22484 38892
rect 22764 38948 22820 40684
rect 22764 38882 22820 38892
rect 22428 38782 22430 38834
rect 22482 38782 22484 38834
rect 22428 38770 22484 38782
rect 22316 38050 22372 38062
rect 22316 37998 22318 38050
rect 22370 37998 22372 38050
rect 22316 37940 22372 37998
rect 22316 37874 22372 37884
rect 22540 37828 22596 37838
rect 22876 37828 22932 43148
rect 23100 42756 23156 42766
rect 23156 42700 23268 42756
rect 23100 42690 23156 42700
rect 22988 42532 23044 42542
rect 22988 42438 23044 42476
rect 23100 42530 23156 42542
rect 23100 42478 23102 42530
rect 23154 42478 23156 42530
rect 22988 41970 23044 41982
rect 22988 41918 22990 41970
rect 23042 41918 23044 41970
rect 22988 41860 23044 41918
rect 22988 41794 23044 41804
rect 23100 41188 23156 42478
rect 23212 42082 23268 42700
rect 23324 42754 23380 43596
rect 23324 42702 23326 42754
rect 23378 42702 23380 42754
rect 23324 42690 23380 42702
rect 23436 43650 23604 43652
rect 23436 43598 23438 43650
rect 23490 43598 23604 43650
rect 23436 43596 23604 43598
rect 23660 43652 24164 43708
rect 24332 43652 24388 43662
rect 23660 43650 23716 43652
rect 23660 43598 23662 43650
rect 23714 43598 23716 43650
rect 23436 42756 23492 43596
rect 23660 43586 23716 43598
rect 24108 43650 24388 43652
rect 24108 43598 24334 43650
rect 24386 43598 24388 43650
rect 24108 43596 24388 43598
rect 23996 43540 24052 43550
rect 23436 42690 23492 42700
rect 23548 43426 23604 43438
rect 23548 43374 23550 43426
rect 23602 43374 23604 43426
rect 23212 42030 23214 42082
rect 23266 42030 23268 42082
rect 23212 42018 23268 42030
rect 23548 42082 23604 43374
rect 23996 43092 24052 43484
rect 23996 43026 24052 43036
rect 23884 42756 23940 42766
rect 23884 42662 23940 42700
rect 23772 42644 23828 42654
rect 23772 42550 23828 42588
rect 23660 42530 23716 42542
rect 23660 42478 23662 42530
rect 23714 42478 23716 42530
rect 23660 42308 23716 42478
rect 24220 42532 24276 43596
rect 24332 43586 24388 43596
rect 24332 42868 24388 42878
rect 24332 42754 24388 42812
rect 24332 42702 24334 42754
rect 24386 42702 24388 42754
rect 24332 42690 24388 42702
rect 24220 42466 24276 42476
rect 23660 42252 23828 42308
rect 23548 42030 23550 42082
rect 23602 42030 23604 42082
rect 23548 42018 23604 42030
rect 23660 42082 23716 42094
rect 23660 42030 23662 42082
rect 23714 42030 23716 42082
rect 23660 41972 23716 42030
rect 23660 41906 23716 41916
rect 23660 41748 23716 41758
rect 23100 41122 23156 41132
rect 23324 41746 23716 41748
rect 23324 41694 23662 41746
rect 23714 41694 23716 41746
rect 23324 41692 23716 41694
rect 23324 41186 23380 41692
rect 23660 41682 23716 41692
rect 23772 41524 23828 42252
rect 23324 41134 23326 41186
rect 23378 41134 23380 41186
rect 23324 41122 23380 41134
rect 23548 41468 23828 41524
rect 24108 41972 24164 41982
rect 24108 41860 24164 41916
rect 24220 41860 24276 41870
rect 24108 41858 24276 41860
rect 24108 41806 24222 41858
rect 24274 41806 24276 41858
rect 24108 41804 24276 41806
rect 23548 41186 23604 41468
rect 23996 41300 24052 41310
rect 23548 41134 23550 41186
rect 23602 41134 23604 41186
rect 23548 41122 23604 41134
rect 23772 41186 23828 41198
rect 23772 41134 23774 41186
rect 23826 41134 23828 41186
rect 23212 41076 23268 41086
rect 23212 40292 23268 41020
rect 23436 40962 23492 40974
rect 23436 40910 23438 40962
rect 23490 40910 23492 40962
rect 23436 40516 23492 40910
rect 23436 40450 23492 40460
rect 23212 40226 23268 40236
rect 23772 39956 23828 41134
rect 23996 41186 24052 41244
rect 23996 41134 23998 41186
rect 24050 41134 24052 41186
rect 23996 40404 24052 41134
rect 24108 41076 24164 41804
rect 24220 41794 24276 41804
rect 24444 41636 24500 45164
rect 25004 44660 25060 56590
rect 25564 55468 25620 59200
rect 27356 56084 27412 56094
rect 27132 56082 27412 56084
rect 27132 56030 27358 56082
rect 27410 56030 27412 56082
rect 27132 56028 27412 56030
rect 26796 55858 26852 55870
rect 26796 55806 26798 55858
rect 26850 55806 26852 55858
rect 25564 55412 25844 55468
rect 25676 54740 25732 54750
rect 25228 54684 25620 54740
rect 25228 53732 25284 54684
rect 25564 54626 25620 54684
rect 25676 54646 25732 54684
rect 25564 54574 25566 54626
rect 25618 54574 25620 54626
rect 25564 54562 25620 54574
rect 25116 53676 25284 53732
rect 25452 54514 25508 54526
rect 25452 54462 25454 54514
rect 25506 54462 25508 54514
rect 25116 52612 25172 53676
rect 25340 53620 25396 53630
rect 25116 52546 25172 52556
rect 25228 53284 25284 53294
rect 25228 52388 25284 53228
rect 25340 53170 25396 53564
rect 25340 53118 25342 53170
rect 25394 53118 25396 53170
rect 25340 53106 25396 53118
rect 25452 52946 25508 54462
rect 25676 53060 25732 53098
rect 25676 52994 25732 53004
rect 25452 52894 25454 52946
rect 25506 52894 25508 52946
rect 25228 52162 25284 52332
rect 25340 52834 25396 52846
rect 25340 52782 25342 52834
rect 25394 52782 25396 52834
rect 25340 52276 25396 52782
rect 25452 52724 25508 52894
rect 25452 52658 25508 52668
rect 25788 52388 25844 55412
rect 26348 55410 26404 55422
rect 26348 55358 26350 55410
rect 26402 55358 26404 55410
rect 25900 53508 25956 53518
rect 25900 53058 25956 53452
rect 25900 53006 25902 53058
rect 25954 53006 25956 53058
rect 25900 52994 25956 53006
rect 26348 52612 26404 55358
rect 26796 55412 26852 55806
rect 26796 55346 26852 55356
rect 27020 54626 27076 54638
rect 27020 54574 27022 54626
rect 27074 54574 27076 54626
rect 26572 54516 26628 54526
rect 26572 54514 26740 54516
rect 26572 54462 26574 54514
rect 26626 54462 26740 54514
rect 26572 54460 26740 54462
rect 26572 54450 26628 54460
rect 26572 53842 26628 53854
rect 26572 53790 26574 53842
rect 26626 53790 26628 53842
rect 26572 52724 26628 53790
rect 26684 53508 26740 54460
rect 27020 53732 27076 54574
rect 27020 53666 27076 53676
rect 26684 53442 26740 53452
rect 26572 52658 26628 52668
rect 26908 53172 26964 53182
rect 26908 52946 26964 53116
rect 26908 52894 26910 52946
rect 26962 52894 26964 52946
rect 26348 52546 26404 52556
rect 25788 52322 25844 52332
rect 26796 52388 26852 52398
rect 26796 52294 26852 52332
rect 25340 52210 25396 52220
rect 25228 52110 25230 52162
rect 25282 52110 25284 52162
rect 25228 52098 25284 52110
rect 25452 52164 25508 52174
rect 26236 52164 26292 52174
rect 25508 52108 25620 52164
rect 25452 52098 25508 52108
rect 25452 51938 25508 51950
rect 25452 51886 25454 51938
rect 25506 51886 25508 51938
rect 25340 50482 25396 50494
rect 25340 50430 25342 50482
rect 25394 50430 25396 50482
rect 25340 50034 25396 50430
rect 25340 49982 25342 50034
rect 25394 49982 25396 50034
rect 25340 49970 25396 49982
rect 25452 50260 25508 51886
rect 25452 49812 25508 50204
rect 25452 49746 25508 49756
rect 25228 49700 25284 49710
rect 25228 49606 25284 49644
rect 25452 48468 25508 48478
rect 25564 48468 25620 52108
rect 26236 52070 26292 52108
rect 25676 52052 25732 52062
rect 25676 51378 25732 51996
rect 26908 52052 26964 52894
rect 26908 51986 26964 51996
rect 27020 52164 27076 52174
rect 25676 51326 25678 51378
rect 25730 51326 25732 51378
rect 25676 51314 25732 51326
rect 26348 51268 26404 51278
rect 26796 51268 26852 51278
rect 26236 51266 26404 51268
rect 26236 51214 26350 51266
rect 26402 51214 26404 51266
rect 26236 51212 26404 51214
rect 26236 50148 26292 51212
rect 26348 51202 26404 51212
rect 26684 51212 26796 51268
rect 25788 50092 26292 50148
rect 25788 49810 25844 50092
rect 26460 50036 26516 50046
rect 25788 49758 25790 49810
rect 25842 49758 25844 49810
rect 25788 49746 25844 49758
rect 25900 50034 26516 50036
rect 25900 49982 26462 50034
rect 26514 49982 26516 50034
rect 25900 49980 26516 49982
rect 25676 49698 25732 49710
rect 25676 49646 25678 49698
rect 25730 49646 25732 49698
rect 25676 49588 25732 49646
rect 25900 49588 25956 49980
rect 26460 49970 26516 49980
rect 26572 49924 26628 49934
rect 26572 49830 26628 49868
rect 26124 49812 26180 49822
rect 26124 49718 26180 49756
rect 26348 49810 26404 49822
rect 26348 49758 26350 49810
rect 26402 49758 26404 49810
rect 25676 49532 25956 49588
rect 26348 49588 26404 49758
rect 26684 49588 26740 51212
rect 26796 51202 26852 51212
rect 27020 50428 27076 52108
rect 26908 50372 27076 50428
rect 26348 49532 26740 49588
rect 26796 50148 26852 50158
rect 26796 49810 26852 50092
rect 26796 49758 26798 49810
rect 26850 49758 26852 49810
rect 25788 49140 25844 49150
rect 25564 48412 25732 48468
rect 25452 48374 25508 48412
rect 25004 44594 25060 44604
rect 25116 48244 25172 48254
rect 24556 44546 24612 44558
rect 24556 44494 24558 44546
rect 24610 44494 24612 44546
rect 24556 44434 24612 44494
rect 24556 44382 24558 44434
rect 24610 44382 24612 44434
rect 24556 43652 24612 44382
rect 25004 44436 25060 44446
rect 25004 44342 25060 44380
rect 25116 43708 25172 48188
rect 25228 48242 25284 48254
rect 25228 48190 25230 48242
rect 25282 48190 25284 48242
rect 25228 47908 25284 48190
rect 25564 48242 25620 48254
rect 25564 48190 25566 48242
rect 25618 48190 25620 48242
rect 25564 48132 25620 48190
rect 25340 47908 25396 47918
rect 25228 47852 25340 47908
rect 25340 47842 25396 47852
rect 25564 47796 25620 48076
rect 25564 47730 25620 47740
rect 25676 47460 25732 48412
rect 25340 47346 25396 47358
rect 25340 47294 25342 47346
rect 25394 47294 25396 47346
rect 25340 46900 25396 47294
rect 25340 46834 25396 46844
rect 25676 46674 25732 47404
rect 25676 46622 25678 46674
rect 25730 46622 25732 46674
rect 25676 46610 25732 46622
rect 25788 48354 25844 49084
rect 26796 48916 26852 49758
rect 25788 48302 25790 48354
rect 25842 48302 25844 48354
rect 25340 46562 25396 46574
rect 25340 46510 25342 46562
rect 25394 46510 25396 46562
rect 25340 45556 25396 46510
rect 25340 45490 25396 45500
rect 25340 45332 25396 45342
rect 25340 45238 25396 45276
rect 24556 43586 24612 43596
rect 25004 43652 25172 43708
rect 25228 45220 25284 45230
rect 25788 45220 25844 48302
rect 26684 48860 26852 48916
rect 26572 47908 26628 47918
rect 26460 47460 26516 47470
rect 26236 47236 26292 47246
rect 26236 46786 26292 47180
rect 26348 47234 26404 47246
rect 26348 47182 26350 47234
rect 26402 47182 26404 47234
rect 26348 47012 26404 47182
rect 26348 46946 26404 46956
rect 26236 46734 26238 46786
rect 26290 46734 26292 46786
rect 26236 46722 26292 46734
rect 26460 46564 26516 47404
rect 26348 46508 26516 46564
rect 26572 46674 26628 47852
rect 26684 47460 26740 48860
rect 26796 48468 26852 48478
rect 26796 47682 26852 48412
rect 26908 48244 26964 50372
rect 27020 49140 27076 49150
rect 27020 49046 27076 49084
rect 26908 48178 26964 48188
rect 27132 48132 27188 56028
rect 27356 56018 27412 56028
rect 27580 55300 27636 59200
rect 28924 55860 28980 59200
rect 29484 56084 29540 56094
rect 29484 55990 29540 56028
rect 28924 55804 29540 55860
rect 27580 55234 27636 55244
rect 28476 55188 28532 55198
rect 28476 55094 28532 55132
rect 29260 55188 29316 55198
rect 28364 55074 28420 55086
rect 28364 55022 28366 55074
rect 28418 55022 28420 55074
rect 28364 54626 28420 55022
rect 28364 54574 28366 54626
rect 28418 54574 28420 54626
rect 28364 54562 28420 54574
rect 27692 54516 27748 54526
rect 27692 54514 28084 54516
rect 27692 54462 27694 54514
rect 27746 54462 28084 54514
rect 27692 54460 28084 54462
rect 27692 54450 27748 54460
rect 27244 53900 27860 53956
rect 27244 53842 27300 53900
rect 27244 53790 27246 53842
rect 27298 53790 27300 53842
rect 27244 53778 27300 53790
rect 27804 53842 27860 53900
rect 27804 53790 27806 53842
rect 27858 53790 27860 53842
rect 27804 53778 27860 53790
rect 27804 53620 27860 53630
rect 27804 53526 27860 53564
rect 27356 53508 27412 53518
rect 27916 53508 27972 53518
rect 27356 53506 27636 53508
rect 27356 53454 27358 53506
rect 27410 53454 27636 53506
rect 27356 53452 27636 53454
rect 27356 53442 27412 53452
rect 27580 53058 27636 53452
rect 27916 53414 27972 53452
rect 28028 53172 28084 54460
rect 29260 53842 29316 55132
rect 29260 53790 29262 53842
rect 29314 53790 29316 53842
rect 29260 53778 29316 53790
rect 28364 53732 28420 53742
rect 28364 53638 28420 53676
rect 29148 53730 29204 53742
rect 29148 53678 29150 53730
rect 29202 53678 29204 53730
rect 29148 53620 29204 53678
rect 29372 53732 29428 53742
rect 29372 53638 29428 53676
rect 29148 53554 29204 53564
rect 29484 53620 29540 55804
rect 29596 55412 29652 59200
rect 29596 55346 29652 55356
rect 29820 54292 29876 54302
rect 29820 53730 29876 54236
rect 29820 53678 29822 53730
rect 29874 53678 29876 53730
rect 29820 53666 29876 53678
rect 29484 53554 29540 53564
rect 28140 53506 28196 53518
rect 28140 53454 28142 53506
rect 28194 53454 28196 53506
rect 28140 53284 28196 53454
rect 28140 53218 28196 53228
rect 29596 53506 29652 53518
rect 29596 53454 29598 53506
rect 29650 53454 29652 53506
rect 29596 53284 29652 53454
rect 28028 53106 28084 53116
rect 27580 53006 27582 53058
rect 27634 53006 27636 53058
rect 27580 52994 27636 53006
rect 29596 52836 29652 53228
rect 29596 52770 29652 52780
rect 29708 53508 29764 53518
rect 29708 52836 29764 53452
rect 30156 53172 30212 53182
rect 29932 53116 30156 53172
rect 29708 52834 29876 52836
rect 29708 52782 29710 52834
rect 29762 52782 29876 52834
rect 29708 52780 29876 52782
rect 29708 52770 29764 52780
rect 29260 52724 29316 52734
rect 28812 52500 28868 52510
rect 28364 51492 28420 51502
rect 27580 50708 27636 50718
rect 27580 50428 27636 50652
rect 27356 50372 27636 50428
rect 28364 50596 28420 51436
rect 28588 51268 28644 51278
rect 28588 51174 28644 51212
rect 28364 50482 28420 50540
rect 28364 50430 28366 50482
rect 28418 50430 28420 50482
rect 28364 50418 28420 50430
rect 28476 50484 28532 50522
rect 28476 50418 28532 50428
rect 28588 50482 28644 50494
rect 28588 50430 28590 50482
rect 28642 50430 28644 50482
rect 28588 50428 28644 50430
rect 28588 50372 28756 50428
rect 27244 50260 27300 50270
rect 27244 50034 27300 50204
rect 27244 49982 27246 50034
rect 27298 49982 27300 50034
rect 27244 49970 27300 49982
rect 27356 50148 27412 50372
rect 27356 50034 27412 50092
rect 27356 49982 27358 50034
rect 27410 49982 27412 50034
rect 27356 49970 27412 49982
rect 27580 49924 27636 49934
rect 27468 49700 27524 49710
rect 27468 49606 27524 49644
rect 27580 49138 27636 49868
rect 27580 49086 27582 49138
rect 27634 49086 27636 49138
rect 27580 49074 27636 49086
rect 27692 49810 27748 49822
rect 27692 49758 27694 49810
rect 27746 49758 27748 49810
rect 27692 49700 27748 49758
rect 28252 49700 28308 49710
rect 27692 49698 28308 49700
rect 27692 49646 28254 49698
rect 28306 49646 28308 49698
rect 27692 49644 28308 49646
rect 27244 48132 27300 48142
rect 27132 48130 27300 48132
rect 27132 48078 27246 48130
rect 27298 48078 27300 48130
rect 27132 48076 27300 48078
rect 27244 48066 27300 48076
rect 27580 48132 27636 48142
rect 27692 48132 27748 49644
rect 28252 49634 28308 49644
rect 28700 49588 28756 50372
rect 28812 49812 28868 52444
rect 29148 51604 29204 51614
rect 29148 50594 29204 51548
rect 29260 51268 29316 52668
rect 29484 52612 29540 52622
rect 29372 52500 29428 52510
rect 29372 52162 29428 52444
rect 29372 52110 29374 52162
rect 29426 52110 29428 52162
rect 29372 52098 29428 52110
rect 29260 51212 29428 51268
rect 29148 50542 29150 50594
rect 29202 50542 29204 50594
rect 29148 50428 29204 50542
rect 29148 50372 29316 50428
rect 29260 50036 29316 50372
rect 29260 49970 29316 49980
rect 28812 49718 28868 49756
rect 29260 49812 29316 49822
rect 29372 49812 29428 51212
rect 29484 50428 29540 52556
rect 29708 52276 29764 52286
rect 29596 52220 29708 52276
rect 29596 52162 29652 52220
rect 29708 52210 29764 52220
rect 29596 52110 29598 52162
rect 29650 52110 29652 52162
rect 29596 52098 29652 52110
rect 29820 52162 29876 52780
rect 29820 52110 29822 52162
rect 29874 52110 29876 52162
rect 29820 52098 29876 52110
rect 29932 51940 29988 53116
rect 30156 53078 30212 53116
rect 30268 52388 30324 59200
rect 30604 56084 30660 56094
rect 30492 54402 30548 54414
rect 30492 54350 30494 54402
rect 30546 54350 30548 54402
rect 30492 53732 30548 54350
rect 30492 53060 30548 53676
rect 30604 53508 30660 56028
rect 30940 55970 30996 59200
rect 31612 56308 31668 59200
rect 31612 56242 31668 56252
rect 30940 55918 30942 55970
rect 30994 55918 30996 55970
rect 30940 55906 30996 55918
rect 30940 55298 30996 55310
rect 30940 55246 30942 55298
rect 30994 55246 30996 55298
rect 30940 54402 30996 55246
rect 31612 55186 31668 55198
rect 31612 55134 31614 55186
rect 31666 55134 31668 55186
rect 31388 54740 31444 54750
rect 30940 54350 30942 54402
rect 30994 54350 30996 54402
rect 30716 53732 30772 53742
rect 30940 53732 30996 54350
rect 30716 53730 30996 53732
rect 30716 53678 30718 53730
rect 30770 53678 30996 53730
rect 30716 53676 30996 53678
rect 30716 53666 30772 53676
rect 30604 53452 30884 53508
rect 30492 52994 30548 53004
rect 30716 53284 30772 53294
rect 30716 53170 30772 53228
rect 30716 53118 30718 53170
rect 30770 53118 30772 53170
rect 30604 52834 30660 52846
rect 30604 52782 30606 52834
rect 30658 52782 30660 52834
rect 30268 52322 30324 52332
rect 30492 52722 30548 52734
rect 30492 52670 30494 52722
rect 30546 52670 30548 52722
rect 30492 52276 30548 52670
rect 30492 52210 30548 52220
rect 30380 52164 30436 52174
rect 30268 52162 30436 52164
rect 30268 52110 30382 52162
rect 30434 52110 30436 52162
rect 30268 52108 30436 52110
rect 30044 52052 30100 52062
rect 30044 51958 30100 51996
rect 29708 51884 29988 51940
rect 29708 51604 29764 51884
rect 29708 51378 29764 51548
rect 29708 51326 29710 51378
rect 29762 51326 29764 51378
rect 29708 51314 29764 51326
rect 30268 50596 30324 52108
rect 30380 52098 30436 52108
rect 30380 51492 30436 51502
rect 30604 51492 30660 52782
rect 30380 51490 30660 51492
rect 30380 51438 30382 51490
rect 30434 51438 30660 51490
rect 30380 51436 30660 51438
rect 30380 51426 30436 51436
rect 30156 50540 30324 50596
rect 30716 50596 30772 53118
rect 29932 50484 29988 50522
rect 29484 50372 29652 50428
rect 29932 50418 29988 50428
rect 29484 49924 29540 49934
rect 29484 49830 29540 49868
rect 29260 49810 29428 49812
rect 29260 49758 29262 49810
rect 29314 49758 29428 49810
rect 29260 49756 29428 49758
rect 29260 49746 29316 49756
rect 29036 49698 29092 49710
rect 29036 49646 29038 49698
rect 29090 49646 29092 49698
rect 29036 49588 29092 49646
rect 28700 49532 29092 49588
rect 28588 49140 28644 49150
rect 27636 48076 27748 48132
rect 27804 48132 27860 48142
rect 27580 48066 27636 48076
rect 26796 47630 26798 47682
rect 26850 47630 26852 47682
rect 26796 47618 26852 47630
rect 26908 48020 26964 48030
rect 26908 47570 26964 47964
rect 26908 47518 26910 47570
rect 26962 47518 26964 47570
rect 26908 47506 26964 47518
rect 27804 47570 27860 48076
rect 27804 47518 27806 47570
rect 27858 47518 27860 47570
rect 27804 47506 27860 47518
rect 27020 47460 27076 47470
rect 26684 47404 26852 47460
rect 26572 46622 26574 46674
rect 26626 46622 26628 46674
rect 24556 43428 24612 43438
rect 24556 42756 24612 43372
rect 24556 42662 24612 42700
rect 24780 42532 24836 42542
rect 24780 42438 24836 42476
rect 24892 42530 24948 42542
rect 24892 42478 24894 42530
rect 24946 42478 24948 42530
rect 24668 41860 24724 41870
rect 24668 41766 24724 41804
rect 24108 41010 24164 41020
rect 24220 41580 24500 41636
rect 23996 40338 24052 40348
rect 23772 39890 23828 39900
rect 24108 40180 24164 40190
rect 23772 38164 23828 38174
rect 23772 38070 23828 38108
rect 23212 37828 23268 37838
rect 22540 37826 23268 37828
rect 22540 37774 22542 37826
rect 22594 37774 23214 37826
rect 23266 37774 23268 37826
rect 22540 37772 23268 37774
rect 22316 37268 22372 37278
rect 22316 37174 22372 37212
rect 22204 36484 22260 36494
rect 22540 36484 22596 37772
rect 23212 37762 23268 37772
rect 23436 37436 23716 37492
rect 23100 37156 23156 37166
rect 23100 36706 23156 37100
rect 23100 36654 23102 36706
rect 23154 36654 23156 36706
rect 23100 36642 23156 36654
rect 22204 36482 22596 36484
rect 22204 36430 22206 36482
rect 22258 36430 22596 36482
rect 22204 36428 22596 36430
rect 23100 36484 23156 36494
rect 23436 36484 23492 37436
rect 23100 36482 23492 36484
rect 23100 36430 23102 36482
rect 23154 36430 23492 36482
rect 23100 36428 23492 36430
rect 23548 37268 23604 37278
rect 23548 36706 23604 37212
rect 23660 37266 23716 37436
rect 23660 37214 23662 37266
rect 23714 37214 23716 37266
rect 23660 37202 23716 37214
rect 23548 36654 23550 36706
rect 23602 36654 23604 36706
rect 22204 36418 22260 36428
rect 22652 36370 22708 36382
rect 22652 36318 22654 36370
rect 22706 36318 22708 36370
rect 22652 35364 22708 36318
rect 22988 36370 23044 36382
rect 22988 36318 22990 36370
rect 23042 36318 23044 36370
rect 22988 36260 23044 36318
rect 22988 36194 23044 36204
rect 23100 36036 23156 36428
rect 22652 35298 22708 35308
rect 22988 35980 23156 36036
rect 23324 36148 23380 36158
rect 22988 35140 23044 35980
rect 23324 35922 23380 36092
rect 23324 35870 23326 35922
rect 23378 35870 23380 35922
rect 23324 35858 23380 35870
rect 22092 35138 23044 35140
rect 22092 35086 22990 35138
rect 23042 35086 23044 35138
rect 22092 35084 23044 35086
rect 22092 31108 22148 35084
rect 22988 35074 23044 35084
rect 23436 35588 23492 35598
rect 23436 35138 23492 35532
rect 23548 35476 23604 36654
rect 23996 37154 24052 37166
rect 23996 37102 23998 37154
rect 24050 37102 24052 37154
rect 23772 36484 23828 36494
rect 23660 36482 23828 36484
rect 23660 36430 23774 36482
rect 23826 36430 23828 36482
rect 23660 36428 23828 36430
rect 23660 35700 23716 36428
rect 23772 36418 23828 36428
rect 23772 35924 23828 35934
rect 23996 35924 24052 37102
rect 23772 35922 24052 35924
rect 23772 35870 23774 35922
rect 23826 35870 24052 35922
rect 23772 35868 24052 35870
rect 24108 35924 24164 40124
rect 24220 39730 24276 41580
rect 24892 41412 24948 42478
rect 25004 42532 25060 43652
rect 25116 42756 25172 42766
rect 25116 42662 25172 42700
rect 25004 42476 25172 42532
rect 24892 41346 24948 41356
rect 24332 41188 24388 41198
rect 24332 41094 24388 41132
rect 24444 41076 24500 41086
rect 24668 41076 24724 41086
rect 24444 40964 24500 41020
rect 24332 40962 24500 40964
rect 24332 40910 24446 40962
rect 24498 40910 24500 40962
rect 24332 40908 24500 40910
rect 24332 40068 24388 40908
rect 24444 40898 24500 40908
rect 24556 41074 24724 41076
rect 24556 41022 24670 41074
rect 24722 41022 24724 41074
rect 24556 41020 24724 41022
rect 24556 40964 24612 41020
rect 24668 41010 24724 41020
rect 25004 41076 25060 41086
rect 25004 40982 25060 41020
rect 24556 40898 24612 40908
rect 25116 40740 25172 42476
rect 24668 40684 25172 40740
rect 24332 40002 24388 40012
rect 24444 40628 24500 40638
rect 24220 39678 24222 39730
rect 24274 39678 24276 39730
rect 24220 39666 24276 39678
rect 24332 39396 24388 39406
rect 24332 37378 24388 39340
rect 24332 37326 24334 37378
rect 24386 37326 24388 37378
rect 24332 37314 24388 37326
rect 24444 39058 24500 40572
rect 24668 40290 24724 40684
rect 25228 40628 25284 45164
rect 25564 45164 25844 45220
rect 26012 46002 26068 46014
rect 26012 45950 26014 46002
rect 26066 45950 26068 46002
rect 25564 44548 25620 45164
rect 26012 45106 26068 45950
rect 26348 45890 26404 46508
rect 26460 46004 26516 46014
rect 26460 45910 26516 45948
rect 26348 45838 26350 45890
rect 26402 45838 26404 45890
rect 26348 45826 26404 45838
rect 26236 45218 26292 45230
rect 26236 45166 26238 45218
rect 26290 45166 26292 45218
rect 26236 45108 26292 45166
rect 26012 45054 26014 45106
rect 26066 45054 26068 45106
rect 26012 44996 26068 45054
rect 25564 44482 25620 44492
rect 25676 44940 26068 44996
rect 26124 45052 26236 45108
rect 25676 44434 25732 44940
rect 26124 44772 26180 45052
rect 26236 45042 26292 45052
rect 26460 44884 26516 44894
rect 26572 44884 26628 46622
rect 26796 46674 26852 47404
rect 27020 47346 27076 47404
rect 27020 47294 27022 47346
rect 27074 47294 27076 47346
rect 27020 47282 27076 47294
rect 28364 47458 28420 47470
rect 28364 47406 28366 47458
rect 28418 47406 28420 47458
rect 27692 47236 27748 47246
rect 27692 47142 27748 47180
rect 27916 47236 27972 47246
rect 27804 47124 27860 47134
rect 26796 46622 26798 46674
rect 26850 46622 26852 46674
rect 26796 46610 26852 46622
rect 27020 46674 27076 46686
rect 27020 46622 27022 46674
rect 27074 46622 27076 46674
rect 26684 46562 26740 46574
rect 26684 46510 26686 46562
rect 26738 46510 26740 46562
rect 26684 46114 26740 46510
rect 26684 46062 26686 46114
rect 26738 46062 26740 46114
rect 26684 46050 26740 46062
rect 27020 45330 27076 46622
rect 27580 46676 27636 46686
rect 27580 46582 27636 46620
rect 27804 46452 27860 47068
rect 27580 46396 27860 46452
rect 27020 45278 27022 45330
rect 27074 45278 27076 45330
rect 26516 44828 26628 44884
rect 26796 45106 26852 45118
rect 26796 45054 26798 45106
rect 26850 45054 26852 45106
rect 26460 44818 26516 44828
rect 26012 44716 26180 44772
rect 25676 44382 25678 44434
rect 25730 44382 25732 44434
rect 25676 44370 25732 44382
rect 25900 44548 25956 44558
rect 25900 44324 25956 44492
rect 25900 44258 25956 44268
rect 25676 43652 25732 43662
rect 25676 42868 25732 43596
rect 25788 43538 25844 43550
rect 25788 43486 25790 43538
rect 25842 43486 25844 43538
rect 25788 42980 25844 43486
rect 25788 42914 25844 42924
rect 25676 42754 25732 42812
rect 25676 42702 25678 42754
rect 25730 42702 25732 42754
rect 25676 42690 25732 42702
rect 26012 42756 26068 44716
rect 26124 44548 26180 44558
rect 26124 44322 26180 44492
rect 26796 44548 26852 45054
rect 27020 45108 27076 45278
rect 27132 45666 27188 45678
rect 27132 45614 27134 45666
rect 27186 45614 27188 45666
rect 27132 45220 27188 45614
rect 27132 45154 27188 45164
rect 27020 45042 27076 45052
rect 27468 45106 27524 45118
rect 27468 45054 27470 45106
rect 27522 45054 27524 45106
rect 26908 44994 26964 45006
rect 26908 44942 26910 44994
rect 26962 44942 26964 44994
rect 26908 44660 26964 44942
rect 26908 44604 27300 44660
rect 26796 44482 26852 44492
rect 27244 44434 27300 44604
rect 27244 44382 27246 44434
rect 27298 44382 27300 44434
rect 27244 44370 27300 44382
rect 26124 44270 26126 44322
rect 26178 44270 26180 44322
rect 26124 42868 26180 44270
rect 27132 44324 27188 44334
rect 27132 44230 27188 44268
rect 26572 44098 26628 44110
rect 26572 44046 26574 44098
rect 26626 44046 26628 44098
rect 26572 43652 26628 44046
rect 27468 43764 27524 45054
rect 27468 43670 27524 43708
rect 26572 43586 26628 43596
rect 27020 43652 27076 43662
rect 27020 43558 27076 43596
rect 27244 43538 27300 43550
rect 27244 43486 27246 43538
rect 27298 43486 27300 43538
rect 26460 43428 26516 43438
rect 26460 43334 26516 43372
rect 27132 43428 27188 43438
rect 27132 43334 27188 43372
rect 26572 43316 26628 43326
rect 26572 43222 26628 43260
rect 26124 42812 26740 42868
rect 26012 42700 26404 42756
rect 25340 42644 25396 42654
rect 25340 42550 25396 42588
rect 25564 42530 25620 42542
rect 25564 42478 25566 42530
rect 25618 42478 25620 42530
rect 25340 40628 25396 40638
rect 25284 40626 25396 40628
rect 25284 40574 25342 40626
rect 25394 40574 25396 40626
rect 25284 40572 25396 40574
rect 25228 40562 25284 40572
rect 25340 40562 25396 40572
rect 24668 40238 24670 40290
rect 24722 40238 24724 40290
rect 24668 40226 24724 40238
rect 24780 40516 24836 40526
rect 24780 39730 24836 40460
rect 24780 39678 24782 39730
rect 24834 39678 24836 39730
rect 24780 39666 24836 39678
rect 25228 40404 25284 40414
rect 24444 39006 24446 39058
rect 24498 39006 24500 39058
rect 24332 36482 24388 36494
rect 24332 36430 24334 36482
rect 24386 36430 24388 36482
rect 24332 36148 24388 36430
rect 24332 36082 24388 36092
rect 23772 35858 23828 35868
rect 24108 35830 24164 35868
rect 23660 35606 23716 35644
rect 23884 35698 23940 35710
rect 23884 35646 23886 35698
rect 23938 35646 23940 35698
rect 23884 35476 23940 35646
rect 23548 35420 23940 35476
rect 23436 35086 23438 35138
rect 23490 35086 23492 35138
rect 23436 35074 23492 35086
rect 23548 35252 23604 35262
rect 22204 34914 22260 34926
rect 22204 34862 22206 34914
rect 22258 34862 22260 34914
rect 22204 34020 22260 34862
rect 23212 34916 23268 34926
rect 22764 34802 22820 34814
rect 22764 34750 22766 34802
rect 22818 34750 22820 34802
rect 22428 34692 22484 34702
rect 22316 34020 22372 34030
rect 22204 34018 22372 34020
rect 22204 33966 22318 34018
rect 22370 33966 22372 34018
rect 22204 33964 22372 33966
rect 22316 33346 22372 33964
rect 22316 33294 22318 33346
rect 22370 33294 22372 33346
rect 22316 33282 22372 33294
rect 22428 33124 22484 34636
rect 22764 33796 22820 34750
rect 22876 34804 22932 34814
rect 22876 34354 22932 34748
rect 23212 34692 23268 34860
rect 23212 34626 23268 34636
rect 22876 34302 22878 34354
rect 22930 34302 22932 34354
rect 22876 34290 22932 34302
rect 23548 34244 23604 35196
rect 23436 34242 23604 34244
rect 23436 34190 23550 34242
rect 23602 34190 23604 34242
rect 23436 34188 23604 34190
rect 22764 33730 22820 33740
rect 23212 33906 23268 33918
rect 23212 33854 23214 33906
rect 23266 33854 23268 33906
rect 22988 33348 23044 33358
rect 22988 33254 23044 33292
rect 22540 33236 22596 33246
rect 22540 33142 22596 33180
rect 22316 33068 22484 33124
rect 22316 31220 22372 33068
rect 22540 32788 22596 32798
rect 22540 31890 22596 32732
rect 23212 32116 23268 33854
rect 23212 32050 23268 32060
rect 22540 31838 22542 31890
rect 22594 31838 22596 31890
rect 22540 31826 22596 31838
rect 22764 31836 23268 31892
rect 22652 31780 22708 31790
rect 22764 31780 22820 31836
rect 22652 31778 22820 31780
rect 22652 31726 22654 31778
rect 22706 31726 22820 31778
rect 22652 31724 22820 31726
rect 23212 31778 23268 31836
rect 23212 31726 23214 31778
rect 23266 31726 23268 31778
rect 22652 31714 22708 31724
rect 23212 31714 23268 31726
rect 22876 31668 22932 31678
rect 22540 31332 22596 31342
rect 22316 31154 22372 31164
rect 22428 31276 22540 31332
rect 22204 31108 22260 31118
rect 22092 31106 22260 31108
rect 22092 31054 22206 31106
rect 22258 31054 22260 31106
rect 22092 31052 22260 31054
rect 21868 30716 22036 30772
rect 21532 30370 21588 30380
rect 21756 30548 21812 30558
rect 21644 30098 21700 30110
rect 21644 30046 21646 30098
rect 21698 30046 21700 30098
rect 21308 29988 21364 29998
rect 21196 29986 21364 29988
rect 21196 29934 21310 29986
rect 21362 29934 21364 29986
rect 21196 29932 21364 29934
rect 21196 29538 21252 29932
rect 21308 29922 21364 29932
rect 21644 29652 21700 30046
rect 21644 29586 21700 29596
rect 21196 29486 21198 29538
rect 21250 29486 21252 29538
rect 21196 29474 21252 29486
rect 20636 26126 20638 26178
rect 20690 26126 20692 26178
rect 20636 25956 20692 26126
rect 20636 25890 20692 25900
rect 20860 26852 21028 26908
rect 21084 27858 21140 27870
rect 21084 27806 21086 27858
rect 21138 27806 21140 27858
rect 21084 26964 21140 27806
rect 21644 27860 21700 27870
rect 21644 27766 21700 27804
rect 19516 25730 19684 25732
rect 19516 25678 19518 25730
rect 19570 25678 19684 25730
rect 19516 25676 19684 25678
rect 19516 25666 19572 25676
rect 19404 25508 19460 25518
rect 19292 25506 19404 25508
rect 19292 25454 19294 25506
rect 19346 25454 19404 25506
rect 19292 25452 19404 25454
rect 19292 25442 19348 25452
rect 17948 25284 18004 25294
rect 17948 25190 18004 25228
rect 19292 25284 19348 25294
rect 18732 25060 18788 25070
rect 18732 24946 18788 25004
rect 18732 24894 18734 24946
rect 18786 24894 18788 24946
rect 18732 24882 18788 24894
rect 19068 24836 19124 24846
rect 18060 24722 18116 24734
rect 18060 24670 18062 24722
rect 18114 24670 18116 24722
rect 17724 24052 17780 24062
rect 17780 23996 17892 24052
rect 17724 23958 17780 23996
rect 17612 23102 17614 23154
rect 17666 23102 17668 23154
rect 17052 22594 17108 22606
rect 17052 22542 17054 22594
rect 17106 22542 17108 22594
rect 17052 22482 17108 22542
rect 17612 22596 17668 23102
rect 17612 22594 17780 22596
rect 17612 22542 17614 22594
rect 17666 22542 17780 22594
rect 17612 22540 17780 22542
rect 17612 22530 17668 22540
rect 17052 22430 17054 22482
rect 17106 22430 17108 22482
rect 17052 22418 17108 22430
rect 17500 22146 17556 22158
rect 17500 22094 17502 22146
rect 17554 22094 17556 22146
rect 17500 21924 17556 22094
rect 17500 21858 17556 21868
rect 17612 21812 17668 21822
rect 17612 21718 17668 21756
rect 17500 21700 17556 21710
rect 17500 21606 17556 21644
rect 17388 21588 17444 21598
rect 17388 21494 17444 21532
rect 17724 20804 17780 22540
rect 17836 22260 17892 23996
rect 18060 23938 18116 24670
rect 18956 24164 19012 24174
rect 18060 23886 18062 23938
rect 18114 23886 18116 23938
rect 18060 23380 18116 23886
rect 18620 23938 18676 23950
rect 18620 23886 18622 23938
rect 18674 23886 18676 23938
rect 18172 23380 18228 23390
rect 18116 23378 18228 23380
rect 18116 23326 18174 23378
rect 18226 23326 18228 23378
rect 18116 23324 18228 23326
rect 18060 23286 18116 23324
rect 18172 23314 18228 23324
rect 17948 22484 18004 22494
rect 17948 22390 18004 22428
rect 18620 22260 18676 23886
rect 18732 23044 18788 23054
rect 18956 23044 19012 24108
rect 19068 24050 19124 24780
rect 19292 24724 19348 25228
rect 19404 25060 19460 25452
rect 20300 25508 20356 25518
rect 20300 25414 20356 25452
rect 19404 24994 19460 25004
rect 19516 25396 19572 25406
rect 19068 23998 19070 24050
rect 19122 23998 19124 24050
rect 19068 23828 19124 23998
rect 19068 23762 19124 23772
rect 19180 24722 19348 24724
rect 19180 24670 19294 24722
rect 19346 24670 19348 24722
rect 19180 24668 19348 24670
rect 18732 23042 18900 23044
rect 18732 22990 18734 23042
rect 18786 22990 18900 23042
rect 18732 22988 18900 22990
rect 18732 22978 18788 22988
rect 18732 22260 18788 22270
rect 17836 22204 18452 22260
rect 18284 22036 18340 22046
rect 18172 21698 18228 21710
rect 18172 21646 18174 21698
rect 18226 21646 18228 21698
rect 18060 21588 18116 21598
rect 18172 21588 18228 21646
rect 18060 21586 18228 21588
rect 18060 21534 18062 21586
rect 18114 21534 18228 21586
rect 18060 21532 18228 21534
rect 18060 21522 18116 21532
rect 17724 20244 17780 20748
rect 18172 21364 18228 21374
rect 18172 20914 18228 21308
rect 18172 20862 18174 20914
rect 18226 20862 18228 20914
rect 17724 20188 18004 20244
rect 17948 20132 18004 20188
rect 17948 20130 18116 20132
rect 17948 20078 17950 20130
rect 18002 20078 18116 20130
rect 17948 20076 18116 20078
rect 17948 20066 18004 20076
rect 17612 19346 17668 19358
rect 17612 19294 17614 19346
rect 17666 19294 17668 19346
rect 17612 19236 17668 19294
rect 17948 19236 18004 19246
rect 17612 19234 18004 19236
rect 17612 19182 17950 19234
rect 18002 19182 18004 19234
rect 17612 19180 18004 19182
rect 17948 19170 18004 19180
rect 17276 19124 17332 19134
rect 17276 19030 17332 19068
rect 17500 19012 17556 19022
rect 17388 19010 17556 19012
rect 17388 18958 17502 19010
rect 17554 18958 17556 19010
rect 17388 18956 17556 18958
rect 17388 18676 17444 18956
rect 17500 18946 17556 18956
rect 18060 18676 18116 20076
rect 16940 18498 16996 18508
rect 17052 18620 17444 18676
rect 17948 18620 18116 18676
rect 18172 19234 18228 20862
rect 18284 20132 18340 21980
rect 18396 21698 18452 22204
rect 18396 21646 18398 21698
rect 18450 21646 18452 21698
rect 18396 20356 18452 21646
rect 18508 22204 18732 22260
rect 18508 21698 18564 22204
rect 18732 22166 18788 22204
rect 18508 21646 18510 21698
rect 18562 21646 18564 21698
rect 18508 21634 18564 21646
rect 18844 21588 18900 22988
rect 18844 21522 18900 21532
rect 18956 21586 19012 22988
rect 19180 23154 19236 24668
rect 19292 24658 19348 24668
rect 19516 23938 19572 25340
rect 19852 25284 19908 25322
rect 19852 25218 19908 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20076 24612 20132 24622
rect 20076 24610 20692 24612
rect 20076 24558 20078 24610
rect 20130 24558 20692 24610
rect 20076 24556 20692 24558
rect 20076 24546 20132 24556
rect 20300 24388 20356 24398
rect 20188 24332 20300 24388
rect 19964 24052 20020 24062
rect 19964 23958 20020 23996
rect 19516 23886 19518 23938
rect 19570 23886 19572 23938
rect 19516 23548 19572 23886
rect 19836 23548 20100 23558
rect 19516 23492 19684 23548
rect 19180 23102 19182 23154
rect 19234 23102 19236 23154
rect 19180 22484 19236 23102
rect 19180 22418 19236 22428
rect 19292 22148 19348 22158
rect 18956 21534 18958 21586
rect 19010 21534 19012 21586
rect 18956 21522 19012 21534
rect 19180 22146 19348 22148
rect 19180 22094 19294 22146
rect 19346 22094 19348 22146
rect 19180 22092 19348 22094
rect 19180 21812 19236 22092
rect 19292 22082 19348 22092
rect 18508 21252 18564 21262
rect 18564 21196 18676 21252
rect 18508 21186 18564 21196
rect 18508 20804 18564 20814
rect 18508 20710 18564 20748
rect 18396 20300 18564 20356
rect 18396 20132 18452 20142
rect 18284 20130 18452 20132
rect 18284 20078 18398 20130
rect 18450 20078 18452 20130
rect 18284 20076 18452 20078
rect 18396 20066 18452 20076
rect 18508 19908 18564 20300
rect 18172 19182 18174 19234
rect 18226 19182 18228 19234
rect 16492 17778 16660 17780
rect 16492 17726 16494 17778
rect 16546 17726 16660 17778
rect 16492 17724 16660 17726
rect 16492 17714 16548 17724
rect 16268 17500 16548 17556
rect 14476 17490 14532 17500
rect 15596 17444 15652 17454
rect 15596 17350 15652 17388
rect 14364 17052 14532 17108
rect 14028 15586 14084 15596
rect 14140 15708 14308 15764
rect 14364 16882 14420 16894
rect 14364 16830 14366 16882
rect 14418 16830 14420 16882
rect 14364 16212 14420 16830
rect 13804 15316 13860 15326
rect 13804 14642 13860 15260
rect 14028 15314 14084 15326
rect 14028 15262 14030 15314
rect 14082 15262 14084 15314
rect 14028 15148 14084 15262
rect 13804 14590 13806 14642
rect 13858 14590 13860 14642
rect 13804 14578 13860 14590
rect 13916 15092 14084 15148
rect 13916 14532 13972 15092
rect 13916 14438 13972 14476
rect 13804 13748 13860 13758
rect 13804 13654 13860 13692
rect 13916 13300 13972 13310
rect 13972 13244 14084 13300
rect 13916 13234 13972 13244
rect 13692 12908 13972 12964
rect 13580 12738 13636 12750
rect 13580 12686 13582 12738
rect 13634 12686 13636 12738
rect 13580 12516 13636 12686
rect 13692 12740 13748 12750
rect 13692 12646 13748 12684
rect 13580 12450 13636 12460
rect 13132 12404 13188 12414
rect 13132 12310 13188 12348
rect 13020 12226 13076 12236
rect 13692 12292 13748 12302
rect 13748 12236 13860 12292
rect 13692 12226 13748 12236
rect 12908 12178 12964 12190
rect 12908 12126 12910 12178
rect 12962 12126 12964 12178
rect 12908 11620 12964 12126
rect 13244 12180 13300 12190
rect 13300 12124 13412 12180
rect 13244 12086 13300 12124
rect 12908 11554 12964 11564
rect 13020 11956 13076 11966
rect 12796 11394 12852 11452
rect 12796 11342 12798 11394
rect 12850 11342 12852 11394
rect 12796 11330 12852 11342
rect 12796 10724 12852 10734
rect 12684 10668 12796 10724
rect 12796 10658 12852 10668
rect 12908 9828 12964 9838
rect 13020 9828 13076 11900
rect 13356 11788 13412 12124
rect 13132 11732 13412 11788
rect 13580 12178 13636 12190
rect 13580 12126 13582 12178
rect 13634 12126 13636 12178
rect 13580 11844 13636 12126
rect 13580 11778 13636 11788
rect 13692 12066 13748 12078
rect 13692 12014 13694 12066
rect 13746 12014 13748 12066
rect 13132 11060 13188 11732
rect 13692 11620 13748 12014
rect 13468 11564 13748 11620
rect 13132 11004 13412 11060
rect 13244 10836 13300 10846
rect 13244 10742 13300 10780
rect 12908 9826 13076 9828
rect 12908 9774 12910 9826
rect 12962 9774 13076 9826
rect 12908 9772 13076 9774
rect 13356 9826 13412 11004
rect 13356 9774 13358 9826
rect 13410 9774 13412 9826
rect 12908 9762 12964 9772
rect 13356 9762 13412 9774
rect 12684 9714 12740 9726
rect 12684 9662 12686 9714
rect 12738 9662 12740 9714
rect 12684 9380 12740 9662
rect 13020 9492 13076 9502
rect 13020 9380 13076 9436
rect 12684 9324 13076 9380
rect 12572 9266 12964 9268
rect 12572 9214 12574 9266
rect 12626 9214 12964 9266
rect 12572 9212 12964 9214
rect 12572 9202 12628 9212
rect 12684 9042 12740 9054
rect 12684 8990 12686 9042
rect 12738 8990 12740 9042
rect 11228 8372 11284 8428
rect 12012 8764 12516 8820
rect 12572 8818 12628 8830
rect 12572 8766 12574 8818
rect 12626 8766 12628 8818
rect 11228 8370 11508 8372
rect 11228 8318 11230 8370
rect 11282 8318 11508 8370
rect 11228 8316 11508 8318
rect 11228 8306 11284 8316
rect 10780 8206 10782 8258
rect 10834 8206 10836 8258
rect 10780 8194 10836 8206
rect 10220 8082 10276 8092
rect 10668 8148 10724 8158
rect 10668 8054 10724 8092
rect 9772 7474 9828 7644
rect 10556 8036 10612 8046
rect 10556 7586 10612 7980
rect 10556 7534 10558 7586
rect 10610 7534 10612 7586
rect 10556 7522 10612 7534
rect 9772 7422 9774 7474
rect 9826 7422 9828 7474
rect 9772 7410 9828 7422
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 11452 6132 11508 8316
rect 12012 8258 12068 8764
rect 12012 8206 12014 8258
rect 12066 8206 12068 8258
rect 12012 8194 12068 8206
rect 12236 8260 12292 8270
rect 12236 8166 12292 8204
rect 12572 8258 12628 8766
rect 12684 8484 12740 8990
rect 12684 8418 12740 8428
rect 12908 8260 12964 9212
rect 12572 8206 12574 8258
rect 12626 8206 12628 8258
rect 12572 8194 12628 8206
rect 12684 8204 12964 8260
rect 12124 8036 12180 8046
rect 12124 7942 12180 7980
rect 12572 8036 12628 8046
rect 11452 6130 11844 6132
rect 11452 6078 11454 6130
rect 11506 6078 11844 6130
rect 11452 6076 11844 6078
rect 11452 6066 11508 6076
rect 11788 5906 11844 6076
rect 12572 6018 12628 7980
rect 12684 7362 12740 8204
rect 12684 7310 12686 7362
rect 12738 7310 12740 7362
rect 12684 7298 12740 7310
rect 13020 7362 13076 9324
rect 13468 8258 13524 11564
rect 13580 11394 13636 11406
rect 13580 11342 13582 11394
rect 13634 11342 13636 11394
rect 13580 9938 13636 11342
rect 13692 11396 13748 11406
rect 13804 11396 13860 12236
rect 13916 12290 13972 12908
rect 13916 12238 13918 12290
rect 13970 12238 13972 12290
rect 13916 11732 13972 12238
rect 13916 11666 13972 11676
rect 13692 11394 13860 11396
rect 13692 11342 13694 11394
rect 13746 11342 13860 11394
rect 13692 11340 13860 11342
rect 14028 11396 14084 13244
rect 14140 12404 14196 15708
rect 14364 15316 14420 16156
rect 14364 15222 14420 15260
rect 14252 15202 14308 15214
rect 14252 15150 14254 15202
rect 14306 15150 14308 15202
rect 14252 13746 14308 15150
rect 14476 15148 14532 17052
rect 14700 16996 14756 17006
rect 14700 16210 14756 16940
rect 15036 16996 15092 17006
rect 14700 16158 14702 16210
rect 14754 16158 14756 16210
rect 14700 16146 14756 16158
rect 14812 16882 14868 16894
rect 14812 16830 14814 16882
rect 14866 16830 14868 16882
rect 14812 16660 14868 16830
rect 14588 16098 14644 16110
rect 14588 16046 14590 16098
rect 14642 16046 14644 16098
rect 14588 15652 14644 16046
rect 14812 16100 14868 16604
rect 14924 16770 14980 16782
rect 14924 16718 14926 16770
rect 14978 16718 14980 16770
rect 14924 16212 14980 16718
rect 15036 16436 15092 16940
rect 16268 16996 16324 17006
rect 16268 16994 16436 16996
rect 16268 16942 16270 16994
rect 16322 16942 16436 16994
rect 16268 16940 16436 16942
rect 16268 16930 16324 16940
rect 16156 16882 16212 16894
rect 16156 16830 16158 16882
rect 16210 16830 16212 16882
rect 15708 16660 15764 16670
rect 15036 16380 15204 16436
rect 15036 16212 15092 16222
rect 14924 16210 15092 16212
rect 14924 16158 15038 16210
rect 15090 16158 15092 16210
rect 14924 16156 15092 16158
rect 15036 16146 15092 16156
rect 14812 16044 14980 16100
rect 14588 15596 14868 15652
rect 14700 15428 14756 15438
rect 14700 15314 14756 15372
rect 14700 15262 14702 15314
rect 14754 15262 14756 15314
rect 14700 15250 14756 15262
rect 14812 15148 14868 15596
rect 14924 15314 14980 16044
rect 14924 15262 14926 15314
rect 14978 15262 14980 15314
rect 14924 15250 14980 15262
rect 15148 15314 15204 16380
rect 15260 16098 15316 16110
rect 15260 16046 15262 16098
rect 15314 16046 15316 16098
rect 15260 15652 15316 16046
rect 15260 15586 15316 15596
rect 15148 15262 15150 15314
rect 15202 15262 15204 15314
rect 15148 15250 15204 15262
rect 15596 15202 15652 15214
rect 15596 15150 15598 15202
rect 15650 15150 15652 15202
rect 14476 15092 14756 15148
rect 14812 15092 14980 15148
rect 14252 13694 14254 13746
rect 14306 13694 14308 13746
rect 14252 13682 14308 13694
rect 14140 12338 14196 12348
rect 14476 13634 14532 13646
rect 14476 13582 14478 13634
rect 14530 13582 14532 13634
rect 14476 12290 14532 13582
rect 14700 13188 14756 15092
rect 14924 14642 14980 15092
rect 15596 15092 15652 15150
rect 15596 15026 15652 15036
rect 14924 14590 14926 14642
rect 14978 14590 14980 14642
rect 14924 14578 14980 14590
rect 14812 14532 14868 14542
rect 14812 14438 14868 14476
rect 15036 14306 15092 14318
rect 15036 14254 15038 14306
rect 15090 14254 15092 14306
rect 15036 13748 15092 14254
rect 15036 13682 15092 13692
rect 14700 13132 14868 13188
rect 14700 12740 14756 12750
rect 14700 12404 14756 12684
rect 14700 12310 14756 12348
rect 14476 12238 14478 12290
rect 14530 12238 14532 12290
rect 14476 12226 14532 12238
rect 14140 12180 14196 12190
rect 14140 12178 14420 12180
rect 14140 12126 14142 12178
rect 14194 12126 14420 12178
rect 14140 12124 14420 12126
rect 14140 12114 14196 12124
rect 14364 12068 14420 12124
rect 14588 12068 14644 12078
rect 14364 12066 14644 12068
rect 14364 12014 14590 12066
rect 14642 12014 14644 12066
rect 14364 12012 14644 12014
rect 14588 12002 14644 12012
rect 14812 11618 14868 13132
rect 15484 12404 15540 12414
rect 15484 12178 15540 12348
rect 15484 12126 15486 12178
rect 15538 12126 15540 12178
rect 15484 12114 15540 12126
rect 15596 12066 15652 12078
rect 15596 12014 15598 12066
rect 15650 12014 15652 12066
rect 14812 11566 14814 11618
rect 14866 11566 14868 11618
rect 14812 11554 14868 11566
rect 15372 11732 15428 11742
rect 13692 11330 13748 11340
rect 14028 11302 14084 11340
rect 14700 11394 14756 11406
rect 14700 11342 14702 11394
rect 14754 11342 14756 11394
rect 13804 11172 13860 11182
rect 13580 9886 13582 9938
rect 13634 9886 13636 9938
rect 13580 9874 13636 9886
rect 13692 11170 13860 11172
rect 13692 11118 13806 11170
rect 13858 11118 13860 11170
rect 13692 11116 13860 11118
rect 13692 9716 13748 11116
rect 13804 11106 13860 11116
rect 13916 11170 13972 11182
rect 13916 11118 13918 11170
rect 13970 11118 13972 11170
rect 13804 10948 13860 10958
rect 13916 10948 13972 11118
rect 14700 11172 14756 11342
rect 14700 11106 14756 11116
rect 15036 11394 15092 11406
rect 15036 11342 15038 11394
rect 15090 11342 15092 11394
rect 13916 10892 14420 10948
rect 13804 10722 13860 10892
rect 13804 10670 13806 10722
rect 13858 10670 13860 10722
rect 13804 10658 13860 10670
rect 13916 10724 13972 10734
rect 13692 9650 13748 9660
rect 13804 10164 13860 10174
rect 13804 9714 13860 10108
rect 13916 9826 13972 10668
rect 14364 10050 14420 10892
rect 14364 9998 14366 10050
rect 14418 9998 14420 10050
rect 14364 9986 14420 9998
rect 14476 10610 14532 10622
rect 14476 10558 14478 10610
rect 14530 10558 14532 10610
rect 13916 9774 13918 9826
rect 13970 9774 13972 9826
rect 13916 9762 13972 9774
rect 13804 9662 13806 9714
rect 13858 9662 13860 9714
rect 13468 8206 13470 8258
rect 13522 8206 13524 8258
rect 13468 8194 13524 8206
rect 13692 8260 13748 8270
rect 13692 8166 13748 8204
rect 13580 8036 13636 8046
rect 13804 8036 13860 9662
rect 14476 9714 14532 10558
rect 14812 10610 14868 10622
rect 14812 10558 14814 10610
rect 14866 10558 14868 10610
rect 14812 10164 14868 10558
rect 15036 10498 15092 11342
rect 15372 10722 15428 11676
rect 15372 10670 15374 10722
rect 15426 10670 15428 10722
rect 15372 10658 15428 10670
rect 15596 10612 15652 12014
rect 15708 12068 15764 16604
rect 16156 16548 16212 16830
rect 16156 16482 16212 16492
rect 16268 16658 16324 16670
rect 16268 16606 16270 16658
rect 16322 16606 16324 16658
rect 15932 15986 15988 15998
rect 15932 15934 15934 15986
rect 15986 15934 15988 15986
rect 15820 12292 15876 12302
rect 15932 12292 15988 15934
rect 16156 15316 16212 15326
rect 16156 15222 16212 15260
rect 15820 12290 15988 12292
rect 15820 12238 15822 12290
rect 15874 12238 15988 12290
rect 15820 12236 15988 12238
rect 16156 14980 16212 14990
rect 15820 12226 15876 12236
rect 15708 12012 15876 12068
rect 15708 11394 15764 11406
rect 15708 11342 15710 11394
rect 15762 11342 15764 11394
rect 15708 10836 15764 11342
rect 15820 11282 15876 12012
rect 15820 11230 15822 11282
rect 15874 11230 15876 11282
rect 15820 11218 15876 11230
rect 16156 10836 16212 14924
rect 16268 14642 16324 16606
rect 16380 15092 16436 16940
rect 16492 15148 16548 17500
rect 17052 17554 17108 18620
rect 17276 18450 17332 18462
rect 17276 18398 17278 18450
rect 17330 18398 17332 18450
rect 17052 17502 17054 17554
rect 17106 17502 17108 17554
rect 16716 17444 16772 17454
rect 16716 17350 16772 17388
rect 16716 16548 16772 16558
rect 16716 16098 16772 16492
rect 17052 16324 17108 17502
rect 17052 16258 17108 16268
rect 17164 18004 17220 18014
rect 17164 16322 17220 17948
rect 17276 16660 17332 18398
rect 17948 18452 18004 18620
rect 17948 18386 18004 18396
rect 18060 18452 18116 18462
rect 18172 18452 18228 19182
rect 18284 19852 18564 19908
rect 18284 18676 18340 19852
rect 18620 19460 18676 21196
rect 18844 20804 18900 20814
rect 18844 20690 18900 20748
rect 19180 20692 19236 21756
rect 19404 21586 19460 21598
rect 19404 21534 19406 21586
rect 19458 21534 19460 21586
rect 19404 20804 19460 21534
rect 19404 20710 19460 20748
rect 19628 20692 19684 23492
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19852 23044 19908 23054
rect 19852 22950 19908 22988
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19964 20804 20020 20814
rect 19964 20710 20020 20748
rect 18844 20638 18846 20690
rect 18898 20638 18900 20690
rect 18844 20626 18900 20638
rect 19068 20636 19236 20692
rect 19516 20690 19684 20692
rect 19516 20638 19630 20690
rect 19682 20638 19684 20690
rect 19516 20636 19684 20638
rect 18956 19908 19012 19918
rect 19068 19908 19124 20636
rect 19404 20244 19460 20254
rect 19516 20244 19572 20636
rect 19628 20626 19684 20636
rect 19404 20242 19572 20244
rect 19404 20190 19406 20242
rect 19458 20190 19572 20242
rect 19404 20188 19572 20190
rect 19628 20468 19684 20478
rect 19628 20244 19684 20412
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19740 20244 19796 20254
rect 19628 20242 19796 20244
rect 19628 20190 19742 20242
rect 19794 20190 19796 20242
rect 19628 20188 19796 20190
rect 19404 20178 19460 20188
rect 19516 20020 19572 20188
rect 19740 20178 19796 20188
rect 19516 19964 20020 20020
rect 18956 19906 19236 19908
rect 18956 19854 18958 19906
rect 19010 19854 19236 19906
rect 18956 19852 19236 19854
rect 18956 19842 19012 19852
rect 18508 19404 18676 19460
rect 18396 19010 18452 19022
rect 18396 18958 18398 19010
rect 18450 18958 18452 19010
rect 18396 18788 18452 18958
rect 18508 19012 18564 19404
rect 18620 19236 18676 19246
rect 18620 19142 18676 19180
rect 19180 19124 19236 19852
rect 19628 19236 19684 19246
rect 19180 19068 19348 19124
rect 18956 19012 19012 19022
rect 18508 19010 19236 19012
rect 18508 18958 18958 19010
rect 19010 18958 19236 19010
rect 18508 18956 19236 18958
rect 18956 18946 19012 18956
rect 18396 18732 19012 18788
rect 18284 18620 18452 18676
rect 18060 18450 18228 18452
rect 18060 18398 18062 18450
rect 18114 18398 18228 18450
rect 18060 18396 18228 18398
rect 18284 18450 18340 18462
rect 18284 18398 18286 18450
rect 18338 18398 18340 18450
rect 18060 18386 18116 18396
rect 17388 17780 17444 17790
rect 17388 17686 17444 17724
rect 18284 17780 18340 18398
rect 18396 18338 18452 18620
rect 18956 18674 19012 18732
rect 18956 18622 18958 18674
rect 19010 18622 19012 18674
rect 18956 18610 19012 18622
rect 19180 18674 19236 18956
rect 19180 18622 19182 18674
rect 19234 18622 19236 18674
rect 19180 18610 19236 18622
rect 18396 18286 18398 18338
rect 18450 18286 18452 18338
rect 18396 18274 18452 18286
rect 18844 18564 18900 18574
rect 18284 17108 18340 17724
rect 18844 17220 18900 18508
rect 19292 18452 19348 19068
rect 19404 19010 19460 19022
rect 19404 18958 19406 19010
rect 19458 18958 19460 19010
rect 19404 18788 19460 18958
rect 19404 18722 19460 18732
rect 19628 19012 19684 19180
rect 19964 19234 20020 19964
rect 19964 19182 19966 19234
rect 20018 19182 20020 19234
rect 19964 19170 20020 19182
rect 19740 19012 19796 19022
rect 19628 19010 19796 19012
rect 19628 18958 19742 19010
rect 19794 18958 19796 19010
rect 19628 18956 19796 18958
rect 19628 18676 19684 18956
rect 19740 18946 19796 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18620 19796 18676
rect 19292 18386 19348 18396
rect 19628 18450 19684 18462
rect 19628 18398 19630 18450
rect 19682 18398 19684 18450
rect 19068 18338 19124 18350
rect 19068 18286 19070 18338
rect 19122 18286 19124 18338
rect 19068 18004 19124 18286
rect 19068 17948 19572 18004
rect 19516 17778 19572 17948
rect 19516 17726 19518 17778
rect 19570 17726 19572 17778
rect 19516 17714 19572 17726
rect 19628 17556 19684 18398
rect 19068 17500 19684 17556
rect 19740 18228 19796 18620
rect 18844 17164 19012 17220
rect 18956 17108 19012 17164
rect 18284 17052 18900 17108
rect 18844 16994 18900 17052
rect 18956 17042 19012 17052
rect 19068 17106 19124 17500
rect 19740 17444 19796 18172
rect 19628 17388 19796 17444
rect 19068 17054 19070 17106
rect 19122 17054 19124 17106
rect 19068 17042 19124 17054
rect 19404 17108 19460 17118
rect 18844 16942 18846 16994
rect 18898 16942 18900 16994
rect 17276 16594 17332 16604
rect 18732 16882 18788 16894
rect 18732 16830 18734 16882
rect 18786 16830 18788 16882
rect 17164 16270 17166 16322
rect 17218 16270 17220 16322
rect 17164 16258 17220 16270
rect 18396 16324 18452 16334
rect 17612 16100 17668 16110
rect 16716 16046 16718 16098
rect 16770 16046 16772 16098
rect 16716 16034 16772 16046
rect 16828 16098 17668 16100
rect 16828 16046 17614 16098
rect 17666 16046 17668 16098
rect 16828 16044 17668 16046
rect 16828 15986 16884 16044
rect 17612 16034 17668 16044
rect 17836 16098 17892 16110
rect 18060 16100 18116 16110
rect 17836 16046 17838 16098
rect 17890 16046 17892 16098
rect 16828 15934 16830 15986
rect 16882 15934 16884 15986
rect 16828 15538 16884 15934
rect 16828 15486 16830 15538
rect 16882 15486 16884 15538
rect 16604 15316 16660 15354
rect 16604 15250 16660 15260
rect 16716 15204 16772 15242
rect 16492 15092 16660 15148
rect 16716 15138 16772 15148
rect 16380 14756 16436 15036
rect 16380 14700 16548 14756
rect 16268 14590 16270 14642
rect 16322 14590 16324 14642
rect 16268 14578 16324 14590
rect 16380 14530 16436 14542
rect 16380 14478 16382 14530
rect 16434 14478 16436 14530
rect 16380 13636 16436 14478
rect 16380 13570 16436 13580
rect 16492 13524 16548 14700
rect 16492 13458 16548 13468
rect 16604 13076 16660 15092
rect 16828 13972 16884 15486
rect 17052 15874 17108 15886
rect 17052 15822 17054 15874
rect 17106 15822 17108 15874
rect 17052 15148 17108 15822
rect 17836 15314 17892 16046
rect 17836 15262 17838 15314
rect 17890 15262 17892 15314
rect 17612 15204 17668 15242
rect 17052 15092 17556 15148
rect 17612 15138 17668 15148
rect 17500 14642 17556 15092
rect 17500 14590 17502 14642
rect 17554 14590 17556 14642
rect 17500 14578 17556 14590
rect 17052 14420 17108 14430
rect 17052 14326 17108 14364
rect 17836 14308 17892 15262
rect 16828 13906 16884 13916
rect 17500 14252 17892 14308
rect 17948 16098 18116 16100
rect 17948 16046 18062 16098
rect 18114 16046 18116 16098
rect 17948 16044 18116 16046
rect 17948 15316 18004 16044
rect 18060 16034 18116 16044
rect 17948 14530 18004 15260
rect 18396 15204 18452 16268
rect 17948 14478 17950 14530
rect 18002 14478 18004 14530
rect 17276 13636 17332 13646
rect 17388 13636 17444 13646
rect 17332 13634 17444 13636
rect 17332 13582 17390 13634
rect 17442 13582 17444 13634
rect 17332 13580 17444 13582
rect 16828 13076 16884 13086
rect 16380 13074 16884 13076
rect 16380 13022 16830 13074
rect 16882 13022 16884 13074
rect 16380 13020 16884 13022
rect 16380 12178 16436 13020
rect 16828 13010 16884 13020
rect 16380 12126 16382 12178
rect 16434 12126 16436 12178
rect 16380 12114 16436 12126
rect 16604 12290 16660 12302
rect 16604 12238 16606 12290
rect 16658 12238 16660 12290
rect 16604 11844 16660 12238
rect 16660 11788 16884 11844
rect 16604 11778 16660 11788
rect 16604 11396 16660 11406
rect 16156 10780 16436 10836
rect 15708 10770 15764 10780
rect 16268 10612 16324 10622
rect 15596 10610 16324 10612
rect 15596 10558 16270 10610
rect 16322 10558 16324 10610
rect 15596 10556 16324 10558
rect 16268 10546 16324 10556
rect 15036 10446 15038 10498
rect 15090 10446 15092 10498
rect 15036 10434 15092 10446
rect 16268 10388 16324 10398
rect 14812 10098 14868 10108
rect 16044 10164 16100 10174
rect 14476 9662 14478 9714
rect 14530 9662 14532 9714
rect 14476 9492 14532 9662
rect 14476 9426 14532 9436
rect 15148 9716 15204 9726
rect 14588 8372 14644 8382
rect 14028 8260 14084 8270
rect 14252 8260 14308 8270
rect 14028 8258 14308 8260
rect 14028 8206 14030 8258
rect 14082 8206 14254 8258
rect 14306 8206 14308 8258
rect 14028 8204 14308 8206
rect 14028 8194 14084 8204
rect 14252 8194 14308 8204
rect 14588 8258 14644 8316
rect 14588 8206 14590 8258
rect 14642 8206 14644 8258
rect 14588 8194 14644 8206
rect 14476 8036 14532 8046
rect 13804 8034 14532 8036
rect 13804 7982 14478 8034
rect 14530 7982 14532 8034
rect 13804 7980 14532 7982
rect 13580 7942 13636 7980
rect 13020 7310 13022 7362
rect 13074 7310 13076 7362
rect 13020 7298 13076 7310
rect 12572 5966 12574 6018
rect 12626 5966 12628 6018
rect 12572 5954 12628 5966
rect 11788 5854 11790 5906
rect 11842 5854 11844 5906
rect 11788 5842 11844 5854
rect 14476 5796 14532 7980
rect 15148 7586 15204 9660
rect 16044 9268 16100 10108
rect 16268 9826 16324 10332
rect 16268 9774 16270 9826
rect 16322 9774 16324 9826
rect 16268 9762 16324 9774
rect 16380 9940 16436 10780
rect 16604 10612 16660 11340
rect 16828 10722 16884 11788
rect 17052 11620 17108 11630
rect 16940 11396 16996 11406
rect 16940 11302 16996 11340
rect 16828 10670 16830 10722
rect 16882 10670 16884 10722
rect 16828 10658 16884 10670
rect 17052 11282 17108 11564
rect 17052 11230 17054 11282
rect 17106 11230 17108 11282
rect 16604 10518 16660 10556
rect 16380 9380 16436 9884
rect 16716 10498 16772 10510
rect 16716 10446 16718 10498
rect 16770 10446 16772 10498
rect 16716 9828 16772 10446
rect 17052 10164 17108 11230
rect 17164 11172 17220 11182
rect 17164 11078 17220 11116
rect 17052 10098 17108 10108
rect 16828 9940 16884 9950
rect 16828 9846 16884 9884
rect 16716 9762 16772 9772
rect 17052 9826 17108 9838
rect 17052 9774 17054 9826
rect 17106 9774 17108 9826
rect 16380 9314 16436 9324
rect 15596 9266 16100 9268
rect 15596 9214 16046 9266
rect 16098 9214 16100 9266
rect 15596 9212 16100 9214
rect 15596 8370 15652 9212
rect 16044 9202 16100 9212
rect 16268 9268 16324 9278
rect 16268 9174 16324 9212
rect 17052 9268 17108 9774
rect 17052 9202 17108 9212
rect 15932 9042 15988 9054
rect 15932 8990 15934 9042
rect 15986 8990 15988 9042
rect 15932 8484 15988 8990
rect 15932 8418 15988 8428
rect 15596 8318 15598 8370
rect 15650 8318 15652 8370
rect 15596 8306 15652 8318
rect 15148 7534 15150 7586
rect 15202 7534 15204 7586
rect 15148 7522 15204 7534
rect 15932 7476 15988 7486
rect 16380 7476 16436 7486
rect 15932 7474 16380 7476
rect 15932 7422 15934 7474
rect 15986 7422 16380 7474
rect 15932 7420 16380 7422
rect 15932 7410 15988 7420
rect 16380 7382 16436 7420
rect 14700 5796 14756 5806
rect 14476 5794 14756 5796
rect 14476 5742 14702 5794
rect 14754 5742 14756 5794
rect 14476 5740 14756 5742
rect 14700 5730 14756 5740
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 16492 3444 16548 3454
rect 17052 3444 17108 3454
rect 16492 3442 17108 3444
rect 16492 3390 16494 3442
rect 16546 3390 17054 3442
rect 17106 3390 17108 3442
rect 16492 3388 17108 3390
rect 17276 3444 17332 13580
rect 17388 13570 17444 13580
rect 17388 12178 17444 12190
rect 17388 12126 17390 12178
rect 17442 12126 17444 12178
rect 17388 11844 17444 12126
rect 17388 11778 17444 11788
rect 17500 11788 17556 14252
rect 17836 13972 17892 13982
rect 17948 13972 18004 14478
rect 18284 15092 18452 15148
rect 18508 15204 18564 15214
rect 18508 15202 18676 15204
rect 18508 15150 18510 15202
rect 18562 15150 18676 15202
rect 18508 15148 18676 15150
rect 18508 15138 18564 15148
rect 18060 14420 18116 14430
rect 18060 14084 18116 14364
rect 18284 14196 18340 15092
rect 18620 14868 18676 15148
rect 18508 14812 18676 14868
rect 18508 14532 18564 14812
rect 18732 14756 18788 16830
rect 18844 16884 18900 16942
rect 18844 16828 19236 16884
rect 19180 15428 19236 16828
rect 19292 15428 19348 15438
rect 19180 15426 19348 15428
rect 19180 15374 19294 15426
rect 19346 15374 19348 15426
rect 19180 15372 19348 15374
rect 19292 15362 19348 15372
rect 19068 15314 19124 15326
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 18508 14466 18564 14476
rect 18620 14700 18788 14756
rect 18956 15204 19012 15214
rect 18396 14420 18452 14430
rect 18396 14326 18452 14364
rect 18284 14140 18564 14196
rect 18060 14028 18340 14084
rect 17948 13916 18228 13972
rect 17836 13636 17892 13916
rect 17948 13636 18004 13646
rect 17836 13634 18004 13636
rect 17836 13582 17950 13634
rect 18002 13582 18004 13634
rect 17836 13580 18004 13582
rect 17948 13570 18004 13580
rect 18060 13636 18116 13646
rect 17612 13524 17668 13534
rect 17612 13430 17668 13468
rect 17612 12404 17668 12414
rect 17612 12402 17892 12404
rect 17612 12350 17614 12402
rect 17666 12350 17892 12402
rect 17612 12348 17892 12350
rect 17612 12338 17668 12348
rect 17724 12178 17780 12190
rect 17724 12126 17726 12178
rect 17778 12126 17780 12178
rect 17500 11732 17668 11788
rect 17388 10612 17444 10622
rect 17388 8930 17444 10556
rect 17612 10052 17668 11732
rect 17724 11732 17780 12126
rect 17724 11666 17780 11676
rect 17836 10836 17892 12348
rect 17948 12292 18004 12302
rect 18060 12292 18116 13580
rect 17948 12290 18116 12292
rect 17948 12238 17950 12290
rect 18002 12238 18116 12290
rect 17948 12236 18116 12238
rect 17948 12226 18004 12236
rect 18172 11788 18228 13916
rect 18284 13858 18340 14028
rect 18508 13970 18564 14140
rect 18508 13918 18510 13970
rect 18562 13918 18564 13970
rect 18508 13906 18564 13918
rect 18284 13806 18286 13858
rect 18338 13806 18340 13858
rect 18284 13794 18340 13806
rect 18396 13636 18452 13646
rect 18396 13542 18452 13580
rect 18620 12402 18676 14700
rect 18844 14644 18900 14654
rect 18732 14532 18788 14542
rect 18732 14438 18788 14476
rect 18844 12962 18900 14588
rect 18956 14418 19012 15148
rect 19068 14754 19124 15262
rect 19404 15148 19460 17052
rect 19628 15426 19684 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20076 17108 20132 17118
rect 20076 17014 20132 17052
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19628 15374 19630 15426
rect 19682 15374 19684 15426
rect 19068 14702 19070 14754
rect 19122 14702 19124 14754
rect 19068 14690 19124 14702
rect 19180 15092 19460 15148
rect 19516 15202 19572 15214
rect 19516 15150 19518 15202
rect 19570 15150 19572 15202
rect 18956 14366 18958 14418
rect 19010 14366 19012 14418
rect 18956 14354 19012 14366
rect 19180 13076 19236 15092
rect 19516 14532 19572 15150
rect 19628 14644 19684 15374
rect 19628 14578 19684 14588
rect 19740 15204 19796 15214
rect 19516 14466 19572 14476
rect 19740 14530 19796 15148
rect 19740 14478 19742 14530
rect 19794 14478 19796 14530
rect 19740 14466 19796 14478
rect 19404 14420 19460 14430
rect 19404 14326 19460 14364
rect 19516 14306 19572 14318
rect 19516 14254 19518 14306
rect 19570 14254 19572 14306
rect 19404 13636 19460 13646
rect 18844 12910 18846 12962
rect 18898 12910 18900 12962
rect 18844 12898 18900 12910
rect 18956 13020 19236 13076
rect 19292 13634 19460 13636
rect 19292 13582 19406 13634
rect 19458 13582 19460 13634
rect 19292 13580 19460 13582
rect 18620 12350 18622 12402
rect 18674 12350 18676 12402
rect 18620 12292 18676 12350
rect 18396 12178 18452 12190
rect 18396 12126 18398 12178
rect 18450 12126 18452 12178
rect 18172 11732 18340 11788
rect 17948 10836 18004 10846
rect 17836 10834 18004 10836
rect 17836 10782 17950 10834
rect 18002 10782 18004 10834
rect 17836 10780 18004 10782
rect 17948 10770 18004 10780
rect 18172 10610 18228 10622
rect 18172 10558 18174 10610
rect 18226 10558 18228 10610
rect 18060 10498 18116 10510
rect 18060 10446 18062 10498
rect 18114 10446 18116 10498
rect 17612 9996 17892 10052
rect 17724 9828 17780 9838
rect 17724 9734 17780 9772
rect 17500 9716 17556 9726
rect 17500 9622 17556 9660
rect 17388 8878 17390 8930
rect 17442 8878 17444 8930
rect 17388 8866 17444 8878
rect 17612 9602 17668 9614
rect 17612 9550 17614 9602
rect 17666 9550 17668 9602
rect 17612 8372 17668 9550
rect 17724 8372 17780 8382
rect 17612 8370 17780 8372
rect 17612 8318 17726 8370
rect 17778 8318 17780 8370
rect 17612 8316 17780 8318
rect 17724 8306 17780 8316
rect 17612 4226 17668 4238
rect 17612 4174 17614 4226
rect 17666 4174 17668 4226
rect 17388 3444 17444 3454
rect 17276 3442 17444 3444
rect 17276 3390 17390 3442
rect 17442 3390 17444 3442
rect 17276 3388 17444 3390
rect 16492 3378 16548 3388
rect 16828 800 16884 3388
rect 17052 3378 17108 3388
rect 17388 3378 17444 3388
rect 17612 3332 17668 4174
rect 17836 4004 17892 9996
rect 18060 9156 18116 10446
rect 18172 9716 18228 10558
rect 18172 9650 18228 9660
rect 18060 9090 18116 9100
rect 18284 6580 18340 11732
rect 18396 10836 18452 12126
rect 18396 10770 18452 10780
rect 18396 10612 18452 10622
rect 18396 9716 18452 10556
rect 18508 10610 18564 10622
rect 18508 10558 18510 10610
rect 18562 10558 18564 10610
rect 18508 10050 18564 10558
rect 18508 9998 18510 10050
rect 18562 9998 18564 10050
rect 18508 9986 18564 9998
rect 18620 9826 18676 12236
rect 18620 9774 18622 9826
rect 18674 9774 18676 9826
rect 18620 9762 18676 9774
rect 18956 9828 19012 13020
rect 19180 12852 19236 12862
rect 19292 12852 19348 13580
rect 19404 13570 19460 13580
rect 19404 12964 19460 12974
rect 19516 12964 19572 14254
rect 20188 14196 20244 24332
rect 20300 24322 20356 24332
rect 20636 24162 20692 24556
rect 20860 24388 20916 26852
rect 21084 26514 21140 26908
rect 21084 26462 21086 26514
rect 21138 26462 21140 26514
rect 21084 26450 21140 26462
rect 21196 27746 21252 27758
rect 21196 27694 21198 27746
rect 21250 27694 21252 27746
rect 21196 26516 21252 27694
rect 21420 27748 21476 27758
rect 21420 27186 21476 27692
rect 21756 27636 21812 30492
rect 21420 27134 21422 27186
rect 21474 27134 21476 27186
rect 21420 27122 21476 27134
rect 21644 27580 21812 27636
rect 21308 27076 21364 27086
rect 21308 26982 21364 27020
rect 21532 26964 21588 27002
rect 21532 26898 21588 26908
rect 21196 26450 21252 26460
rect 21308 25396 21364 25406
rect 21308 25302 21364 25340
rect 20860 24322 20916 24332
rect 20636 24110 20638 24162
rect 20690 24110 20692 24162
rect 20636 24098 20692 24110
rect 20748 24052 20804 24062
rect 21420 24052 21476 24062
rect 20748 24050 21476 24052
rect 20748 23998 20750 24050
rect 20802 23998 21422 24050
rect 21474 23998 21476 24050
rect 20748 23996 21476 23998
rect 20748 23986 20804 23996
rect 21420 23986 21476 23996
rect 21532 23940 21588 23950
rect 21532 23846 21588 23884
rect 21308 23828 21364 23838
rect 21364 23772 21476 23828
rect 21308 23762 21364 23772
rect 21420 23714 21476 23772
rect 21420 23662 21422 23714
rect 21474 23662 21476 23714
rect 21420 23650 21476 23662
rect 20636 23044 20692 23054
rect 20636 22594 20692 22988
rect 20636 22542 20638 22594
rect 20690 22542 20692 22594
rect 20636 22530 20692 22542
rect 20748 22260 20804 22270
rect 20748 22258 21140 22260
rect 20748 22206 20750 22258
rect 20802 22206 21140 22258
rect 20748 22204 21140 22206
rect 20748 22194 20804 22204
rect 20972 22036 21028 22046
rect 20972 21810 21028 21980
rect 20972 21758 20974 21810
rect 21026 21758 21028 21810
rect 20972 21746 21028 21758
rect 21084 21810 21140 22204
rect 21084 21758 21086 21810
rect 21138 21758 21140 21810
rect 21084 21746 21140 21758
rect 21196 21812 21252 21822
rect 21196 21718 21252 21756
rect 21420 21700 21476 21710
rect 21420 21606 21476 21644
rect 20860 21586 20916 21598
rect 20860 21534 20862 21586
rect 20914 21534 20916 21586
rect 20524 20802 20580 20814
rect 20524 20750 20526 20802
rect 20578 20750 20580 20802
rect 20524 20356 20580 20750
rect 20860 20804 20916 21534
rect 20860 20738 20916 20748
rect 20524 20290 20580 20300
rect 20748 20692 20804 20702
rect 20300 19906 20356 19918
rect 20300 19854 20302 19906
rect 20354 19854 20356 19906
rect 20300 18116 20356 19854
rect 20748 19122 20804 20636
rect 21196 20020 21252 20030
rect 21644 20020 21700 27580
rect 21868 26908 21924 30716
rect 22204 29540 22260 31052
rect 22428 30660 22484 31276
rect 22540 31266 22596 31276
rect 22876 30996 22932 31612
rect 22988 31666 23044 31678
rect 22988 31614 22990 31666
rect 23042 31614 23044 31666
rect 22988 31220 23044 31614
rect 22988 31154 23044 31164
rect 23212 31554 23268 31566
rect 23212 31502 23214 31554
rect 23266 31502 23268 31554
rect 22988 30996 23044 31006
rect 22876 30994 23044 30996
rect 22876 30942 22990 30994
rect 23042 30942 23044 30994
rect 22876 30940 23044 30942
rect 22540 30884 22596 30894
rect 22540 30882 22708 30884
rect 22540 30830 22542 30882
rect 22594 30830 22708 30882
rect 22540 30828 22708 30830
rect 22540 30818 22596 30828
rect 22428 30604 22596 30660
rect 22316 30436 22372 30446
rect 22316 30100 22372 30380
rect 22428 30434 22484 30446
rect 22428 30382 22430 30434
rect 22482 30382 22484 30434
rect 22428 30324 22484 30382
rect 22428 30258 22484 30268
rect 22540 30210 22596 30604
rect 22540 30158 22542 30210
rect 22594 30158 22596 30210
rect 22540 30146 22596 30158
rect 22428 30100 22484 30110
rect 22316 30098 22484 30100
rect 22316 30046 22430 30098
rect 22482 30046 22484 30098
rect 22316 30044 22484 30046
rect 22428 30034 22484 30044
rect 22652 29764 22708 30828
rect 22876 30436 22932 30446
rect 22876 30342 22932 30380
rect 22988 30100 23044 30940
rect 23100 30996 23156 31006
rect 23100 30322 23156 30940
rect 23212 30884 23268 31502
rect 23324 30884 23380 30894
rect 23212 30882 23380 30884
rect 23212 30830 23326 30882
rect 23378 30830 23380 30882
rect 23212 30828 23380 30830
rect 23324 30818 23380 30828
rect 23100 30270 23102 30322
rect 23154 30270 23156 30322
rect 23100 30258 23156 30270
rect 23100 30100 23156 30110
rect 22988 30098 23156 30100
rect 22988 30046 23102 30098
rect 23154 30046 23156 30098
rect 22988 30044 23156 30046
rect 23100 30034 23156 30044
rect 22652 29708 23044 29764
rect 22428 29652 22484 29662
rect 22428 29558 22484 29596
rect 22316 29540 22372 29550
rect 22204 29484 22316 29540
rect 22316 29474 22372 29484
rect 21980 29428 22036 29438
rect 21980 29426 22260 29428
rect 21980 29374 21982 29426
rect 22034 29374 22260 29426
rect 21980 29372 22260 29374
rect 21980 29362 22036 29372
rect 21980 29204 22036 29214
rect 21980 28420 22036 29148
rect 22204 28756 22260 29372
rect 22764 29204 22820 29214
rect 22204 28662 22260 28700
rect 22316 29202 22820 29204
rect 22316 29150 22766 29202
rect 22818 29150 22820 29202
rect 22316 29148 22820 29150
rect 21980 27636 22036 28364
rect 22092 28084 22148 28094
rect 22316 28084 22372 29148
rect 22764 29138 22820 29148
rect 22092 28082 22372 28084
rect 22092 28030 22094 28082
rect 22146 28030 22372 28082
rect 22092 28028 22372 28030
rect 22092 28018 22148 28028
rect 22988 27970 23044 29708
rect 23436 29652 23492 34188
rect 23548 34178 23604 34188
rect 23772 34692 23828 35420
rect 24108 34916 24164 34926
rect 24444 34916 24500 39006
rect 25116 39284 25172 39294
rect 25116 38500 25172 39228
rect 25228 38834 25284 40348
rect 25340 40292 25396 40302
rect 25396 40236 25508 40292
rect 25340 40226 25396 40236
rect 25452 38948 25508 40236
rect 25564 39060 25620 42478
rect 25900 42532 25956 42542
rect 25900 42194 25956 42476
rect 25900 42142 25902 42194
rect 25954 42142 25956 42194
rect 25900 42130 25956 42142
rect 26124 42194 26180 42700
rect 26348 42642 26404 42700
rect 26348 42590 26350 42642
rect 26402 42590 26404 42642
rect 26348 42578 26404 42590
rect 26124 42142 26126 42194
rect 26178 42142 26180 42194
rect 26124 42130 26180 42142
rect 26236 42532 26292 42542
rect 26236 41972 26292 42476
rect 26460 42420 26516 42812
rect 26684 42756 26740 42812
rect 26908 42756 26964 42766
rect 26684 42754 26964 42756
rect 26684 42702 26910 42754
rect 26962 42702 26964 42754
rect 26684 42700 26964 42702
rect 26908 42690 26964 42700
rect 27244 42756 27300 43486
rect 27244 42690 27300 42700
rect 26348 42364 26516 42420
rect 26572 42644 26628 42654
rect 26572 42420 26628 42588
rect 26348 42082 26404 42364
rect 26572 42354 26628 42364
rect 26684 42530 26740 42542
rect 26684 42478 26686 42530
rect 26738 42478 26740 42530
rect 26684 42196 26740 42478
rect 26684 42130 26740 42140
rect 26348 42030 26350 42082
rect 26402 42030 26404 42082
rect 26348 42018 26404 42030
rect 26796 42084 26852 42094
rect 26796 42082 26964 42084
rect 26796 42030 26798 42082
rect 26850 42030 26964 42082
rect 26796 42028 26964 42030
rect 26796 42018 26852 42028
rect 26124 41916 26292 41972
rect 26684 41970 26740 41982
rect 26684 41918 26686 41970
rect 26738 41918 26740 41970
rect 25676 41412 25732 41422
rect 25676 40514 25732 41356
rect 25788 41186 25844 41198
rect 25788 41134 25790 41186
rect 25842 41134 25844 41186
rect 25788 40740 25844 41134
rect 25788 40674 25844 40684
rect 25676 40462 25678 40514
rect 25730 40462 25732 40514
rect 25676 40450 25732 40462
rect 25788 40516 25844 40526
rect 26124 40516 26180 41916
rect 26236 41748 26292 41758
rect 26684 41748 26740 41918
rect 26908 41860 26964 42028
rect 27356 41860 27412 41870
rect 26908 41804 27356 41860
rect 26236 41746 26740 41748
rect 26236 41694 26238 41746
rect 26290 41694 26740 41746
rect 26236 41692 26740 41694
rect 26796 41748 26852 41758
rect 26796 41746 26964 41748
rect 26796 41694 26798 41746
rect 26850 41694 26964 41746
rect 26796 41692 26964 41694
rect 26236 41682 26292 41692
rect 26796 41682 26852 41692
rect 26460 41076 26516 41086
rect 26460 41074 26852 41076
rect 26460 41022 26462 41074
rect 26514 41022 26852 41074
rect 26460 41020 26852 41022
rect 26460 41010 26516 41020
rect 26684 40628 26740 40638
rect 26684 40534 26740 40572
rect 26796 40626 26852 41020
rect 26796 40574 26798 40626
rect 26850 40574 26852 40626
rect 26796 40562 26852 40574
rect 26908 40626 26964 41692
rect 27020 41076 27076 41804
rect 27356 41766 27412 41804
rect 27020 41010 27076 41020
rect 26908 40574 26910 40626
rect 26962 40574 26964 40626
rect 26908 40562 26964 40574
rect 25788 40514 26068 40516
rect 25788 40462 25790 40514
rect 25842 40462 26068 40514
rect 25788 40460 26068 40462
rect 26124 40460 26404 40516
rect 25788 40450 25844 40460
rect 25788 40180 25844 40190
rect 25788 40178 25956 40180
rect 25788 40126 25790 40178
rect 25842 40126 25956 40178
rect 25788 40124 25956 40126
rect 25788 40114 25844 40124
rect 25676 39060 25732 39070
rect 25564 39058 25732 39060
rect 25564 39006 25678 39058
rect 25730 39006 25732 39058
rect 25564 39004 25732 39006
rect 25676 38994 25732 39004
rect 25900 39058 25956 40124
rect 25900 39006 25902 39058
rect 25954 39006 25956 39058
rect 25900 38994 25956 39006
rect 25452 38892 25620 38948
rect 25228 38782 25230 38834
rect 25282 38782 25284 38834
rect 25228 38770 25284 38782
rect 25452 38722 25508 38734
rect 25452 38670 25454 38722
rect 25506 38670 25508 38722
rect 25452 38668 25508 38670
rect 25116 38434 25172 38444
rect 25228 38612 25508 38668
rect 25228 37378 25284 38612
rect 25564 37380 25620 38892
rect 25788 38836 25844 38846
rect 25788 38742 25844 38780
rect 25676 38164 25732 38174
rect 25732 38108 25844 38164
rect 25676 38098 25732 38108
rect 25228 37326 25230 37378
rect 25282 37326 25284 37378
rect 25228 37314 25284 37326
rect 25340 37324 25620 37380
rect 24780 36820 24836 36830
rect 24780 36594 24836 36764
rect 24780 36542 24782 36594
rect 24834 36542 24836 36594
rect 24780 36530 24836 36542
rect 24780 36372 24836 36382
rect 24668 35924 24724 35934
rect 24668 35830 24724 35868
rect 24108 34822 24164 34860
rect 24220 34860 24500 34916
rect 23884 34804 23940 34814
rect 23884 34710 23940 34748
rect 23772 34242 23828 34636
rect 23772 34190 23774 34242
rect 23826 34190 23828 34242
rect 23772 34178 23828 34190
rect 23548 34020 23604 34030
rect 23548 33124 23604 33964
rect 24108 33460 24164 33470
rect 24220 33460 24276 34860
rect 24444 34692 24500 34702
rect 24444 34598 24500 34636
rect 24780 34356 24836 36316
rect 25116 36148 25172 36158
rect 25116 35026 25172 36092
rect 25228 35812 25284 35822
rect 25340 35812 25396 37324
rect 25676 37268 25732 37278
rect 25676 37174 25732 37212
rect 25564 37154 25620 37166
rect 25564 37102 25566 37154
rect 25618 37102 25620 37154
rect 25564 36706 25620 37102
rect 25564 36654 25566 36706
rect 25618 36654 25620 36706
rect 25564 36642 25620 36654
rect 25228 35810 25396 35812
rect 25228 35758 25230 35810
rect 25282 35758 25396 35810
rect 25228 35756 25396 35758
rect 25452 36370 25508 36382
rect 25452 36318 25454 36370
rect 25506 36318 25508 36370
rect 25228 35746 25284 35756
rect 25452 35588 25508 36318
rect 25564 36260 25620 36270
rect 25564 36166 25620 36204
rect 25452 35522 25508 35532
rect 25116 34974 25118 35026
rect 25170 34974 25172 35026
rect 25116 34962 25172 34974
rect 25228 34356 25284 34366
rect 24780 34354 25284 34356
rect 24780 34302 24782 34354
rect 24834 34302 25230 34354
rect 25282 34302 25284 34354
rect 24780 34300 25284 34302
rect 24780 34290 24836 34300
rect 25228 34290 25284 34300
rect 25564 34244 25620 34254
rect 24108 33458 24276 33460
rect 24108 33406 24110 33458
rect 24162 33406 24276 33458
rect 24108 33404 24276 33406
rect 24108 33394 24164 33404
rect 24220 33348 24276 33404
rect 25452 34242 25620 34244
rect 25452 34190 25566 34242
rect 25618 34190 25620 34242
rect 25452 34188 25620 34190
rect 24220 33282 24276 33292
rect 24892 33348 24948 33358
rect 24892 33254 24948 33292
rect 25340 33348 25396 33358
rect 23548 33058 23604 33068
rect 24444 33234 24500 33246
rect 24444 33182 24446 33234
rect 24498 33182 24500 33234
rect 24444 32788 24500 33182
rect 24556 33236 24612 33246
rect 24556 33142 24612 33180
rect 24444 32722 24500 32732
rect 25228 32676 25284 32686
rect 25228 32582 25284 32620
rect 23660 32116 23716 32126
rect 23716 32060 23828 32116
rect 23660 32050 23716 32060
rect 23548 31668 23604 31678
rect 23548 31666 23716 31668
rect 23548 31614 23550 31666
rect 23602 31614 23716 31666
rect 23548 31612 23716 31614
rect 23548 31602 23604 31612
rect 23660 30884 23716 31612
rect 23772 31332 23828 32060
rect 23996 31892 24052 31902
rect 23996 31798 24052 31836
rect 24668 31892 24724 31902
rect 25340 31892 25396 33292
rect 25452 32564 25508 34188
rect 25564 34178 25620 34188
rect 25676 33236 25732 33246
rect 25676 33142 25732 33180
rect 25676 32900 25732 32910
rect 25564 32788 25620 32798
rect 25564 32694 25620 32732
rect 25676 32786 25732 32844
rect 25676 32734 25678 32786
rect 25730 32734 25732 32786
rect 25676 32722 25732 32734
rect 25452 32470 25508 32508
rect 25452 31892 25508 31902
rect 25340 31890 25732 31892
rect 25340 31838 25454 31890
rect 25506 31838 25732 31890
rect 25340 31836 25732 31838
rect 24220 31780 24276 31790
rect 24220 31778 24388 31780
rect 24220 31726 24222 31778
rect 24274 31726 24388 31778
rect 24220 31724 24388 31726
rect 24220 31714 24276 31724
rect 23884 31668 23940 31678
rect 23884 31574 23940 31612
rect 24332 31332 24388 31724
rect 24556 31668 24612 31678
rect 23772 31276 24164 31332
rect 23772 30996 23828 31006
rect 23772 30902 23828 30940
rect 23548 30324 23604 30334
rect 23660 30324 23716 30828
rect 23772 30324 23828 30334
rect 23660 30322 23828 30324
rect 23660 30270 23774 30322
rect 23826 30270 23828 30322
rect 23660 30268 23828 30270
rect 23548 30230 23604 30268
rect 23772 30258 23828 30268
rect 24108 30322 24164 31276
rect 24108 30270 24110 30322
rect 24162 30270 24164 30322
rect 24108 30258 24164 30270
rect 24220 31276 24388 31332
rect 24444 31554 24500 31566
rect 24444 31502 24446 31554
rect 24498 31502 24500 31554
rect 24444 31332 24500 31502
rect 24220 30994 24276 31276
rect 24444 31266 24500 31276
rect 24220 30942 24222 30994
rect 24274 30942 24276 30994
rect 24220 30212 24276 30942
rect 24444 30996 24500 31006
rect 24556 30996 24612 31612
rect 24668 31554 24724 31836
rect 25452 31826 25508 31836
rect 25676 31778 25732 31836
rect 25676 31726 25678 31778
rect 25730 31726 25732 31778
rect 25676 31714 25732 31726
rect 24668 31502 24670 31554
rect 24722 31502 24724 31554
rect 24668 31220 24724 31502
rect 24780 31666 24836 31678
rect 24780 31614 24782 31666
rect 24834 31614 24836 31666
rect 24780 31556 24836 31614
rect 24836 31500 25284 31556
rect 24780 31490 24836 31500
rect 24668 31154 24724 31164
rect 25228 31106 25284 31500
rect 25452 31220 25508 31230
rect 25452 31126 25508 31164
rect 25228 31054 25230 31106
rect 25282 31054 25284 31106
rect 25228 31042 25284 31054
rect 24500 30940 24612 30996
rect 24444 30902 24500 30940
rect 24332 30882 24388 30894
rect 24332 30830 24334 30882
rect 24386 30830 24388 30882
rect 24332 30772 24388 30830
rect 25340 30884 25396 30894
rect 25340 30790 25396 30828
rect 24332 30706 24388 30716
rect 25788 30436 25844 38108
rect 26012 37828 26068 40460
rect 26236 40292 26292 40302
rect 26236 40198 26292 40236
rect 26236 39956 26292 39966
rect 26124 39732 26180 39742
rect 26124 38164 26180 39676
rect 26124 38098 26180 38108
rect 26012 37762 26068 37772
rect 26236 36594 26292 39900
rect 26348 36708 26404 40460
rect 26460 40292 26516 40302
rect 26460 40290 26628 40292
rect 26460 40238 26462 40290
rect 26514 40238 26628 40290
rect 26460 40236 26628 40238
rect 26460 40226 26516 40236
rect 26460 39620 26516 39630
rect 26460 38834 26516 39564
rect 26460 38782 26462 38834
rect 26514 38782 26516 38834
rect 26460 38770 26516 38782
rect 26572 38052 26628 40236
rect 27580 39732 27636 46396
rect 27916 45444 27972 47180
rect 28252 46562 28308 46574
rect 28252 46510 28254 46562
rect 28306 46510 28308 46562
rect 28252 46004 28308 46510
rect 28140 45948 28308 46004
rect 28140 45890 28196 45948
rect 28140 45838 28142 45890
rect 28194 45838 28196 45890
rect 28140 45826 28196 45838
rect 28028 45668 28084 45678
rect 28028 45574 28084 45612
rect 28252 45666 28308 45678
rect 28252 45614 28254 45666
rect 28306 45614 28308 45666
rect 28252 45444 28308 45614
rect 27916 45388 28308 45444
rect 27916 44434 27972 44446
rect 27916 44382 27918 44434
rect 27970 44382 27972 44434
rect 27916 43652 27972 44382
rect 28364 43876 28420 47406
rect 28364 43810 28420 43820
rect 27916 43586 27972 43596
rect 28140 43316 28196 43326
rect 28140 42754 28196 43260
rect 28140 42702 28142 42754
rect 28194 42702 28196 42754
rect 28140 42690 28196 42702
rect 28252 42644 28308 42654
rect 28252 42550 28308 42588
rect 28476 42530 28532 42542
rect 28476 42478 28478 42530
rect 28530 42478 28532 42530
rect 27916 41188 27972 41198
rect 27916 40740 27972 41132
rect 28476 40964 28532 42478
rect 28588 41298 28644 49084
rect 28924 48916 28980 48926
rect 28700 45892 28756 45902
rect 28700 45890 28868 45892
rect 28700 45838 28702 45890
rect 28754 45838 28868 45890
rect 28700 45836 28868 45838
rect 28700 45826 28756 45836
rect 28812 45668 28868 45836
rect 28700 43426 28756 43438
rect 28700 43374 28702 43426
rect 28754 43374 28756 43426
rect 28700 42644 28756 43374
rect 28700 42578 28756 42588
rect 28812 42420 28868 45612
rect 28588 41246 28590 41298
rect 28642 41246 28644 41298
rect 28588 41234 28644 41246
rect 28700 42364 28868 42420
rect 28476 40908 28644 40964
rect 27916 40628 27972 40684
rect 27580 39666 27636 39676
rect 27692 40626 27972 40628
rect 27692 40574 27918 40626
rect 27970 40574 27972 40626
rect 27692 40572 27972 40574
rect 27692 39620 27748 40572
rect 27916 40562 27972 40572
rect 28476 40740 28532 40750
rect 26908 39506 26964 39518
rect 26908 39454 26910 39506
rect 26962 39454 26964 39506
rect 26908 38836 26964 39454
rect 27132 39060 27188 39070
rect 27132 38946 27188 39004
rect 27132 38894 27134 38946
rect 27186 38894 27188 38946
rect 27132 38882 27188 38894
rect 26908 38770 26964 38780
rect 27692 38724 27748 39564
rect 28252 39732 28308 39742
rect 28252 39618 28308 39676
rect 28252 39566 28254 39618
rect 28306 39566 28308 39618
rect 28252 39554 28308 39566
rect 28028 39396 28084 39406
rect 28028 39302 28084 39340
rect 28140 39394 28196 39406
rect 28140 39342 28142 39394
rect 28194 39342 28196 39394
rect 28140 39060 28196 39342
rect 28140 38994 28196 39004
rect 27692 38658 27748 38668
rect 26572 37996 27300 38052
rect 26908 37378 26964 37390
rect 26908 37326 26910 37378
rect 26962 37326 26964 37378
rect 26684 37268 26740 37278
rect 26348 36642 26404 36652
rect 26460 37266 26740 37268
rect 26460 37214 26686 37266
rect 26738 37214 26740 37266
rect 26460 37212 26740 37214
rect 26236 36542 26238 36594
rect 26290 36542 26292 36594
rect 26236 36530 26292 36542
rect 26460 36482 26516 37212
rect 26684 37202 26740 37212
rect 26908 36708 26964 37326
rect 26460 36430 26462 36482
rect 26514 36430 26516 36482
rect 26460 36418 26516 36430
rect 26572 36652 26964 36708
rect 26572 36260 26628 36652
rect 26796 36484 26852 36494
rect 26796 36390 26852 36428
rect 26572 35924 26628 36204
rect 26908 36260 26964 36652
rect 26908 36194 26964 36204
rect 27020 37266 27076 37278
rect 27020 37214 27022 37266
rect 27074 37214 27076 37266
rect 27020 36932 27076 37214
rect 26684 35924 26740 35934
rect 26572 35922 26740 35924
rect 26572 35870 26686 35922
rect 26738 35870 26740 35922
rect 26572 35868 26740 35870
rect 26684 35858 26740 35868
rect 25900 35698 25956 35710
rect 25900 35646 25902 35698
rect 25954 35646 25956 35698
rect 25900 34692 25956 35646
rect 26124 35700 26180 35710
rect 26460 35700 26516 35710
rect 26124 35698 26516 35700
rect 26124 35646 26126 35698
rect 26178 35646 26462 35698
rect 26514 35646 26516 35698
rect 26124 35644 26516 35646
rect 26124 35634 26180 35644
rect 26460 35634 26516 35644
rect 26796 35698 26852 35710
rect 26796 35646 26798 35698
rect 26850 35646 26852 35698
rect 26796 35588 26852 35646
rect 26572 35532 26852 35588
rect 26572 35308 26628 35532
rect 27020 35476 27076 36876
rect 27244 35810 27300 37996
rect 27804 37828 27860 37838
rect 27244 35758 27246 35810
rect 27298 35758 27300 35810
rect 27244 35746 27300 35758
rect 27580 37266 27636 37278
rect 27580 37214 27582 37266
rect 27634 37214 27636 37266
rect 27580 36820 27636 37214
rect 27580 36484 27636 36764
rect 27804 36708 27860 37772
rect 28364 37492 28420 37502
rect 28476 37492 28532 40684
rect 28588 39618 28644 40908
rect 28588 39566 28590 39618
rect 28642 39566 28644 39618
rect 28588 39554 28644 39566
rect 28588 37828 28644 37838
rect 28588 37734 28644 37772
rect 28700 37604 28756 42364
rect 28812 41188 28868 41198
rect 28812 40626 28868 41132
rect 28812 40574 28814 40626
rect 28866 40574 28868 40626
rect 28812 40562 28868 40574
rect 28924 38724 28980 48860
rect 29372 48804 29428 48814
rect 29148 48802 29428 48804
rect 29148 48750 29374 48802
rect 29426 48750 29428 48802
rect 29148 48748 29428 48750
rect 29148 47346 29204 48748
rect 29372 48738 29428 48748
rect 29260 48244 29316 48254
rect 29260 47682 29316 48188
rect 29372 48132 29428 48142
rect 29372 48038 29428 48076
rect 29260 47630 29262 47682
rect 29314 47630 29316 47682
rect 29260 47618 29316 47630
rect 29596 47460 29652 50372
rect 30156 50260 30212 50540
rect 30716 50530 30772 50540
rect 30828 50428 30884 53452
rect 30940 53172 30996 53676
rect 31276 54684 31388 54740
rect 31276 53284 31332 54684
rect 31388 54646 31444 54684
rect 31612 54516 31668 55134
rect 31612 54450 31668 54460
rect 32172 54626 32228 54638
rect 32172 54574 32174 54626
rect 32226 54574 32228 54626
rect 31388 54402 31444 54414
rect 31388 54350 31390 54402
rect 31442 54350 31444 54402
rect 31388 53842 31444 54350
rect 31388 53790 31390 53842
rect 31442 53790 31444 53842
rect 31388 53778 31444 53790
rect 31612 54290 31668 54302
rect 31612 54238 31614 54290
rect 31666 54238 31668 54290
rect 31276 53218 31332 53228
rect 30940 53106 30996 53116
rect 31612 53170 31668 54238
rect 31612 53118 31614 53170
rect 31666 53118 31668 53170
rect 31612 53106 31668 53118
rect 31836 53060 31892 53070
rect 31836 52966 31892 53004
rect 31500 52948 31556 52958
rect 31500 52854 31556 52892
rect 31948 52948 32004 52958
rect 32172 52948 32228 54574
rect 32284 53508 32340 59200
rect 33180 56308 33236 56318
rect 33180 56214 33236 56252
rect 32284 53442 32340 53452
rect 32396 56082 32452 56094
rect 32396 56030 32398 56082
rect 32450 56030 32452 56082
rect 31948 52946 32228 52948
rect 31948 52894 31950 52946
rect 32002 52894 32228 52946
rect 31948 52892 32228 52894
rect 31388 52388 31444 52398
rect 31388 52294 31444 52332
rect 29932 50204 30212 50260
rect 30268 50372 30884 50428
rect 31724 52052 31780 52062
rect 29932 48916 29988 50204
rect 29932 48850 29988 48860
rect 30044 50036 30100 50046
rect 29148 47294 29150 47346
rect 29202 47294 29204 47346
rect 29148 47124 29204 47294
rect 29260 47404 29652 47460
rect 30044 48804 30100 49980
rect 30156 49922 30212 49934
rect 30156 49870 30158 49922
rect 30210 49870 30212 49922
rect 30156 49812 30212 49870
rect 30156 49746 30212 49756
rect 30044 48242 30100 48748
rect 30044 48190 30046 48242
rect 30098 48190 30100 48242
rect 30044 47458 30100 48190
rect 30044 47406 30046 47458
rect 30098 47406 30100 47458
rect 29260 47346 29316 47404
rect 30044 47394 30100 47406
rect 29260 47294 29262 47346
rect 29314 47294 29316 47346
rect 29260 47282 29316 47294
rect 29148 47058 29204 47068
rect 30156 47124 30212 47134
rect 30156 46788 30212 47068
rect 30156 46722 30212 46732
rect 29148 46676 29204 46686
rect 29148 44324 29204 46620
rect 30268 46564 30324 50372
rect 30492 50148 30548 50158
rect 30492 50034 30548 50092
rect 30492 49982 30494 50034
rect 30546 49982 30548 50034
rect 30492 49970 30548 49982
rect 30940 50148 30996 50158
rect 30716 49026 30772 49038
rect 30716 48974 30718 49026
rect 30770 48974 30772 49026
rect 30380 48804 30436 48814
rect 30716 48804 30772 48974
rect 30940 48914 30996 50092
rect 30940 48862 30942 48914
rect 30994 48862 30996 48914
rect 30940 48850 30996 48862
rect 31500 49812 31556 49822
rect 30380 48802 30772 48804
rect 30380 48750 30382 48802
rect 30434 48750 30772 48802
rect 30380 48748 30772 48750
rect 30380 48738 30436 48748
rect 30716 48692 30772 48748
rect 31388 48804 31444 48814
rect 31388 48710 31444 48748
rect 30716 48636 31332 48692
rect 30716 48466 30772 48478
rect 30716 48414 30718 48466
rect 30770 48414 30772 48466
rect 30380 48244 30436 48254
rect 30380 48150 30436 48188
rect 30716 47570 30772 48414
rect 30940 48356 30996 48366
rect 30716 47518 30718 47570
rect 30770 47518 30772 47570
rect 30716 47506 30772 47518
rect 30828 48242 30884 48254
rect 30828 48190 30830 48242
rect 30882 48190 30884 48242
rect 30828 46788 30884 48190
rect 30940 48242 30996 48300
rect 30940 48190 30942 48242
rect 30994 48190 30996 48242
rect 30940 48178 30996 48190
rect 30828 46722 30884 46732
rect 30940 46676 30996 46686
rect 30940 46582 30996 46620
rect 30380 46564 30436 46574
rect 30268 46562 30436 46564
rect 30268 46510 30382 46562
rect 30434 46510 30436 46562
rect 30268 46508 30436 46510
rect 30380 46498 30436 46508
rect 29260 45668 29316 45678
rect 29260 45574 29316 45612
rect 30604 45220 30660 45230
rect 30492 45218 30996 45220
rect 30492 45166 30606 45218
rect 30658 45166 30996 45218
rect 30492 45164 30996 45166
rect 29484 45108 29540 45118
rect 29484 45014 29540 45052
rect 30380 45108 30436 45118
rect 29932 44994 29988 45006
rect 29932 44942 29934 44994
rect 29986 44942 29988 44994
rect 29932 44772 29988 44942
rect 29932 44706 29988 44716
rect 29148 44230 29204 44268
rect 29932 44212 29988 44222
rect 29708 44210 29988 44212
rect 29708 44158 29934 44210
rect 29986 44158 29988 44210
rect 29708 44156 29988 44158
rect 29708 43762 29764 44156
rect 29932 44146 29988 44156
rect 29708 43710 29710 43762
rect 29762 43710 29764 43762
rect 29708 43698 29764 43710
rect 30380 43764 30436 45052
rect 29036 43652 29092 43662
rect 29036 43558 29092 43596
rect 29148 43652 29204 43662
rect 29148 43650 29316 43652
rect 29148 43598 29150 43650
rect 29202 43598 29316 43650
rect 29148 43596 29316 43598
rect 29148 43586 29204 43596
rect 29148 43314 29204 43326
rect 29148 43262 29150 43314
rect 29202 43262 29204 43314
rect 29036 41970 29092 41982
rect 29036 41918 29038 41970
rect 29090 41918 29092 41970
rect 29036 41748 29092 41918
rect 29036 40740 29092 41692
rect 29148 41188 29204 43262
rect 29260 42644 29316 43596
rect 29596 43540 29652 43550
rect 29596 43446 29652 43484
rect 29820 43538 29876 43550
rect 29820 43486 29822 43538
rect 29874 43486 29876 43538
rect 29820 42868 29876 43486
rect 29820 42802 29876 42812
rect 30156 43538 30212 43550
rect 30156 43486 30158 43538
rect 30210 43486 30212 43538
rect 29260 42550 29316 42588
rect 29372 42420 29428 42430
rect 29372 42196 29428 42364
rect 29372 42194 29876 42196
rect 29372 42142 29374 42194
rect 29426 42142 29876 42194
rect 29372 42140 29876 42142
rect 29372 42130 29428 42140
rect 29148 41132 29764 41188
rect 29484 40962 29540 40974
rect 29484 40910 29486 40962
rect 29538 40910 29540 40962
rect 29148 40740 29204 40750
rect 29036 40684 29148 40740
rect 29148 40674 29204 40684
rect 29484 40740 29540 40910
rect 29484 40674 29540 40684
rect 29260 40292 29316 40302
rect 29260 39732 29316 40236
rect 29260 39638 29316 39676
rect 29596 38822 29652 38834
rect 29596 38770 29598 38822
rect 29650 38770 29652 38822
rect 29260 38724 29316 38734
rect 28924 38722 29316 38724
rect 28924 38670 29262 38722
rect 29314 38670 29316 38722
rect 28924 38668 29316 38670
rect 29596 38724 29652 38770
rect 29260 38658 29316 38668
rect 29484 38612 29652 38668
rect 28364 37490 28532 37492
rect 28364 37438 28366 37490
rect 28418 37438 28532 37490
rect 28364 37436 28532 37438
rect 28588 37548 28756 37604
rect 28924 38500 28980 38510
rect 28364 37426 28420 37436
rect 27916 37266 27972 37278
rect 27916 37214 27918 37266
rect 27970 37214 27972 37266
rect 27916 36932 27972 37214
rect 28028 37268 28084 37278
rect 28028 37174 28084 37212
rect 28140 37266 28196 37278
rect 28140 37214 28142 37266
rect 28194 37214 28196 37266
rect 27916 36866 27972 36876
rect 28140 36820 28196 37214
rect 28140 36754 28196 36764
rect 28476 37044 28532 37054
rect 27804 36652 27972 36708
rect 26460 35252 26628 35308
rect 26796 35420 27076 35476
rect 26460 34914 26516 35252
rect 26796 35138 26852 35420
rect 26796 35086 26798 35138
rect 26850 35086 26852 35138
rect 26796 35074 26852 35086
rect 26460 34862 26462 34914
rect 26514 34862 26516 34914
rect 26236 34802 26292 34814
rect 26236 34750 26238 34802
rect 26290 34750 26292 34802
rect 26236 34692 26292 34750
rect 25900 34690 26292 34692
rect 25900 34638 25902 34690
rect 25954 34638 26292 34690
rect 25900 34636 26292 34638
rect 25900 34626 25956 34636
rect 26236 34020 26292 34636
rect 26460 34692 26516 34862
rect 27580 34916 27636 36428
rect 27804 36372 27860 36382
rect 27804 35812 27860 36316
rect 27916 36148 27972 36652
rect 28476 36594 28532 36988
rect 28476 36542 28478 36594
rect 28530 36542 28532 36594
rect 28476 36530 28532 36542
rect 28028 36372 28084 36382
rect 28028 36278 28084 36316
rect 28252 36370 28308 36382
rect 28252 36318 28254 36370
rect 28306 36318 28308 36370
rect 28252 36148 28308 36318
rect 27916 36092 28308 36148
rect 27804 35746 27860 35756
rect 27580 34850 27636 34860
rect 27916 35698 27972 35710
rect 27916 35646 27918 35698
rect 27970 35646 27972 35698
rect 26460 34626 26516 34636
rect 27244 34692 27300 34702
rect 27692 34692 27748 34702
rect 27300 34690 27748 34692
rect 27300 34638 27694 34690
rect 27746 34638 27748 34690
rect 27300 34636 27748 34638
rect 26460 34020 26516 34030
rect 26236 34018 26516 34020
rect 26236 33966 26462 34018
rect 26514 33966 26516 34018
rect 26236 33964 26516 33966
rect 25900 33572 25956 33582
rect 25900 32676 25956 33516
rect 26460 33236 26516 33964
rect 25900 32562 25956 32620
rect 25900 32510 25902 32562
rect 25954 32510 25956 32562
rect 25900 32498 25956 32510
rect 26236 33180 26516 33236
rect 24220 30146 24276 30156
rect 25340 30380 25844 30436
rect 26012 31668 26068 31678
rect 23996 29988 24052 29998
rect 23996 29894 24052 29932
rect 24220 29986 24276 29998
rect 24220 29934 24222 29986
rect 24274 29934 24276 29986
rect 23324 29540 23380 29550
rect 23324 29446 23380 29484
rect 23436 29426 23492 29596
rect 23436 29374 23438 29426
rect 23490 29374 23492 29426
rect 23436 29362 23492 29374
rect 24220 28868 24276 29934
rect 24892 29988 24948 29998
rect 24892 29316 24948 29932
rect 25340 29650 25396 30380
rect 25340 29598 25342 29650
rect 25394 29598 25396 29650
rect 25340 29586 25396 29598
rect 24892 29250 24948 29260
rect 25676 28980 25732 30380
rect 25228 28868 25284 28878
rect 23772 28812 24276 28868
rect 25116 28812 25228 28868
rect 23660 28420 23716 28430
rect 22988 27918 22990 27970
rect 23042 27918 23044 27970
rect 22988 27906 23044 27918
rect 23212 28418 23716 28420
rect 23212 28366 23662 28418
rect 23714 28366 23716 28418
rect 23212 28364 23716 28366
rect 22428 27860 22484 27870
rect 22428 27766 22484 27804
rect 23212 27858 23268 28364
rect 23660 28354 23716 28364
rect 23660 27972 23716 27982
rect 23772 27972 23828 28812
rect 24668 28756 24724 28766
rect 24724 28700 24836 28756
rect 24668 28690 24724 28700
rect 24220 28532 24276 28542
rect 23660 27970 23828 27972
rect 23660 27918 23662 27970
rect 23714 27918 23828 27970
rect 23660 27916 23828 27918
rect 23996 28420 24052 28430
rect 23660 27906 23716 27916
rect 23212 27806 23214 27858
rect 23266 27806 23268 27858
rect 21980 27580 22484 27636
rect 22428 27186 22484 27580
rect 22428 27134 22430 27186
rect 22482 27134 22484 27186
rect 22428 27122 22484 27134
rect 22764 27412 22820 27422
rect 22764 27074 22820 27356
rect 23212 27186 23268 27806
rect 23996 27860 24052 28364
rect 24108 27860 24164 27870
rect 23996 27858 24164 27860
rect 23996 27806 24110 27858
rect 24162 27806 24164 27858
rect 23996 27804 24164 27806
rect 23996 27300 24052 27804
rect 24108 27794 24164 27804
rect 24108 27300 24164 27310
rect 23996 27298 24164 27300
rect 23996 27246 24110 27298
rect 24162 27246 24164 27298
rect 23996 27244 24164 27246
rect 24108 27234 24164 27244
rect 23212 27134 23214 27186
rect 23266 27134 23268 27186
rect 22764 27022 22766 27074
rect 22818 27022 22820 27074
rect 22764 27010 22820 27022
rect 23100 27076 23156 27086
rect 21756 26850 21812 26862
rect 21868 26852 22148 26908
rect 21756 26798 21758 26850
rect 21810 26798 21812 26850
rect 21756 26292 21812 26798
rect 21756 26198 21812 26236
rect 21980 26290 22036 26302
rect 21980 26238 21982 26290
rect 22034 26238 22036 26290
rect 21980 25956 22036 26238
rect 21980 25890 22036 25900
rect 21756 25732 21812 25742
rect 21756 25618 21812 25676
rect 21756 25566 21758 25618
rect 21810 25566 21812 25618
rect 21756 25554 21812 25566
rect 21980 23826 22036 23838
rect 21980 23774 21982 23826
rect 22034 23774 22036 23826
rect 21756 23714 21812 23726
rect 21756 23662 21758 23714
rect 21810 23662 21812 23714
rect 21756 21812 21812 23662
rect 21980 23268 22036 23774
rect 21756 20692 21812 21756
rect 21756 20626 21812 20636
rect 21868 23044 21924 23054
rect 21868 22484 21924 22988
rect 21868 21586 21924 22428
rect 21980 23042 22036 23212
rect 21980 22990 21982 23042
rect 22034 22990 22036 23042
rect 21980 22036 22036 22990
rect 22092 22708 22148 26852
rect 22764 26516 22820 26526
rect 22764 26422 22820 26460
rect 22428 26404 22484 26414
rect 22428 26178 22484 26348
rect 22428 26126 22430 26178
rect 22482 26126 22484 26178
rect 22428 26114 22484 26126
rect 22988 26402 23044 26414
rect 22988 26350 22990 26402
rect 23042 26350 23044 26402
rect 22988 26068 23044 26350
rect 23100 26402 23156 27020
rect 23212 26908 23268 27134
rect 23436 27076 23492 27114
rect 23436 27010 23492 27020
rect 23884 27076 23940 27086
rect 23884 26982 23940 27020
rect 23212 26852 23492 26908
rect 23100 26350 23102 26402
rect 23154 26350 23156 26402
rect 23100 26338 23156 26350
rect 22652 26012 22988 26068
rect 22428 25506 22484 25518
rect 22428 25454 22430 25506
rect 22482 25454 22484 25506
rect 22428 25284 22484 25454
rect 22652 25394 22708 26012
rect 22988 26002 23044 26012
rect 23324 26180 23380 26190
rect 22652 25342 22654 25394
rect 22706 25342 22708 25394
rect 22652 25330 22708 25342
rect 22876 25508 22932 25518
rect 22428 25060 22484 25228
rect 22428 24994 22484 25004
rect 22876 24946 22932 25452
rect 22876 24894 22878 24946
rect 22930 24894 22932 24946
rect 22876 24882 22932 24894
rect 22764 24722 22820 24734
rect 22764 24670 22766 24722
rect 22818 24670 22820 24722
rect 22204 24612 22260 24622
rect 22764 24612 22820 24670
rect 22204 24610 22820 24612
rect 22204 24558 22206 24610
rect 22258 24558 22820 24610
rect 22204 24556 22820 24558
rect 23324 24610 23380 26124
rect 23324 24558 23326 24610
rect 23378 24558 23380 24610
rect 22204 23940 22260 24556
rect 22204 23874 22260 23884
rect 22764 23940 22820 23950
rect 23324 23940 23380 24558
rect 22764 23938 23380 23940
rect 22764 23886 22766 23938
rect 22818 23886 23380 23938
rect 22764 23884 23380 23886
rect 22428 23716 22484 23726
rect 22764 23716 22820 23884
rect 22428 23714 22820 23716
rect 22428 23662 22430 23714
rect 22482 23662 22820 23714
rect 22428 23660 22820 23662
rect 22428 23044 22484 23660
rect 22988 23156 23044 23166
rect 23436 23156 23492 26852
rect 23548 26178 23604 26190
rect 23548 26126 23550 26178
rect 23602 26126 23604 26178
rect 23548 26068 23604 26126
rect 24108 26180 24164 26190
rect 24108 26086 24164 26124
rect 23548 26002 23604 26012
rect 24108 25618 24164 25630
rect 24108 25566 24110 25618
rect 24162 25566 24164 25618
rect 23660 24834 23716 24846
rect 23660 24782 23662 24834
rect 23714 24782 23716 24834
rect 23548 24052 23604 24062
rect 23660 24052 23716 24782
rect 23996 24836 24052 24846
rect 23996 24742 24052 24780
rect 23548 24050 23716 24052
rect 23548 23998 23550 24050
rect 23602 23998 23716 24050
rect 23548 23996 23716 23998
rect 23548 23986 23604 23996
rect 22988 23154 23492 23156
rect 22988 23102 22990 23154
rect 23042 23102 23438 23154
rect 23490 23102 23492 23154
rect 22988 23100 23492 23102
rect 22988 23090 23044 23100
rect 23436 23044 23492 23100
rect 23884 23044 23940 23054
rect 23436 22988 23828 23044
rect 22428 22950 22484 22988
rect 22092 22652 23044 22708
rect 21980 21970 22036 21980
rect 22316 22258 22372 22270
rect 22316 22206 22318 22258
rect 22370 22206 22372 22258
rect 21868 21534 21870 21586
rect 21922 21534 21924 21586
rect 21868 20916 21924 21534
rect 21084 19236 21140 19246
rect 20748 19070 20750 19122
rect 20802 19070 20804 19122
rect 20748 19058 20804 19070
rect 20972 19180 21084 19236
rect 20412 19012 20468 19022
rect 20412 18918 20468 18956
rect 20860 19012 20916 19022
rect 20860 18674 20916 18956
rect 20860 18622 20862 18674
rect 20914 18622 20916 18674
rect 20860 18610 20916 18622
rect 20300 18050 20356 18060
rect 20300 17836 20692 17892
rect 20300 17666 20356 17836
rect 20636 17780 20692 17836
rect 20860 17780 20916 17790
rect 20972 17780 21028 19180
rect 21084 19170 21140 19180
rect 21196 19124 21252 19964
rect 21084 19012 21140 19022
rect 21084 18674 21140 18956
rect 21084 18622 21086 18674
rect 21138 18622 21140 18674
rect 21084 18610 21140 18622
rect 20636 17778 21028 17780
rect 20636 17726 20862 17778
rect 20914 17726 21028 17778
rect 20636 17724 21028 17726
rect 20860 17714 20916 17724
rect 20300 17614 20302 17666
rect 20354 17614 20356 17666
rect 20300 17602 20356 17614
rect 20524 17668 20580 17678
rect 20412 17108 20468 17118
rect 20412 17014 20468 17052
rect 20524 15314 20580 17612
rect 20748 17108 20804 17118
rect 20748 17014 20804 17052
rect 21196 16882 21252 19068
rect 21196 16830 21198 16882
rect 21250 16830 21252 16882
rect 21196 16818 21252 16830
rect 21308 19964 21700 20020
rect 21308 16660 21364 19964
rect 21868 19908 21924 20860
rect 22092 21700 22148 21710
rect 21980 20804 22036 20814
rect 21980 20710 22036 20748
rect 22092 20802 22148 21644
rect 22204 20916 22260 20926
rect 22316 20916 22372 22206
rect 22428 22146 22484 22158
rect 22428 22094 22430 22146
rect 22482 22094 22484 22146
rect 22428 21700 22484 22094
rect 22540 21700 22596 21710
rect 22428 21698 22596 21700
rect 22428 21646 22542 21698
rect 22594 21646 22596 21698
rect 22428 21644 22596 21646
rect 22540 21634 22596 21644
rect 22204 20914 22372 20916
rect 22204 20862 22206 20914
rect 22258 20862 22372 20914
rect 22204 20860 22372 20862
rect 22204 20850 22260 20860
rect 22092 20750 22094 20802
rect 22146 20750 22148 20802
rect 22092 20738 22148 20750
rect 22428 20804 22484 20814
rect 22316 20692 22372 20702
rect 22204 20636 22316 20692
rect 22204 20356 22260 20636
rect 22316 20598 22372 20636
rect 21644 19906 21924 19908
rect 21644 19854 21870 19906
rect 21922 19854 21924 19906
rect 21644 19852 21924 19854
rect 21644 19236 21700 19852
rect 21868 19842 21924 19852
rect 22092 20300 22260 20356
rect 21644 19142 21700 19180
rect 22092 18674 22148 20300
rect 22092 18622 22094 18674
rect 22146 18622 22148 18674
rect 22092 18610 22148 18622
rect 22204 19908 22260 19918
rect 21420 18562 21476 18574
rect 21420 18510 21422 18562
rect 21474 18510 21476 18562
rect 21420 17892 21476 18510
rect 21980 18450 22036 18462
rect 21980 18398 21982 18450
rect 22034 18398 22036 18450
rect 21420 17836 21588 17892
rect 21420 17668 21476 17678
rect 21420 17574 21476 17612
rect 20524 15262 20526 15314
rect 20578 15262 20580 15314
rect 20524 15250 20580 15262
rect 21084 16604 21364 16660
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20188 14130 20244 14140
rect 20300 14532 20356 14542
rect 19836 14074 20100 14084
rect 20188 13636 20244 13646
rect 20188 13074 20244 13580
rect 20188 13022 20190 13074
rect 20242 13022 20244 13074
rect 20188 13010 20244 13022
rect 19404 12962 19572 12964
rect 19404 12910 19406 12962
rect 19458 12910 19572 12962
rect 19404 12908 19572 12910
rect 19628 12962 19684 12974
rect 19628 12910 19630 12962
rect 19682 12910 19684 12962
rect 19404 12898 19460 12908
rect 19180 12850 19348 12852
rect 19180 12798 19182 12850
rect 19234 12798 19348 12850
rect 19180 12796 19348 12798
rect 19180 12786 19236 12796
rect 19068 12738 19124 12750
rect 19068 12686 19070 12738
rect 19122 12686 19124 12738
rect 19068 12628 19124 12686
rect 19068 12562 19124 12572
rect 19180 12292 19236 12302
rect 19180 12198 19236 12236
rect 19292 12290 19348 12796
rect 19628 12628 19684 12910
rect 20300 12962 20356 14476
rect 20300 12910 20302 12962
rect 20354 12910 20356 12962
rect 20300 12898 20356 12910
rect 20076 12740 20132 12750
rect 20076 12738 20244 12740
rect 20076 12686 20078 12738
rect 20130 12686 20244 12738
rect 20076 12684 20244 12686
rect 20076 12674 20132 12684
rect 19292 12238 19294 12290
rect 19346 12238 19348 12290
rect 19292 11284 19348 12238
rect 19516 12572 19684 12628
rect 19836 12572 20100 12582
rect 19516 12290 19572 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19740 12404 19796 12414
rect 19740 12310 19796 12348
rect 19964 12404 20020 12414
rect 20188 12404 20244 12684
rect 19964 12402 20244 12404
rect 19964 12350 19966 12402
rect 20018 12350 20244 12402
rect 19964 12348 20244 12350
rect 19964 12338 20020 12348
rect 19516 12238 19518 12290
rect 19570 12238 19572 12290
rect 19516 12226 19572 12238
rect 19852 12066 19908 12078
rect 19852 12014 19854 12066
rect 19906 12014 19908 12066
rect 19516 11284 19572 11294
rect 19292 11282 19572 11284
rect 19292 11230 19518 11282
rect 19570 11230 19572 11282
rect 19292 11228 19572 11230
rect 19516 11218 19572 11228
rect 19852 11172 19908 12014
rect 19628 11116 19908 11172
rect 20076 11172 20132 12348
rect 20636 12292 20692 12302
rect 20636 12198 20692 12236
rect 20748 12292 20804 12302
rect 20748 12290 20916 12292
rect 20748 12238 20750 12290
rect 20802 12238 20916 12290
rect 20748 12236 20916 12238
rect 20748 12226 20804 12236
rect 20412 12178 20468 12190
rect 20412 12126 20414 12178
rect 20466 12126 20468 12178
rect 20412 11956 20468 12126
rect 20748 11956 20804 11966
rect 20412 11954 20804 11956
rect 20412 11902 20750 11954
rect 20802 11902 20804 11954
rect 20412 11900 20804 11902
rect 20748 11890 20804 11900
rect 20860 11732 20916 12236
rect 20748 11396 20804 11406
rect 20860 11396 20916 11676
rect 20748 11394 20916 11396
rect 20748 11342 20750 11394
rect 20802 11342 20916 11394
rect 20748 11340 20916 11342
rect 20076 11116 20244 11172
rect 19628 10724 19684 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20188 10836 20244 11116
rect 20076 10780 20244 10836
rect 19964 10724 20020 10734
rect 19628 10722 20020 10724
rect 19628 10670 19966 10722
rect 20018 10670 20020 10722
rect 19628 10668 20020 10670
rect 19964 10658 20020 10668
rect 19292 10610 19348 10622
rect 19292 10558 19294 10610
rect 19346 10558 19348 10610
rect 19068 9828 19124 9838
rect 18956 9772 19068 9828
rect 19068 9734 19124 9772
rect 18508 9716 18564 9726
rect 18396 9714 18564 9716
rect 18396 9662 18510 9714
rect 18562 9662 18564 9714
rect 18396 9660 18564 9662
rect 18508 9650 18564 9660
rect 18508 8260 18564 8270
rect 18956 8260 19012 8270
rect 18508 8258 18956 8260
rect 18508 8206 18510 8258
rect 18562 8206 18956 8258
rect 18508 8204 18956 8206
rect 18508 7476 18564 8204
rect 18956 8166 19012 8204
rect 19292 8260 19348 10558
rect 19852 9828 19908 9838
rect 19852 9734 19908 9772
rect 19404 9716 19460 9726
rect 19404 9622 19460 9660
rect 20076 9716 20132 10780
rect 20748 10500 20804 11340
rect 20748 10434 20804 10444
rect 20076 9650 20132 9660
rect 20748 9604 20804 9614
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19516 9156 19572 9166
rect 19516 9062 19572 9100
rect 20188 9044 20244 9054
rect 20748 9044 20804 9548
rect 21084 9380 21140 16604
rect 21532 16100 21588 17836
rect 21532 16034 21588 16044
rect 21756 17108 21812 17118
rect 21756 15876 21812 17052
rect 21980 16884 22036 18398
rect 22204 18450 22260 19852
rect 22316 19796 22372 19806
rect 22316 19346 22372 19740
rect 22316 19294 22318 19346
rect 22370 19294 22372 19346
rect 22316 19282 22372 19294
rect 22316 19124 22372 19134
rect 22316 18674 22372 19068
rect 22316 18622 22318 18674
rect 22370 18622 22372 18674
rect 22316 18610 22372 18622
rect 22204 18398 22206 18450
rect 22258 18398 22260 18450
rect 22204 18386 22260 18398
rect 22428 18450 22484 20748
rect 22540 20690 22596 20702
rect 22540 20638 22542 20690
rect 22594 20638 22596 20690
rect 22540 19236 22596 20638
rect 22540 19170 22596 19180
rect 22428 18398 22430 18450
rect 22482 18398 22484 18450
rect 22092 17892 22148 17902
rect 22092 17778 22148 17836
rect 22092 17726 22094 17778
rect 22146 17726 22148 17778
rect 22092 17714 22148 17726
rect 22428 17108 22484 18398
rect 22428 17042 22484 17052
rect 22876 18340 22932 18350
rect 22876 17668 22932 18284
rect 22876 16996 22932 17612
rect 21980 16098 22036 16828
rect 22540 16994 22932 16996
rect 22540 16942 22878 16994
rect 22930 16942 22932 16994
rect 22540 16940 22932 16942
rect 21980 16046 21982 16098
rect 22034 16046 22036 16098
rect 21980 16034 22036 16046
rect 22204 16100 22260 16110
rect 22204 16006 22260 16044
rect 22428 15986 22484 15998
rect 22428 15934 22430 15986
rect 22482 15934 22484 15986
rect 21868 15876 21924 15886
rect 21756 15874 21924 15876
rect 21756 15822 21870 15874
rect 21922 15822 21924 15874
rect 21756 15820 21924 15822
rect 21868 15810 21924 15820
rect 22092 15874 22148 15886
rect 22092 15822 22094 15874
rect 22146 15822 22148 15874
rect 21196 15202 21252 15214
rect 21196 15150 21198 15202
rect 21250 15150 21252 15202
rect 21196 15148 21252 15150
rect 22092 15148 22148 15822
rect 22428 15316 22484 15934
rect 22428 15250 22484 15260
rect 22540 15148 22596 16940
rect 22876 16930 22932 16940
rect 22764 16772 22820 16782
rect 22988 16772 23044 22652
rect 23436 20916 23492 20926
rect 23436 20822 23492 20860
rect 23660 19908 23716 19918
rect 23660 19814 23716 19852
rect 23548 19796 23604 19806
rect 23772 19796 23828 22988
rect 23884 22950 23940 22988
rect 23884 20916 23940 20926
rect 23884 20802 23940 20860
rect 23884 20750 23886 20802
rect 23938 20750 23940 20802
rect 23884 20738 23940 20750
rect 24108 20356 24164 25566
rect 23996 20300 24164 20356
rect 23884 19796 23940 19806
rect 23772 19740 23884 19796
rect 23548 19702 23604 19740
rect 23884 19730 23940 19740
rect 23996 18452 24052 20300
rect 24108 20132 24164 20142
rect 24220 20132 24276 28476
rect 24668 28418 24724 28430
rect 24668 28366 24670 28418
rect 24722 28366 24724 28418
rect 24556 27746 24612 27758
rect 24556 27694 24558 27746
rect 24610 27694 24612 27746
rect 24332 27074 24388 27086
rect 24332 27022 24334 27074
rect 24386 27022 24388 27074
rect 24332 26180 24388 27022
rect 24556 26516 24612 27694
rect 24556 26450 24612 26460
rect 24668 26404 24724 28366
rect 24556 26180 24612 26190
rect 24332 26178 24612 26180
rect 24332 26126 24558 26178
rect 24610 26126 24612 26178
rect 24332 26124 24612 26126
rect 24556 25844 24612 26124
rect 24556 25778 24612 25788
rect 24556 25508 24612 25518
rect 24668 25508 24724 26348
rect 24780 27074 24836 28700
rect 25116 28754 25172 28812
rect 25228 28802 25284 28812
rect 25676 28866 25732 28924
rect 25676 28814 25678 28866
rect 25730 28814 25732 28866
rect 25676 28802 25732 28814
rect 25116 28702 25118 28754
rect 25170 28702 25172 28754
rect 25116 28690 25172 28702
rect 25900 28644 25956 28654
rect 25900 28530 25956 28588
rect 25900 28478 25902 28530
rect 25954 28478 25956 28530
rect 25900 28466 25956 28478
rect 26012 28532 26068 31612
rect 26012 28466 26068 28476
rect 25788 28418 25844 28430
rect 25788 28366 25790 28418
rect 25842 28366 25844 28418
rect 25788 28084 25844 28366
rect 25788 28028 26068 28084
rect 25564 27916 25844 27972
rect 25564 27858 25620 27916
rect 25564 27806 25566 27858
rect 25618 27806 25620 27858
rect 25564 27794 25620 27806
rect 25676 27746 25732 27758
rect 25676 27694 25678 27746
rect 25730 27694 25732 27746
rect 25676 27300 25732 27694
rect 25452 27244 25732 27300
rect 25452 27186 25508 27244
rect 25452 27134 25454 27186
rect 25506 27134 25508 27186
rect 25452 27122 25508 27134
rect 24780 27022 24782 27074
rect 24834 27022 24836 27074
rect 24780 26180 24836 27022
rect 25228 27076 25284 27086
rect 25228 26514 25284 27020
rect 25788 26908 25844 27916
rect 25900 27860 25956 27870
rect 25900 27766 25956 27804
rect 26012 27858 26068 28028
rect 26012 27806 26014 27858
rect 26066 27806 26068 27858
rect 26012 27794 26068 27806
rect 26236 26908 26292 33180
rect 27244 32788 27300 34636
rect 27692 34626 27748 34636
rect 27916 34356 27972 35646
rect 27916 34290 27972 34300
rect 28028 34244 28084 36092
rect 28140 35700 28196 35710
rect 28476 35700 28532 35710
rect 28140 35698 28532 35700
rect 28140 35646 28142 35698
rect 28194 35646 28478 35698
rect 28530 35646 28532 35698
rect 28140 35644 28532 35646
rect 28140 35634 28196 35644
rect 28476 35634 28532 35644
rect 28140 34916 28196 34926
rect 28140 34822 28196 34860
rect 28028 34178 28084 34188
rect 27804 33458 27860 33470
rect 27804 33406 27806 33458
rect 27858 33406 27860 33458
rect 27804 32900 27860 33406
rect 28588 33460 28644 37548
rect 28924 37490 28980 38444
rect 29484 38162 29540 38612
rect 29484 38110 29486 38162
rect 29538 38110 29540 38162
rect 29484 38098 29540 38110
rect 29708 38050 29764 41132
rect 29820 40514 29876 42140
rect 30044 42084 30100 42094
rect 29932 42028 30044 42084
rect 29932 40626 29988 42028
rect 30044 42018 30100 42028
rect 30044 41524 30100 41534
rect 30044 41188 30100 41468
rect 30156 41300 30212 43486
rect 30268 42868 30324 42878
rect 30268 41970 30324 42812
rect 30380 42642 30436 43708
rect 30380 42590 30382 42642
rect 30434 42590 30436 42642
rect 30380 42578 30436 42590
rect 30492 42420 30548 45164
rect 30604 45154 30660 45164
rect 30940 45108 30996 45164
rect 31164 45108 31220 45118
rect 30940 45106 31220 45108
rect 30940 45054 31166 45106
rect 31218 45054 31220 45106
rect 30940 45052 31220 45054
rect 31164 45042 31220 45052
rect 31276 44772 31332 48636
rect 31500 48354 31556 49756
rect 31500 48302 31502 48354
rect 31554 48302 31556 48354
rect 31500 48290 31556 48302
rect 31724 48244 31780 51996
rect 31836 49698 31892 49710
rect 31836 49646 31838 49698
rect 31890 49646 31892 49698
rect 31836 48804 31892 49646
rect 31836 48738 31892 48748
rect 31612 48242 31780 48244
rect 31612 48190 31726 48242
rect 31778 48190 31780 48242
rect 31612 48188 31780 48190
rect 31388 45332 31444 45342
rect 31388 45218 31444 45276
rect 31388 45166 31390 45218
rect 31442 45166 31444 45218
rect 31388 45154 31444 45166
rect 31612 45108 31668 48188
rect 31724 48178 31780 48188
rect 31948 48242 32004 52892
rect 32060 50708 32116 50718
rect 32060 50706 32228 50708
rect 32060 50654 32062 50706
rect 32114 50654 32228 50706
rect 32060 50652 32228 50654
rect 32060 50642 32116 50652
rect 32172 50372 32228 50652
rect 32172 49812 32228 50316
rect 32172 49718 32228 49756
rect 31948 48190 31950 48242
rect 32002 48190 32004 48242
rect 31948 47796 32004 48190
rect 32172 48020 32228 48030
rect 31948 47730 32004 47740
rect 32060 48018 32228 48020
rect 32060 47966 32174 48018
rect 32226 47966 32228 48018
rect 32060 47964 32228 47966
rect 31836 47012 31892 47022
rect 31836 46898 31892 46956
rect 31836 46846 31838 46898
rect 31890 46846 31892 46898
rect 31836 46834 31892 46846
rect 32060 46564 32116 47964
rect 32172 47954 32228 47964
rect 32172 47012 32228 47022
rect 32172 46786 32228 46956
rect 32172 46734 32174 46786
rect 32226 46734 32228 46786
rect 32172 46722 32228 46734
rect 32284 46788 32340 46798
rect 32284 46694 32340 46732
rect 31948 46508 32340 46564
rect 31724 46116 31780 46126
rect 31724 46004 31780 46060
rect 31724 46002 31892 46004
rect 31724 45950 31726 46002
rect 31778 45950 31892 46002
rect 31724 45948 31892 45950
rect 31724 45938 31780 45948
rect 31724 45108 31780 45118
rect 31612 45052 31724 45108
rect 31724 45014 31780 45052
rect 31500 44996 31556 45006
rect 31500 44902 31556 44940
rect 31276 44716 31780 44772
rect 30716 42644 30772 42654
rect 31276 42644 31332 42654
rect 30716 42642 31332 42644
rect 30716 42590 30718 42642
rect 30770 42590 31278 42642
rect 31330 42590 31332 42642
rect 30716 42588 31332 42590
rect 30716 42578 30772 42588
rect 30268 41918 30270 41970
rect 30322 41918 30324 41970
rect 30268 41906 30324 41918
rect 30380 42364 30548 42420
rect 30268 41748 30324 41758
rect 30380 41748 30436 42364
rect 30716 42084 30772 42094
rect 30716 41990 30772 42028
rect 31276 42084 31332 42588
rect 31276 42018 31332 42028
rect 30492 41972 30548 41982
rect 30492 41878 30548 41916
rect 30940 41972 30996 41982
rect 30940 41878 30996 41916
rect 30828 41858 30884 41870
rect 30828 41806 30830 41858
rect 30882 41806 30884 41858
rect 30324 41692 30436 41748
rect 30716 41748 30772 41758
rect 30268 41682 30324 41692
rect 30156 41244 30324 41300
rect 30044 41186 30212 41188
rect 30044 41134 30046 41186
rect 30098 41134 30212 41186
rect 30044 41132 30212 41134
rect 30044 41122 30100 41132
rect 29932 40574 29934 40626
rect 29986 40574 29988 40626
rect 29932 40562 29988 40574
rect 30044 40852 30100 40862
rect 29820 40462 29822 40514
rect 29874 40462 29876 40514
rect 29820 40450 29876 40462
rect 30044 40402 30100 40796
rect 30044 40350 30046 40402
rect 30098 40350 30100 40402
rect 30044 40338 30100 40350
rect 29932 40292 29988 40302
rect 29932 38668 29988 40236
rect 30156 39956 30212 41132
rect 30156 39890 30212 39900
rect 30268 39732 30324 41244
rect 30716 41188 30772 41692
rect 30828 41412 30884 41806
rect 31388 41860 31444 41870
rect 31388 41766 31444 41804
rect 30828 41356 31444 41412
rect 31388 41298 31444 41356
rect 31388 41246 31390 41298
rect 31442 41246 31444 41298
rect 31388 41234 31444 41246
rect 30716 41094 30772 41132
rect 30940 40852 30996 40862
rect 30940 40628 30996 40796
rect 30828 40626 30996 40628
rect 30828 40574 30942 40626
rect 30994 40574 30996 40626
rect 30828 40572 30996 40574
rect 30716 40514 30772 40526
rect 30716 40462 30718 40514
rect 30770 40462 30772 40514
rect 30268 39666 30324 39676
rect 30380 40404 30436 40414
rect 30716 40404 30772 40462
rect 30380 40402 30772 40404
rect 30380 40350 30382 40402
rect 30434 40350 30772 40402
rect 30380 40348 30772 40350
rect 30268 39060 30324 39070
rect 30380 39060 30436 40348
rect 30828 39844 30884 40572
rect 30940 40562 30996 40572
rect 31612 40852 31668 40862
rect 31612 40626 31668 40796
rect 31612 40574 31614 40626
rect 31666 40574 31668 40626
rect 31612 40562 31668 40574
rect 31276 40402 31332 40414
rect 31276 40350 31278 40402
rect 31330 40350 31332 40402
rect 31052 40180 31108 40190
rect 31052 40086 31108 40124
rect 30604 39788 30828 39844
rect 30604 39730 30660 39788
rect 30828 39750 30884 39788
rect 30604 39678 30606 39730
rect 30658 39678 30660 39730
rect 30604 39666 30660 39678
rect 31164 39732 31220 39742
rect 30324 39004 30436 39060
rect 30268 38994 30324 39004
rect 30380 38722 30436 38734
rect 30380 38670 30382 38722
rect 30434 38670 30436 38722
rect 30380 38668 30436 38670
rect 29932 38612 30212 38668
rect 29708 37998 29710 38050
rect 29762 37998 29764 38050
rect 29708 37986 29764 37998
rect 30156 38164 30212 38612
rect 30156 38050 30212 38108
rect 30268 38612 30436 38668
rect 30268 38162 30324 38612
rect 31164 38276 31220 39676
rect 30940 38220 31220 38276
rect 30268 38110 30270 38162
rect 30322 38110 30324 38162
rect 30268 38098 30324 38110
rect 30828 38164 30884 38174
rect 30828 38070 30884 38108
rect 30156 37998 30158 38050
rect 30210 37998 30212 38050
rect 30156 37986 30212 37998
rect 30716 38052 30772 38062
rect 30492 37940 30548 37950
rect 28924 37438 28926 37490
rect 28978 37438 28980 37490
rect 28924 37426 28980 37438
rect 29036 37828 29092 37838
rect 30380 37828 30436 37838
rect 29036 37490 29092 37772
rect 29036 37438 29038 37490
rect 29090 37438 29092 37490
rect 29036 37426 29092 37438
rect 30268 37826 30436 37828
rect 30268 37774 30382 37826
rect 30434 37774 30436 37826
rect 30268 37772 30436 37774
rect 29148 37380 29204 37390
rect 28812 37268 28868 37278
rect 28700 36484 28756 36494
rect 28812 36484 28868 37212
rect 28700 36482 28868 36484
rect 28700 36430 28702 36482
rect 28754 36430 28868 36482
rect 28700 36428 28868 36430
rect 28700 36418 28756 36428
rect 28700 36260 28756 36270
rect 29148 36260 29204 37324
rect 29260 37378 29316 37390
rect 29260 37326 29262 37378
rect 29314 37326 29316 37378
rect 29260 37044 29316 37326
rect 30268 37044 30324 37772
rect 30380 37762 30436 37772
rect 30380 37492 30436 37502
rect 30492 37492 30548 37884
rect 30380 37490 30548 37492
rect 30380 37438 30382 37490
rect 30434 37438 30548 37490
rect 30380 37436 30548 37438
rect 30716 37490 30772 37996
rect 30716 37438 30718 37490
rect 30770 37438 30772 37490
rect 30380 37426 30436 37436
rect 29260 36978 29316 36988
rect 30156 36988 30324 37044
rect 30044 36932 30100 36942
rect 30044 36370 30100 36876
rect 30044 36318 30046 36370
rect 30098 36318 30100 36370
rect 28756 36204 29204 36260
rect 29708 36260 29764 36270
rect 28700 35922 28756 36204
rect 28700 35870 28702 35922
rect 28754 35870 28756 35922
rect 28700 35858 28756 35870
rect 28812 35698 28868 35710
rect 28812 35646 28814 35698
rect 28866 35646 28868 35698
rect 28812 34692 28868 35646
rect 29036 35588 29092 35598
rect 28812 34626 28868 34636
rect 28924 35364 28980 35374
rect 28588 33404 28756 33460
rect 27804 32834 27860 32844
rect 28476 33234 28532 33246
rect 28476 33182 28478 33234
rect 28530 33182 28532 33234
rect 27020 32732 27300 32788
rect 28476 32788 28532 33182
rect 28588 33236 28644 33246
rect 28588 33142 28644 33180
rect 26460 32674 26516 32686
rect 26460 32622 26462 32674
rect 26514 32622 26516 32674
rect 26460 31890 26516 32622
rect 26796 32562 26852 32574
rect 26796 32510 26798 32562
rect 26850 32510 26852 32562
rect 26460 31838 26462 31890
rect 26514 31838 26516 31890
rect 26460 31826 26516 31838
rect 26684 32004 26740 32014
rect 26572 29426 26628 29438
rect 26572 29374 26574 29426
rect 26626 29374 26628 29426
rect 26348 29316 26404 29326
rect 26572 29316 26628 29374
rect 26348 29314 26628 29316
rect 26348 29262 26350 29314
rect 26402 29262 26628 29314
rect 26348 29260 26628 29262
rect 26348 28756 26404 29260
rect 26684 28868 26740 31948
rect 26796 31218 26852 32510
rect 26796 31166 26798 31218
rect 26850 31166 26852 31218
rect 26796 31154 26852 31166
rect 26348 28690 26404 28700
rect 26572 28756 26628 28766
rect 26460 28644 26516 28654
rect 26572 28644 26628 28700
rect 26516 28588 26628 28644
rect 26460 28550 26516 28588
rect 26684 28082 26740 28812
rect 26684 28030 26686 28082
rect 26738 28030 26740 28082
rect 26684 27860 26740 28030
rect 26684 27794 26740 27804
rect 26796 28980 26852 28990
rect 26796 26908 26852 28924
rect 27020 28756 27076 32732
rect 28476 32722 28532 32732
rect 27244 32450 27300 32462
rect 27244 32398 27246 32450
rect 27298 32398 27300 32450
rect 27244 32340 27300 32398
rect 27244 32274 27300 32284
rect 28588 31892 28644 31902
rect 28588 31798 28644 31836
rect 27804 31106 27860 31118
rect 27804 31054 27806 31106
rect 27858 31054 27860 31106
rect 27132 30772 27188 30782
rect 27132 30770 27300 30772
rect 27132 30718 27134 30770
rect 27186 30718 27300 30770
rect 27132 30716 27300 30718
rect 27132 30706 27188 30716
rect 27132 30210 27188 30222
rect 27132 30158 27134 30210
rect 27186 30158 27188 30210
rect 27132 28868 27188 30158
rect 27244 29540 27300 30716
rect 27804 30660 27860 31054
rect 27804 30594 27860 30604
rect 27916 30994 27972 31006
rect 27916 30942 27918 30994
rect 27970 30942 27972 30994
rect 27244 29474 27300 29484
rect 27356 29986 27412 29998
rect 27356 29934 27358 29986
rect 27410 29934 27412 29986
rect 27356 29538 27412 29934
rect 27356 29486 27358 29538
rect 27410 29486 27412 29538
rect 27356 29474 27412 29486
rect 27916 29652 27972 30942
rect 27244 28868 27300 28878
rect 27132 28866 27300 28868
rect 27132 28814 27246 28866
rect 27298 28814 27300 28866
rect 27132 28812 27300 28814
rect 27244 28802 27300 28812
rect 27020 28700 27188 28756
rect 25676 26852 25844 26908
rect 26012 26852 26292 26908
rect 26348 26852 26852 26908
rect 25452 26740 25508 26750
rect 25228 26462 25230 26514
rect 25282 26462 25284 26514
rect 25228 26450 25284 26462
rect 25340 26516 25396 26526
rect 25340 26422 25396 26460
rect 24780 26114 24836 26124
rect 25452 26290 25508 26684
rect 25452 26238 25454 26290
rect 25506 26238 25508 26290
rect 24556 25506 24724 25508
rect 24556 25454 24558 25506
rect 24610 25454 24724 25506
rect 24556 25452 24724 25454
rect 24892 25844 24948 25854
rect 24556 25442 24612 25452
rect 24892 25284 24948 25788
rect 25452 25844 25508 26238
rect 25452 25778 25508 25788
rect 25004 25284 25060 25294
rect 24892 25282 25060 25284
rect 24892 25230 25006 25282
rect 25058 25230 25060 25282
rect 24892 25228 25060 25230
rect 24668 24612 24724 24622
rect 24780 24612 24836 24622
rect 24668 24610 24780 24612
rect 24668 24558 24670 24610
rect 24722 24558 24780 24610
rect 24668 24556 24780 24558
rect 24668 24546 24724 24556
rect 24780 23044 24836 24556
rect 24668 21476 24724 21486
rect 24668 21382 24724 21420
rect 24668 20916 24724 20926
rect 24556 20692 24612 20702
rect 24556 20598 24612 20636
rect 24108 20130 24612 20132
rect 24108 20078 24110 20130
rect 24162 20078 24612 20130
rect 24108 20076 24612 20078
rect 24108 20020 24164 20076
rect 24108 19954 24164 19964
rect 24444 19348 24500 19358
rect 24444 19254 24500 19292
rect 24220 18452 24276 18462
rect 23996 18450 24276 18452
rect 23996 18398 24222 18450
rect 24274 18398 24276 18450
rect 23996 18396 24276 18398
rect 23884 18340 23940 18350
rect 23884 18246 23940 18284
rect 24220 18004 24276 18396
rect 22764 15986 22820 16716
rect 22764 15934 22766 15986
rect 22818 15934 22820 15986
rect 22764 15922 22820 15934
rect 22876 16716 23044 16772
rect 24108 17948 24220 18004
rect 21196 15092 21588 15148
rect 21532 14754 21588 15092
rect 21532 14702 21534 14754
rect 21586 14702 21588 14754
rect 21532 14690 21588 14702
rect 21644 15092 22148 15148
rect 22428 15092 22596 15148
rect 21644 14642 21700 15092
rect 21644 14590 21646 14642
rect 21698 14590 21700 14642
rect 21644 14578 21700 14590
rect 22428 14530 22484 15092
rect 22428 14478 22430 14530
rect 22482 14478 22484 14530
rect 22092 14308 22148 14318
rect 22092 14306 22260 14308
rect 22092 14254 22094 14306
rect 22146 14254 22260 14306
rect 22092 14252 22260 14254
rect 22092 14242 22148 14252
rect 22204 13746 22260 14252
rect 22204 13694 22206 13746
rect 22258 13694 22260 13746
rect 21532 13636 21588 13646
rect 21532 13542 21588 13580
rect 22204 13636 22260 13694
rect 22428 13636 22484 14478
rect 22876 13972 22932 16716
rect 23996 16660 24052 16670
rect 22988 16100 23044 16110
rect 22988 15204 23044 16044
rect 23660 16100 23716 16110
rect 23660 16006 23716 16044
rect 23772 15988 23828 15998
rect 22988 15138 23044 15148
rect 23100 15876 23156 15886
rect 23100 14084 23156 15820
rect 23660 15428 23716 15438
rect 23212 15426 23716 15428
rect 23212 15374 23662 15426
rect 23714 15374 23716 15426
rect 23212 15372 23716 15374
rect 23212 14642 23268 15372
rect 23660 15362 23716 15372
rect 23324 15204 23380 15242
rect 23324 15138 23380 15148
rect 23212 14590 23214 14642
rect 23266 14590 23268 14642
rect 23212 14578 23268 14590
rect 23100 14018 23156 14028
rect 22876 13906 22932 13916
rect 22764 13636 22820 13646
rect 22204 13634 22820 13636
rect 22204 13582 22766 13634
rect 22818 13582 22820 13634
rect 22204 13580 22820 13582
rect 21868 12180 21924 12190
rect 22204 12180 22260 13580
rect 22764 13570 22820 13580
rect 22540 12740 22596 12750
rect 22540 12290 22596 12684
rect 22540 12238 22542 12290
rect 22594 12238 22596 12290
rect 22540 12226 22596 12238
rect 21868 12178 22260 12180
rect 21868 12126 21870 12178
rect 21922 12126 22260 12178
rect 21868 12124 22260 12126
rect 21868 9604 21924 12124
rect 23772 10612 23828 15932
rect 23996 15426 24052 16604
rect 23996 15374 23998 15426
rect 24050 15374 24052 15426
rect 23996 15362 24052 15374
rect 24108 15148 24164 17948
rect 24220 17938 24276 17948
rect 24444 18340 24500 18350
rect 24220 17780 24276 17790
rect 24220 17778 24388 17780
rect 24220 17726 24222 17778
rect 24274 17726 24388 17778
rect 24220 17724 24388 17726
rect 24220 17714 24276 17724
rect 24332 16882 24388 17724
rect 24332 16830 24334 16882
rect 24386 16830 24388 16882
rect 24332 16210 24388 16830
rect 24332 16158 24334 16210
rect 24386 16158 24388 16210
rect 24332 16146 24388 16158
rect 24444 15538 24500 18284
rect 24556 16324 24612 20076
rect 24668 18450 24724 20860
rect 24668 18398 24670 18450
rect 24722 18398 24724 18450
rect 24668 18386 24724 18398
rect 24780 17556 24836 22988
rect 24780 17490 24836 17500
rect 24668 16994 24724 17006
rect 24668 16942 24670 16994
rect 24722 16942 24724 16994
rect 24668 16772 24724 16942
rect 24668 16706 24724 16716
rect 24668 16324 24724 16334
rect 24556 16322 24724 16324
rect 24556 16270 24670 16322
rect 24722 16270 24724 16322
rect 24556 16268 24724 16270
rect 24668 16258 24724 16268
rect 24556 15988 24612 15998
rect 24556 15894 24612 15932
rect 24444 15486 24446 15538
rect 24498 15486 24500 15538
rect 24444 15474 24500 15486
rect 23884 15092 24164 15148
rect 23884 13076 23940 15092
rect 24668 13972 24724 13982
rect 24668 13878 24724 13916
rect 23884 13074 24388 13076
rect 23884 13022 23886 13074
rect 23938 13022 24388 13074
rect 23884 13020 24388 13022
rect 23884 13010 23940 13020
rect 24332 12962 24388 13020
rect 24332 12910 24334 12962
rect 24386 12910 24388 12962
rect 24332 12898 24388 12910
rect 24108 12852 24164 12862
rect 24108 12758 24164 12796
rect 24668 12852 24724 12862
rect 24668 12758 24724 12796
rect 24220 12740 24276 12750
rect 24220 12646 24276 12684
rect 24668 12066 24724 12078
rect 24668 12014 24670 12066
rect 24722 12014 24724 12066
rect 24668 11508 24724 12014
rect 24668 11442 24724 11452
rect 24892 11396 24948 25228
rect 25004 25218 25060 25228
rect 25676 24946 25732 26852
rect 25900 26292 25956 26302
rect 25900 25844 25956 26236
rect 25900 25778 25956 25788
rect 25676 24894 25678 24946
rect 25730 24894 25732 24946
rect 25676 24882 25732 24894
rect 25452 24722 25508 24734
rect 25452 24670 25454 24722
rect 25506 24670 25508 24722
rect 25452 24612 25508 24670
rect 25452 24546 25508 24556
rect 25900 24722 25956 24734
rect 25900 24670 25902 24722
rect 25954 24670 25956 24722
rect 25900 24276 25956 24670
rect 25900 24210 25956 24220
rect 25676 24050 25732 24062
rect 25676 23998 25678 24050
rect 25730 23998 25732 24050
rect 25676 23940 25732 23998
rect 26012 24052 26068 26852
rect 26236 26178 26292 26190
rect 26236 26126 26238 26178
rect 26290 26126 26292 26178
rect 26236 25844 26292 26126
rect 26236 25778 26292 25788
rect 26236 25508 26292 25518
rect 26236 25414 26292 25452
rect 26124 25284 26180 25294
rect 26124 24834 26180 25228
rect 26124 24782 26126 24834
rect 26178 24782 26180 24834
rect 26124 24770 26180 24782
rect 26236 24388 26292 24398
rect 26012 23996 26180 24052
rect 25676 23874 25732 23884
rect 26012 23826 26068 23838
rect 26012 23774 26014 23826
rect 26066 23774 26068 23826
rect 25340 22482 25396 22494
rect 25340 22430 25342 22482
rect 25394 22430 25396 22482
rect 25340 21924 25396 22430
rect 25340 21858 25396 21868
rect 25788 22146 25844 22158
rect 25788 22094 25790 22146
rect 25842 22094 25844 22146
rect 25788 21588 25844 22094
rect 26012 21812 26068 23774
rect 26012 21746 26068 21756
rect 26012 21588 26068 21598
rect 25788 21586 26068 21588
rect 25788 21534 26014 21586
rect 26066 21534 26068 21586
rect 25788 21532 26068 21534
rect 25340 21474 25396 21486
rect 25340 21422 25342 21474
rect 25394 21422 25396 21474
rect 25340 20916 25396 21422
rect 26012 21476 26068 21532
rect 26012 21410 26068 21420
rect 25340 20850 25396 20860
rect 25564 21364 25620 21374
rect 25228 19346 25284 19358
rect 25228 19294 25230 19346
rect 25282 19294 25284 19346
rect 25228 19236 25284 19294
rect 25228 19170 25284 19180
rect 25228 18452 25284 18462
rect 25228 18358 25284 18396
rect 25452 18450 25508 18462
rect 25452 18398 25454 18450
rect 25506 18398 25508 18450
rect 25340 18338 25396 18350
rect 25340 18286 25342 18338
rect 25394 18286 25396 18338
rect 25340 18228 25396 18286
rect 25004 18172 25396 18228
rect 25004 17892 25060 18172
rect 25228 18004 25284 18014
rect 25452 18004 25508 18398
rect 25284 17948 25508 18004
rect 25228 17938 25284 17948
rect 25564 17892 25620 21308
rect 25788 20020 25844 20030
rect 25676 20018 25844 20020
rect 25676 19966 25790 20018
rect 25842 19966 25844 20018
rect 25676 19964 25844 19966
rect 25676 19348 25732 19964
rect 25788 19954 25844 19964
rect 26012 19348 26068 19358
rect 25676 19234 25732 19292
rect 25676 19182 25678 19234
rect 25730 19182 25732 19234
rect 25676 19170 25732 19182
rect 25788 19346 26068 19348
rect 25788 19294 26014 19346
rect 26066 19294 26068 19346
rect 25788 19292 26068 19294
rect 25788 18562 25844 19292
rect 26012 19282 26068 19292
rect 26124 19124 26180 23996
rect 26236 23938 26292 24332
rect 26236 23886 26238 23938
rect 26290 23886 26292 23938
rect 26236 21476 26292 23886
rect 26236 21410 26292 21420
rect 26348 19460 26404 26852
rect 26796 25508 26852 25518
rect 26684 25452 26796 25508
rect 26684 24162 26740 25452
rect 26796 25414 26852 25452
rect 26908 25396 26964 25406
rect 26908 25302 26964 25340
rect 27132 25172 27188 28700
rect 27580 28642 27636 28654
rect 27580 28590 27582 28642
rect 27634 28590 27636 28642
rect 27580 27860 27636 28590
rect 27916 28644 27972 29596
rect 28028 28644 28084 28654
rect 27916 28642 28084 28644
rect 27916 28590 28030 28642
rect 28082 28590 28084 28642
rect 27916 28588 28084 28590
rect 28028 28578 28084 28588
rect 28364 28644 28420 28654
rect 28364 28530 28420 28588
rect 28364 28478 28366 28530
rect 28418 28478 28420 28530
rect 28364 28466 28420 28478
rect 28364 28084 28420 28094
rect 28364 27990 28420 28028
rect 28588 27972 28644 27982
rect 28588 27878 28644 27916
rect 27580 27794 27636 27804
rect 28700 27858 28756 33404
rect 28924 31668 28980 35308
rect 29036 35138 29092 35532
rect 29708 35364 29764 36204
rect 30044 36148 30100 36318
rect 30044 36082 30100 36092
rect 30156 35812 30212 36988
rect 30716 36932 30772 37438
rect 30716 36866 30772 36876
rect 30940 36594 30996 38220
rect 31276 36932 31332 40350
rect 31612 39508 31668 39518
rect 31388 39506 31668 39508
rect 31388 39454 31614 39506
rect 31666 39454 31668 39506
rect 31388 39452 31668 39454
rect 31388 39394 31444 39452
rect 31612 39442 31668 39452
rect 31388 39342 31390 39394
rect 31442 39342 31444 39394
rect 31388 38388 31444 39342
rect 31388 38322 31444 38332
rect 31388 37940 31444 37950
rect 31724 37940 31780 44716
rect 31836 44436 31892 45948
rect 31948 45220 32004 46508
rect 32284 46450 32340 46508
rect 32284 46398 32286 46450
rect 32338 46398 32340 46450
rect 32284 46386 32340 46398
rect 32060 46116 32116 46126
rect 32396 46116 32452 56030
rect 33180 55412 33236 55422
rect 32508 54516 32564 54526
rect 32508 54514 32676 54516
rect 32508 54462 32510 54514
rect 32562 54462 32676 54514
rect 32508 54460 32676 54462
rect 32508 54450 32564 54460
rect 32620 53284 32676 54460
rect 33180 54514 33236 55356
rect 33628 55188 33684 59200
rect 35980 56082 36036 56094
rect 35980 56030 35982 56082
rect 36034 56030 36036 56082
rect 35308 55972 35364 55982
rect 35980 55972 36036 56030
rect 35308 55970 36036 55972
rect 35308 55918 35310 55970
rect 35362 55918 36036 55970
rect 35308 55916 36036 55918
rect 35308 55860 35364 55916
rect 35084 55804 35364 55860
rect 33740 55412 33796 55422
rect 35084 55412 35140 55804
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35756 55524 35812 55534
rect 35756 55430 35812 55468
rect 33740 55318 33796 55356
rect 34972 55356 35140 55412
rect 35980 55412 36036 55916
rect 36316 55412 36372 59200
rect 36764 55970 36820 55982
rect 36764 55918 36766 55970
rect 36818 55918 36820 55970
rect 36764 55524 36820 55918
rect 36764 55458 36820 55468
rect 36316 55356 36484 55412
rect 33628 55132 33796 55188
rect 33628 54852 33684 54862
rect 33180 54462 33182 54514
rect 33234 54462 33236 54514
rect 33180 53844 33236 54462
rect 33292 54628 33348 54638
rect 33292 54514 33348 54572
rect 33628 54626 33684 54796
rect 33628 54574 33630 54626
rect 33682 54574 33684 54626
rect 33628 54562 33684 54574
rect 33292 54462 33294 54514
rect 33346 54462 33348 54514
rect 33292 54292 33348 54462
rect 33516 54404 33572 54414
rect 33516 54310 33572 54348
rect 33740 54292 33796 55132
rect 34188 55076 34244 55086
rect 34076 55074 34244 55076
rect 34076 55022 34190 55074
rect 34242 55022 34244 55074
rect 34076 55020 34244 55022
rect 33964 54404 34020 54414
rect 33964 54310 34020 54348
rect 33292 54226 33348 54236
rect 33628 54236 33796 54292
rect 33180 53778 33236 53788
rect 33516 53842 33572 53854
rect 33516 53790 33518 53842
rect 33570 53790 33572 53842
rect 32732 53284 32788 53294
rect 32620 53228 32732 53284
rect 32732 53218 32788 53228
rect 33516 53284 33572 53790
rect 33628 53732 33684 54236
rect 33852 53732 33908 53742
rect 34076 53732 34132 55020
rect 34188 55010 34244 55020
rect 34636 55076 34692 55086
rect 34412 54852 34468 54862
rect 34188 54740 34244 54750
rect 34188 54646 34244 54684
rect 34188 54404 34244 54414
rect 34188 54310 34244 54348
rect 33628 53666 33684 53676
rect 33740 53730 34132 53732
rect 33740 53678 33854 53730
rect 33906 53678 34132 53730
rect 33740 53676 34132 53678
rect 34188 53844 34244 53854
rect 33516 53218 33572 53228
rect 32508 53172 32564 53182
rect 32508 53078 32564 53116
rect 33292 53172 33348 53182
rect 33292 52162 33348 53116
rect 33292 52110 33294 52162
rect 33346 52110 33348 52162
rect 33292 52098 33348 52110
rect 33516 52946 33572 52958
rect 33516 52894 33518 52946
rect 33570 52894 33572 52946
rect 33068 52052 33124 52062
rect 33068 51602 33124 51996
rect 33068 51550 33070 51602
rect 33122 51550 33124 51602
rect 33068 51538 33124 51550
rect 33292 51378 33348 51390
rect 33292 51326 33294 51378
rect 33346 51326 33348 51378
rect 32508 51268 32564 51278
rect 33292 51268 33348 51326
rect 32508 51266 33348 51268
rect 32508 51214 32510 51266
rect 32562 51214 33348 51266
rect 32508 51212 33348 51214
rect 32508 50596 32564 51212
rect 32620 50596 32676 50606
rect 32508 50594 32676 50596
rect 32508 50542 32622 50594
rect 32674 50542 32676 50594
rect 32508 50540 32676 50542
rect 32620 50530 32676 50540
rect 32732 50482 32788 50494
rect 32732 50430 32734 50482
rect 32786 50430 32788 50482
rect 32732 50372 32788 50430
rect 32732 50306 32788 50316
rect 32060 45778 32116 46060
rect 32060 45726 32062 45778
rect 32114 45726 32116 45778
rect 32060 45714 32116 45726
rect 32172 46060 32452 46116
rect 32508 49924 32564 49934
rect 31948 45106 32004 45164
rect 31948 45054 31950 45106
rect 32002 45054 32004 45106
rect 31948 45042 32004 45054
rect 31836 44370 31892 44380
rect 32060 44436 32116 44446
rect 32172 44436 32228 46060
rect 32508 46004 32564 49868
rect 33292 49698 33348 49710
rect 33292 49646 33294 49698
rect 33346 49646 33348 49698
rect 32956 49026 33012 49038
rect 32956 48974 32958 49026
rect 33010 48974 33012 49026
rect 32956 48916 33012 48974
rect 33068 48916 33124 48926
rect 32956 48860 33068 48916
rect 33068 48850 33124 48860
rect 33180 48692 33236 48702
rect 33180 48242 33236 48636
rect 33180 48190 33182 48242
rect 33234 48190 33236 48242
rect 33180 48178 33236 48190
rect 32620 48020 32676 48030
rect 32620 48018 33236 48020
rect 32620 47966 32622 48018
rect 32674 47966 33236 48018
rect 32620 47964 33236 47966
rect 32620 47954 32676 47964
rect 32844 47796 32900 47806
rect 32900 47740 33012 47796
rect 32844 47730 32900 47740
rect 32844 47570 32900 47582
rect 32844 47518 32846 47570
rect 32898 47518 32900 47570
rect 32844 46452 32900 47518
rect 32844 46386 32900 46396
rect 32284 45948 32564 46004
rect 32284 45890 32340 45948
rect 32284 45838 32286 45890
rect 32338 45838 32340 45890
rect 32284 45332 32340 45838
rect 32284 45266 32340 45276
rect 32396 45666 32452 45678
rect 32396 45614 32398 45666
rect 32450 45614 32452 45666
rect 32396 44996 32452 45614
rect 32508 45666 32564 45678
rect 32508 45614 32510 45666
rect 32562 45614 32564 45666
rect 32508 45220 32564 45614
rect 32508 45154 32564 45164
rect 32956 45108 33012 47740
rect 33180 47458 33236 47964
rect 33292 47682 33348 49646
rect 33292 47630 33294 47682
rect 33346 47630 33348 47682
rect 33292 47618 33348 47630
rect 33404 48916 33460 48926
rect 33180 47406 33182 47458
rect 33234 47406 33236 47458
rect 33180 47394 33236 47406
rect 33292 47234 33348 47246
rect 33292 47182 33294 47234
rect 33346 47182 33348 47234
rect 33180 46564 33236 46574
rect 33292 46564 33348 47182
rect 33180 46562 33348 46564
rect 33180 46510 33182 46562
rect 33234 46510 33348 46562
rect 33180 46508 33348 46510
rect 33180 46498 33236 46508
rect 33180 45108 33236 45118
rect 32956 45052 33124 45108
rect 32396 44940 33012 44996
rect 32060 44434 32228 44436
rect 32060 44382 32062 44434
rect 32114 44382 32228 44434
rect 32060 44380 32228 44382
rect 32956 44434 33012 44940
rect 32956 44382 32958 44434
rect 33010 44382 33012 44434
rect 32060 44370 32116 44380
rect 32956 44370 33012 44382
rect 32508 44324 32564 44334
rect 32508 44230 32564 44268
rect 33068 43764 33124 45052
rect 33180 44322 33236 45052
rect 33292 44772 33348 46508
rect 33404 45892 33460 48860
rect 33404 45556 33460 45836
rect 33404 45490 33460 45500
rect 33404 45332 33460 45342
rect 33404 45106 33460 45276
rect 33404 45054 33406 45106
rect 33458 45054 33460 45106
rect 33404 45042 33460 45054
rect 33292 44706 33348 44716
rect 33516 44548 33572 52894
rect 33628 50484 33684 50494
rect 33628 49810 33684 50428
rect 33740 50428 33796 53676
rect 33852 53666 33908 53676
rect 34076 53508 34132 53518
rect 34076 53170 34132 53452
rect 34076 53118 34078 53170
rect 34130 53118 34132 53170
rect 34076 53106 34132 53118
rect 34076 52050 34132 52062
rect 34076 51998 34078 52050
rect 34130 51998 34132 52050
rect 33964 51604 34020 51614
rect 33852 51548 33964 51604
rect 33852 51490 33908 51548
rect 33964 51538 34020 51548
rect 33852 51438 33854 51490
rect 33906 51438 33908 51490
rect 33852 51426 33908 51438
rect 33964 51380 34020 51390
rect 34076 51380 34132 51998
rect 33964 51378 34132 51380
rect 33964 51326 33966 51378
rect 34018 51326 34132 51378
rect 33964 51324 34132 51326
rect 33964 51314 34020 51324
rect 34076 50484 34132 50494
rect 34188 50484 34244 53788
rect 34412 52948 34468 54796
rect 34636 54516 34692 55020
rect 34748 54516 34804 54526
rect 34636 54514 34804 54516
rect 34636 54462 34750 54514
rect 34802 54462 34804 54514
rect 34636 54460 34804 54462
rect 34636 53172 34692 54460
rect 34748 54450 34804 54460
rect 34636 53106 34692 53116
rect 34412 52052 34468 52892
rect 34132 50428 34244 50484
rect 34300 51378 34356 51390
rect 34300 51326 34302 51378
rect 34354 51326 34356 51378
rect 33740 50372 34020 50428
rect 34076 50418 34132 50428
rect 33628 49758 33630 49810
rect 33682 49758 33684 49810
rect 33628 49746 33684 49758
rect 33740 49138 33796 49150
rect 33740 49086 33742 49138
rect 33794 49086 33796 49138
rect 33740 48692 33796 49086
rect 33964 49140 34020 50372
rect 34300 50260 34356 51326
rect 34300 50036 34356 50204
rect 34300 49970 34356 49980
rect 34412 50034 34468 51996
rect 34860 52948 34916 52958
rect 34636 51604 34692 51614
rect 34636 51510 34692 51548
rect 34524 51380 34580 51390
rect 34524 51286 34580 51324
rect 34748 51378 34804 51390
rect 34748 51326 34750 51378
rect 34802 51326 34804 51378
rect 34748 51268 34804 51326
rect 34748 51202 34804 51212
rect 34860 51156 34916 52892
rect 34972 52164 35028 55356
rect 35980 55346 36036 55356
rect 35644 55188 35700 55198
rect 35644 55094 35700 55132
rect 36316 55186 36372 55198
rect 36316 55134 36318 55186
rect 36370 55134 36372 55186
rect 35084 55076 35140 55086
rect 36204 55076 36260 55086
rect 35084 54982 35140 55020
rect 35868 55074 36260 55076
rect 35868 55022 36206 55074
rect 36258 55022 36260 55074
rect 35868 55020 36260 55022
rect 35868 54740 35924 55020
rect 36204 55010 36260 55020
rect 35532 54684 35924 54740
rect 35532 54626 35588 54684
rect 35532 54574 35534 54626
rect 35586 54574 35588 54626
rect 35532 54562 35588 54574
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 36316 53844 36372 55134
rect 36428 55076 36484 55356
rect 36988 55300 37044 59200
rect 37660 55636 37716 59200
rect 38332 55972 38388 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 42812 56082 42868 56094
rect 42812 56030 42814 56082
rect 42866 56030 42868 56082
rect 38332 55906 38388 55916
rect 39004 55970 39060 55982
rect 39004 55918 39006 55970
rect 39058 55918 39060 55970
rect 37660 55580 37940 55636
rect 37100 55412 37156 55422
rect 37100 55318 37156 55356
rect 37660 55412 37716 55422
rect 36988 55234 37044 55244
rect 37660 55300 37716 55356
rect 37660 55298 37828 55300
rect 37660 55246 37662 55298
rect 37714 55246 37828 55298
rect 37660 55244 37828 55246
rect 37660 55234 37716 55244
rect 36428 55010 36484 55020
rect 37660 54402 37716 54414
rect 37660 54350 37662 54402
rect 37714 54350 37716 54402
rect 37660 54068 37716 54350
rect 37772 54292 37828 55244
rect 37884 54740 37940 55580
rect 39004 55468 39060 55918
rect 40012 55970 40068 55982
rect 42140 55972 42196 55982
rect 40012 55918 40014 55970
rect 40066 55918 40068 55970
rect 40012 55468 40068 55918
rect 42028 55970 42196 55972
rect 42028 55918 42142 55970
rect 42194 55918 42196 55970
rect 42028 55916 42196 55918
rect 39004 55412 39172 55468
rect 40012 55412 40180 55468
rect 37884 54674 37940 54684
rect 38332 55188 38388 55198
rect 38332 54738 38388 55132
rect 38444 55188 38500 55198
rect 38444 55186 39060 55188
rect 38444 55134 38446 55186
rect 38498 55134 39060 55186
rect 38444 55132 39060 55134
rect 38444 55122 38500 55132
rect 38332 54686 38334 54738
rect 38386 54686 38388 54738
rect 38332 54674 38388 54686
rect 38780 54964 38836 54974
rect 38220 54628 38276 54638
rect 38220 54534 38276 54572
rect 37996 54516 38052 54526
rect 37772 54226 37828 54236
rect 37884 54514 38052 54516
rect 37884 54462 37998 54514
rect 38050 54462 38052 54514
rect 37884 54460 38052 54462
rect 37884 54404 37940 54460
rect 37996 54450 38052 54460
rect 38444 54514 38500 54526
rect 38444 54462 38446 54514
rect 38498 54462 38500 54514
rect 37716 54012 37828 54068
rect 37660 54002 37716 54012
rect 36316 53778 36372 53788
rect 37660 53844 37716 53854
rect 37660 53750 37716 53788
rect 36988 53732 37044 53742
rect 35420 53620 35476 53630
rect 35420 53526 35476 53564
rect 35868 53284 35924 53294
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 34972 52108 35364 52164
rect 34972 51492 35028 51502
rect 34972 51398 35028 51436
rect 35308 51380 35364 52108
rect 35420 51380 35476 51390
rect 35308 51378 35588 51380
rect 35308 51326 35422 51378
rect 35474 51326 35588 51378
rect 35308 51324 35588 51326
rect 35420 51314 35476 51324
rect 34860 51100 35028 51156
rect 34860 50370 34916 50382
rect 34860 50318 34862 50370
rect 34914 50318 34916 50370
rect 34412 49982 34414 50034
rect 34466 49982 34468 50034
rect 34412 49970 34468 49982
rect 34748 50148 34804 50158
rect 34748 50034 34804 50092
rect 34748 49982 34750 50034
rect 34802 49982 34804 50034
rect 34748 49970 34804 49982
rect 33964 49074 34020 49084
rect 34076 49698 34132 49710
rect 34076 49646 34078 49698
rect 34130 49646 34132 49698
rect 33740 46898 33796 48636
rect 33964 48130 34020 48142
rect 33964 48078 33966 48130
rect 34018 48078 34020 48130
rect 33964 47236 34020 48078
rect 34076 47458 34132 49646
rect 34860 48020 34916 50318
rect 34860 47954 34916 47964
rect 34972 47684 35028 51100
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35308 50484 35364 50522
rect 35308 50418 35364 50428
rect 35196 49700 35252 49710
rect 35532 49700 35588 51324
rect 35868 50428 35924 53228
rect 36988 53170 37044 53676
rect 37772 53730 37828 54012
rect 37772 53678 37774 53730
rect 37826 53678 37828 53730
rect 37772 53666 37828 53678
rect 36988 53118 36990 53170
rect 37042 53118 37044 53170
rect 36988 53106 37044 53118
rect 37212 53506 37268 53518
rect 37212 53454 37214 53506
rect 37266 53454 37268 53506
rect 35980 52948 36036 52958
rect 35980 52854 36036 52892
rect 36316 51938 36372 51950
rect 36316 51886 36318 51938
rect 36370 51886 36372 51938
rect 36316 51492 36372 51886
rect 37212 51828 37268 53454
rect 37660 53508 37716 53518
rect 37884 53508 37940 54348
rect 37660 53506 37940 53508
rect 37660 53454 37662 53506
rect 37714 53454 37940 53506
rect 37660 53452 37940 53454
rect 37996 54180 38052 54190
rect 37996 53506 38052 54124
rect 38444 54180 38500 54462
rect 38444 54114 38500 54124
rect 38556 54514 38612 54526
rect 38556 54462 38558 54514
rect 38610 54462 38612 54514
rect 38556 54068 38612 54462
rect 38780 54516 38836 54908
rect 39004 54738 39060 55132
rect 39116 54964 39172 55412
rect 39116 54898 39172 54908
rect 39788 54740 39844 54750
rect 39004 54686 39006 54738
rect 39058 54686 39060 54738
rect 39004 54674 39060 54686
rect 39116 54738 39844 54740
rect 39116 54686 39790 54738
rect 39842 54686 39844 54738
rect 39116 54684 39844 54686
rect 39116 54626 39172 54684
rect 39788 54674 39844 54684
rect 39116 54574 39118 54626
rect 39170 54574 39172 54626
rect 39116 54562 39172 54574
rect 40124 54628 40180 55412
rect 40124 54534 40180 54572
rect 40572 55410 40628 55422
rect 40572 55358 40574 55410
rect 40626 55358 40628 55410
rect 38556 53844 38612 54012
rect 38556 53778 38612 53788
rect 38668 54292 38724 54302
rect 38220 53620 38276 53630
rect 38220 53526 38276 53564
rect 37996 53454 37998 53506
rect 38050 53454 38052 53506
rect 37324 53060 37380 53070
rect 37324 52162 37380 53004
rect 37324 52110 37326 52162
rect 37378 52110 37380 52162
rect 37324 52098 37380 52110
rect 37660 52050 37716 53452
rect 37996 52836 38052 53454
rect 38668 53506 38724 54236
rect 38668 53454 38670 53506
rect 38722 53454 38724 53506
rect 38668 53172 38724 53454
rect 38668 53106 38724 53116
rect 37996 52770 38052 52780
rect 37660 51998 37662 52050
rect 37714 51998 37716 52050
rect 37660 51986 37716 51998
rect 38556 52052 38612 52062
rect 38780 52052 38836 54460
rect 39564 54514 39620 54526
rect 39564 54462 39566 54514
rect 39618 54462 39620 54514
rect 39564 54404 39620 54462
rect 39564 54338 39620 54348
rect 39676 54514 39732 54526
rect 39676 54462 39678 54514
rect 39730 54462 39732 54514
rect 39676 54068 39732 54462
rect 39900 54516 39956 54526
rect 39900 54422 39956 54460
rect 40572 54068 40628 55358
rect 40908 55300 40964 55310
rect 39676 54012 40628 54068
rect 40796 55298 40964 55300
rect 40796 55246 40910 55298
rect 40962 55246 40964 55298
rect 40796 55244 40964 55246
rect 39900 53844 39956 53854
rect 39116 53732 39172 53742
rect 39116 53638 39172 53676
rect 39788 53620 39844 53630
rect 39340 53618 39844 53620
rect 39340 53566 39790 53618
rect 39842 53566 39844 53618
rect 39340 53564 39844 53566
rect 39340 53172 39396 53564
rect 39788 53554 39844 53564
rect 39900 53396 39956 53788
rect 38556 52050 38836 52052
rect 38556 51998 38558 52050
rect 38610 51998 38836 52050
rect 38556 51996 38836 51998
rect 39116 53116 39396 53172
rect 39676 53340 39956 53396
rect 40012 53620 40068 54012
rect 38556 51986 38612 51996
rect 35980 51436 36372 51492
rect 36988 51492 37044 51502
rect 35980 51380 36036 51436
rect 35980 50596 36036 51324
rect 36092 51268 36148 51278
rect 36092 51266 36932 51268
rect 36092 51214 36094 51266
rect 36146 51214 36932 51266
rect 36092 51212 36932 51214
rect 36092 51202 36148 51212
rect 35980 50530 36036 50540
rect 36428 50594 36484 50606
rect 36428 50542 36430 50594
rect 36482 50542 36484 50594
rect 36428 50428 36484 50542
rect 35868 50372 36484 50428
rect 36540 50596 36596 50606
rect 35980 50036 36036 50046
rect 35980 49942 36036 49980
rect 36316 50036 36372 50046
rect 36316 49942 36372 49980
rect 36092 49812 36148 49822
rect 36092 49718 36148 49756
rect 36540 49812 36596 50540
rect 36876 50034 36932 51212
rect 36876 49982 36878 50034
rect 36930 49982 36932 50034
rect 36876 49970 36932 49982
rect 36988 50594 37044 51436
rect 37212 51268 37268 51772
rect 39116 51716 39172 53116
rect 39228 52946 39284 52958
rect 39228 52894 39230 52946
rect 39282 52894 39284 52946
rect 39228 52052 39284 52894
rect 39564 52948 39620 52958
rect 39676 52948 39732 53340
rect 39564 52946 39732 52948
rect 39564 52894 39566 52946
rect 39618 52894 39732 52946
rect 39564 52892 39732 52894
rect 39788 52948 39844 52958
rect 39788 52946 39956 52948
rect 39788 52894 39790 52946
rect 39842 52894 39956 52946
rect 39788 52892 39956 52894
rect 39228 51986 39284 51996
rect 39340 52834 39396 52846
rect 39340 52782 39342 52834
rect 39394 52782 39396 52834
rect 39004 51660 39172 51716
rect 39004 51602 39060 51660
rect 39004 51550 39006 51602
rect 39058 51550 39060 51602
rect 39004 51538 39060 51550
rect 39116 51492 39172 51502
rect 39340 51492 39396 52782
rect 39564 52162 39620 52892
rect 39788 52276 39844 52892
rect 39900 52834 39956 52892
rect 39900 52782 39902 52834
rect 39954 52782 39956 52834
rect 39900 52770 39956 52782
rect 39564 52110 39566 52162
rect 39618 52110 39620 52162
rect 39564 52098 39620 52110
rect 39676 52220 39844 52276
rect 39116 51490 39396 51492
rect 39116 51438 39118 51490
rect 39170 51438 39396 51490
rect 39116 51436 39396 51438
rect 39452 52052 39508 52062
rect 39452 51490 39508 51996
rect 39452 51438 39454 51490
rect 39506 51438 39508 51490
rect 39116 51426 39172 51436
rect 39452 51426 39508 51438
rect 38780 51380 38836 51390
rect 38780 51286 38836 51324
rect 36988 50542 36990 50594
rect 37042 50542 37044 50594
rect 36988 49924 37044 50542
rect 37100 50708 37156 50718
rect 37100 50482 37156 50652
rect 37100 50430 37102 50482
rect 37154 50430 37156 50482
rect 37100 50418 37156 50430
rect 37212 50036 37268 51212
rect 38332 51266 38388 51278
rect 38332 51214 38334 51266
rect 38386 51214 38388 51266
rect 36988 49868 37156 49924
rect 36540 49810 36708 49812
rect 36540 49758 36542 49810
rect 36594 49758 36708 49810
rect 36540 49756 36708 49758
rect 36540 49746 36596 49756
rect 35084 49698 35588 49700
rect 35084 49646 35198 49698
rect 35250 49646 35588 49698
rect 35084 49644 35588 49646
rect 36204 49700 36260 49710
rect 35084 48692 35140 49644
rect 35196 49634 35252 49644
rect 36204 49606 36260 49644
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35532 48804 35588 48814
rect 36316 48804 36372 48814
rect 35532 48802 35700 48804
rect 35532 48750 35534 48802
rect 35586 48750 35700 48802
rect 35532 48748 35700 48750
rect 35532 48738 35588 48748
rect 35084 48626 35140 48636
rect 35644 48244 35700 48748
rect 36372 48748 36596 48804
rect 36316 48710 36372 48748
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 34076 47406 34078 47458
rect 34130 47406 34132 47458
rect 34076 47394 34132 47406
rect 34748 47628 35028 47684
rect 35532 47684 35588 47694
rect 34188 47236 34244 47246
rect 33964 47234 34244 47236
rect 33964 47182 34190 47234
rect 34242 47182 34244 47234
rect 33964 47180 34244 47182
rect 34188 47170 34244 47180
rect 34300 47236 34356 47246
rect 33740 46846 33742 46898
rect 33794 46846 33796 46898
rect 33740 46834 33796 46846
rect 34076 46788 34132 46798
rect 34076 46694 34132 46732
rect 33964 46674 34020 46686
rect 33964 46622 33966 46674
rect 34018 46622 34020 46674
rect 33964 46452 34020 46622
rect 33964 46386 34020 46396
rect 33964 46004 34020 46014
rect 33852 45332 33908 45342
rect 33740 45276 33852 45332
rect 33180 44270 33182 44322
rect 33234 44270 33236 44322
rect 33180 44258 33236 44270
rect 33292 44492 33572 44548
rect 33628 44996 33684 45006
rect 33068 43698 33124 43708
rect 32956 43540 33012 43550
rect 32508 43538 33012 43540
rect 32508 43486 32958 43538
rect 33010 43486 33012 43538
rect 32508 43484 33012 43486
rect 32508 42756 32564 43484
rect 32956 43474 33012 43484
rect 33292 43316 33348 44492
rect 33628 44100 33684 44940
rect 33404 43764 33460 43774
rect 33404 43650 33460 43708
rect 33628 43762 33684 44044
rect 33628 43710 33630 43762
rect 33682 43710 33684 43762
rect 33628 43698 33684 43710
rect 33404 43598 33406 43650
rect 33458 43598 33460 43650
rect 33404 43586 33460 43598
rect 33516 43652 33572 43662
rect 33516 43558 33572 43596
rect 33740 43540 33796 45276
rect 33852 45266 33908 45276
rect 33852 45106 33908 45118
rect 33852 45054 33854 45106
rect 33906 45054 33908 45106
rect 33852 44996 33908 45054
rect 33852 44930 33908 44940
rect 33964 44324 34020 45948
rect 34300 45444 34356 47180
rect 34524 47236 34580 47246
rect 34524 47142 34580 47180
rect 34300 45388 34692 45444
rect 34412 45220 34468 45230
rect 34412 45126 34468 45164
rect 34524 45218 34580 45230
rect 34524 45166 34526 45218
rect 34578 45166 34580 45218
rect 34524 45108 34580 45166
rect 34076 44996 34132 45006
rect 34524 44996 34580 45052
rect 34076 44994 34356 44996
rect 34076 44942 34078 44994
rect 34130 44942 34356 44994
rect 34076 44940 34356 44942
rect 34076 44930 34132 44940
rect 33964 44258 34020 44268
rect 34076 44660 34132 44670
rect 33852 44212 33908 44222
rect 33852 44118 33908 44156
rect 33628 43484 33796 43540
rect 33628 43428 33684 43484
rect 31948 42754 32564 42756
rect 31948 42702 32510 42754
rect 32562 42702 32564 42754
rect 31948 42700 32564 42702
rect 31948 42194 32004 42700
rect 32508 42690 32564 42700
rect 32620 43260 33348 43316
rect 33516 43372 33684 43428
rect 31948 42142 31950 42194
rect 32002 42142 32004 42194
rect 31948 40626 32004 42142
rect 31948 40574 31950 40626
rect 32002 40574 32004 40626
rect 31948 39506 32004 40574
rect 32396 41972 32452 41982
rect 32284 40180 32340 40190
rect 32284 39618 32340 40124
rect 32396 39842 32452 41916
rect 32508 41076 32564 41086
rect 32508 40404 32564 41020
rect 32508 40310 32564 40348
rect 32396 39790 32398 39842
rect 32450 39790 32452 39842
rect 32396 39778 32452 39790
rect 32284 39566 32286 39618
rect 32338 39566 32340 39618
rect 32284 39554 32340 39566
rect 32508 39620 32564 39630
rect 31948 39454 31950 39506
rect 32002 39454 32004 39506
rect 31948 39442 32004 39454
rect 32396 39396 32452 39406
rect 32396 39302 32452 39340
rect 32508 39284 32564 39564
rect 32508 39218 32564 39228
rect 32508 38724 32564 38734
rect 32620 38724 32676 43260
rect 32732 42644 32788 42654
rect 32732 42550 32788 42588
rect 32508 38722 32676 38724
rect 32508 38670 32510 38722
rect 32562 38670 32676 38722
rect 32508 38668 32676 38670
rect 32844 42084 32900 42094
rect 32844 39732 32900 42028
rect 33516 41298 33572 43372
rect 34076 43316 34132 44604
rect 34188 44210 34244 44222
rect 34188 44158 34190 44210
rect 34242 44158 34244 44210
rect 34188 43652 34244 44158
rect 34188 43586 34244 43596
rect 33516 41246 33518 41298
rect 33570 41246 33572 41298
rect 33516 41234 33572 41246
rect 33628 43260 34132 43316
rect 33628 40516 33684 43260
rect 33740 42868 33796 42878
rect 33740 42642 33796 42812
rect 33740 42590 33742 42642
rect 33794 42590 33796 42642
rect 33740 42578 33796 42590
rect 34076 42642 34132 42654
rect 34076 42590 34078 42642
rect 34130 42590 34132 42642
rect 34076 42532 34132 42590
rect 34188 42532 34244 42542
rect 34076 42476 34188 42532
rect 34188 42466 34244 42476
rect 33740 42196 33796 42206
rect 33740 41748 33796 42140
rect 33796 41692 33908 41748
rect 33740 41682 33796 41692
rect 33628 40460 33796 40516
rect 32508 38658 32564 38668
rect 31836 38388 31892 38398
rect 31836 38164 31892 38332
rect 31836 38162 32228 38164
rect 31836 38110 31838 38162
rect 31890 38110 32228 38162
rect 31836 38108 32228 38110
rect 31836 38098 31892 38108
rect 32172 38050 32228 38108
rect 32172 37998 32174 38050
rect 32226 37998 32228 38050
rect 32172 37986 32228 37998
rect 31444 37884 31780 37940
rect 31388 37490 31444 37884
rect 31388 37438 31390 37490
rect 31442 37438 31444 37490
rect 31388 37426 31444 37438
rect 32508 37826 32564 37838
rect 32508 37774 32510 37826
rect 32562 37774 32564 37826
rect 31836 37156 31892 37166
rect 31724 37154 31892 37156
rect 31724 37102 31838 37154
rect 31890 37102 31892 37154
rect 31724 37100 31892 37102
rect 31276 36876 31556 36932
rect 30940 36542 30942 36594
rect 30994 36542 30996 36594
rect 30940 36530 30996 36542
rect 30380 36484 30436 36494
rect 30828 36484 30884 36494
rect 30380 36482 30884 36484
rect 30380 36430 30382 36482
rect 30434 36430 30830 36482
rect 30882 36430 30884 36482
rect 30380 36428 30884 36430
rect 31500 36484 31556 36876
rect 31612 36484 31668 36494
rect 31500 36428 31612 36484
rect 30380 36418 30436 36428
rect 30268 36258 30324 36270
rect 30268 36206 30270 36258
rect 30322 36206 30324 36258
rect 30268 36148 30324 36206
rect 30268 36082 30324 36092
rect 30492 36258 30548 36270
rect 30492 36206 30494 36258
rect 30546 36206 30548 36258
rect 30492 36036 30548 36206
rect 30492 35970 30548 35980
rect 30268 35812 30324 35822
rect 30156 35810 30324 35812
rect 30156 35758 30270 35810
rect 30322 35758 30324 35810
rect 30156 35756 30324 35758
rect 30268 35746 30324 35756
rect 30604 35810 30660 36428
rect 30828 36418 30884 36428
rect 31612 36418 31668 36428
rect 31052 36260 31108 36270
rect 31052 36166 31108 36204
rect 31276 36258 31332 36270
rect 31276 36206 31278 36258
rect 31330 36206 31332 36258
rect 30604 35758 30606 35810
rect 30658 35758 30660 35810
rect 30604 35746 30660 35758
rect 30716 36148 30772 36158
rect 29708 35298 29764 35308
rect 29820 35698 29876 35710
rect 29820 35646 29822 35698
rect 29874 35646 29876 35698
rect 29036 35086 29038 35138
rect 29090 35086 29092 35138
rect 29036 35074 29092 35086
rect 29820 35028 29876 35646
rect 30044 35700 30100 35710
rect 30044 35698 30212 35700
rect 30044 35646 30046 35698
rect 30098 35646 30212 35698
rect 30044 35644 30212 35646
rect 30044 35634 30100 35644
rect 29932 35028 29988 35038
rect 30156 35028 30212 35644
rect 30604 35588 30660 35598
rect 30492 35476 30548 35486
rect 30492 35308 30548 35420
rect 30268 35196 30548 35308
rect 30380 35028 30436 35038
rect 29820 35026 30100 35028
rect 29820 34974 29934 35026
rect 29986 34974 30100 35026
rect 29820 34972 30100 34974
rect 30156 35026 30436 35028
rect 30156 34974 30382 35026
rect 30434 34974 30436 35026
rect 30156 34972 30436 34974
rect 29932 34962 29988 34972
rect 29484 34914 29540 34926
rect 29484 34862 29486 34914
rect 29538 34862 29540 34914
rect 29484 34692 29540 34862
rect 29484 34626 29540 34636
rect 29708 34914 29764 34926
rect 29708 34862 29710 34914
rect 29762 34862 29764 34914
rect 29596 34132 29652 34142
rect 29708 34132 29764 34862
rect 29932 34244 29988 34254
rect 29932 34150 29988 34188
rect 29596 34130 29764 34132
rect 29596 34078 29598 34130
rect 29650 34078 29764 34130
rect 29596 34076 29764 34078
rect 29596 33684 29652 34076
rect 29036 33628 29652 33684
rect 29036 31892 29092 33628
rect 29148 33458 29204 33470
rect 29148 33406 29150 33458
rect 29202 33406 29204 33458
rect 29148 33124 29204 33406
rect 29148 33068 29988 33124
rect 29484 32900 29540 32910
rect 29484 32676 29540 32844
rect 29820 32788 29876 32798
rect 29820 32694 29876 32732
rect 29484 32674 29652 32676
rect 29484 32622 29486 32674
rect 29538 32622 29652 32674
rect 29484 32620 29652 32622
rect 29484 32610 29540 32620
rect 29148 32450 29204 32462
rect 29148 32398 29150 32450
rect 29202 32398 29204 32450
rect 29148 32340 29204 32398
rect 29148 32274 29204 32284
rect 29260 32452 29316 32462
rect 29148 31892 29204 31902
rect 29036 31836 29148 31892
rect 29148 31826 29204 31836
rect 28924 31612 29204 31668
rect 28700 27806 28702 27858
rect 28754 27806 28756 27858
rect 28700 27794 28756 27806
rect 28812 27858 28868 27870
rect 28812 27806 28814 27858
rect 28866 27806 28868 27858
rect 28812 27748 28868 27806
rect 29036 27858 29092 27870
rect 29036 27806 29038 27858
rect 29090 27806 29092 27858
rect 29036 27748 29092 27806
rect 28812 27692 29092 27748
rect 27580 27186 27636 27198
rect 27580 27134 27582 27186
rect 27634 27134 27636 27186
rect 27580 26516 27636 27134
rect 28476 26740 28532 26750
rect 27580 26450 27636 26460
rect 28140 26516 28196 26526
rect 28476 26516 28532 26684
rect 27692 26292 27748 26302
rect 27580 26236 27692 26292
rect 27244 25396 27300 25406
rect 27244 25302 27300 25340
rect 27468 25396 27524 25406
rect 27468 25302 27524 25340
rect 27356 25284 27412 25294
rect 27356 25190 27412 25228
rect 27132 25116 27300 25172
rect 27020 25060 27076 25070
rect 26684 24110 26686 24162
rect 26738 24110 26740 24162
rect 26684 24098 26740 24110
rect 26908 24722 26964 24734
rect 26908 24670 26910 24722
rect 26962 24670 26964 24722
rect 26460 23940 26516 23950
rect 26460 23846 26516 23884
rect 26908 23268 26964 24670
rect 26908 23202 26964 23212
rect 26572 21812 26628 21822
rect 26572 20916 26628 21756
rect 26908 21700 26964 21710
rect 26908 21606 26964 21644
rect 26684 21476 26740 21486
rect 26684 21382 26740 21420
rect 27020 21140 27076 25004
rect 27132 23714 27188 23726
rect 27132 23662 27134 23714
rect 27186 23662 27188 23714
rect 27132 23548 27188 23662
rect 27244 23548 27300 25116
rect 27580 24948 27636 26236
rect 27692 26226 27748 26236
rect 28140 26290 28196 26460
rect 28140 26238 28142 26290
rect 28194 26238 28196 26290
rect 27804 26178 27860 26190
rect 27804 26126 27806 26178
rect 27858 26126 27860 26178
rect 27356 24892 27580 24948
rect 27356 24722 27412 24892
rect 27580 24882 27636 24892
rect 27692 25394 27748 25406
rect 27692 25342 27694 25394
rect 27746 25342 27748 25394
rect 27356 24670 27358 24722
rect 27410 24670 27412 24722
rect 27356 24658 27412 24670
rect 27580 24724 27636 24734
rect 27692 24724 27748 25342
rect 27804 25396 27860 26126
rect 27804 25060 27860 25340
rect 28028 25506 28084 25518
rect 28028 25454 28030 25506
rect 28082 25454 28084 25506
rect 28028 25394 28084 25454
rect 28140 25508 28196 26238
rect 28252 26514 28532 26516
rect 28252 26462 28478 26514
rect 28530 26462 28532 26514
rect 28252 26460 28532 26462
rect 28252 25730 28308 26460
rect 28476 26450 28532 26460
rect 28812 26514 28868 27692
rect 29148 26908 29204 31612
rect 29260 29092 29316 32396
rect 29596 31892 29652 32620
rect 29708 32562 29764 32574
rect 29708 32510 29710 32562
rect 29762 32510 29764 32562
rect 29708 32340 29764 32510
rect 29708 32274 29764 32284
rect 29932 32562 29988 33068
rect 30044 32900 30100 34972
rect 30380 34962 30436 34972
rect 30492 34916 30548 35196
rect 30604 35028 30660 35532
rect 30716 35140 30772 36092
rect 31276 36036 31332 36206
rect 30828 35980 31332 36036
rect 30828 35922 30884 35980
rect 30828 35870 30830 35922
rect 30882 35870 30884 35922
rect 30828 35858 30884 35870
rect 31164 35812 31220 35822
rect 31052 35756 31164 35812
rect 30828 35698 30884 35710
rect 30828 35646 30830 35698
rect 30882 35646 30884 35698
rect 30828 35364 30884 35646
rect 30828 35298 30884 35308
rect 30716 35084 30996 35140
rect 30604 34972 30884 35028
rect 30492 34860 30660 34916
rect 30268 34692 30324 34702
rect 30268 34598 30324 34636
rect 30492 34690 30548 34702
rect 30492 34638 30494 34690
rect 30546 34638 30548 34690
rect 30492 34244 30548 34638
rect 30044 32844 30212 32900
rect 30044 32676 30100 32686
rect 30044 32582 30100 32620
rect 29932 32510 29934 32562
rect 29986 32510 29988 32562
rect 29708 31892 29764 31902
rect 29596 31890 29764 31892
rect 29596 31838 29710 31890
rect 29762 31838 29764 31890
rect 29596 31836 29764 31838
rect 29708 31826 29764 31836
rect 29484 31780 29540 31790
rect 29484 31686 29540 31724
rect 29820 31556 29876 31566
rect 29820 31462 29876 31500
rect 29932 31220 29988 32510
rect 30156 32004 30212 32844
rect 29932 31154 29988 31164
rect 30044 31948 30212 32004
rect 29708 31106 29764 31118
rect 29708 31054 29710 31106
rect 29762 31054 29764 31106
rect 29484 30996 29540 31006
rect 29484 30902 29540 30940
rect 29708 30324 29764 31054
rect 29820 30996 29876 31006
rect 29820 30902 29876 30940
rect 29708 30258 29764 30268
rect 30044 30212 30100 31948
rect 30380 31892 30436 31902
rect 30156 31780 30212 31790
rect 30156 31686 30212 31724
rect 30268 31556 30324 31566
rect 30268 31108 30324 31500
rect 30156 30324 30212 30334
rect 30156 30230 30212 30268
rect 29820 30210 30100 30212
rect 29820 30158 30046 30210
rect 30098 30158 30100 30210
rect 29820 30156 30100 30158
rect 29484 29428 29540 29438
rect 29484 29314 29540 29372
rect 29484 29262 29486 29314
rect 29538 29262 29540 29314
rect 29484 29250 29540 29262
rect 29820 29092 29876 30156
rect 30044 30146 30100 30156
rect 30268 30098 30324 31052
rect 30268 30046 30270 30098
rect 30322 30046 30324 30098
rect 29260 29036 29540 29092
rect 29260 28084 29316 28094
rect 29260 27990 29316 28028
rect 29036 26852 29204 26908
rect 29372 27972 29428 27982
rect 29372 27858 29428 27916
rect 29372 27806 29374 27858
rect 29426 27806 29428 27858
rect 29372 26908 29428 27806
rect 29484 27636 29540 29036
rect 29596 29036 29876 29092
rect 29932 29428 29988 29438
rect 30268 29428 30324 30046
rect 30380 30882 30436 31836
rect 30380 30830 30382 30882
rect 30434 30830 30436 30882
rect 30380 30098 30436 30830
rect 30492 30660 30548 34188
rect 30492 30594 30548 30604
rect 30380 30046 30382 30098
rect 30434 30046 30436 30098
rect 30380 30034 30436 30046
rect 30380 29428 30436 29438
rect 30268 29426 30436 29428
rect 30268 29374 30382 29426
rect 30434 29374 30436 29426
rect 30268 29372 30436 29374
rect 29596 28644 29652 29036
rect 29596 28530 29652 28588
rect 29932 28642 29988 29372
rect 30380 29362 30436 29372
rect 29932 28590 29934 28642
rect 29986 28590 29988 28642
rect 29932 28578 29988 28590
rect 30380 28644 30436 28654
rect 30604 28644 30660 34860
rect 30716 31220 30772 31230
rect 30716 30994 30772 31164
rect 30716 30942 30718 30994
rect 30770 30942 30772 30994
rect 30716 30930 30772 30942
rect 30828 30436 30884 34972
rect 30940 35026 30996 35084
rect 30940 34974 30942 35026
rect 30994 34974 30996 35026
rect 30940 34914 30996 34974
rect 30940 34862 30942 34914
rect 30994 34862 30996 34914
rect 30940 34850 30996 34862
rect 31052 33572 31108 35756
rect 31164 35718 31220 35756
rect 31612 35812 31668 35822
rect 31612 35718 31668 35756
rect 31276 35700 31332 35710
rect 31164 34914 31220 34926
rect 31164 34862 31166 34914
rect 31218 34862 31220 34914
rect 31164 34354 31220 34862
rect 31164 34302 31166 34354
rect 31218 34302 31220 34354
rect 31164 34290 31220 34302
rect 31052 33506 31108 33516
rect 30380 28642 30660 28644
rect 30380 28590 30382 28642
rect 30434 28590 30660 28642
rect 30380 28588 30660 28590
rect 30380 28578 30436 28588
rect 29596 28478 29598 28530
rect 29650 28478 29652 28530
rect 29596 28466 29652 28478
rect 29708 28084 29764 28094
rect 29708 27970 29764 28028
rect 30268 28084 30324 28094
rect 30268 27990 30324 28028
rect 29708 27918 29710 27970
rect 29762 27918 29764 27970
rect 29708 27906 29764 27918
rect 30492 27636 30548 27646
rect 29484 27580 29764 27636
rect 29372 26852 29652 26908
rect 28812 26462 28814 26514
rect 28866 26462 28868 26514
rect 28812 26450 28868 26462
rect 28924 26740 28980 26750
rect 28924 26290 28980 26684
rect 28924 26238 28926 26290
rect 28978 26238 28980 26290
rect 28924 26226 28980 26238
rect 28252 25678 28254 25730
rect 28306 25678 28308 25730
rect 28252 25666 28308 25678
rect 28476 25620 28532 25630
rect 28196 25452 28420 25508
rect 28140 25414 28196 25452
rect 28028 25342 28030 25394
rect 28082 25342 28084 25394
rect 28028 25330 28084 25342
rect 27804 24994 27860 25004
rect 28028 24948 28084 24958
rect 27804 24724 27860 24734
rect 27580 24722 27860 24724
rect 27580 24670 27582 24722
rect 27634 24670 27806 24722
rect 27858 24670 27860 24722
rect 27580 24668 27860 24670
rect 27580 24658 27636 24668
rect 27804 24658 27860 24668
rect 27356 23940 27412 23950
rect 27356 23846 27412 23884
rect 27580 23940 27636 23950
rect 28028 23940 28084 24892
rect 28364 24612 28420 25452
rect 28476 25172 28532 25564
rect 28588 25396 28644 25406
rect 28588 25394 28756 25396
rect 28588 25342 28590 25394
rect 28642 25342 28756 25394
rect 28588 25340 28756 25342
rect 28588 25330 28644 25340
rect 28476 25116 28644 25172
rect 28588 24722 28644 25116
rect 28588 24670 28590 24722
rect 28642 24670 28644 24722
rect 28588 24658 28644 24670
rect 28476 24612 28532 24622
rect 28364 24610 28532 24612
rect 28364 24558 28478 24610
rect 28530 24558 28532 24610
rect 28364 24556 28532 24558
rect 28476 24546 28532 24556
rect 28700 24612 28756 25340
rect 29036 24948 29092 26852
rect 29148 26292 29204 26302
rect 29484 26292 29540 26302
rect 29148 26198 29204 26236
rect 29372 26290 29540 26292
rect 29372 26238 29486 26290
rect 29538 26238 29540 26290
rect 29372 26236 29540 26238
rect 28700 24546 28756 24556
rect 28812 24892 29092 24948
rect 28812 23940 28868 24892
rect 27132 23492 27300 23548
rect 27580 23492 27636 23884
rect 27692 23938 28084 23940
rect 27692 23886 28030 23938
rect 28082 23886 28084 23938
rect 27692 23884 28084 23886
rect 27692 23826 27748 23884
rect 28028 23874 28084 23884
rect 28252 23884 28868 23940
rect 29148 24834 29204 24846
rect 29148 24782 29150 24834
rect 29202 24782 29204 24834
rect 27692 23774 27694 23826
rect 27746 23774 27748 23826
rect 27692 23762 27748 23774
rect 28140 23714 28196 23726
rect 28140 23662 28142 23714
rect 28194 23662 28196 23714
rect 28140 23492 28196 23662
rect 27020 21074 27076 21084
rect 26684 20916 26740 20926
rect 26460 20914 26964 20916
rect 26460 20862 26686 20914
rect 26738 20862 26964 20914
rect 26460 20860 26964 20862
rect 26460 20018 26516 20860
rect 26684 20850 26740 20860
rect 26908 20692 26964 20860
rect 27020 20692 27076 20702
rect 26908 20690 27076 20692
rect 26908 20638 27022 20690
rect 27074 20638 27076 20690
rect 26908 20636 27076 20638
rect 27020 20626 27076 20636
rect 26684 20580 26740 20590
rect 26684 20130 26740 20524
rect 26684 20078 26686 20130
rect 26738 20078 26740 20130
rect 26684 20066 26740 20078
rect 27132 20578 27188 20590
rect 27132 20526 27134 20578
rect 27186 20526 27188 20578
rect 27132 20132 27188 20526
rect 27132 20066 27188 20076
rect 26460 19966 26462 20018
rect 26514 19966 26516 20018
rect 26460 19954 26516 19966
rect 26348 19458 26964 19460
rect 26348 19406 26350 19458
rect 26402 19406 26964 19458
rect 26348 19404 26964 19406
rect 26348 19394 26404 19404
rect 26908 19346 26964 19404
rect 26908 19294 26910 19346
rect 26962 19294 26964 19346
rect 26908 19282 26964 19294
rect 27244 19236 27300 23492
rect 27468 23436 27636 23492
rect 27692 23436 28196 23492
rect 27244 19180 27412 19236
rect 26124 19030 26180 19068
rect 27132 19124 27188 19134
rect 27188 19068 27300 19124
rect 27132 19058 27188 19068
rect 26796 19012 26852 19022
rect 26572 18788 26628 18798
rect 25788 18510 25790 18562
rect 25842 18510 25844 18562
rect 25788 18498 25844 18510
rect 26460 18732 26572 18788
rect 26348 18450 26404 18462
rect 26348 18398 26350 18450
rect 26402 18398 26404 18450
rect 26348 18228 26404 18398
rect 26348 18162 26404 18172
rect 25004 17826 25060 17836
rect 25452 17836 25620 17892
rect 25228 17666 25284 17678
rect 25228 17614 25230 17666
rect 25282 17614 25284 17666
rect 25228 16884 25284 17614
rect 25228 16818 25284 16828
rect 25340 17556 25396 17566
rect 25116 16322 25172 16334
rect 25116 16270 25118 16322
rect 25170 16270 25172 16322
rect 25116 16210 25172 16270
rect 25116 16158 25118 16210
rect 25170 16158 25172 16210
rect 25116 16146 25172 16158
rect 25228 15316 25284 15326
rect 25004 13972 25060 13982
rect 25004 13300 25060 13916
rect 25004 13186 25060 13244
rect 25004 13134 25006 13186
rect 25058 13134 25060 13186
rect 25004 13122 25060 13134
rect 25116 12852 25172 12862
rect 25116 12758 25172 12796
rect 25228 11396 25284 15260
rect 25340 15148 25396 17500
rect 25452 16436 25508 17836
rect 26460 17780 26516 18732
rect 26572 18722 26628 18732
rect 26796 18674 26852 18956
rect 27244 19010 27300 19068
rect 27244 18958 27246 19010
rect 27298 18958 27300 19010
rect 27244 18946 27300 18958
rect 26796 18622 26798 18674
rect 26850 18622 26852 18674
rect 26796 18610 26852 18622
rect 27132 18788 27188 18798
rect 26572 18450 26628 18462
rect 26572 18398 26574 18450
rect 26626 18398 26628 18450
rect 26572 18228 26628 18398
rect 26684 18452 26740 18462
rect 26684 18358 26740 18396
rect 27020 18450 27076 18462
rect 27020 18398 27022 18450
rect 27074 18398 27076 18450
rect 27020 18340 27076 18398
rect 27020 18274 27076 18284
rect 26572 18172 26852 18228
rect 26796 17780 26852 18172
rect 27020 17780 27076 17790
rect 26460 17724 26628 17780
rect 26796 17778 27076 17780
rect 26796 17726 27022 17778
rect 27074 17726 27076 17778
rect 26796 17724 27076 17726
rect 25452 16370 25508 16380
rect 25564 17666 25620 17678
rect 25564 17614 25566 17666
rect 25618 17614 25620 17666
rect 25564 16882 25620 17614
rect 25676 17668 25732 17678
rect 26124 17668 26180 17678
rect 25676 17666 26516 17668
rect 25676 17614 25678 17666
rect 25730 17614 26126 17666
rect 26178 17614 26516 17666
rect 25676 17612 26516 17614
rect 25676 17602 25732 17612
rect 26124 17602 26180 17612
rect 26012 17444 26068 17454
rect 25900 17388 26012 17444
rect 25788 17108 25844 17118
rect 25788 17014 25844 17052
rect 25564 16830 25566 16882
rect 25618 16830 25620 16882
rect 25564 16772 25620 16830
rect 25564 16100 25620 16716
rect 25676 16884 25732 16894
rect 25676 16210 25732 16828
rect 25788 16324 25844 16334
rect 25900 16324 25956 17388
rect 26012 17378 26068 17388
rect 26460 17332 26516 17612
rect 26572 17666 26628 17724
rect 27020 17714 27076 17724
rect 26572 17614 26574 17666
rect 26626 17614 26628 17666
rect 26572 17602 26628 17614
rect 26908 17556 26964 17566
rect 26460 17276 26740 17332
rect 26684 17106 26740 17276
rect 26684 17054 26686 17106
rect 26738 17054 26740 17106
rect 26684 17042 26740 17054
rect 26796 17108 26852 17118
rect 26908 17108 26964 17500
rect 26796 17106 26964 17108
rect 26796 17054 26798 17106
rect 26850 17054 26964 17106
rect 26796 17052 26964 17054
rect 26796 17042 26852 17052
rect 26908 16884 26964 16894
rect 27132 16884 27188 18732
rect 26908 16882 27188 16884
rect 26908 16830 26910 16882
rect 26962 16830 27188 16882
rect 26908 16828 27188 16830
rect 26908 16818 26964 16828
rect 26796 16772 26852 16782
rect 25788 16322 26292 16324
rect 25788 16270 25790 16322
rect 25842 16270 26292 16322
rect 25788 16268 26292 16270
rect 25788 16258 25844 16268
rect 25676 16158 25678 16210
rect 25730 16158 25732 16210
rect 25676 16146 25732 16158
rect 25564 16034 25620 16044
rect 26124 15986 26180 15998
rect 26124 15934 26126 15986
rect 26178 15934 26180 15986
rect 25900 15316 25956 15326
rect 25340 15092 25620 15148
rect 25340 14868 25396 14878
rect 25340 14642 25396 14812
rect 25340 14590 25342 14642
rect 25394 14590 25396 14642
rect 25340 14578 25396 14590
rect 25564 13972 25620 15092
rect 25900 14642 25956 15260
rect 25900 14590 25902 14642
rect 25954 14590 25956 14642
rect 25900 14578 25956 14590
rect 26012 14420 26068 14430
rect 26012 14326 26068 14364
rect 26012 14196 26068 14206
rect 26012 13972 26068 14140
rect 25564 13878 25620 13916
rect 25900 13970 26068 13972
rect 25900 13918 26014 13970
rect 26066 13918 26068 13970
rect 25900 13916 26068 13918
rect 25340 13748 25396 13758
rect 25340 12962 25396 13692
rect 25340 12910 25342 12962
rect 25394 12910 25396 12962
rect 25340 12178 25396 12910
rect 25340 12126 25342 12178
rect 25394 12126 25396 12178
rect 25340 11788 25396 12126
rect 25788 12178 25844 12190
rect 25788 12126 25790 12178
rect 25842 12126 25844 12178
rect 25340 11732 25620 11788
rect 24892 11340 25060 11396
rect 24892 11170 24948 11182
rect 24892 11118 24894 11170
rect 24946 11118 24948 11170
rect 23772 10556 23940 10612
rect 22092 10500 22148 10510
rect 22092 10406 22148 10444
rect 22540 10498 22596 10510
rect 22540 10446 22542 10498
rect 22594 10446 22596 10498
rect 22204 9828 22260 9838
rect 22540 9828 22596 10446
rect 23548 10500 23604 10510
rect 23548 10498 23828 10500
rect 23548 10446 23550 10498
rect 23602 10446 23828 10498
rect 23548 10444 23828 10446
rect 23548 10434 23604 10444
rect 23436 10388 23492 10398
rect 22988 10386 23492 10388
rect 22988 10334 23438 10386
rect 23490 10334 23492 10386
rect 22988 10332 23492 10334
rect 22988 9938 23044 10332
rect 23436 10322 23492 10332
rect 22988 9886 22990 9938
rect 23042 9886 23044 9938
rect 22988 9874 23044 9886
rect 23660 10164 23716 10174
rect 22204 9826 22596 9828
rect 22204 9774 22206 9826
rect 22258 9774 22596 9826
rect 22204 9772 22596 9774
rect 22652 9828 22708 9838
rect 22204 9604 22260 9772
rect 21924 9548 22260 9604
rect 21868 9510 21924 9548
rect 21084 9314 21140 9324
rect 22428 9268 22484 9278
rect 22652 9268 22708 9772
rect 22428 9266 22708 9268
rect 22428 9214 22430 9266
rect 22482 9214 22654 9266
rect 22706 9214 22708 9266
rect 22428 9212 22708 9214
rect 22428 9202 22484 9212
rect 22652 9202 22708 9212
rect 22988 9268 23044 9278
rect 22988 9174 23044 9212
rect 23436 9268 23492 9278
rect 19292 8194 19348 8204
rect 20076 9042 20804 9044
rect 20076 8990 20190 9042
rect 20242 8990 20750 9042
rect 20802 8990 20804 9042
rect 20076 8988 20804 8990
rect 20076 8260 20132 8988
rect 20188 8978 20244 8988
rect 20748 8978 20804 8988
rect 23436 9042 23492 9212
rect 23660 9266 23716 10108
rect 23660 9214 23662 9266
rect 23714 9214 23716 9266
rect 23660 9202 23716 9214
rect 23772 9266 23828 10444
rect 23772 9214 23774 9266
rect 23826 9214 23828 9266
rect 23772 9202 23828 9214
rect 23884 9828 23940 10556
rect 23884 9266 23940 9772
rect 23884 9214 23886 9266
rect 23938 9214 23940 9266
rect 23884 9202 23940 9214
rect 24668 9604 24724 9614
rect 24892 9604 24948 11118
rect 24724 9548 24948 9604
rect 24668 9266 24724 9548
rect 24668 9214 24670 9266
rect 24722 9214 24724 9266
rect 24668 9202 24724 9214
rect 24108 9156 24164 9166
rect 24108 9062 24164 9100
rect 23436 8990 23438 9042
rect 23490 8990 23492 9042
rect 23436 8978 23492 8990
rect 20076 8194 20132 8204
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 18508 7410 18564 7420
rect 18284 6514 18340 6524
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 18172 4228 18228 4238
rect 18172 4226 18676 4228
rect 18172 4174 18174 4226
rect 18226 4174 18676 4226
rect 18172 4172 18676 4174
rect 18172 4162 18228 4172
rect 17836 3938 17892 3948
rect 18396 4004 18452 4014
rect 18060 3780 18116 3790
rect 17724 3442 17780 3454
rect 17724 3390 17726 3442
rect 17778 3390 17780 3442
rect 17724 3332 17780 3390
rect 18060 3442 18116 3724
rect 18060 3390 18062 3442
rect 18114 3390 18116 3442
rect 18060 3378 18116 3390
rect 18172 3444 18228 3454
rect 17500 3276 17780 3332
rect 17500 800 17556 3276
rect 18172 800 18228 3388
rect 18396 3442 18452 3948
rect 18396 3390 18398 3442
rect 18450 3390 18452 3442
rect 18396 3378 18452 3390
rect 18620 3554 18676 4172
rect 25004 3666 25060 11340
rect 25116 11340 25284 11396
rect 25340 11508 25396 11518
rect 25340 11394 25396 11452
rect 25340 11342 25342 11394
rect 25394 11342 25396 11394
rect 25116 10164 25172 11340
rect 25340 11330 25396 11342
rect 25564 11282 25620 11732
rect 25564 11230 25566 11282
rect 25618 11230 25620 11282
rect 25564 11218 25620 11230
rect 25788 11172 25844 12126
rect 25900 11732 25956 13916
rect 26012 13906 26068 13916
rect 26012 13748 26068 13758
rect 26124 13748 26180 15934
rect 26236 14532 26292 16268
rect 26796 16322 26852 16716
rect 26796 16270 26798 16322
rect 26850 16270 26852 16322
rect 26796 16258 26852 16270
rect 27132 16212 27188 16828
rect 27244 17554 27300 17566
rect 27244 17502 27246 17554
rect 27298 17502 27300 17554
rect 27244 16882 27300 17502
rect 27244 16830 27246 16882
rect 27298 16830 27300 16882
rect 27244 16818 27300 16830
rect 27356 16772 27412 19180
rect 27468 18564 27524 23436
rect 27692 23378 27748 23436
rect 27692 23326 27694 23378
rect 27746 23326 27748 23378
rect 27692 23314 27748 23326
rect 27580 23268 27636 23278
rect 27580 23174 27636 23212
rect 27692 23156 27748 23166
rect 27692 19012 27748 23100
rect 28252 22820 28308 23884
rect 29148 23826 29204 24782
rect 29372 24388 29428 26236
rect 29484 26226 29540 26236
rect 29484 25282 29540 25294
rect 29484 25230 29486 25282
rect 29538 25230 29540 25282
rect 29484 25060 29540 25230
rect 29484 24994 29540 25004
rect 29596 24724 29652 26852
rect 29708 26404 29764 27580
rect 30380 27580 30492 27636
rect 30156 26962 30212 26974
rect 30156 26910 30158 26962
rect 30210 26910 30212 26962
rect 30156 26908 30212 26910
rect 30380 26908 30436 27580
rect 30492 27570 30548 27580
rect 30156 26852 30436 26908
rect 30492 27412 30548 27422
rect 30492 27074 30548 27356
rect 30492 27022 30494 27074
rect 30546 27022 30548 27074
rect 30156 26404 30212 26414
rect 29708 26402 30212 26404
rect 29708 26350 29710 26402
rect 29762 26350 30158 26402
rect 30210 26350 30212 26402
rect 29708 26348 30212 26350
rect 29708 26338 29764 26348
rect 30156 26338 30212 26348
rect 29708 25732 29764 25742
rect 29708 25284 29764 25676
rect 29820 25508 29876 25518
rect 29820 25506 29988 25508
rect 29820 25454 29822 25506
rect 29874 25454 29988 25506
rect 29820 25452 29988 25454
rect 29820 25442 29876 25452
rect 29820 25284 29876 25294
rect 29708 25228 29820 25284
rect 29820 24836 29876 25228
rect 29932 24948 29988 25452
rect 30156 24948 30212 24958
rect 29932 24946 30212 24948
rect 29932 24894 30158 24946
rect 30210 24894 30212 24946
rect 29932 24892 30212 24894
rect 30268 24948 30324 26852
rect 30492 26516 30548 27022
rect 30604 26740 30660 28588
rect 30716 30380 30884 30436
rect 30940 33460 30996 33470
rect 30716 28308 30772 30380
rect 30828 30210 30884 30222
rect 30828 30158 30830 30210
rect 30882 30158 30884 30210
rect 30828 30100 30884 30158
rect 30828 30034 30884 30044
rect 30940 29876 30996 33404
rect 31276 33460 31332 35644
rect 31500 35252 31556 35262
rect 31388 34804 31444 34814
rect 31388 34710 31444 34748
rect 31500 34802 31556 35196
rect 31724 35140 31780 37100
rect 31836 37090 31892 37100
rect 32508 37044 32564 37774
rect 32508 36978 32564 36988
rect 32732 36708 32788 36718
rect 32732 36594 32788 36652
rect 32732 36542 32734 36594
rect 32786 36542 32788 36594
rect 32172 36484 32228 36494
rect 31836 36260 31892 36270
rect 31836 36166 31892 36204
rect 32172 35922 32228 36428
rect 32172 35870 32174 35922
rect 32226 35870 32228 35922
rect 32172 35858 32228 35870
rect 32508 35698 32564 35710
rect 32508 35646 32510 35698
rect 32562 35646 32564 35698
rect 32508 35252 32564 35646
rect 32732 35700 32788 36542
rect 32844 35812 32900 39676
rect 33180 40292 33236 40302
rect 33180 39058 33236 40236
rect 33740 40068 33796 40460
rect 33852 40404 33908 41692
rect 34188 41188 34244 41198
rect 33852 40338 33908 40348
rect 33964 41186 34244 41188
rect 33964 41134 34190 41186
rect 34242 41134 34244 41186
rect 33964 41132 34244 41134
rect 33964 40180 34020 41132
rect 34188 41122 34244 41132
rect 34300 41076 34356 44940
rect 34412 44940 34580 44996
rect 34412 44660 34468 44940
rect 34412 44594 34468 44604
rect 34636 44548 34692 45388
rect 34748 45332 34804 47628
rect 34972 47460 35028 47470
rect 34972 47346 35028 47404
rect 34972 47294 34974 47346
rect 35026 47294 35028 47346
rect 34972 47282 35028 47294
rect 35196 47458 35252 47470
rect 35196 47406 35198 47458
rect 35250 47406 35252 47458
rect 35196 47124 35252 47406
rect 35196 47058 35252 47068
rect 35532 46898 35588 47628
rect 35532 46846 35534 46898
rect 35586 46846 35588 46898
rect 35532 46834 35588 46846
rect 35196 46674 35252 46686
rect 35196 46622 35198 46674
rect 35250 46622 35252 46674
rect 34860 46564 34916 46574
rect 35196 46564 35252 46622
rect 34860 46562 35252 46564
rect 34860 46510 34862 46562
rect 34914 46510 35252 46562
rect 34860 46508 35252 46510
rect 34860 45668 34916 46508
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35644 45892 35700 48188
rect 36092 48580 36148 48590
rect 36092 48130 36148 48524
rect 36540 48468 36596 48748
rect 36652 48692 36708 49756
rect 36988 49700 37044 49710
rect 36988 49606 37044 49644
rect 36764 48692 36820 48702
rect 36652 48636 36764 48692
rect 36764 48626 36820 48636
rect 36540 48466 36820 48468
rect 36540 48414 36542 48466
rect 36594 48414 36820 48466
rect 36540 48412 36820 48414
rect 36540 48402 36596 48412
rect 36092 48078 36094 48130
rect 36146 48078 36148 48130
rect 36092 48066 36148 48078
rect 36428 48132 36484 48142
rect 36428 47682 36484 48076
rect 36428 47630 36430 47682
rect 36482 47630 36484 47682
rect 36428 47618 36484 47630
rect 35756 47572 35812 47582
rect 35756 47234 35812 47516
rect 36092 47460 36148 47470
rect 36092 47366 36148 47404
rect 36428 47460 36484 47470
rect 36764 47460 36820 48412
rect 36876 48356 36932 48366
rect 36876 48242 36932 48300
rect 36876 48190 36878 48242
rect 36930 48190 36932 48242
rect 36876 47684 36932 48190
rect 37100 48242 37156 49868
rect 37212 49138 37268 49980
rect 37548 50708 37604 50718
rect 37212 49086 37214 49138
rect 37266 49086 37268 49138
rect 37212 49074 37268 49086
rect 37436 49810 37492 49822
rect 37436 49758 37438 49810
rect 37490 49758 37492 49810
rect 37436 48804 37492 49758
rect 37548 49812 37604 50652
rect 38332 50708 38388 51214
rect 39564 51268 39620 51278
rect 39564 51174 39620 51212
rect 39004 51156 39060 51166
rect 38332 50642 38388 50652
rect 38892 50820 38948 50830
rect 38220 50484 38276 50494
rect 38220 49922 38276 50428
rect 38220 49870 38222 49922
rect 38274 49870 38276 49922
rect 38220 49858 38276 49870
rect 37548 49138 37604 49756
rect 37548 49086 37550 49138
rect 37602 49086 37604 49138
rect 37548 49074 37604 49086
rect 38332 49588 38388 49598
rect 38108 49028 38164 49038
rect 38108 48934 38164 48972
rect 37436 48738 37492 48748
rect 37996 48692 38052 48702
rect 37660 48356 37716 48366
rect 37100 48190 37102 48242
rect 37154 48190 37156 48242
rect 37100 48178 37156 48190
rect 37436 48242 37492 48254
rect 37436 48190 37438 48242
rect 37490 48190 37492 48242
rect 36988 48132 37044 48142
rect 36988 48038 37044 48076
rect 36876 47618 36932 47628
rect 37436 47684 37492 48190
rect 37660 48242 37716 48300
rect 37660 48190 37662 48242
rect 37714 48190 37716 48242
rect 37660 48178 37716 48190
rect 37996 48242 38052 48636
rect 38332 48580 38388 49532
rect 38444 48804 38500 48814
rect 38444 48692 38500 48748
rect 38444 48636 38836 48692
rect 38332 48524 38500 48580
rect 37996 48190 37998 48242
rect 38050 48190 38052 48242
rect 37996 48178 38052 48190
rect 38332 48242 38388 48254
rect 38332 48190 38334 48242
rect 38386 48190 38388 48242
rect 37436 47618 37492 47628
rect 37884 48130 37940 48142
rect 37884 48078 37886 48130
rect 37938 48078 37940 48130
rect 36988 47460 37044 47470
rect 36484 47404 36596 47460
rect 36764 47458 37044 47460
rect 36764 47406 36990 47458
rect 37042 47406 37044 47458
rect 36764 47404 37044 47406
rect 36428 47394 36484 47404
rect 36316 47348 36372 47358
rect 36316 47254 36372 47292
rect 35756 47182 35758 47234
rect 35810 47182 35812 47234
rect 35756 47124 35812 47182
rect 35756 47058 35812 47068
rect 36092 47236 36148 47246
rect 35868 45892 35924 45902
rect 35644 45836 35868 45892
rect 35532 45780 35588 45790
rect 35588 45724 35812 45780
rect 35532 45714 35588 45724
rect 34860 45602 34916 45612
rect 34748 45266 34804 45276
rect 34748 45106 34804 45118
rect 34748 45054 34750 45106
rect 34802 45054 34804 45106
rect 34748 44996 34804 45054
rect 35084 45108 35140 45118
rect 35084 45014 35140 45052
rect 35756 45106 35812 45724
rect 35868 45668 35924 45836
rect 35868 45666 36036 45668
rect 35868 45614 35870 45666
rect 35922 45614 36036 45666
rect 35868 45612 36036 45614
rect 35868 45602 35924 45612
rect 35756 45054 35758 45106
rect 35810 45054 35812 45106
rect 34748 44930 34804 44940
rect 35756 44772 35812 45054
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35756 44706 35812 44716
rect 35196 44650 35460 44660
rect 34636 44492 35364 44548
rect 34524 44324 34580 44334
rect 34412 44210 34468 44222
rect 34412 44158 34414 44210
rect 34466 44158 34468 44210
rect 34412 43764 34468 44158
rect 34412 43698 34468 43708
rect 34412 43540 34468 43550
rect 34412 42642 34468 43484
rect 34412 42590 34414 42642
rect 34466 42590 34468 42642
rect 34412 42578 34468 42590
rect 34524 43538 34580 44268
rect 35308 44322 35364 44492
rect 35308 44270 35310 44322
rect 35362 44270 35364 44322
rect 34748 44210 34804 44222
rect 34748 44158 34750 44210
rect 34802 44158 34804 44210
rect 34636 44098 34692 44110
rect 34636 44046 34638 44098
rect 34690 44046 34692 44098
rect 34636 43652 34692 44046
rect 34748 44100 34804 44158
rect 34860 44212 34916 44222
rect 35084 44212 35140 44222
rect 34916 44210 35140 44212
rect 34916 44158 35086 44210
rect 35138 44158 35140 44210
rect 34916 44156 35140 44158
rect 34860 44146 34916 44156
rect 35084 44146 35140 44156
rect 34748 44034 34804 44044
rect 35196 44098 35252 44110
rect 35196 44046 35198 44098
rect 35250 44046 35252 44098
rect 34636 43596 34804 43652
rect 34524 43486 34526 43538
rect 34578 43486 34580 43538
rect 34524 42196 34580 43486
rect 34748 42756 34804 43596
rect 35196 43650 35252 44046
rect 35308 43764 35364 44270
rect 35308 43698 35364 43708
rect 35644 44322 35700 44334
rect 35644 44270 35646 44322
rect 35698 44270 35700 44322
rect 35196 43598 35198 43650
rect 35250 43598 35252 43650
rect 35196 43586 35252 43598
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35532 42868 35588 42878
rect 34748 42690 34804 42700
rect 35420 42756 35476 42766
rect 35420 42662 35476 42700
rect 35532 42754 35588 42812
rect 35532 42702 35534 42754
rect 35586 42702 35588 42754
rect 35532 42690 35588 42702
rect 34748 42532 34804 42542
rect 34804 42476 34916 42532
rect 34748 42438 34804 42476
rect 34748 42196 34804 42206
rect 34580 42194 34804 42196
rect 34580 42142 34750 42194
rect 34802 42142 34804 42194
rect 34580 42140 34804 42142
rect 34524 42130 34580 42140
rect 34748 42130 34804 42140
rect 34300 41020 34692 41076
rect 34524 40292 34580 40302
rect 33628 40012 33796 40068
rect 33852 40124 34020 40180
rect 34076 40290 34580 40292
rect 34076 40238 34526 40290
rect 34578 40238 34580 40290
rect 34076 40236 34580 40238
rect 33180 39006 33182 39058
rect 33234 39006 33236 39058
rect 33180 38994 33236 39006
rect 33516 39956 33572 39966
rect 33516 38052 33572 39900
rect 33628 38668 33684 40012
rect 33740 39394 33796 39406
rect 33740 39342 33742 39394
rect 33794 39342 33796 39394
rect 33740 39284 33796 39342
rect 33852 39284 33908 40124
rect 34076 39730 34132 40236
rect 34524 40226 34580 40236
rect 34076 39678 34078 39730
rect 34130 39678 34132 39730
rect 34076 39666 34132 39678
rect 34524 39618 34580 39630
rect 34524 39566 34526 39618
rect 34578 39566 34580 39618
rect 33964 39508 34020 39518
rect 33964 39414 34020 39452
rect 34188 39394 34244 39406
rect 34188 39342 34190 39394
rect 34242 39342 34244 39394
rect 34188 39284 34244 39342
rect 33740 39228 34244 39284
rect 34188 39172 34244 39228
rect 34188 39106 34244 39116
rect 33964 39060 34020 39070
rect 33964 38966 34020 39004
rect 34300 39060 34356 39070
rect 34300 38966 34356 39004
rect 34524 39058 34580 39566
rect 34524 39006 34526 39058
rect 34578 39006 34580 39058
rect 34524 38994 34580 39006
rect 34188 38834 34244 38846
rect 34188 38782 34190 38834
rect 34242 38782 34244 38834
rect 33628 38612 34132 38668
rect 33516 37986 33572 37996
rect 33180 37828 33236 37838
rect 33628 37828 33684 37838
rect 33964 37828 34020 37838
rect 33180 37826 33964 37828
rect 33180 37774 33182 37826
rect 33234 37774 33630 37826
rect 33682 37774 33964 37826
rect 33180 37772 33964 37774
rect 33068 37604 33124 37614
rect 33068 36370 33124 37548
rect 33180 37492 33236 37772
rect 33628 37762 33684 37772
rect 33964 37734 34020 37772
rect 33180 37426 33236 37436
rect 33404 37604 33460 37614
rect 33404 37490 33460 37548
rect 33404 37438 33406 37490
rect 33458 37438 33460 37490
rect 33404 37426 33460 37438
rect 33852 37604 33908 37614
rect 33852 37154 33908 37548
rect 33852 37102 33854 37154
rect 33906 37102 33908 37154
rect 33292 37044 33348 37054
rect 33852 37044 33908 37102
rect 33292 36482 33348 36988
rect 33516 36988 33908 37044
rect 33404 36596 33460 36606
rect 33516 36596 33572 36988
rect 34076 36932 34132 38612
rect 33460 36540 33572 36596
rect 33852 36876 34132 36932
rect 33404 36530 33460 36540
rect 33292 36430 33294 36482
rect 33346 36430 33348 36482
rect 33292 36418 33348 36430
rect 33068 36318 33070 36370
rect 33122 36318 33124 36370
rect 33068 36306 33124 36318
rect 33068 35812 33124 35822
rect 32844 35810 33348 35812
rect 32844 35758 33070 35810
rect 33122 35758 33348 35810
rect 32844 35756 33348 35758
rect 33068 35746 33124 35756
rect 32732 35634 32788 35644
rect 32508 35186 32564 35196
rect 32956 35588 33012 35598
rect 33292 35588 33348 35756
rect 33404 35810 33460 35822
rect 33404 35758 33406 35810
rect 33458 35758 33460 35810
rect 33404 35700 33460 35758
rect 33404 35644 33796 35700
rect 33292 35532 33684 35588
rect 31724 35074 31780 35084
rect 32956 35026 33012 35532
rect 32956 34974 32958 35026
rect 33010 34974 33012 35026
rect 32956 34962 33012 34974
rect 33628 35026 33684 35532
rect 33628 34974 33630 35026
rect 33682 34974 33684 35026
rect 33628 34962 33684 34974
rect 33740 35252 33796 35644
rect 31724 34916 31780 34926
rect 32060 34916 32116 34926
rect 31724 34914 32116 34916
rect 31724 34862 31726 34914
rect 31778 34862 32062 34914
rect 32114 34862 32116 34914
rect 31724 34860 32116 34862
rect 31724 34850 31780 34860
rect 32060 34850 32116 34860
rect 32284 34914 32340 34926
rect 32284 34862 32286 34914
rect 32338 34862 32340 34914
rect 31500 34750 31502 34802
rect 31554 34750 31556 34802
rect 31500 34738 31556 34750
rect 31612 34020 31668 34030
rect 31612 33926 31668 33964
rect 32284 34020 32340 34862
rect 33740 34692 33796 35196
rect 33740 34626 33796 34636
rect 33740 34020 33796 34030
rect 32284 33954 32340 33964
rect 33628 34018 33796 34020
rect 33628 33966 33742 34018
rect 33794 33966 33796 34018
rect 33628 33964 33796 33966
rect 31276 33394 31332 33404
rect 33628 33908 33684 33964
rect 33740 33954 33796 33964
rect 32060 33346 32116 33358
rect 32060 33294 32062 33346
rect 32114 33294 32116 33346
rect 31276 33236 31332 33246
rect 31276 33142 31332 33180
rect 31724 33236 31780 33246
rect 31724 32786 31780 33180
rect 32060 33124 32116 33294
rect 32508 33236 32564 33246
rect 32508 33142 32564 33180
rect 32396 33124 32452 33134
rect 32060 33058 32116 33068
rect 32284 33122 32452 33124
rect 32284 33070 32398 33122
rect 32450 33070 32452 33122
rect 32284 33068 32452 33070
rect 31724 32734 31726 32786
rect 31778 32734 31780 32786
rect 31724 32722 31780 32734
rect 31388 32676 31444 32686
rect 31388 32562 31444 32620
rect 31388 32510 31390 32562
rect 31442 32510 31444 32562
rect 31388 32498 31444 32510
rect 31612 32562 31668 32574
rect 31612 32510 31614 32562
rect 31666 32510 31668 32562
rect 31052 32450 31108 32462
rect 31052 32398 31054 32450
rect 31106 32398 31108 32450
rect 31052 32340 31108 32398
rect 31052 32274 31108 32284
rect 30828 29820 30996 29876
rect 31052 31052 31332 31108
rect 30828 28756 30884 29820
rect 31052 29540 31108 31052
rect 31276 30996 31332 31052
rect 31500 30996 31556 31006
rect 31276 30994 31556 30996
rect 31276 30942 31502 30994
rect 31554 30942 31556 30994
rect 31276 30940 31556 30942
rect 31500 30930 31556 30940
rect 31164 30884 31220 30894
rect 31164 30790 31220 30828
rect 30940 29484 31108 29540
rect 31500 30660 31556 30670
rect 30940 29428 30996 29484
rect 30940 29334 30996 29372
rect 31052 29316 31108 29326
rect 31052 29222 31108 29260
rect 30828 28662 30884 28700
rect 31500 28642 31556 30604
rect 31612 30436 31668 32510
rect 31836 32562 31892 32574
rect 31836 32510 31838 32562
rect 31890 32510 31892 32562
rect 31836 32340 31892 32510
rect 31836 32274 31892 32284
rect 31948 32562 32004 32574
rect 31948 32510 31950 32562
rect 32002 32510 32004 32562
rect 31948 31220 32004 32510
rect 32172 31668 32228 31678
rect 32172 31574 32228 31612
rect 31948 31154 32004 31164
rect 31724 31108 31780 31118
rect 31724 31014 31780 31052
rect 31836 30996 31892 31006
rect 31836 30902 31892 30940
rect 31948 30994 32004 31006
rect 31948 30942 31950 30994
rect 32002 30942 32004 30994
rect 31948 30772 32004 30942
rect 31948 30706 32004 30716
rect 32172 30994 32228 31006
rect 32172 30942 32174 30994
rect 32226 30942 32228 30994
rect 31612 30370 31668 30380
rect 31612 30212 31668 30222
rect 31612 30118 31668 30156
rect 31836 30100 31892 30110
rect 31724 30044 31836 30100
rect 31612 29314 31668 29326
rect 31612 29262 31614 29314
rect 31666 29262 31668 29314
rect 31612 28754 31668 29262
rect 31612 28702 31614 28754
rect 31666 28702 31668 28754
rect 31612 28690 31668 28702
rect 31500 28590 31502 28642
rect 31554 28590 31556 28642
rect 31500 28578 31556 28590
rect 31724 28642 31780 30044
rect 31836 30034 31892 30044
rect 32172 29764 32228 30942
rect 32284 30210 32340 33068
rect 32396 33058 32452 33068
rect 32956 33124 33012 33134
rect 32956 32564 33012 33068
rect 32956 32498 33012 32508
rect 33180 31220 33236 31230
rect 33180 31106 33236 31164
rect 33180 31054 33182 31106
rect 33234 31054 33236 31106
rect 33180 31042 33236 31054
rect 33516 30996 33572 31006
rect 33292 30994 33572 30996
rect 33292 30942 33518 30994
rect 33570 30942 33572 30994
rect 33292 30940 33572 30942
rect 33292 30884 33348 30940
rect 33516 30930 33572 30940
rect 33180 30828 33348 30884
rect 32284 30158 32286 30210
rect 32338 30158 32340 30210
rect 32284 30146 32340 30158
rect 33068 30770 33124 30782
rect 33068 30718 33070 30770
rect 33122 30718 33124 30770
rect 33068 30100 33124 30718
rect 33068 30034 33124 30044
rect 33180 29764 33236 30828
rect 33516 30772 33572 30782
rect 33516 29876 33572 30716
rect 33628 29988 33684 33852
rect 33852 33124 33908 36876
rect 34076 36596 34132 36606
rect 33964 36370 34020 36382
rect 33964 36318 33966 36370
rect 34018 36318 34020 36370
rect 33964 35698 34020 36318
rect 34076 36370 34132 36540
rect 34076 36318 34078 36370
rect 34130 36318 34132 36370
rect 34076 36306 34132 36318
rect 34188 35924 34244 38782
rect 34636 38668 34692 41020
rect 34748 40964 34804 40974
rect 34860 40964 34916 42476
rect 35084 42196 35140 42206
rect 35084 41972 35140 42140
rect 35084 41878 35140 41916
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35644 41412 35700 44270
rect 35868 42642 35924 42654
rect 35868 42590 35870 42642
rect 35922 42590 35924 42642
rect 35756 42530 35812 42542
rect 35756 42478 35758 42530
rect 35810 42478 35812 42530
rect 35756 42084 35812 42478
rect 35868 42308 35924 42590
rect 35868 42242 35924 42252
rect 35868 42084 35924 42094
rect 35756 42082 35924 42084
rect 35756 42030 35870 42082
rect 35922 42030 35924 42082
rect 35756 42028 35924 42030
rect 35868 42018 35924 42028
rect 35644 41356 35812 41412
rect 34748 40962 34916 40964
rect 34748 40910 34750 40962
rect 34802 40910 34916 40962
rect 34748 40908 34916 40910
rect 34748 40898 34804 40908
rect 34860 39396 34916 40908
rect 35644 40964 35700 40974
rect 35644 40870 35700 40908
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35084 39620 35140 39630
rect 34860 39302 34916 39340
rect 34972 39618 35140 39620
rect 34972 39566 35086 39618
rect 35138 39566 35140 39618
rect 34972 39564 35140 39566
rect 34636 38612 34916 38668
rect 34300 37940 34356 37950
rect 34300 37846 34356 37884
rect 34636 37828 34692 37838
rect 34636 37734 34692 37772
rect 34412 37492 34468 37502
rect 34468 37436 34580 37492
rect 34412 37398 34468 37436
rect 34412 37044 34468 37054
rect 34300 36372 34356 36382
rect 34300 36278 34356 36316
rect 33964 35646 33966 35698
rect 34018 35646 34020 35698
rect 33964 34580 34020 35646
rect 34076 35868 34244 35924
rect 34076 35588 34132 35868
rect 34412 35810 34468 36988
rect 34524 36708 34580 37436
rect 34748 37380 34804 37390
rect 34524 36642 34580 36652
rect 34636 37378 34804 37380
rect 34636 37326 34750 37378
rect 34802 37326 34804 37378
rect 34636 37324 34804 37326
rect 34636 36484 34692 37324
rect 34748 37314 34804 37324
rect 34636 36390 34692 36428
rect 34748 36484 34804 36494
rect 34860 36484 34916 38612
rect 34972 38388 35028 39564
rect 35084 39554 35140 39564
rect 35308 39396 35364 39406
rect 35308 38948 35364 39340
rect 35756 39058 35812 41356
rect 35868 40964 35924 40974
rect 35868 39620 35924 40908
rect 35868 39526 35924 39564
rect 35980 39396 36036 45612
rect 36092 40628 36148 47180
rect 36540 46898 36596 47404
rect 36988 47394 37044 47404
rect 37436 47460 37492 47470
rect 36540 46846 36542 46898
rect 36594 46846 36596 46898
rect 36540 46834 36596 46846
rect 36764 47236 36820 47246
rect 36764 46786 36820 47180
rect 36764 46734 36766 46786
rect 36818 46734 36820 46786
rect 36764 46722 36820 46734
rect 36652 46676 36708 46686
rect 36652 46582 36708 46620
rect 37100 46674 37156 46686
rect 37100 46622 37102 46674
rect 37154 46622 37156 46674
rect 36204 46564 36260 46574
rect 36204 46004 36260 46508
rect 37100 46564 37156 46622
rect 37100 46498 37156 46508
rect 36204 45938 36260 45948
rect 37324 46452 37380 46462
rect 36316 45106 36372 45118
rect 36316 45054 36318 45106
rect 36370 45054 36372 45106
rect 36316 43540 36372 45054
rect 37324 45106 37380 46396
rect 37324 45054 37326 45106
rect 37378 45054 37380 45106
rect 37324 45042 37380 45054
rect 36316 43474 36372 43484
rect 37324 43428 37380 43438
rect 37436 43428 37492 47404
rect 37772 47348 37828 47358
rect 37772 47254 37828 47292
rect 37884 47236 37940 48078
rect 37884 47170 37940 47180
rect 37996 47012 38052 47022
rect 37884 46676 37940 46686
rect 37884 46582 37940 46620
rect 37996 46116 38052 46956
rect 38332 46564 38388 48190
rect 38332 46498 38388 46508
rect 37996 46002 38052 46060
rect 37996 45950 37998 46002
rect 38050 45950 38052 46002
rect 37996 45938 38052 45950
rect 38332 45330 38388 45342
rect 38332 45278 38334 45330
rect 38386 45278 38388 45330
rect 38332 45220 38388 45278
rect 37884 45164 38388 45220
rect 37884 45106 37940 45164
rect 37884 45054 37886 45106
rect 37938 45054 37940 45106
rect 37884 45042 37940 45054
rect 37996 44994 38052 45006
rect 37996 44942 37998 44994
rect 38050 44942 38052 44994
rect 37772 43764 37828 43774
rect 37772 43650 37828 43708
rect 37772 43598 37774 43650
rect 37826 43598 37828 43650
rect 37772 43586 37828 43598
rect 37324 43426 37492 43428
rect 37324 43374 37326 43426
rect 37378 43374 37492 43426
rect 37324 43372 37492 43374
rect 37660 43540 37716 43550
rect 37324 43362 37380 43372
rect 36428 41972 36484 41982
rect 36428 41300 36484 41916
rect 37436 41412 37492 41422
rect 36428 41298 36708 41300
rect 36428 41246 36430 41298
rect 36482 41246 36708 41298
rect 36428 41244 36708 41246
rect 36428 41234 36484 41244
rect 36092 40562 36148 40572
rect 36204 40964 36260 40974
rect 35756 39006 35758 39058
rect 35810 39006 35812 39058
rect 35756 38994 35812 39006
rect 35868 39340 36036 39396
rect 36204 39394 36260 40908
rect 36652 40852 36708 41244
rect 37436 41298 37492 41356
rect 37436 41246 37438 41298
rect 37490 41246 37492 41298
rect 37436 41234 37492 41246
rect 36988 40964 37044 40974
rect 36988 40870 37044 40908
rect 37660 40964 37716 43484
rect 37996 42084 38052 44942
rect 38108 44548 38164 44558
rect 38108 44454 38164 44492
rect 38444 44324 38500 48524
rect 38780 48466 38836 48636
rect 38780 48414 38782 48466
rect 38834 48414 38836 48466
rect 38780 48402 38836 48414
rect 38780 47684 38836 47694
rect 38668 46116 38724 46126
rect 38668 45106 38724 46060
rect 38668 45054 38670 45106
rect 38722 45054 38724 45106
rect 38668 45042 38724 45054
rect 38668 44548 38724 44558
rect 37660 40898 37716 40908
rect 37884 42028 38052 42084
rect 38108 44268 38500 44324
rect 38556 44324 38612 44334
rect 36652 40786 36708 40796
rect 37100 40852 37156 40862
rect 37100 40404 37156 40796
rect 36652 40290 36708 40302
rect 36652 40238 36654 40290
rect 36706 40238 36708 40290
rect 36652 40068 36708 40238
rect 36652 40002 36708 40012
rect 36204 39342 36206 39394
rect 36258 39342 36260 39394
rect 35252 38892 35364 38948
rect 35420 38948 35476 38958
rect 35084 38722 35140 38734
rect 35084 38670 35086 38722
rect 35138 38670 35140 38722
rect 35084 38668 35140 38670
rect 35252 38668 35308 38892
rect 35420 38854 35476 38892
rect 35532 38836 35588 38846
rect 35532 38834 35812 38836
rect 35532 38782 35534 38834
rect 35586 38782 35812 38834
rect 35532 38780 35812 38782
rect 35532 38770 35588 38780
rect 35084 38612 35308 38668
rect 35420 38724 35476 38734
rect 35420 38610 35476 38668
rect 35420 38558 35422 38610
rect 35474 38558 35476 38610
rect 35420 38546 35476 38558
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 34972 38332 35140 38388
rect 35196 38378 35460 38388
rect 35644 38388 35700 38398
rect 34972 38164 35028 38174
rect 34972 37938 35028 38108
rect 34972 37886 34974 37938
rect 35026 37886 35028 37938
rect 34972 37874 35028 37886
rect 35084 37940 35140 38332
rect 35644 38050 35700 38332
rect 35644 37998 35646 38050
rect 35698 37998 35700 38050
rect 35644 37986 35700 37998
rect 35084 37492 35140 37884
rect 35308 37826 35364 37838
rect 35308 37774 35310 37826
rect 35362 37774 35364 37826
rect 35196 37492 35252 37502
rect 35084 37436 35196 37492
rect 35196 37426 35252 37436
rect 35308 37380 35364 37774
rect 35756 37380 35812 38780
rect 35308 37314 35364 37324
rect 35644 37324 35812 37380
rect 35308 37154 35364 37166
rect 35308 37102 35310 37154
rect 35362 37102 35364 37154
rect 35308 37044 35364 37102
rect 35308 36978 35364 36988
rect 35644 37044 35700 37324
rect 35644 36978 35700 36988
rect 35756 37154 35812 37166
rect 35756 37102 35758 37154
rect 35810 37102 35812 37154
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35756 36708 35812 37102
rect 35868 36820 35924 39340
rect 35980 38948 36036 38958
rect 35980 38164 36036 38892
rect 35980 38098 36036 38108
rect 36092 38834 36148 38846
rect 36092 38782 36094 38834
rect 36146 38782 36148 38834
rect 35980 37938 36036 37950
rect 35980 37886 35982 37938
rect 36034 37886 36036 37938
rect 35980 37380 36036 37886
rect 36092 37380 36148 38782
rect 36204 38388 36260 39342
rect 36540 39396 36596 39406
rect 36540 38500 36596 39340
rect 36652 38948 36708 38958
rect 36652 38854 36708 38892
rect 36988 38948 37044 38958
rect 36988 38854 37044 38892
rect 36204 38322 36260 38332
rect 36428 38444 36596 38500
rect 36876 38834 36932 38846
rect 36876 38782 36878 38834
rect 36930 38782 36932 38834
rect 36428 37938 36484 38444
rect 36876 38388 36932 38782
rect 37100 38668 37156 40348
rect 37772 40402 37828 40414
rect 37772 40350 37774 40402
rect 37826 40350 37828 40402
rect 37436 40292 37492 40302
rect 37324 40290 37492 40292
rect 37324 40238 37438 40290
rect 37490 40238 37492 40290
rect 37324 40236 37492 40238
rect 37212 39620 37268 39630
rect 37212 39526 37268 39564
rect 37324 38948 37380 40236
rect 37436 40226 37492 40236
rect 37548 39732 37604 39742
rect 37548 39506 37604 39676
rect 37772 39620 37828 40350
rect 37884 40404 37940 42028
rect 37996 41860 38052 41870
rect 38108 41860 38164 44268
rect 38556 44230 38612 44268
rect 38668 43764 38724 44492
rect 38668 43698 38724 43708
rect 38780 44546 38836 47628
rect 38892 47460 38948 50764
rect 39004 48580 39060 51100
rect 39116 50596 39172 50606
rect 39116 50502 39172 50540
rect 39004 48514 39060 48524
rect 38892 47394 38948 47404
rect 39676 47012 39732 52220
rect 40012 52164 40068 53564
rect 40124 53844 40180 53854
rect 40124 52834 40180 53788
rect 40124 52782 40126 52834
rect 40178 52782 40180 52834
rect 40124 52770 40180 52782
rect 40236 53060 40292 53070
rect 40236 52276 40292 53004
rect 40236 52210 40292 52220
rect 39788 52162 40068 52164
rect 39788 52110 40014 52162
rect 40066 52110 40068 52162
rect 39788 52108 40068 52110
rect 39788 51490 39844 52108
rect 40012 52098 40068 52108
rect 39788 51438 39790 51490
rect 39842 51438 39844 51490
rect 39788 51426 39844 51438
rect 40236 51938 40292 51950
rect 40236 51886 40238 51938
rect 40290 51886 40292 51938
rect 40012 51380 40068 51390
rect 40012 51378 40180 51380
rect 40012 51326 40014 51378
rect 40066 51326 40180 51378
rect 40012 51324 40180 51326
rect 40012 51314 40068 51324
rect 39788 50370 39844 50382
rect 39788 50318 39790 50370
rect 39842 50318 39844 50370
rect 39788 49026 39844 50318
rect 40124 49700 40180 51324
rect 40236 50428 40292 51886
rect 40796 51156 40852 55244
rect 40908 55234 40964 55244
rect 41244 54740 41300 54750
rect 41244 54738 41972 54740
rect 41244 54686 41246 54738
rect 41298 54686 41972 54738
rect 41244 54684 41972 54686
rect 41244 54674 41300 54684
rect 41132 54628 41188 54638
rect 40908 54514 40964 54526
rect 40908 54462 40910 54514
rect 40962 54462 40964 54514
rect 40908 54404 40964 54462
rect 40908 54338 40964 54348
rect 41132 54514 41188 54572
rect 41916 54626 41972 54684
rect 42028 54738 42084 55916
rect 42140 55906 42196 55916
rect 42812 55468 42868 56030
rect 42140 55410 42196 55422
rect 42140 55358 42142 55410
rect 42194 55358 42196 55410
rect 42140 55300 42196 55358
rect 42140 55234 42196 55244
rect 42588 55412 42868 55468
rect 43260 56084 43316 56094
rect 46172 56084 46228 56094
rect 46620 56084 46676 56094
rect 42028 54686 42030 54738
rect 42082 54686 42084 54738
rect 42028 54674 42084 54686
rect 42476 54740 42532 54750
rect 41916 54574 41918 54626
rect 41970 54574 41972 54626
rect 41916 54562 41972 54574
rect 41132 54462 41134 54514
rect 41186 54462 41188 54514
rect 41020 53172 41076 53182
rect 41020 53078 41076 53116
rect 41132 52052 41188 54462
rect 41356 54516 41412 54526
rect 41356 54422 41412 54460
rect 41580 54514 41636 54526
rect 41580 54462 41582 54514
rect 41634 54462 41636 54514
rect 41468 53732 41524 53742
rect 41468 53170 41524 53676
rect 41468 53118 41470 53170
rect 41522 53118 41524 53170
rect 41468 53106 41524 53118
rect 41580 53172 41636 54462
rect 42252 54180 42308 54190
rect 41916 53844 41972 53854
rect 41916 53750 41972 53788
rect 42252 53618 42308 54124
rect 42252 53566 42254 53618
rect 42306 53566 42308 53618
rect 42252 53554 42308 53566
rect 41916 53172 41972 53182
rect 41580 53170 42084 53172
rect 41580 53118 41918 53170
rect 41970 53118 42084 53170
rect 41580 53116 42084 53118
rect 41916 53106 41972 53116
rect 42028 53060 42084 53116
rect 42028 52994 42084 53004
rect 41804 52052 41860 52062
rect 41132 52050 41860 52052
rect 41132 51998 41806 52050
rect 41858 51998 41860 52050
rect 41132 51996 41860 51998
rect 40796 51090 40852 51100
rect 40908 51378 40964 51390
rect 40908 51326 40910 51378
rect 40962 51326 40964 51378
rect 40908 50820 40964 51326
rect 41356 51380 41412 51390
rect 40908 50754 40964 50764
rect 41132 51268 41188 51278
rect 41132 50818 41188 51212
rect 41132 50766 41134 50818
rect 41186 50766 41188 50818
rect 41132 50754 41188 50766
rect 40796 50596 40852 50606
rect 40796 50482 40852 50540
rect 40796 50430 40798 50482
rect 40850 50430 40852 50482
rect 40236 50372 40628 50428
rect 40796 50418 40852 50430
rect 41244 50484 41300 50494
rect 41244 50390 41300 50428
rect 41356 50482 41412 51324
rect 41356 50430 41358 50482
rect 41410 50430 41412 50482
rect 40348 49700 40404 49710
rect 40124 49644 40348 49700
rect 40348 49606 40404 49644
rect 39788 48974 39790 49026
rect 39842 48974 39844 49026
rect 39788 48962 39844 48974
rect 39900 49140 39956 49150
rect 39900 48914 39956 49084
rect 39900 48862 39902 48914
rect 39954 48862 39956 48914
rect 39900 48850 39956 48862
rect 40572 48914 40628 50372
rect 40572 48862 40574 48914
rect 40626 48862 40628 48914
rect 40572 48850 40628 48862
rect 41020 49700 41076 49710
rect 40012 48130 40068 48142
rect 40012 48078 40014 48130
rect 40066 48078 40068 48130
rect 39900 47684 39956 47694
rect 39900 47570 39956 47628
rect 39900 47518 39902 47570
rect 39954 47518 39956 47570
rect 39900 47506 39956 47518
rect 40012 47236 40068 48078
rect 40348 48132 40404 48142
rect 40460 48132 40516 48142
rect 40348 48130 40460 48132
rect 40348 48078 40350 48130
rect 40402 48078 40460 48130
rect 40348 48076 40460 48078
rect 40348 48066 40404 48076
rect 40124 48020 40180 48030
rect 40124 47460 40180 47964
rect 40124 47366 40180 47404
rect 40348 47570 40404 47582
rect 40348 47518 40350 47570
rect 40402 47518 40404 47570
rect 40012 47170 40068 47180
rect 39676 46956 40180 47012
rect 39004 46564 39060 46574
rect 38892 44994 38948 45006
rect 38892 44942 38894 44994
rect 38946 44942 38948 44994
rect 38892 44660 38948 44942
rect 38892 44594 38948 44604
rect 38780 44494 38782 44546
rect 38834 44494 38836 44546
rect 38780 43540 38836 44494
rect 39004 44436 39060 46508
rect 40012 46564 40068 46574
rect 40012 46470 40068 46508
rect 40124 45892 40180 46956
rect 40236 46004 40292 46014
rect 40236 45910 40292 45948
rect 40124 45798 40180 45836
rect 39564 45668 39620 45678
rect 39900 45668 39956 45678
rect 39564 45666 39900 45668
rect 39564 45614 39566 45666
rect 39618 45614 39900 45666
rect 39564 45612 39900 45614
rect 39564 45602 39620 45612
rect 39900 45574 39956 45612
rect 40348 45668 40404 47518
rect 40460 47572 40516 48076
rect 40460 47506 40516 47516
rect 40460 47236 40516 47246
rect 40460 46676 40516 47180
rect 40684 47234 40740 47246
rect 40684 47182 40686 47234
rect 40738 47182 40740 47234
rect 40684 46788 40740 47182
rect 40908 46788 40964 46798
rect 40684 46732 40908 46788
rect 40460 46116 40516 46620
rect 40908 46674 40964 46732
rect 40908 46622 40910 46674
rect 40962 46622 40964 46674
rect 40908 46610 40964 46622
rect 40460 46050 40516 46060
rect 41020 46340 41076 49644
rect 41132 48468 41188 48478
rect 41356 48468 41412 50430
rect 41804 50428 41860 51996
rect 42476 51490 42532 54684
rect 42588 54516 42644 55412
rect 42588 53844 42644 54460
rect 42588 53778 42644 53788
rect 42924 54404 42980 54414
rect 42924 54068 42980 54348
rect 42924 53618 42980 54012
rect 42924 53566 42926 53618
rect 42978 53566 42980 53618
rect 42924 53554 42980 53566
rect 43148 53730 43204 53742
rect 43148 53678 43150 53730
rect 43202 53678 43204 53730
rect 42476 51438 42478 51490
rect 42530 51438 42532 51490
rect 42476 51426 42532 51438
rect 42588 53508 42644 53518
rect 42588 51380 42644 53452
rect 43148 53508 43204 53678
rect 43148 53442 43204 53452
rect 41916 50596 41972 50606
rect 41916 50502 41972 50540
rect 42252 50482 42308 50494
rect 42252 50430 42254 50482
rect 42306 50430 42308 50482
rect 41468 50372 41524 50382
rect 41804 50372 42084 50428
rect 41468 49026 41524 50316
rect 41692 49812 41748 49822
rect 41692 49718 41748 49756
rect 41468 48974 41470 49026
rect 41522 48974 41524 49026
rect 41468 48962 41524 48974
rect 42028 48916 42084 50372
rect 42028 48850 42084 48860
rect 42252 50260 42308 50430
rect 42588 50482 42644 51324
rect 42588 50430 42590 50482
rect 42642 50430 42644 50482
rect 42588 50418 42644 50430
rect 43036 50482 43092 50494
rect 43036 50430 43038 50482
rect 43090 50430 43092 50482
rect 43036 50260 43092 50430
rect 42252 50204 43092 50260
rect 41804 48804 41860 48814
rect 41804 48468 41860 48748
rect 41132 48466 41860 48468
rect 41132 48414 41134 48466
rect 41186 48414 41860 48466
rect 41132 48412 41860 48414
rect 41132 48402 41188 48412
rect 41356 48242 41412 48254
rect 41356 48190 41358 48242
rect 41410 48190 41412 48242
rect 41356 48132 41412 48190
rect 41804 48242 41860 48412
rect 42140 48468 42196 48478
rect 42140 48354 42196 48412
rect 42140 48302 42142 48354
rect 42194 48302 42196 48354
rect 42140 48290 42196 48302
rect 41804 48190 41806 48242
rect 41858 48190 41860 48242
rect 41804 48178 41860 48190
rect 41356 48066 41412 48076
rect 42028 48130 42084 48142
rect 42028 48078 42030 48130
rect 42082 48078 42084 48130
rect 42028 47572 42084 48078
rect 42140 47572 42196 47582
rect 42028 47570 42196 47572
rect 42028 47518 42142 47570
rect 42194 47518 42196 47570
rect 42028 47516 42196 47518
rect 42140 47506 42196 47516
rect 41244 47460 41300 47470
rect 41244 46786 41300 47404
rect 41468 47458 41524 47470
rect 41468 47406 41470 47458
rect 41522 47406 41524 47458
rect 41468 47236 41524 47406
rect 41468 47170 41524 47180
rect 42252 47012 42308 50204
rect 42364 49698 42420 49710
rect 42364 49646 42366 49698
rect 42418 49646 42420 49698
rect 42364 49250 42420 49646
rect 43260 49588 43316 56028
rect 45388 56082 46676 56084
rect 45388 56030 46174 56082
rect 46226 56030 46622 56082
rect 46674 56030 46676 56082
rect 45388 56028 46676 56030
rect 43820 55858 43876 55870
rect 43820 55806 43822 55858
rect 43874 55806 43876 55858
rect 43820 55524 43876 55806
rect 45388 55468 45444 56028
rect 46172 56018 46228 56028
rect 46620 56018 46676 56028
rect 49532 56084 49588 56094
rect 49532 55990 49588 56028
rect 50428 56084 50484 56094
rect 50428 55990 50484 56028
rect 47628 55972 47684 55982
rect 47628 55878 47684 55916
rect 43820 55458 43876 55468
rect 45276 55412 45444 55468
rect 45500 55412 45556 55422
rect 49644 55412 49700 55422
rect 43932 55188 43988 55198
rect 43932 55094 43988 55132
rect 43820 55076 43876 55086
rect 43372 55074 43876 55076
rect 43372 55022 43822 55074
rect 43874 55022 43876 55074
rect 43372 55020 43876 55022
rect 43372 54626 43428 55020
rect 43820 55010 43876 55020
rect 44940 55076 44996 55086
rect 44940 55074 45108 55076
rect 44940 55022 44942 55074
rect 44994 55022 45108 55074
rect 44940 55020 45108 55022
rect 44940 55010 44996 55020
rect 43372 54574 43374 54626
rect 43426 54574 43428 54626
rect 43372 54562 43428 54574
rect 45052 54516 45108 55020
rect 43820 54068 43876 54078
rect 43596 53732 43652 53742
rect 43596 53638 43652 53676
rect 43820 53730 43876 54012
rect 44156 53844 44212 53854
rect 44940 53844 44996 53854
rect 44156 53842 44996 53844
rect 44156 53790 44158 53842
rect 44210 53790 44942 53842
rect 44994 53790 44996 53842
rect 44156 53788 44996 53790
rect 44156 53778 44212 53788
rect 44940 53778 44996 53788
rect 43820 53678 43822 53730
rect 43874 53678 43876 53730
rect 43820 53666 43876 53678
rect 45052 53732 45108 54460
rect 44156 53620 44212 53630
rect 44156 53526 44212 53564
rect 44044 53506 44100 53518
rect 44828 53508 44884 53518
rect 44044 53454 44046 53506
rect 44098 53454 44100 53506
rect 43708 53060 43764 53070
rect 43708 52164 43764 53004
rect 44044 53060 44100 53454
rect 44268 53506 44884 53508
rect 44268 53454 44830 53506
rect 44882 53454 44884 53506
rect 44268 53452 44884 53454
rect 44044 52994 44100 53004
rect 44156 53060 44212 53070
rect 44268 53060 44324 53452
rect 44828 53442 44884 53452
rect 44156 53058 44324 53060
rect 44156 53006 44158 53058
rect 44210 53006 44324 53058
rect 44156 53004 44324 53006
rect 44156 52994 44212 53004
rect 43484 52108 43764 52164
rect 44940 52948 44996 52958
rect 45052 52948 45108 53676
rect 44940 52946 45108 52948
rect 44940 52894 44942 52946
rect 44994 52894 45108 52946
rect 44940 52892 45108 52894
rect 44940 52164 44996 52892
rect 45164 52164 45220 52174
rect 44940 52162 45220 52164
rect 44940 52110 45166 52162
rect 45218 52110 45220 52162
rect 44940 52108 45220 52110
rect 43260 49522 43316 49532
rect 43372 50484 43428 50494
rect 43484 50484 43540 52108
rect 44156 51828 44212 51838
rect 44156 51602 44212 51772
rect 44156 51550 44158 51602
rect 44210 51550 44212 51602
rect 44156 51538 44212 51550
rect 43820 51380 43876 51390
rect 45052 51380 45108 51390
rect 43820 51286 43876 51324
rect 44716 51378 45108 51380
rect 44716 51326 45054 51378
rect 45106 51326 45108 51378
rect 44716 51324 45108 51326
rect 43428 50428 43540 50484
rect 42364 49198 42366 49250
rect 42418 49198 42420 49250
rect 42364 49186 42420 49198
rect 42700 49140 42756 49150
rect 43148 49140 43204 49150
rect 42700 49138 43204 49140
rect 42700 49086 42702 49138
rect 42754 49086 43150 49138
rect 43202 49086 43204 49138
rect 42700 49084 43204 49086
rect 42700 49074 42756 49084
rect 43148 49074 43204 49084
rect 43372 49026 43428 50428
rect 44716 50148 44772 51324
rect 45052 51314 45108 51324
rect 44940 50484 44996 50494
rect 44940 50390 44996 50428
rect 45052 50372 45108 50382
rect 45052 50278 45108 50316
rect 44772 50092 44884 50148
rect 44716 50082 44772 50092
rect 44604 50036 44660 50046
rect 43372 48974 43374 49026
rect 43426 48974 43428 49026
rect 43372 48962 43428 48974
rect 44492 49698 44548 49710
rect 44492 49646 44494 49698
rect 44546 49646 44548 49698
rect 42924 48916 42980 48926
rect 42476 48804 42532 48814
rect 42476 48710 42532 48748
rect 42812 48468 42868 48506
rect 42812 48402 42868 48412
rect 42588 48244 42644 48254
rect 42812 48244 42868 48254
rect 42924 48244 42980 48860
rect 43036 48914 43092 48926
rect 43036 48862 43038 48914
rect 43090 48862 43092 48914
rect 43036 48804 43092 48862
rect 43596 48916 43652 48926
rect 43596 48822 43652 48860
rect 44492 48916 44548 49646
rect 43036 48354 43092 48748
rect 43036 48302 43038 48354
rect 43090 48302 43092 48354
rect 43036 48290 43092 48302
rect 43596 48354 43652 48366
rect 43596 48302 43598 48354
rect 43650 48302 43652 48354
rect 42588 48242 42756 48244
rect 42588 48190 42590 48242
rect 42642 48190 42756 48242
rect 42588 48188 42756 48190
rect 42588 48178 42644 48188
rect 42700 48020 42756 48188
rect 42812 48242 42980 48244
rect 42812 48190 42814 48242
rect 42866 48190 42980 48242
rect 42812 48188 42980 48190
rect 42812 48178 42868 48188
rect 43596 48020 43652 48302
rect 43932 48244 43988 48254
rect 43932 48242 44324 48244
rect 43932 48190 43934 48242
rect 43986 48190 44324 48242
rect 43932 48188 44324 48190
rect 43932 48178 43988 48188
rect 42700 47964 43652 48020
rect 42252 46956 42532 47012
rect 41244 46734 41246 46786
rect 41298 46734 41300 46786
rect 41244 46722 41300 46734
rect 42364 46786 42420 46798
rect 42364 46734 42366 46786
rect 42418 46734 42420 46786
rect 41132 46676 41188 46686
rect 41132 46582 41188 46620
rect 41692 46676 41748 46686
rect 42252 46676 42308 46686
rect 41692 46674 42308 46676
rect 41692 46622 41694 46674
rect 41746 46622 42254 46674
rect 42306 46622 42308 46674
rect 41692 46620 42308 46622
rect 41692 46610 41748 46620
rect 42252 46610 42308 46620
rect 41916 46452 41972 46462
rect 41916 46358 41972 46396
rect 42140 46450 42196 46462
rect 42140 46398 42142 46450
rect 42194 46398 42196 46450
rect 40796 46004 40852 46014
rect 40796 45910 40852 45948
rect 41020 45890 41076 46284
rect 42140 46340 42196 46398
rect 42140 46274 42196 46284
rect 42140 46116 42196 46126
rect 42140 46002 42196 46060
rect 42140 45950 42142 46002
rect 42194 45950 42196 46002
rect 42140 45938 42196 45950
rect 41020 45838 41022 45890
rect 41074 45838 41076 45890
rect 41020 45826 41076 45838
rect 41580 45892 41636 45902
rect 40348 45666 41524 45668
rect 40348 45614 40350 45666
rect 40402 45614 41524 45666
rect 40348 45612 41524 45614
rect 40348 45602 40404 45612
rect 39004 44434 39620 44436
rect 39004 44382 39006 44434
rect 39058 44382 39620 44434
rect 39004 44380 39620 44382
rect 39004 44370 39060 44380
rect 39564 44324 39620 44380
rect 39564 44322 39732 44324
rect 39564 44270 39566 44322
rect 39618 44270 39732 44322
rect 39564 44268 39732 44270
rect 39564 44258 39620 44268
rect 39340 44212 39396 44222
rect 39340 44118 39396 44156
rect 39452 44098 39508 44110
rect 39452 44046 39454 44098
rect 39506 44046 39508 44098
rect 39452 43764 39508 44046
rect 39340 43708 39508 43764
rect 39004 43540 39060 43550
rect 38780 43538 39060 43540
rect 38780 43486 39006 43538
rect 39058 43486 39060 43538
rect 38780 43484 39060 43486
rect 39004 43474 39060 43484
rect 37996 41858 38164 41860
rect 37996 41806 37998 41858
rect 38050 41806 38164 41858
rect 37996 41804 38164 41806
rect 38220 43426 38276 43438
rect 38220 43374 38222 43426
rect 38274 43374 38276 43426
rect 38220 41860 38276 43374
rect 39340 43426 39396 43708
rect 39340 43374 39342 43426
rect 39394 43374 39396 43426
rect 39340 43362 39396 43374
rect 39004 43314 39060 43326
rect 39004 43262 39006 43314
rect 39058 43262 39060 43314
rect 39004 42754 39060 43262
rect 39004 42702 39006 42754
rect 39058 42702 39060 42754
rect 39004 42690 39060 42702
rect 39676 42754 39732 44268
rect 39676 42702 39678 42754
rect 39730 42702 39732 42754
rect 39676 42690 39732 42702
rect 40012 44322 40068 44334
rect 40012 44270 40014 44322
rect 40066 44270 40068 44322
rect 38444 42532 38500 42542
rect 38444 42438 38500 42476
rect 38668 42532 38724 42542
rect 38892 42532 38948 42542
rect 38668 42530 38836 42532
rect 38668 42478 38670 42530
rect 38722 42478 38836 42530
rect 38668 42476 38836 42478
rect 38668 42466 38724 42476
rect 38780 42084 38836 42476
rect 38892 42438 38948 42476
rect 40012 42196 40068 44270
rect 41468 44322 41524 45612
rect 41580 45106 41636 45836
rect 42364 45892 42420 46734
rect 42364 45826 42420 45836
rect 41580 45054 41582 45106
rect 41634 45054 41636 45106
rect 41580 45042 41636 45054
rect 41692 45778 41748 45790
rect 41692 45726 41694 45778
rect 41746 45726 41748 45778
rect 41468 44270 41470 44322
rect 41522 44270 41524 44322
rect 41468 44258 41524 44270
rect 40236 44212 40292 44222
rect 40124 43652 40180 43662
rect 40124 43558 40180 43596
rect 40236 43650 40292 44156
rect 41580 44098 41636 44110
rect 41580 44046 41582 44098
rect 41634 44046 41636 44098
rect 40236 43598 40238 43650
rect 40290 43598 40292 43650
rect 40236 43586 40292 43598
rect 41020 43652 41076 43662
rect 41020 43426 41076 43596
rect 41020 43374 41022 43426
rect 41074 43374 41076 43426
rect 40124 43314 40180 43326
rect 40124 43262 40126 43314
rect 40178 43262 40180 43314
rect 40124 42754 40180 43262
rect 40124 42702 40126 42754
rect 40178 42702 40180 42754
rect 40124 42690 40180 42702
rect 40348 42644 40404 42654
rect 40236 42642 40404 42644
rect 40236 42590 40350 42642
rect 40402 42590 40404 42642
rect 40236 42588 40404 42590
rect 40124 42196 40180 42206
rect 40012 42140 40124 42196
rect 38780 42028 39284 42084
rect 39228 41970 39284 42028
rect 39228 41918 39230 41970
rect 39282 41918 39284 41970
rect 39228 41906 39284 41918
rect 39676 42082 39732 42094
rect 39676 42030 39678 42082
rect 39730 42030 39732 42082
rect 38444 41860 38500 41870
rect 37996 41794 38052 41804
rect 38220 41794 38276 41804
rect 38332 41858 38500 41860
rect 38332 41806 38446 41858
rect 38498 41806 38500 41858
rect 38332 41804 38500 41806
rect 38220 41188 38276 41198
rect 38332 41188 38388 41804
rect 38444 41794 38500 41804
rect 38780 41860 38836 41870
rect 38892 41860 38948 41870
rect 38836 41858 38948 41860
rect 38836 41806 38894 41858
rect 38946 41806 38948 41858
rect 38836 41804 38948 41806
rect 38220 41186 38388 41188
rect 38220 41134 38222 41186
rect 38274 41134 38388 41186
rect 38220 41132 38388 41134
rect 38444 41636 38500 41646
rect 38108 40740 38164 40750
rect 38108 40626 38164 40684
rect 38108 40574 38110 40626
rect 38162 40574 38164 40626
rect 38108 40562 38164 40574
rect 38220 40516 38276 41132
rect 38444 41074 38500 41580
rect 38444 41022 38446 41074
rect 38498 41022 38500 41074
rect 38444 41010 38500 41022
rect 38780 41186 38836 41804
rect 38892 41794 38948 41804
rect 39676 41636 39732 42030
rect 39900 41970 39956 41982
rect 39900 41918 39902 41970
rect 39954 41918 39956 41970
rect 39676 41570 39732 41580
rect 39788 41858 39844 41870
rect 39788 41806 39790 41858
rect 39842 41806 39844 41858
rect 39788 41412 39844 41806
rect 39564 41356 39844 41412
rect 39564 41298 39620 41356
rect 39564 41246 39566 41298
rect 39618 41246 39620 41298
rect 39564 41234 39620 41246
rect 38780 41134 38782 41186
rect 38834 41134 38836 41186
rect 38668 40740 38724 40750
rect 38668 40626 38724 40684
rect 38668 40574 38670 40626
rect 38722 40574 38724 40626
rect 38668 40562 38724 40574
rect 38220 40460 38612 40516
rect 37884 40348 38388 40404
rect 37772 39554 37828 39564
rect 37548 39454 37550 39506
rect 37602 39454 37604 39506
rect 37548 39442 37604 39454
rect 37324 38882 37380 38892
rect 37996 39394 38052 39406
rect 37996 39342 37998 39394
rect 38050 39342 38052 39394
rect 37436 38836 37492 38846
rect 37996 38836 38052 39342
rect 37436 38834 38052 38836
rect 37436 38782 37438 38834
rect 37490 38782 38052 38834
rect 37436 38780 38052 38782
rect 37436 38668 37492 38780
rect 38220 38722 38276 38734
rect 38220 38670 38222 38722
rect 38274 38670 38276 38722
rect 38220 38668 38276 38670
rect 36540 38332 36932 38388
rect 36988 38610 37044 38622
rect 37100 38612 37716 38668
rect 36988 38558 36990 38610
rect 37042 38558 37044 38610
rect 36540 38274 36596 38332
rect 36540 38222 36542 38274
rect 36594 38222 36596 38274
rect 36540 38210 36596 38222
rect 36988 38276 37044 38558
rect 37324 38276 37380 38286
rect 36988 38274 37380 38276
rect 36988 38222 37326 38274
rect 37378 38222 37380 38274
rect 36988 38220 37380 38222
rect 37324 38210 37380 38220
rect 36428 37886 36430 37938
rect 36482 37886 36484 37938
rect 36204 37826 36260 37838
rect 36204 37774 36206 37826
rect 36258 37774 36260 37826
rect 36204 37716 36260 37774
rect 36204 37650 36260 37660
rect 36092 37324 36260 37380
rect 35980 37314 36036 37324
rect 36092 37154 36148 37166
rect 36092 37102 36094 37154
rect 36146 37102 36148 37154
rect 36092 37042 36148 37102
rect 36092 36990 36094 37042
rect 36146 36990 36148 37042
rect 36092 36978 36148 36990
rect 35868 36764 36036 36820
rect 35756 36652 35924 36708
rect 35084 36596 35140 36606
rect 35084 36594 35476 36596
rect 35084 36542 35086 36594
rect 35138 36542 35476 36594
rect 35084 36540 35476 36542
rect 35084 36530 35140 36540
rect 34748 36482 34916 36484
rect 34748 36430 34750 36482
rect 34802 36430 34916 36482
rect 34748 36428 34916 36430
rect 34748 36418 34804 36428
rect 34972 36260 35028 36270
rect 34636 36258 35028 36260
rect 34636 36206 34974 36258
rect 35026 36206 35028 36258
rect 34636 36204 35028 36206
rect 34524 35924 34580 35934
rect 34636 35924 34692 36204
rect 34972 36194 35028 36204
rect 35084 36260 35140 36270
rect 35084 36166 35140 36204
rect 34524 35922 34692 35924
rect 34524 35870 34526 35922
rect 34578 35870 34692 35922
rect 34524 35868 34692 35870
rect 34524 35858 34580 35868
rect 34412 35758 34414 35810
rect 34466 35758 34468 35810
rect 34188 35700 34244 35710
rect 34188 35606 34244 35644
rect 34076 35522 34132 35532
rect 34300 34692 34356 34702
rect 34300 34598 34356 34636
rect 33964 34514 34020 34524
rect 34412 34356 34468 35758
rect 35420 35812 35476 36540
rect 35532 36372 35588 36382
rect 35532 36278 35588 36316
rect 35756 36372 35812 36382
rect 35644 36260 35700 36270
rect 35644 36166 35700 36204
rect 35532 35812 35588 35822
rect 35420 35810 35588 35812
rect 35420 35758 35534 35810
rect 35586 35758 35588 35810
rect 35420 35756 35588 35758
rect 35532 35746 35588 35756
rect 34860 35698 34916 35710
rect 34860 35646 34862 35698
rect 34914 35646 34916 35698
rect 34860 35588 34916 35646
rect 35196 35588 35252 35598
rect 34860 35532 35196 35588
rect 35196 35522 35252 35532
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34412 34290 34468 34300
rect 34524 35028 34580 35038
rect 34524 34690 34580 34972
rect 34636 34916 34692 34926
rect 35196 34916 35252 34926
rect 34636 34914 35252 34916
rect 34636 34862 34638 34914
rect 34690 34862 35198 34914
rect 35250 34862 35252 34914
rect 34636 34860 35252 34862
rect 34636 34850 34692 34860
rect 35196 34850 35252 34860
rect 35644 34914 35700 34926
rect 35644 34862 35646 34914
rect 35698 34862 35700 34914
rect 34524 34638 34526 34690
rect 34578 34638 34580 34690
rect 34412 34132 34468 34142
rect 34300 34076 34412 34132
rect 34188 34020 34244 34030
rect 34188 33926 34244 33964
rect 34300 33796 34356 34076
rect 34412 34066 34468 34076
rect 34188 33740 34356 33796
rect 34188 33348 34244 33740
rect 34524 33684 34580 34638
rect 34748 34690 34804 34702
rect 34748 34638 34750 34690
rect 34802 34638 34804 34690
rect 34748 34580 34804 34638
rect 34748 34514 34804 34524
rect 35532 34692 35588 34702
rect 34972 34468 35028 34478
rect 34748 34020 34804 34030
rect 34748 33926 34804 33964
rect 34972 33908 35028 34412
rect 35532 34130 35588 34636
rect 35532 34078 35534 34130
rect 35586 34078 35588 34130
rect 35532 34066 35588 34078
rect 34972 33814 35028 33852
rect 35308 33908 35364 33918
rect 35308 33906 35588 33908
rect 35308 33854 35310 33906
rect 35362 33854 35588 33906
rect 35308 33852 35588 33854
rect 35308 33842 35364 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 34524 33628 35140 33684
rect 35196 33674 35460 33684
rect 34300 33570 34356 33582
rect 34300 33518 34302 33570
rect 34354 33518 34356 33570
rect 34300 33460 34356 33518
rect 34860 33460 34916 33470
rect 34300 33458 34916 33460
rect 34300 33406 34862 33458
rect 34914 33406 34916 33458
rect 34300 33404 34916 33406
rect 34860 33394 34916 33404
rect 34188 33292 34468 33348
rect 34412 33236 34468 33292
rect 34412 33234 35028 33236
rect 34412 33182 34414 33234
rect 34466 33182 35028 33234
rect 34412 33180 35028 33182
rect 34412 33170 34468 33180
rect 33740 32564 33796 32574
rect 33740 30212 33796 32508
rect 33852 32452 33908 33068
rect 34300 33124 34356 33134
rect 34300 33030 34356 33068
rect 34748 32564 34804 32574
rect 34636 32562 34804 32564
rect 34636 32510 34750 32562
rect 34802 32510 34804 32562
rect 34636 32508 34804 32510
rect 33852 32386 33908 32396
rect 33964 32450 34020 32462
rect 33964 32398 33966 32450
rect 34018 32398 34020 32450
rect 33964 31444 34020 32398
rect 34636 32338 34692 32508
rect 34748 32498 34804 32508
rect 34636 32286 34638 32338
rect 34690 32286 34692 32338
rect 33964 31378 34020 31388
rect 34300 31444 34356 31454
rect 34300 31218 34356 31388
rect 34300 31166 34302 31218
rect 34354 31166 34356 31218
rect 34300 31154 34356 31166
rect 34188 30996 34244 31006
rect 34188 30902 34244 30940
rect 33740 30146 33796 30156
rect 33852 30884 33908 30894
rect 33628 29932 33796 29988
rect 33516 29820 33684 29876
rect 32172 29698 32228 29708
rect 32508 29708 33236 29764
rect 31836 29426 31892 29438
rect 31836 29374 31838 29426
rect 31890 29374 31892 29426
rect 31836 29316 31892 29374
rect 32396 29316 32452 29326
rect 31836 28756 31892 29260
rect 31836 28690 31892 28700
rect 31948 29314 32452 29316
rect 31948 29262 32398 29314
rect 32450 29262 32452 29314
rect 31948 29260 32452 29262
rect 31724 28590 31726 28642
rect 31778 28590 31780 28642
rect 31724 28578 31780 28590
rect 30716 28252 31332 28308
rect 31052 27748 31108 27758
rect 30940 27746 31108 27748
rect 30940 27694 31054 27746
rect 31106 27694 31108 27746
rect 30940 27692 31108 27694
rect 30940 26964 30996 27692
rect 31052 27682 31108 27692
rect 31164 27076 31220 27086
rect 31164 26982 31220 27020
rect 30940 26898 30996 26908
rect 30604 26674 30660 26684
rect 30604 26516 30660 26526
rect 31276 26516 31332 28252
rect 31836 28084 31892 28094
rect 31948 28084 32004 29260
rect 32396 29250 32452 29260
rect 32508 28866 32564 29708
rect 33292 29540 33348 29550
rect 33292 29446 33348 29484
rect 33180 29428 33236 29438
rect 33068 29426 33236 29428
rect 33068 29374 33182 29426
rect 33234 29374 33236 29426
rect 33068 29372 33236 29374
rect 32508 28814 32510 28866
rect 32562 28814 32564 28866
rect 32508 28802 32564 28814
rect 32956 29092 33012 29102
rect 32396 28756 32452 28766
rect 32396 28662 32452 28700
rect 32060 28644 32116 28654
rect 32060 28550 32116 28588
rect 31836 28082 32004 28084
rect 31836 28030 31838 28082
rect 31890 28030 32004 28082
rect 31836 28028 32004 28030
rect 31836 28018 31892 28028
rect 31948 27860 32004 27870
rect 31948 27766 32004 27804
rect 32060 27858 32116 27870
rect 32060 27806 32062 27858
rect 32114 27806 32116 27858
rect 32060 27524 32116 27806
rect 32284 27748 32340 27758
rect 32956 27748 33012 29036
rect 33068 28196 33124 29372
rect 33180 29362 33236 29372
rect 33404 29426 33460 29438
rect 33404 29374 33406 29426
rect 33458 29374 33460 29426
rect 33292 29316 33348 29326
rect 33292 29204 33348 29260
rect 33180 29148 33348 29204
rect 33404 29204 33460 29374
rect 33180 28530 33236 29148
rect 33404 29138 33460 29148
rect 33516 29426 33572 29438
rect 33516 29374 33518 29426
rect 33570 29374 33572 29426
rect 33516 28980 33572 29374
rect 33292 28924 33572 28980
rect 33292 28754 33348 28924
rect 33292 28702 33294 28754
rect 33346 28702 33348 28754
rect 33292 28644 33348 28702
rect 33404 28756 33460 28766
rect 33404 28662 33460 28700
rect 33292 28578 33348 28588
rect 33180 28478 33182 28530
rect 33234 28478 33236 28530
rect 33180 28466 33236 28478
rect 33628 28532 33684 29820
rect 33628 28466 33684 28476
rect 33068 28140 33348 28196
rect 33292 27970 33348 28140
rect 33292 27918 33294 27970
rect 33346 27918 33348 27970
rect 33292 27906 33348 27918
rect 32284 27746 32452 27748
rect 32284 27694 32286 27746
rect 32338 27694 32452 27746
rect 32284 27692 32452 27694
rect 32956 27692 33236 27748
rect 32284 27682 32340 27692
rect 32060 27458 32116 27468
rect 32396 27188 32452 27692
rect 32508 27636 32564 27646
rect 32508 27634 33124 27636
rect 32508 27582 32510 27634
rect 32562 27582 33124 27634
rect 32508 27580 33124 27582
rect 32508 27570 32564 27580
rect 33068 27298 33124 27580
rect 33068 27246 33070 27298
rect 33122 27246 33124 27298
rect 33068 27234 33124 27246
rect 33180 27300 33236 27692
rect 32508 27188 32564 27198
rect 32396 27186 32564 27188
rect 32396 27134 32510 27186
rect 32562 27134 32564 27186
rect 32396 27132 32564 27134
rect 32508 27122 32564 27132
rect 32620 27188 32676 27198
rect 31612 27076 31668 27086
rect 31612 26964 31668 27020
rect 32060 27076 32116 27086
rect 31724 26964 31780 26974
rect 31612 26962 31780 26964
rect 31612 26910 31726 26962
rect 31778 26910 31780 26962
rect 31612 26908 31780 26910
rect 31724 26898 31780 26908
rect 31836 26964 31892 27002
rect 32060 26982 32116 27020
rect 32284 27076 32340 27086
rect 31836 26898 31892 26908
rect 32284 26962 32340 27020
rect 32620 27074 32676 27132
rect 32620 27022 32622 27074
rect 32674 27022 32676 27074
rect 32620 27010 32676 27022
rect 32284 26910 32286 26962
rect 32338 26910 32340 26962
rect 32284 26898 32340 26910
rect 32956 26964 33012 27002
rect 32956 26898 33012 26908
rect 33068 26964 33124 26974
rect 33180 26964 33236 27244
rect 33628 27188 33684 27198
rect 33628 27094 33684 27132
rect 33068 26962 33236 26964
rect 33068 26910 33070 26962
rect 33122 26910 33236 26962
rect 33068 26908 33236 26910
rect 33740 26908 33796 29932
rect 33852 29652 33908 30828
rect 34300 30770 34356 30782
rect 34300 30718 34302 30770
rect 34354 30718 34356 30770
rect 34300 30548 34356 30718
rect 33852 29586 33908 29596
rect 33964 30492 34356 30548
rect 34636 30548 34692 32286
rect 34972 31218 35028 33180
rect 35084 32338 35140 33628
rect 35308 33346 35364 33358
rect 35308 33294 35310 33346
rect 35362 33294 35364 33346
rect 35308 33124 35364 33294
rect 35308 33058 35364 33068
rect 35420 32676 35476 32686
rect 35308 32620 35420 32676
rect 35308 32562 35364 32620
rect 35420 32610 35476 32620
rect 35308 32510 35310 32562
rect 35362 32510 35364 32562
rect 35308 32498 35364 32510
rect 35084 32286 35086 32338
rect 35138 32286 35140 32338
rect 35084 32274 35140 32286
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34972 31166 34974 31218
rect 35026 31166 35028 31218
rect 34972 31154 35028 31166
rect 35420 30996 35476 31006
rect 35532 30996 35588 33852
rect 35644 33684 35700 34862
rect 35644 33618 35700 33628
rect 35756 33458 35812 36316
rect 35868 36370 35924 36652
rect 35868 36318 35870 36370
rect 35922 36318 35924 36370
rect 35868 35028 35924 36318
rect 35868 34962 35924 34972
rect 35980 34804 36036 36764
rect 36092 36708 36148 36718
rect 36092 36482 36148 36652
rect 36092 36430 36094 36482
rect 36146 36430 36148 36482
rect 36092 36418 36148 36430
rect 36092 35028 36148 35038
rect 36204 35028 36260 37324
rect 36092 35026 36260 35028
rect 36092 34974 36094 35026
rect 36146 34974 36260 35026
rect 36092 34972 36260 34974
rect 36316 37044 36372 37054
rect 36092 34962 36148 34972
rect 35756 33406 35758 33458
rect 35810 33406 35812 33458
rect 35756 33394 35812 33406
rect 35868 34748 36036 34804
rect 35868 31668 35924 34748
rect 35980 34130 36036 34142
rect 35980 34078 35982 34130
rect 36034 34078 36036 34130
rect 35980 33124 36036 34078
rect 36204 34132 36260 34142
rect 36204 34038 36260 34076
rect 36092 34018 36148 34030
rect 36092 33966 36094 34018
rect 36146 33966 36148 34018
rect 36092 33460 36148 33966
rect 36092 33404 36260 33460
rect 35980 33058 36036 33068
rect 36092 33234 36148 33246
rect 36092 33182 36094 33234
rect 36146 33182 36148 33234
rect 35980 32562 36036 32574
rect 35980 32510 35982 32562
rect 36034 32510 36036 32562
rect 35980 32452 36036 32510
rect 35980 32386 36036 32396
rect 35868 31602 35924 31612
rect 36092 31444 36148 33182
rect 36204 32562 36260 33404
rect 36316 32676 36372 36988
rect 36428 37042 36484 37886
rect 37100 38052 37156 38062
rect 37548 38052 37604 38062
rect 36988 37716 37044 37726
rect 36428 36990 36430 37042
rect 36482 36990 36484 37042
rect 36428 36978 36484 36990
rect 36540 37380 36596 37390
rect 36540 37154 36596 37324
rect 36540 37102 36542 37154
rect 36594 37102 36596 37154
rect 36428 34580 36484 34590
rect 36428 34020 36484 34524
rect 36540 34468 36596 37102
rect 36876 37266 36932 37278
rect 36876 37214 36878 37266
rect 36930 37214 36932 37266
rect 36764 37044 36820 37054
rect 36876 37044 36932 37214
rect 36764 37042 36932 37044
rect 36764 36990 36766 37042
rect 36818 36990 36932 37042
rect 36764 36988 36932 36990
rect 36764 35308 36820 36988
rect 36988 36708 37044 37660
rect 36988 35924 37044 36652
rect 37100 37378 37156 37996
rect 37324 38050 37604 38052
rect 37324 37998 37550 38050
rect 37602 37998 37604 38050
rect 37324 37996 37604 37998
rect 37324 37490 37380 37996
rect 37548 37986 37604 37996
rect 37660 37828 37716 38612
rect 37884 38612 38276 38668
rect 37772 38164 37828 38174
rect 37772 38050 37828 38108
rect 37884 38162 37940 38612
rect 38332 38276 38388 40348
rect 38444 39620 38500 39630
rect 38444 39396 38500 39564
rect 38444 39330 38500 39340
rect 37884 38110 37886 38162
rect 37938 38110 37940 38162
rect 37884 38098 37940 38110
rect 37996 38220 38388 38276
rect 37772 37998 37774 38050
rect 37826 37998 37828 38050
rect 37772 37986 37828 37998
rect 37996 38050 38052 38220
rect 37996 37998 37998 38050
rect 38050 37998 38052 38050
rect 37996 37986 38052 37998
rect 37324 37438 37326 37490
rect 37378 37438 37380 37490
rect 37324 37426 37380 37438
rect 37548 37772 37716 37828
rect 37100 37326 37102 37378
rect 37154 37326 37156 37378
rect 37100 36596 37156 37326
rect 37436 37380 37492 37390
rect 37436 37286 37492 37324
rect 37100 36502 37156 36540
rect 36988 35858 37044 35868
rect 37548 35588 37604 37772
rect 37772 37268 37828 37278
rect 37772 37174 37828 37212
rect 38220 37266 38276 37278
rect 38220 37214 38222 37266
rect 38274 37214 38276 37266
rect 38220 37156 38276 37214
rect 38556 37268 38612 40460
rect 38780 40404 38836 41134
rect 39900 40628 39956 41918
rect 39788 40572 39956 40628
rect 38780 40338 38836 40348
rect 39564 40514 39620 40526
rect 39564 40462 39566 40514
rect 39618 40462 39620 40514
rect 39116 40290 39172 40302
rect 39116 40238 39118 40290
rect 39170 40238 39172 40290
rect 38892 39396 38948 39406
rect 38892 39302 38948 39340
rect 39116 38668 39172 40238
rect 38556 37202 38612 37212
rect 39004 38612 39172 38668
rect 38220 37090 38276 37100
rect 39004 36148 39060 38612
rect 39228 38500 39284 38510
rect 39004 36082 39060 36092
rect 39116 36482 39172 36494
rect 39116 36430 39118 36482
rect 39170 36430 39172 36482
rect 37548 35522 37604 35532
rect 37660 35586 37716 35598
rect 37660 35534 37662 35586
rect 37714 35534 37716 35586
rect 36540 34402 36596 34412
rect 36652 35252 36820 35308
rect 36540 34020 36596 34030
rect 36428 34018 36596 34020
rect 36428 33966 36542 34018
rect 36594 33966 36596 34018
rect 36428 33964 36596 33966
rect 36428 33234 36484 33964
rect 36540 33954 36596 33964
rect 36652 34020 36708 35252
rect 37660 35140 37716 35534
rect 37660 35074 37716 35084
rect 38108 35588 38164 35598
rect 37100 35028 37156 35038
rect 37100 34934 37156 34972
rect 37660 34692 37716 34702
rect 37436 34690 37716 34692
rect 37436 34638 37662 34690
rect 37714 34638 37716 34690
rect 37436 34636 37716 34638
rect 37100 34356 37156 34366
rect 37100 34262 37156 34300
rect 36428 33182 36430 33234
rect 36482 33182 36484 33234
rect 36428 33170 36484 33182
rect 36540 33684 36596 33694
rect 36540 33012 36596 33628
rect 36316 32610 36372 32620
rect 36428 32956 36596 33012
rect 36204 32510 36206 32562
rect 36258 32510 36260 32562
rect 36204 32498 36260 32510
rect 35756 31388 36148 31444
rect 36204 31554 36260 31566
rect 36204 31502 36206 31554
rect 36258 31502 36260 31554
rect 35756 30996 35812 31388
rect 35420 30994 35812 30996
rect 35420 30942 35422 30994
rect 35474 30942 35812 30994
rect 35420 30940 35812 30942
rect 35420 30930 35476 30940
rect 35868 30884 35924 30894
rect 35868 30790 35924 30828
rect 35644 30772 35700 30782
rect 35644 30678 35700 30716
rect 36204 30660 36260 31502
rect 36316 30660 36372 30670
rect 35196 30604 35460 30614
rect 36204 30604 36316 30660
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 33852 29428 33908 29438
rect 33964 29428 34020 30492
rect 34636 30482 34692 30492
rect 34412 30324 34468 30334
rect 34412 30230 34468 30268
rect 35084 30324 35140 30334
rect 34524 30212 34580 30222
rect 34860 30212 34916 30250
rect 34580 30156 34692 30212
rect 34524 30146 34580 30156
rect 34188 30100 34244 30110
rect 34076 30044 34188 30100
rect 34076 29650 34132 30044
rect 34188 30034 34244 30044
rect 34076 29598 34078 29650
rect 34130 29598 34132 29650
rect 34076 29586 34132 29598
rect 34300 29652 34356 29662
rect 34300 29558 34356 29596
rect 34524 29540 34580 29550
rect 33852 29426 34020 29428
rect 33852 29374 33854 29426
rect 33906 29374 34020 29426
rect 33852 29372 34020 29374
rect 34412 29428 34468 29438
rect 33852 29362 33908 29372
rect 33852 29204 33908 29214
rect 33852 28754 33908 29148
rect 33852 28702 33854 28754
rect 33906 28702 33908 28754
rect 33852 28690 33908 28702
rect 34412 28756 34468 29372
rect 34412 28690 34468 28700
rect 34076 28644 34132 28654
rect 33964 27858 34020 27870
rect 33964 27806 33966 27858
rect 34018 27806 34020 27858
rect 33964 27300 34020 27806
rect 33964 27234 34020 27244
rect 33068 26898 33124 26908
rect 31500 26852 31556 26862
rect 31500 26850 31668 26852
rect 31500 26798 31502 26850
rect 31554 26798 31668 26850
rect 31500 26796 31668 26798
rect 31500 26786 31556 26796
rect 30492 26514 30660 26516
rect 30492 26462 30606 26514
rect 30658 26462 30660 26514
rect 30492 26460 30660 26462
rect 30604 26450 30660 26460
rect 31052 26514 31332 26516
rect 31052 26462 31278 26514
rect 31330 26462 31332 26514
rect 31052 26460 31332 26462
rect 30940 26404 30996 26414
rect 30716 26402 30996 26404
rect 30716 26350 30942 26402
rect 30994 26350 30996 26402
rect 30716 26348 30996 26350
rect 30380 26180 30436 26190
rect 30380 25506 30436 26124
rect 30716 25620 30772 26348
rect 30940 26338 30996 26348
rect 31052 25620 31108 26460
rect 31276 26450 31332 26460
rect 31500 26292 31556 26302
rect 31500 26198 31556 26236
rect 30380 25454 30382 25506
rect 30434 25454 30436 25506
rect 30380 25442 30436 25454
rect 30492 25564 30772 25620
rect 30828 25564 31108 25620
rect 30492 25172 30548 25564
rect 30604 25396 30660 25406
rect 30828 25396 30884 25564
rect 30604 25394 30884 25396
rect 30604 25342 30606 25394
rect 30658 25342 30884 25394
rect 30604 25340 30884 25342
rect 30604 25330 30660 25340
rect 31276 25284 31332 25294
rect 31500 25284 31556 25294
rect 31276 25282 31556 25284
rect 31276 25230 31278 25282
rect 31330 25230 31502 25282
rect 31554 25230 31556 25282
rect 31276 25228 31556 25230
rect 31276 25218 31332 25228
rect 30492 25116 30772 25172
rect 30268 24892 30548 24948
rect 30156 24882 30212 24892
rect 29820 24780 30100 24836
rect 29596 24668 29764 24724
rect 29596 24500 29652 24510
rect 29372 24322 29428 24332
rect 29484 24498 29652 24500
rect 29484 24446 29598 24498
rect 29650 24446 29652 24498
rect 29484 24444 29652 24446
rect 29484 23938 29540 24444
rect 29596 24434 29652 24444
rect 29484 23886 29486 23938
rect 29538 23886 29540 23938
rect 29484 23874 29540 23886
rect 29148 23774 29150 23826
rect 29202 23774 29204 23826
rect 28364 23714 28420 23726
rect 28364 23662 28366 23714
rect 28418 23662 28420 23714
rect 28364 23380 28420 23662
rect 28364 23324 28868 23380
rect 28812 23268 28868 23324
rect 29036 23268 29092 23278
rect 28812 23266 28980 23268
rect 28812 23214 28814 23266
rect 28866 23214 28980 23266
rect 28812 23212 28980 23214
rect 28812 23202 28868 23212
rect 28700 23154 28756 23166
rect 28700 23102 28702 23154
rect 28754 23102 28756 23154
rect 28028 22764 28308 22820
rect 28364 23042 28420 23054
rect 28364 22990 28366 23042
rect 28418 22990 28420 23042
rect 27804 22484 27860 22494
rect 28028 22484 28084 22764
rect 28364 22708 28420 22990
rect 28700 23044 28756 23102
rect 28812 23044 28868 23054
rect 28700 22988 28812 23044
rect 28812 22978 28868 22988
rect 28924 22932 28980 23212
rect 29036 23174 29092 23212
rect 29148 23044 29204 23774
rect 29260 23716 29316 23726
rect 29260 23714 29428 23716
rect 29260 23662 29262 23714
rect 29314 23662 29428 23714
rect 29260 23660 29428 23662
rect 29260 23650 29316 23660
rect 29148 22978 29204 22988
rect 29036 22932 29092 22942
rect 28924 22876 29036 22932
rect 29036 22866 29092 22876
rect 28364 22642 28420 22652
rect 29372 22708 29428 23660
rect 29708 23604 29764 24668
rect 29820 24612 29876 24622
rect 29820 24518 29876 24556
rect 29932 24050 29988 24780
rect 30044 24722 30100 24780
rect 30044 24670 30046 24722
rect 30098 24670 30100 24722
rect 30044 24658 30100 24670
rect 30268 24724 30324 24734
rect 30268 24630 30324 24668
rect 30492 24162 30548 24892
rect 30492 24110 30494 24162
rect 30546 24110 30548 24162
rect 30492 24098 30548 24110
rect 29932 23998 29934 24050
rect 29986 23998 29988 24050
rect 29932 23986 29988 23998
rect 30604 24052 30660 24062
rect 30604 23958 30660 23996
rect 29708 23548 30212 23604
rect 29708 23380 29764 23390
rect 29708 23378 29988 23380
rect 29708 23326 29710 23378
rect 29762 23326 29988 23378
rect 29708 23324 29988 23326
rect 29708 23314 29764 23324
rect 29372 22642 29428 22652
rect 29484 23154 29540 23166
rect 29484 23102 29486 23154
rect 29538 23102 29540 23154
rect 27804 22482 28084 22484
rect 27804 22430 27806 22482
rect 27858 22430 28084 22482
rect 27804 22428 28084 22430
rect 27804 22418 27860 22428
rect 28028 22370 28084 22428
rect 28140 22596 28196 22606
rect 28140 22482 28196 22540
rect 28140 22430 28142 22482
rect 28194 22430 28196 22482
rect 28140 22418 28196 22430
rect 28028 22318 28030 22370
rect 28082 22318 28084 22370
rect 28028 22148 28084 22318
rect 28588 22370 28644 22382
rect 29148 22372 29204 22382
rect 28588 22318 28590 22370
rect 28642 22318 28644 22370
rect 28588 22260 28644 22318
rect 28588 22194 28644 22204
rect 28700 22370 29204 22372
rect 28700 22318 29150 22370
rect 29202 22318 29204 22370
rect 28700 22316 29204 22318
rect 28028 22082 28084 22092
rect 28252 22146 28308 22158
rect 28252 22094 28254 22146
rect 28306 22094 28308 22146
rect 28252 21924 28308 22094
rect 28252 21858 28308 21868
rect 28700 21810 28756 22316
rect 29148 22306 29204 22316
rect 28700 21758 28702 21810
rect 28754 21758 28756 21810
rect 28700 21746 28756 21758
rect 29148 22148 29204 22158
rect 29148 21812 29204 22092
rect 28476 21700 28532 21738
rect 28476 21634 28532 21644
rect 28028 21588 28084 21598
rect 28028 21252 28084 21532
rect 28028 21186 28084 21196
rect 28364 21588 28420 21598
rect 27916 20802 27972 20814
rect 27916 20750 27918 20802
rect 27970 20750 27972 20802
rect 27916 20132 27972 20750
rect 28140 20804 28196 20814
rect 28140 20692 28196 20748
rect 28140 20690 28308 20692
rect 28140 20638 28142 20690
rect 28194 20638 28308 20690
rect 28140 20636 28308 20638
rect 28140 20626 28196 20636
rect 28252 20356 28308 20636
rect 28364 20580 28420 21532
rect 28476 21476 28532 21486
rect 28476 20916 28532 21420
rect 28476 20802 28532 20860
rect 28476 20750 28478 20802
rect 28530 20750 28532 20802
rect 28476 20738 28532 20750
rect 29148 20690 29204 21756
rect 29148 20638 29150 20690
rect 29202 20638 29204 20690
rect 29148 20626 29204 20638
rect 29372 22146 29428 22158
rect 29372 22094 29374 22146
rect 29426 22094 29428 22146
rect 28364 20514 28420 20524
rect 28588 20580 28644 20590
rect 28588 20486 28644 20524
rect 28252 20300 28420 20356
rect 27916 20020 27972 20076
rect 28252 20130 28308 20142
rect 28252 20078 28254 20130
rect 28306 20078 28308 20130
rect 28140 20020 28196 20030
rect 27916 20018 28196 20020
rect 27916 19966 28142 20018
rect 28194 19966 28196 20018
rect 27916 19964 28196 19966
rect 28140 19954 28196 19964
rect 28028 19236 28084 19246
rect 28252 19236 28308 20078
rect 28364 19346 28420 20300
rect 29372 20132 29428 22094
rect 29484 21588 29540 23102
rect 29708 23154 29764 23166
rect 29708 23102 29710 23154
rect 29762 23102 29764 23154
rect 29596 23044 29652 23054
rect 29596 22372 29652 22988
rect 29708 22596 29764 23102
rect 29708 22530 29764 22540
rect 29820 22932 29876 22942
rect 29708 22372 29764 22382
rect 29596 22370 29764 22372
rect 29596 22318 29710 22370
rect 29762 22318 29764 22370
rect 29596 22316 29764 22318
rect 29708 22306 29764 22316
rect 29820 22258 29876 22876
rect 29820 22206 29822 22258
rect 29874 22206 29876 22258
rect 29820 22194 29876 22206
rect 29596 22148 29652 22158
rect 29596 21810 29652 22092
rect 29596 21758 29598 21810
rect 29650 21758 29652 21810
rect 29596 21746 29652 21758
rect 29932 21810 29988 23324
rect 30044 23156 30100 23166
rect 30044 23062 30100 23100
rect 29932 21758 29934 21810
rect 29986 21758 29988 21810
rect 29932 21746 29988 21758
rect 30044 22596 30100 22606
rect 29484 21494 29540 21532
rect 29708 21588 29764 21598
rect 30044 21588 30100 22540
rect 29708 21586 30100 21588
rect 29708 21534 29710 21586
rect 29762 21534 30100 21586
rect 29708 21532 30100 21534
rect 29708 21522 29764 21532
rect 30044 20804 30100 20814
rect 30156 20804 30212 23548
rect 30716 23492 30772 25116
rect 30100 20748 30212 20804
rect 30380 23436 30772 23492
rect 31052 24162 31108 24174
rect 31052 24110 31054 24162
rect 31106 24110 31108 24162
rect 31052 24050 31108 24110
rect 31052 23998 31054 24050
rect 31106 23998 31108 24050
rect 30044 20710 30100 20748
rect 29932 20692 29988 20702
rect 29932 20598 29988 20636
rect 29484 20580 29540 20590
rect 29820 20580 29876 20590
rect 29540 20524 29764 20580
rect 29484 20486 29540 20524
rect 29372 20076 29540 20132
rect 28364 19294 28366 19346
rect 28418 19294 28420 19346
rect 28364 19282 28420 19294
rect 29372 19906 29428 19918
rect 29372 19854 29374 19906
rect 29426 19854 29428 19906
rect 28084 19180 28308 19236
rect 28588 19236 28644 19246
rect 28028 19142 28084 19180
rect 27692 18956 28196 19012
rect 27468 18508 27748 18564
rect 27468 18340 27524 18350
rect 27468 18338 27636 18340
rect 27468 18286 27470 18338
rect 27522 18286 27636 18338
rect 27468 18284 27636 18286
rect 27468 18274 27524 18284
rect 27580 17668 27636 18284
rect 27580 17574 27636 17612
rect 27468 17444 27524 17454
rect 27468 17350 27524 17388
rect 27692 16996 27748 18508
rect 28028 18338 28084 18350
rect 28028 18286 28030 18338
rect 28082 18286 28084 18338
rect 28028 18228 28084 18286
rect 28028 18162 28084 18172
rect 27692 16930 27748 16940
rect 27804 17668 27860 17678
rect 27356 16706 27412 16716
rect 27356 16548 27412 16558
rect 27132 16156 27300 16212
rect 26348 16098 26404 16110
rect 26348 16046 26350 16098
rect 26402 16046 26404 16098
rect 26348 14868 26404 16046
rect 26348 14802 26404 14812
rect 26572 16100 26628 16110
rect 26348 14532 26404 14542
rect 26236 14530 26404 14532
rect 26236 14478 26350 14530
rect 26402 14478 26404 14530
rect 26236 14476 26404 14478
rect 26348 14466 26404 14476
rect 26572 14530 26628 16044
rect 27020 16100 27076 16110
rect 27076 16044 27188 16100
rect 27020 16034 27076 16044
rect 26908 15316 26964 15326
rect 26908 15222 26964 15260
rect 26796 15202 26852 15214
rect 26796 15150 26798 15202
rect 26850 15150 26852 15202
rect 26796 14644 26852 15150
rect 26908 14868 26964 14878
rect 26908 14644 26964 14812
rect 26796 14588 26964 14644
rect 26572 14478 26574 14530
rect 26626 14478 26628 14530
rect 26572 14466 26628 14478
rect 26684 14532 26740 14542
rect 26684 14438 26740 14476
rect 26908 14530 26964 14588
rect 26908 14478 26910 14530
rect 26962 14478 26964 14530
rect 26908 14466 26964 14478
rect 26796 14420 26852 14430
rect 26796 14326 26852 14364
rect 27020 13972 27076 13982
rect 26460 13748 26516 13758
rect 26068 13692 26180 13748
rect 26348 13746 26516 13748
rect 26348 13694 26462 13746
rect 26514 13694 26516 13746
rect 26348 13692 26516 13694
rect 26012 13654 26068 13692
rect 26348 13636 26404 13692
rect 26460 13682 26516 13692
rect 26796 13746 26852 13758
rect 26796 13694 26798 13746
rect 26850 13694 26852 13746
rect 26124 13580 26404 13636
rect 26684 13634 26740 13646
rect 26684 13582 26686 13634
rect 26738 13582 26740 13634
rect 26124 13074 26180 13580
rect 26236 13412 26292 13422
rect 26236 13186 26292 13356
rect 26236 13134 26238 13186
rect 26290 13134 26292 13186
rect 26236 13122 26292 13134
rect 26572 13412 26628 13422
rect 26124 13022 26126 13074
rect 26178 13022 26180 13074
rect 26124 13010 26180 13022
rect 26460 13076 26516 13086
rect 26012 12740 26068 12750
rect 26012 12646 26068 12684
rect 26236 12292 26292 12302
rect 26460 12292 26516 13020
rect 26572 12404 26628 13356
rect 26684 12962 26740 13582
rect 26796 13076 26852 13694
rect 26796 13010 26852 13020
rect 26684 12910 26686 12962
rect 26738 12910 26740 12962
rect 26684 12898 26740 12910
rect 26908 12964 26964 12974
rect 26908 12870 26964 12908
rect 27020 12962 27076 13916
rect 27132 13860 27188 16044
rect 27244 15316 27300 16156
rect 27356 16210 27412 16492
rect 27356 16158 27358 16210
rect 27410 16158 27412 16210
rect 27356 16146 27412 16158
rect 27692 15988 27748 15998
rect 27692 15894 27748 15932
rect 27804 15986 27860 17612
rect 28140 17666 28196 18956
rect 28476 18564 28532 18574
rect 28588 18564 28644 19180
rect 29372 19234 29428 19854
rect 29372 19182 29374 19234
rect 29426 19182 29428 19234
rect 29036 19010 29092 19022
rect 29036 18958 29038 19010
rect 29090 18958 29092 19010
rect 29036 18788 29092 18958
rect 29036 18722 29092 18732
rect 28476 18562 28644 18564
rect 28476 18510 28478 18562
rect 28530 18510 28644 18562
rect 28476 18508 28644 18510
rect 28476 18498 28532 18508
rect 29372 18450 29428 19182
rect 29372 18398 29374 18450
rect 29426 18398 29428 18450
rect 29372 18386 29428 18398
rect 29484 19346 29540 20076
rect 29708 20018 29764 20524
rect 30380 20580 30436 23436
rect 30492 23268 30548 23278
rect 30492 23174 30548 23212
rect 30940 23268 30996 23278
rect 30604 23154 30660 23166
rect 30828 23156 30884 23166
rect 30604 23102 30606 23154
rect 30658 23102 30660 23154
rect 30492 22930 30548 22942
rect 30492 22878 30494 22930
rect 30546 22878 30548 22930
rect 30492 22260 30548 22878
rect 30492 21700 30548 22204
rect 30604 22258 30660 23102
rect 30604 22206 30606 22258
rect 30658 22206 30660 22258
rect 30604 21924 30660 22206
rect 30716 23154 30884 23156
rect 30716 23102 30830 23154
rect 30882 23102 30884 23154
rect 30716 23100 30884 23102
rect 30716 22148 30772 23100
rect 30828 23090 30884 23100
rect 30940 22820 30996 23212
rect 31052 23156 31108 23998
rect 31276 24052 31332 24062
rect 31276 23378 31332 23996
rect 31276 23326 31278 23378
rect 31330 23326 31332 23378
rect 31276 23314 31332 23326
rect 31388 23268 31444 25228
rect 31500 25218 31556 25228
rect 31388 23202 31444 23212
rect 31052 23090 31108 23100
rect 31500 23156 31556 23166
rect 31500 23062 31556 23100
rect 30828 22764 30996 22820
rect 31388 23042 31444 23054
rect 31388 22990 31390 23042
rect 31442 22990 31444 23042
rect 30828 22258 30884 22764
rect 31388 22708 31444 22990
rect 31612 22820 31668 26796
rect 31724 26740 31780 26750
rect 31724 23044 31780 26684
rect 33180 26514 33236 26908
rect 33180 26462 33182 26514
rect 33234 26462 33236 26514
rect 33180 26450 33236 26462
rect 33628 26852 33796 26908
rect 33964 27074 34020 27086
rect 33964 27022 33966 27074
rect 34018 27022 34020 27074
rect 33964 26964 34020 27022
rect 33964 26898 34020 26908
rect 32060 25506 32116 25518
rect 32060 25454 32062 25506
rect 32114 25454 32116 25506
rect 31948 23714 32004 23726
rect 31948 23662 31950 23714
rect 32002 23662 32004 23714
rect 31948 23156 32004 23662
rect 32060 23492 32116 25454
rect 33068 24724 33124 24734
rect 33068 24630 33124 24668
rect 33180 24722 33236 24734
rect 33180 24670 33182 24722
rect 33234 24670 33236 24722
rect 32284 24276 32340 24286
rect 33180 24276 33236 24670
rect 32340 24220 32676 24276
rect 32284 24210 32340 24220
rect 32620 23828 32676 24220
rect 32732 24220 33236 24276
rect 33516 24724 33572 24734
rect 32732 24162 32788 24220
rect 32732 24110 32734 24162
rect 32786 24110 32788 24162
rect 32732 24098 32788 24110
rect 32732 23828 32788 23838
rect 32060 23426 32116 23436
rect 32508 23826 32788 23828
rect 32508 23774 32734 23826
rect 32786 23774 32788 23826
rect 32508 23772 32788 23774
rect 32508 23378 32564 23772
rect 32732 23762 32788 23772
rect 32844 23826 32900 23838
rect 33180 23828 33236 23838
rect 32844 23774 32846 23826
rect 32898 23774 32900 23826
rect 32844 23716 32900 23774
rect 32844 23650 32900 23660
rect 32956 23826 33236 23828
rect 32956 23774 33182 23826
rect 33234 23774 33236 23826
rect 32956 23772 33236 23774
rect 32508 23326 32510 23378
rect 32562 23326 32564 23378
rect 32508 23268 32564 23326
rect 32508 23202 32564 23212
rect 32284 23156 32340 23166
rect 31948 23154 32340 23156
rect 31948 23102 32286 23154
rect 32338 23102 32340 23154
rect 31948 23100 32340 23102
rect 31724 22978 31780 22988
rect 32060 22932 32116 22942
rect 31948 22876 32060 22932
rect 31612 22764 31892 22820
rect 31388 22652 31780 22708
rect 30940 22482 30996 22494
rect 30940 22430 30942 22482
rect 30994 22430 30996 22482
rect 30940 22372 30996 22430
rect 31612 22482 31668 22494
rect 31612 22430 31614 22482
rect 31666 22430 31668 22482
rect 31388 22372 31444 22382
rect 30940 22306 30996 22316
rect 31052 22370 31444 22372
rect 31052 22318 31390 22370
rect 31442 22318 31444 22370
rect 31052 22316 31444 22318
rect 30828 22206 30830 22258
rect 30882 22206 30884 22258
rect 30828 22194 30884 22206
rect 31052 22148 31108 22316
rect 31388 22306 31444 22316
rect 31500 22372 31556 22382
rect 31612 22372 31668 22430
rect 31556 22316 31668 22372
rect 31500 22306 31556 22316
rect 30716 22082 30772 22092
rect 30940 22092 31108 22148
rect 30604 21868 30884 21924
rect 30604 21700 30660 21710
rect 30492 21698 30660 21700
rect 30492 21646 30606 21698
rect 30658 21646 30660 21698
rect 30492 21644 30660 21646
rect 30604 21634 30660 21644
rect 30716 21698 30772 21710
rect 30716 21646 30718 21698
rect 30770 21646 30772 21698
rect 30492 21364 30548 21374
rect 30492 20802 30548 21308
rect 30716 21252 30772 21646
rect 30828 21700 30884 21868
rect 30940 21810 30996 22092
rect 30940 21758 30942 21810
rect 30994 21758 30996 21810
rect 30940 21746 30996 21758
rect 31052 21924 31108 21934
rect 30828 21634 30884 21644
rect 31052 21588 31108 21868
rect 31500 21812 31556 21822
rect 31500 21718 31556 21756
rect 31724 21812 31780 22652
rect 31836 22372 31892 22764
rect 31948 22372 32004 22876
rect 32060 22866 32116 22876
rect 32060 22372 32116 22382
rect 31948 22370 32116 22372
rect 31948 22318 32062 22370
rect 32114 22318 32116 22370
rect 31948 22316 32116 22318
rect 31836 22306 31892 22316
rect 32060 22306 32116 22316
rect 32284 22260 32340 23100
rect 32956 22932 33012 23772
rect 33180 23762 33236 23772
rect 33516 23604 33572 24668
rect 33292 23548 33572 23604
rect 33180 23492 33236 23502
rect 33068 23156 33124 23166
rect 33068 23062 33124 23100
rect 32956 22866 33012 22876
rect 33180 22596 33236 23436
rect 32620 22540 33236 22596
rect 32620 22482 32676 22540
rect 32620 22430 32622 22482
rect 32674 22430 32676 22482
rect 32284 22194 32340 22204
rect 32396 22372 32452 22382
rect 31836 22148 31892 22158
rect 31836 22054 31892 22092
rect 31948 22146 32004 22158
rect 31948 22094 31950 22146
rect 32002 22094 32004 22146
rect 31724 21746 31780 21756
rect 31276 21588 31332 21598
rect 30716 21186 30772 21196
rect 30940 21532 31108 21588
rect 31164 21586 31332 21588
rect 31164 21534 31278 21586
rect 31330 21534 31332 21586
rect 31164 21532 31332 21534
rect 30492 20750 30494 20802
rect 30546 20750 30548 20802
rect 30492 20738 30548 20750
rect 30380 20524 30772 20580
rect 29820 20486 29876 20524
rect 29708 19966 29710 20018
rect 29762 19966 29764 20018
rect 29708 19954 29764 19966
rect 30380 20356 30436 20366
rect 29484 19294 29486 19346
rect 29538 19294 29540 19346
rect 28252 18226 28308 18238
rect 28252 18174 28254 18226
rect 28306 18174 28308 18226
rect 28252 18004 28308 18174
rect 28924 18228 28980 18238
rect 29484 18228 29540 19294
rect 29708 19236 29764 19246
rect 29708 19142 29764 19180
rect 30156 18564 30212 18574
rect 29708 18508 29988 18564
rect 29708 18452 29764 18508
rect 28924 18226 29540 18228
rect 28924 18174 28926 18226
rect 28978 18174 29540 18226
rect 28924 18172 29540 18174
rect 29596 18396 29764 18452
rect 29932 18450 29988 18508
rect 29932 18398 29934 18450
rect 29986 18398 29988 18450
rect 28924 18162 28980 18172
rect 28252 17938 28308 17948
rect 29372 18004 29428 18014
rect 28140 17614 28142 17666
rect 28194 17614 28196 17666
rect 28140 17108 28196 17614
rect 28364 17668 28420 17678
rect 28364 17574 28420 17612
rect 29372 17666 29428 17948
rect 29372 17614 29374 17666
rect 29426 17614 29428 17666
rect 29372 17602 29428 17614
rect 28588 17556 28644 17566
rect 28476 17444 28532 17454
rect 28476 17350 28532 17388
rect 28588 17332 28644 17500
rect 29148 17556 29204 17566
rect 29148 17462 29204 17500
rect 28588 17266 28644 17276
rect 29260 17442 29316 17454
rect 29260 17390 29262 17442
rect 29314 17390 29316 17442
rect 28252 17108 28308 17118
rect 28140 17106 28308 17108
rect 28140 17054 28254 17106
rect 28306 17054 28308 17106
rect 28140 17052 28308 17054
rect 28252 17042 28308 17052
rect 28476 16996 28532 17006
rect 28364 16772 28420 16782
rect 28364 16210 28420 16716
rect 28364 16158 28366 16210
rect 28418 16158 28420 16210
rect 28364 16146 28420 16158
rect 27804 15934 27806 15986
rect 27858 15934 27860 15986
rect 27804 15764 27860 15934
rect 27580 15708 27860 15764
rect 28028 15874 28084 15886
rect 28028 15822 28030 15874
rect 28082 15822 28084 15874
rect 27580 15426 27636 15708
rect 27580 15374 27582 15426
rect 27634 15374 27636 15426
rect 27580 15362 27636 15374
rect 28028 15428 28084 15822
rect 27244 15260 27524 15316
rect 27468 15204 27524 15260
rect 27916 15314 27972 15326
rect 27916 15262 27918 15314
rect 27970 15262 27972 15314
rect 27468 15148 27860 15204
rect 27132 13766 27188 13804
rect 27244 15092 27300 15102
rect 27020 12910 27022 12962
rect 27074 12910 27076 12962
rect 27020 12898 27076 12910
rect 27244 12962 27300 15036
rect 27692 14756 27748 14766
rect 27244 12910 27246 12962
rect 27298 12910 27300 12962
rect 27244 12898 27300 12910
rect 27356 14754 27748 14756
rect 27356 14702 27694 14754
rect 27746 14702 27748 14754
rect 27356 14700 27748 14702
rect 26796 12738 26852 12750
rect 26796 12686 26798 12738
rect 26850 12686 26852 12738
rect 26684 12404 26740 12414
rect 26572 12402 26740 12404
rect 26572 12350 26686 12402
rect 26738 12350 26740 12402
rect 26572 12348 26740 12350
rect 26684 12338 26740 12348
rect 26796 12402 26852 12686
rect 26796 12350 26798 12402
rect 26850 12350 26852 12402
rect 26236 12290 26516 12292
rect 26236 12238 26238 12290
rect 26290 12238 26516 12290
rect 26236 12236 26516 12238
rect 26236 12226 26292 12236
rect 26796 11956 26852 12350
rect 26908 12740 26964 12750
rect 26908 12402 26964 12684
rect 27356 12740 27412 14700
rect 27692 14690 27748 14700
rect 27580 14532 27636 14542
rect 27468 14420 27524 14430
rect 27468 13746 27524 14364
rect 27468 13694 27470 13746
rect 27522 13694 27524 13746
rect 27468 13682 27524 13694
rect 27580 13186 27636 14476
rect 27804 14418 27860 15148
rect 27916 14868 27972 15262
rect 27916 14802 27972 14812
rect 28028 14754 28084 15372
rect 28476 15314 28532 16940
rect 28924 16884 28980 16894
rect 29260 16884 29316 17390
rect 29484 17220 29540 17230
rect 28924 16882 29316 16884
rect 28924 16830 28926 16882
rect 28978 16830 29316 16882
rect 28924 16828 29316 16830
rect 29372 17164 29484 17220
rect 29372 16882 29428 17164
rect 29484 17154 29540 17164
rect 29484 16996 29540 17006
rect 29484 16902 29540 16940
rect 29372 16830 29374 16882
rect 29426 16830 29428 16882
rect 28924 16818 28980 16828
rect 29372 16818 29428 16830
rect 28588 16660 28644 16670
rect 28588 16566 28644 16604
rect 28812 15428 28868 15438
rect 28812 15334 28868 15372
rect 29036 15426 29092 15438
rect 29036 15374 29038 15426
rect 29090 15374 29092 15426
rect 28476 15262 28478 15314
rect 28530 15262 28532 15314
rect 28476 15148 28532 15262
rect 28476 15092 28980 15148
rect 28028 14702 28030 14754
rect 28082 14702 28084 14754
rect 28028 14690 28084 14702
rect 27804 14366 27806 14418
rect 27858 14366 27860 14418
rect 27804 14354 27860 14366
rect 28924 13970 28980 15092
rect 28924 13918 28926 13970
rect 28978 13918 28980 13970
rect 27580 13134 27582 13186
rect 27634 13134 27636 13186
rect 27580 13076 27636 13134
rect 27692 13860 27748 13870
rect 28364 13860 28420 13870
rect 27692 13858 28420 13860
rect 27692 13806 27694 13858
rect 27746 13806 28366 13858
rect 28418 13806 28420 13858
rect 27692 13804 28420 13806
rect 27692 13188 27748 13804
rect 28364 13794 28420 13804
rect 28252 13634 28308 13646
rect 28252 13582 28254 13634
rect 28306 13582 28308 13634
rect 27804 13524 27860 13534
rect 27804 13430 27860 13468
rect 28140 13522 28196 13534
rect 28140 13470 28142 13522
rect 28194 13470 28196 13522
rect 28140 13412 28196 13470
rect 27916 13356 28196 13412
rect 28252 13412 28308 13582
rect 28924 13524 28980 13918
rect 28924 13458 28980 13468
rect 27804 13188 27860 13198
rect 27692 13186 27860 13188
rect 27692 13134 27806 13186
rect 27858 13134 27860 13186
rect 27692 13132 27860 13134
rect 27804 13122 27860 13132
rect 27580 13020 27748 13076
rect 27692 12964 27748 13020
rect 27916 12964 27972 13356
rect 28252 13346 28308 13356
rect 29036 13300 29092 15374
rect 29148 15204 29204 15214
rect 29596 15204 29652 18396
rect 29932 18386 29988 18398
rect 29820 18340 29876 18350
rect 29148 15202 29652 15204
rect 29148 15150 29150 15202
rect 29202 15150 29652 15202
rect 29148 15148 29652 15150
rect 29708 18338 29876 18340
rect 29708 18286 29822 18338
rect 29874 18286 29876 18338
rect 29708 18284 29876 18286
rect 29148 15138 29204 15148
rect 29708 14420 29764 18284
rect 29820 18274 29876 18284
rect 30156 18004 30212 18508
rect 30156 17938 30212 17948
rect 29820 17668 29876 17678
rect 30156 17668 30212 17678
rect 29820 17666 30212 17668
rect 29820 17614 29822 17666
rect 29874 17614 30158 17666
rect 30210 17614 30212 17666
rect 29820 17612 30212 17614
rect 29820 17602 29876 17612
rect 30156 17602 30212 17612
rect 30268 17668 30324 17678
rect 30268 17574 30324 17612
rect 30044 17442 30100 17454
rect 30380 17444 30436 20300
rect 30044 17390 30046 17442
rect 30098 17390 30100 17442
rect 30044 17332 30100 17390
rect 30044 17266 30100 17276
rect 30156 17388 30436 17444
rect 30492 17444 30548 17454
rect 29708 14354 29764 14364
rect 29372 13860 29428 13870
rect 29372 13766 29428 13804
rect 28924 13244 29092 13300
rect 29932 13636 29988 13646
rect 27692 12908 27972 12964
rect 28140 12962 28196 12974
rect 28140 12910 28142 12962
rect 28194 12910 28196 12962
rect 27356 12674 27412 12684
rect 26908 12350 26910 12402
rect 26962 12350 26964 12402
rect 26908 12338 26964 12350
rect 28140 12404 28196 12910
rect 28364 12964 28420 12974
rect 28364 12870 28420 12908
rect 28140 12338 28196 12348
rect 28252 12738 28308 12750
rect 28252 12686 28254 12738
rect 28306 12686 28308 12738
rect 28252 12292 28308 12686
rect 28476 12740 28532 12750
rect 28476 12738 28868 12740
rect 28476 12686 28478 12738
rect 28530 12686 28868 12738
rect 28476 12684 28868 12686
rect 28476 12674 28532 12684
rect 28252 12226 28308 12236
rect 28812 12290 28868 12684
rect 28924 12404 28980 13244
rect 29932 13074 29988 13580
rect 29932 13022 29934 13074
rect 29986 13022 29988 13074
rect 29932 13010 29988 13022
rect 29148 12964 29204 12974
rect 29148 12870 29204 12908
rect 29372 12962 29428 12974
rect 29372 12910 29374 12962
rect 29426 12910 29428 12962
rect 29372 12516 29428 12910
rect 28924 12338 28980 12348
rect 29036 12460 29428 12516
rect 28812 12238 28814 12290
rect 28866 12238 28868 12290
rect 25900 11394 25956 11676
rect 26572 11900 26852 11956
rect 27356 12180 27412 12190
rect 25900 11342 25902 11394
rect 25954 11342 25956 11394
rect 25900 11330 25956 11342
rect 26012 11396 26068 11406
rect 26012 11302 26068 11340
rect 26572 11394 26628 11900
rect 26572 11342 26574 11394
rect 26626 11342 26628 11394
rect 26572 11330 26628 11342
rect 26796 11732 26852 11742
rect 26124 11172 26180 11182
rect 25788 11170 26180 11172
rect 25788 11118 26126 11170
rect 26178 11118 26180 11170
rect 25788 11116 26180 11118
rect 26124 10724 26180 11116
rect 26796 10834 26852 11676
rect 27356 11618 27412 12124
rect 27580 12178 27636 12190
rect 27580 12126 27582 12178
rect 27634 12126 27636 12178
rect 27580 11732 27636 12126
rect 27580 11666 27636 11676
rect 27916 12178 27972 12190
rect 27916 12126 27918 12178
rect 27970 12126 27972 12178
rect 27356 11566 27358 11618
rect 27410 11566 27412 11618
rect 27356 11554 27412 11566
rect 27132 11508 27188 11518
rect 27132 11414 27188 11452
rect 27468 11396 27524 11406
rect 27916 11396 27972 12126
rect 28364 11732 28420 11742
rect 28364 11506 28420 11676
rect 28364 11454 28366 11506
rect 28418 11454 28420 11506
rect 28364 11442 28420 11454
rect 27468 11394 27972 11396
rect 27468 11342 27470 11394
rect 27522 11342 27972 11394
rect 27468 11340 27972 11342
rect 27468 11330 27524 11340
rect 26796 10782 26798 10834
rect 26850 10782 26852 10834
rect 26796 10770 26852 10782
rect 26124 10658 26180 10668
rect 27244 10724 27300 10734
rect 27244 10630 27300 10668
rect 27580 10610 27636 11340
rect 27580 10558 27582 10610
rect 27634 10558 27636 10610
rect 25116 9938 25172 10108
rect 26796 10500 26852 10510
rect 26684 9940 26740 9950
rect 25116 9886 25118 9938
rect 25170 9886 25172 9938
rect 25116 9874 25172 9886
rect 26236 9938 26740 9940
rect 26236 9886 26686 9938
rect 26738 9886 26740 9938
rect 26236 9884 26740 9886
rect 25228 9604 25284 9614
rect 25228 9044 25284 9548
rect 25228 8950 25284 8988
rect 26012 8930 26068 8942
rect 26012 8878 26014 8930
rect 26066 8878 26068 8930
rect 26012 8484 26068 8878
rect 26124 8484 26180 8494
rect 26012 8482 26180 8484
rect 26012 8430 26126 8482
rect 26178 8430 26180 8482
rect 26012 8428 26180 8430
rect 26124 8418 26180 8428
rect 26236 8370 26292 9884
rect 26684 9874 26740 9884
rect 26684 9602 26740 9614
rect 26684 9550 26686 9602
rect 26738 9550 26740 9602
rect 26684 9268 26740 9550
rect 26684 9202 26740 9212
rect 26796 9602 26852 10444
rect 27244 10052 27300 10062
rect 27020 9828 27076 9838
rect 27020 9734 27076 9772
rect 27244 9826 27300 9996
rect 27244 9774 27246 9826
rect 27298 9774 27300 9826
rect 27244 9762 27300 9774
rect 26796 9550 26798 9602
rect 26850 9550 26852 9602
rect 26796 9156 26852 9550
rect 26796 9090 26852 9100
rect 26236 8318 26238 8370
rect 26290 8318 26292 8370
rect 26236 8306 26292 8318
rect 27020 9044 27076 9054
rect 27020 7700 27076 8988
rect 27580 8932 27636 10558
rect 27804 10052 27860 10062
rect 27804 9826 27860 9996
rect 28812 10052 28868 12238
rect 29036 12066 29092 12460
rect 29820 12404 29876 12414
rect 29820 12310 29876 12348
rect 29036 12014 29038 12066
rect 29090 12014 29092 12066
rect 29036 12002 29092 12014
rect 29148 12292 29204 12302
rect 29148 12178 29204 12236
rect 29596 12292 29652 12302
rect 29596 12198 29652 12236
rect 29148 12126 29150 12178
rect 29202 12126 29204 12178
rect 29148 11284 29204 12126
rect 29484 12180 29540 12190
rect 29484 12086 29540 12124
rect 29148 11218 29204 11228
rect 29932 11284 29988 11294
rect 29932 11190 29988 11228
rect 30044 11282 30100 11294
rect 30044 11230 30046 11282
rect 30098 11230 30100 11282
rect 30044 10052 30100 11230
rect 28868 9996 29204 10052
rect 28812 9986 28868 9996
rect 27804 9774 27806 9826
rect 27858 9774 27860 9826
rect 27804 9762 27860 9774
rect 28028 9828 28084 9838
rect 28028 9734 28084 9772
rect 28252 9714 28308 9726
rect 28252 9662 28254 9714
rect 28306 9662 28308 9714
rect 27692 9602 27748 9614
rect 27692 9550 27694 9602
rect 27746 9550 27748 9602
rect 27692 9268 27748 9550
rect 27916 9604 27972 9614
rect 27916 9510 27972 9548
rect 28252 9492 28308 9662
rect 28252 9426 28308 9436
rect 28588 9604 28644 9614
rect 27692 9202 27748 9212
rect 28588 9154 28644 9548
rect 29148 9266 29204 9996
rect 29708 9996 30044 10052
rect 29708 9938 29764 9996
rect 29708 9886 29710 9938
rect 29762 9886 29764 9938
rect 29708 9874 29764 9886
rect 29148 9214 29150 9266
rect 29202 9214 29204 9266
rect 29148 9202 29204 9214
rect 28588 9102 28590 9154
rect 28642 9102 28644 9154
rect 28588 9090 28644 9102
rect 29484 9044 29540 9054
rect 29484 8950 29540 8988
rect 28140 8932 28196 8942
rect 27580 8930 28196 8932
rect 27580 8878 28142 8930
rect 28194 8878 28196 8930
rect 27580 8876 28196 8878
rect 28140 8866 28196 8876
rect 30044 8930 30100 9996
rect 30044 8878 30046 8930
rect 30098 8878 30100 8930
rect 30044 8866 30100 8878
rect 28476 8820 28532 8830
rect 28252 8818 28532 8820
rect 28252 8766 28478 8818
rect 28530 8766 28532 8818
rect 28252 8764 28532 8766
rect 27020 7698 27412 7700
rect 27020 7646 27022 7698
rect 27074 7646 27412 7698
rect 27020 7644 27412 7646
rect 27020 7634 27076 7644
rect 27356 7474 27412 7644
rect 28140 7588 28196 7598
rect 28252 7588 28308 8764
rect 28476 8754 28532 8764
rect 28140 7586 28308 7588
rect 28140 7534 28142 7586
rect 28194 7534 28308 7586
rect 28140 7532 28308 7534
rect 28140 7522 28196 7532
rect 27356 7422 27358 7474
rect 27410 7422 27412 7474
rect 27356 7410 27412 7422
rect 25004 3614 25006 3666
rect 25058 3614 25060 3666
rect 25004 3602 25060 3614
rect 18620 3502 18622 3554
rect 18674 3502 18676 3554
rect 18620 3444 18676 3502
rect 29148 3556 29204 3566
rect 29148 3554 29876 3556
rect 29148 3502 29150 3554
rect 29202 3502 29876 3554
rect 29148 3500 29876 3502
rect 29148 3490 29204 3500
rect 18620 3378 18676 3388
rect 24108 3444 24164 3454
rect 24556 3444 24612 3454
rect 24108 3442 24612 3444
rect 24108 3390 24110 3442
rect 24162 3390 24558 3442
rect 24610 3390 24612 3442
rect 24108 3388 24612 3390
rect 24108 3378 24164 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 24220 800 24276 3388
rect 24556 3378 24612 3388
rect 29820 3442 29876 3500
rect 29820 3390 29822 3442
rect 29874 3390 29876 3442
rect 29596 3332 29652 3342
rect 29596 3238 29652 3276
rect 29820 2324 29876 3390
rect 30156 3442 30212 17388
rect 30492 17350 30548 17388
rect 30268 16996 30324 17006
rect 30268 16902 30324 16940
rect 30716 15148 30772 20524
rect 30940 20020 30996 21532
rect 31052 20916 31108 20926
rect 31052 20822 31108 20860
rect 31164 20580 31220 21532
rect 31276 21522 31332 21532
rect 31388 21586 31444 21598
rect 31388 21534 31390 21586
rect 31442 21534 31444 21586
rect 31388 20916 31444 21534
rect 31836 21586 31892 21598
rect 31836 21534 31838 21586
rect 31890 21534 31892 21586
rect 31388 20850 31444 20860
rect 31500 21476 31556 21486
rect 31052 20020 31108 20030
rect 30940 20018 31108 20020
rect 30940 19966 31054 20018
rect 31106 19966 31108 20018
rect 30940 19964 31108 19966
rect 31052 19954 31108 19964
rect 30940 18452 30996 18462
rect 30940 18116 30996 18396
rect 30940 18050 30996 18060
rect 31052 18004 31108 18014
rect 30940 17780 30996 17790
rect 30940 16996 30996 17724
rect 31052 17666 31108 17948
rect 31052 17614 31054 17666
rect 31106 17614 31108 17666
rect 31052 17220 31108 17614
rect 31052 17154 31108 17164
rect 31164 17444 31220 20524
rect 31500 20468 31556 21420
rect 31276 19348 31332 19358
rect 31276 19254 31332 19292
rect 31388 18452 31444 18462
rect 31500 18452 31556 20412
rect 31836 19908 31892 21534
rect 31948 20130 32004 22094
rect 32396 22036 32452 22316
rect 32620 22148 32676 22430
rect 33180 22372 33236 22382
rect 33292 22372 33348 23548
rect 33628 23380 33684 26852
rect 33740 26178 33796 26190
rect 33964 26180 34020 26190
rect 33740 26126 33742 26178
rect 33794 26126 33796 26178
rect 33740 25956 33796 26126
rect 33740 25890 33796 25900
rect 33852 26124 33964 26180
rect 33852 24164 33908 26124
rect 33964 26086 34020 26124
rect 33964 25282 34020 25294
rect 33964 25230 33966 25282
rect 34018 25230 34020 25282
rect 33964 24724 34020 25230
rect 34076 25284 34132 28588
rect 34188 27748 34244 27758
rect 34188 27746 34468 27748
rect 34188 27694 34190 27746
rect 34242 27694 34468 27746
rect 34188 27692 34468 27694
rect 34188 27682 34244 27692
rect 34188 27300 34244 27310
rect 34188 27186 34244 27244
rect 34188 27134 34190 27186
rect 34242 27134 34244 27186
rect 34188 27122 34244 27134
rect 34412 27074 34468 27692
rect 34412 27022 34414 27074
rect 34466 27022 34468 27074
rect 34412 27010 34468 27022
rect 34412 26290 34468 26302
rect 34412 26238 34414 26290
rect 34466 26238 34468 26290
rect 34412 25956 34468 26238
rect 34412 25890 34468 25900
rect 34076 25218 34132 25228
rect 34188 25844 34244 25854
rect 34188 25618 34244 25788
rect 34188 25566 34190 25618
rect 34242 25566 34244 25618
rect 33964 24658 34020 24668
rect 34188 24164 34244 25566
rect 33516 23324 33628 23380
rect 33404 22596 33460 22606
rect 33404 22502 33460 22540
rect 33516 22372 33572 23324
rect 33628 23314 33684 23324
rect 33740 24108 33908 24164
rect 33964 24108 34244 24164
rect 33180 22370 33348 22372
rect 33180 22318 33182 22370
rect 33234 22318 33348 22370
rect 33180 22316 33348 22318
rect 33404 22316 33572 22372
rect 33628 23154 33684 23166
rect 33628 23102 33630 23154
rect 33682 23102 33684 23154
rect 33628 22372 33684 23102
rect 32620 22082 32676 22092
rect 32956 22260 33012 22270
rect 32172 21812 32228 21822
rect 32172 21754 32228 21756
rect 32172 21702 32174 21754
rect 32226 21702 32228 21754
rect 32172 21690 32228 21702
rect 32284 21698 32340 21710
rect 32284 21646 32286 21698
rect 32338 21646 32340 21698
rect 32284 21588 32340 21646
rect 32172 21532 32340 21588
rect 31948 20078 31950 20130
rect 32002 20078 32004 20130
rect 31948 20066 32004 20078
rect 32060 20132 32116 20142
rect 32172 20132 32228 21532
rect 32284 21364 32340 21374
rect 32284 21270 32340 21308
rect 32060 20130 32228 20132
rect 32060 20078 32062 20130
rect 32114 20078 32228 20130
rect 32060 20076 32228 20078
rect 32060 20066 32116 20076
rect 31836 19852 32116 19908
rect 32060 19794 32116 19852
rect 32060 19742 32062 19794
rect 32114 19742 32116 19794
rect 32060 19730 32116 19742
rect 32172 19572 32228 20076
rect 32060 19516 32228 19572
rect 31612 19348 31668 19358
rect 31612 19234 31668 19292
rect 31612 19182 31614 19234
rect 31666 19182 31668 19234
rect 31612 19170 31668 19182
rect 31836 19010 31892 19022
rect 31836 18958 31838 19010
rect 31890 18958 31892 19010
rect 31836 18900 31892 18958
rect 32060 18900 32116 19516
rect 32396 19460 32452 21980
rect 32956 21476 33012 22204
rect 33180 21924 33236 22316
rect 33180 21858 33236 21868
rect 33180 21476 33236 21486
rect 32956 21474 33236 21476
rect 32956 21422 33182 21474
rect 33234 21422 33236 21474
rect 32956 21420 33236 21422
rect 32956 20356 33012 20366
rect 33068 20356 33124 21420
rect 33180 21410 33236 21420
rect 33180 20916 33236 20926
rect 33180 20822 33236 20860
rect 33012 20300 33124 20356
rect 32956 20290 33012 20300
rect 33292 19796 33348 19806
rect 32172 19404 32452 19460
rect 32508 19404 33124 19460
rect 32172 19012 32228 19404
rect 32508 19348 32564 19404
rect 32284 19292 32564 19348
rect 32284 19234 32340 19292
rect 32284 19182 32286 19234
rect 32338 19182 32340 19234
rect 32284 19170 32340 19182
rect 32844 19236 32900 19246
rect 32844 19142 32900 19180
rect 32396 19122 32452 19134
rect 32396 19070 32398 19122
rect 32450 19070 32452 19122
rect 32396 19012 32452 19070
rect 32172 18956 32452 19012
rect 32508 19010 32564 19022
rect 32508 18958 32510 19010
rect 32562 18958 32564 19010
rect 31836 18844 32228 18900
rect 31388 18450 31556 18452
rect 31388 18398 31390 18450
rect 31442 18398 31556 18450
rect 31388 18396 31556 18398
rect 31612 18562 31668 18574
rect 31612 18510 31614 18562
rect 31666 18510 31668 18562
rect 31388 17780 31444 18396
rect 31612 18228 31668 18510
rect 32060 18562 32116 18574
rect 32060 18510 32062 18562
rect 32114 18510 32116 18562
rect 32060 18452 32116 18510
rect 31948 18340 32004 18350
rect 31948 18246 32004 18284
rect 31388 17714 31444 17724
rect 31500 18172 31612 18228
rect 31276 17444 31332 17454
rect 31164 17442 31332 17444
rect 31164 17390 31278 17442
rect 31330 17390 31332 17442
rect 31164 17388 31332 17390
rect 31052 16996 31108 17006
rect 30940 16994 31108 16996
rect 30940 16942 31054 16994
rect 31106 16942 31108 16994
rect 30940 16940 31108 16942
rect 31164 16996 31220 17388
rect 31276 17378 31332 17388
rect 31164 16940 31444 16996
rect 31052 16930 31108 16940
rect 31276 16324 31332 16334
rect 31164 16268 31276 16324
rect 31052 15428 31108 15438
rect 31052 15314 31108 15372
rect 31052 15262 31054 15314
rect 31106 15262 31108 15314
rect 31052 15250 31108 15262
rect 31164 15202 31220 16268
rect 31276 16258 31332 16268
rect 31164 15150 31166 15202
rect 31218 15150 31220 15202
rect 30604 15092 30660 15102
rect 30716 15092 30996 15148
rect 31164 15138 31220 15150
rect 31276 15428 31332 15438
rect 30604 14998 30660 15036
rect 30716 14418 30772 14430
rect 30716 14366 30718 14418
rect 30770 14366 30772 14418
rect 30716 12964 30772 14366
rect 30940 13970 30996 15092
rect 30940 13918 30942 13970
rect 30994 13918 30996 13970
rect 30940 13412 30996 13918
rect 31164 14530 31220 14542
rect 31164 14478 31166 14530
rect 31218 14478 31220 14530
rect 31164 13972 31220 14478
rect 31164 13906 31220 13916
rect 31052 13860 31108 13870
rect 31052 13748 31108 13804
rect 31164 13748 31220 13758
rect 31052 13746 31220 13748
rect 31052 13694 31166 13746
rect 31218 13694 31220 13746
rect 31052 13692 31220 13694
rect 31164 13682 31220 13692
rect 30940 13346 30996 13356
rect 31276 13300 31332 15372
rect 31052 13244 31332 13300
rect 30940 12964 30996 12974
rect 30716 12898 30772 12908
rect 30828 12962 30996 12964
rect 30828 12910 30942 12962
rect 30994 12910 30996 12962
rect 30828 12908 30996 12910
rect 30828 12740 30884 12908
rect 30940 12898 30996 12908
rect 30380 12684 30884 12740
rect 30380 12402 30436 12684
rect 30380 12350 30382 12402
rect 30434 12350 30436 12402
rect 30380 12338 30436 12350
rect 30940 12404 30996 12414
rect 30492 12292 30548 12302
rect 30716 12292 30772 12302
rect 30268 12178 30324 12190
rect 30268 12126 30270 12178
rect 30322 12126 30324 12178
rect 30268 11396 30324 12126
rect 30268 11302 30324 11340
rect 30492 12178 30548 12236
rect 30492 12126 30494 12178
rect 30546 12126 30548 12178
rect 30492 10948 30548 12126
rect 30604 12290 30772 12292
rect 30604 12238 30718 12290
rect 30770 12238 30772 12290
rect 30604 12236 30772 12238
rect 30604 11170 30660 12236
rect 30716 12226 30772 12236
rect 30940 11394 30996 12348
rect 30940 11342 30942 11394
rect 30994 11342 30996 11394
rect 30604 11118 30606 11170
rect 30658 11118 30660 11170
rect 30604 11106 30660 11118
rect 30716 11284 30772 11294
rect 30716 11282 30884 11284
rect 30716 11230 30718 11282
rect 30770 11230 30884 11282
rect 30716 11228 30884 11230
rect 30716 10948 30772 11228
rect 30492 10892 30772 10948
rect 30268 9044 30324 9054
rect 30268 7362 30324 8988
rect 30828 8930 30884 11228
rect 30940 10386 30996 11342
rect 30940 10334 30942 10386
rect 30994 10334 30996 10386
rect 30940 10322 30996 10334
rect 30828 8878 30830 8930
rect 30882 8878 30884 8930
rect 30828 8866 30884 8878
rect 31052 8708 31108 13244
rect 31388 13188 31444 16940
rect 31164 13132 31444 13188
rect 31164 11396 31220 13132
rect 31500 13076 31556 18172
rect 31612 18162 31668 18172
rect 32060 17780 32116 18396
rect 32060 17714 32116 17724
rect 31724 17556 31780 17566
rect 31724 17462 31780 17500
rect 31836 16100 31892 16110
rect 31836 16098 32004 16100
rect 31836 16046 31838 16098
rect 31890 16046 32004 16098
rect 31836 16044 32004 16046
rect 31836 16034 31892 16044
rect 31836 15540 31892 15550
rect 31836 15314 31892 15484
rect 31948 15428 32004 16044
rect 31948 15362 32004 15372
rect 32060 16098 32116 16110
rect 32060 16046 32062 16098
rect 32114 16046 32116 16098
rect 31836 15262 31838 15314
rect 31890 15262 31892 15314
rect 31836 15250 31892 15262
rect 31612 15204 31668 15214
rect 31612 14642 31668 15148
rect 31612 14590 31614 14642
rect 31666 14590 31668 14642
rect 31612 14578 31668 14590
rect 32060 15092 32116 16046
rect 31612 13972 31668 13982
rect 32060 13972 32116 15036
rect 31668 13916 32116 13972
rect 31612 13524 31668 13916
rect 31724 13748 31780 13758
rect 31724 13746 31892 13748
rect 31724 13694 31726 13746
rect 31778 13694 31892 13746
rect 31724 13692 31892 13694
rect 31724 13682 31780 13692
rect 31612 13468 31780 13524
rect 31276 13020 31556 13076
rect 31276 12852 31332 13020
rect 31612 12964 31668 12974
rect 31612 12870 31668 12908
rect 31388 12852 31444 12862
rect 31276 12796 31388 12852
rect 31388 12758 31444 12796
rect 31500 12738 31556 12750
rect 31500 12686 31502 12738
rect 31554 12686 31556 12738
rect 31500 12628 31556 12686
rect 31500 12562 31556 12572
rect 31612 12404 31668 12414
rect 31612 12178 31668 12348
rect 31612 12126 31614 12178
rect 31666 12126 31668 12178
rect 31612 12114 31668 12126
rect 31276 11396 31332 11406
rect 31164 11340 31276 11396
rect 31276 11302 31332 11340
rect 31500 11284 31556 11294
rect 31500 11190 31556 11228
rect 31388 11170 31444 11182
rect 31388 11118 31390 11170
rect 31442 11118 31444 11170
rect 31276 10498 31332 10510
rect 31276 10446 31278 10498
rect 31330 10446 31332 10498
rect 31276 10386 31332 10446
rect 31276 10334 31278 10386
rect 31330 10334 31332 10386
rect 31276 10322 31332 10334
rect 31388 9716 31444 11118
rect 31724 10500 31780 13468
rect 31836 13412 31892 13692
rect 31836 12404 31892 13356
rect 31948 12850 32004 12862
rect 31948 12798 31950 12850
rect 32002 12798 32004 12850
rect 31948 12628 32004 12798
rect 31948 12562 32004 12572
rect 32060 12852 32116 12862
rect 32172 12852 32228 18844
rect 32508 18676 32564 18958
rect 32956 19012 33012 19022
rect 32956 18918 33012 18956
rect 33068 19012 33124 19404
rect 33292 19234 33348 19740
rect 33292 19182 33294 19234
rect 33346 19182 33348 19234
rect 33292 19170 33348 19182
rect 33068 19010 33348 19012
rect 33068 18958 33070 19010
rect 33122 18958 33348 19010
rect 33068 18956 33348 18958
rect 33068 18946 33124 18956
rect 32284 18620 32564 18676
rect 32284 18562 32340 18620
rect 32284 18510 32286 18562
rect 32338 18510 32340 18562
rect 32284 18498 32340 18510
rect 33068 18452 33124 18462
rect 33068 18358 33124 18396
rect 33292 18450 33348 18956
rect 33292 18398 33294 18450
rect 33346 18398 33348 18450
rect 32620 18340 32676 18350
rect 32620 17778 32676 18284
rect 33180 18340 33236 18350
rect 33180 18246 33236 18284
rect 33292 18116 33348 18398
rect 32620 17726 32622 17778
rect 32674 17726 32676 17778
rect 32620 17714 32676 17726
rect 33180 18060 33348 18116
rect 32396 17668 32452 17678
rect 32396 17574 32452 17612
rect 33068 17668 33124 17678
rect 33180 17668 33236 18060
rect 33068 17666 33236 17668
rect 33068 17614 33070 17666
rect 33122 17614 33236 17666
rect 33068 17612 33236 17614
rect 33292 17668 33348 17678
rect 33068 17220 33124 17612
rect 33292 17574 33348 17612
rect 32844 17164 33124 17220
rect 33180 17444 33236 17454
rect 32508 16884 32564 16894
rect 32284 16100 32340 16110
rect 32508 16100 32564 16828
rect 32284 16098 32564 16100
rect 32284 16046 32286 16098
rect 32338 16046 32564 16098
rect 32284 16044 32564 16046
rect 32284 16034 32340 16044
rect 32508 15538 32564 16044
rect 32732 15988 32788 15998
rect 32732 15894 32788 15932
rect 32508 15486 32510 15538
rect 32562 15486 32564 15538
rect 32508 15474 32564 15486
rect 32620 15540 32676 15550
rect 32844 15540 32900 17164
rect 33180 16884 33236 17388
rect 33068 16324 33124 16334
rect 33068 16230 33124 16268
rect 33180 16100 33236 16828
rect 33292 16548 33348 16558
rect 33404 16548 33460 22316
rect 33628 22278 33684 22316
rect 33628 22148 33684 22158
rect 33516 22092 33628 22148
rect 33516 19236 33572 22092
rect 33628 22082 33684 22092
rect 33740 21700 33796 24108
rect 33852 23938 33908 23950
rect 33852 23886 33854 23938
rect 33906 23886 33908 23938
rect 33852 23268 33908 23886
rect 33964 23380 34020 24108
rect 34076 23940 34132 23950
rect 34076 23938 34356 23940
rect 34076 23886 34078 23938
rect 34130 23886 34356 23938
rect 34076 23884 34356 23886
rect 34076 23874 34132 23884
rect 33964 23324 34244 23380
rect 33852 22596 33908 23212
rect 34076 23156 34132 23166
rect 33964 23044 34020 23054
rect 33964 22950 34020 22988
rect 34076 22708 34132 23100
rect 34076 22642 34132 22652
rect 33852 22530 33908 22540
rect 34076 22148 34132 22158
rect 34076 22054 34132 22092
rect 33740 21634 33796 21644
rect 33964 21924 34020 21934
rect 33964 21476 34020 21868
rect 33740 21474 34020 21476
rect 33740 21422 33966 21474
rect 34018 21422 34020 21474
rect 33740 21420 34020 21422
rect 33516 18452 33572 19180
rect 33516 17890 33572 18396
rect 33516 17838 33518 17890
rect 33570 17838 33572 17890
rect 33516 17826 33572 17838
rect 33628 20132 33684 20142
rect 33628 18450 33684 20076
rect 33628 18398 33630 18450
rect 33682 18398 33684 18450
rect 33628 16772 33684 18398
rect 33628 16706 33684 16716
rect 33348 16492 33460 16548
rect 33292 16482 33348 16492
rect 33180 16098 33572 16100
rect 33180 16046 33182 16098
rect 33234 16046 33572 16098
rect 33180 16044 33572 16046
rect 33180 16034 33236 16044
rect 33068 15988 33124 15998
rect 33068 15894 33124 15932
rect 33292 15876 33348 15886
rect 33348 15820 33460 15876
rect 33292 15810 33348 15820
rect 32284 15428 32340 15438
rect 32284 15334 32340 15372
rect 32396 15204 32452 15242
rect 32396 15138 32452 15148
rect 32620 14642 32676 15484
rect 32620 14590 32622 14642
rect 32674 14590 32676 14642
rect 32620 14578 32676 14590
rect 32732 15484 32900 15540
rect 32060 12850 32228 12852
rect 32060 12798 32062 12850
rect 32114 12798 32228 12850
rect 32060 12796 32228 12798
rect 31836 12338 31892 12348
rect 32060 12404 32116 12796
rect 32284 12740 32340 12750
rect 32060 12338 32116 12348
rect 32172 12738 32340 12740
rect 32172 12686 32286 12738
rect 32338 12686 32340 12738
rect 32172 12684 32340 12686
rect 32060 12068 32116 12078
rect 32060 11974 32116 12012
rect 32172 11844 32228 12684
rect 32284 12674 32340 12684
rect 32508 12740 32564 12750
rect 32508 12292 32564 12684
rect 32508 12198 32564 12236
rect 31836 11788 32228 11844
rect 31836 11394 31892 11788
rect 31836 11342 31838 11394
rect 31890 11342 31892 11394
rect 31836 11330 31892 11342
rect 32172 11396 32228 11406
rect 32172 11302 32228 11340
rect 31388 9650 31444 9660
rect 31500 10444 31780 10500
rect 32284 11170 32340 11182
rect 32284 11118 32286 11170
rect 32338 11118 32340 11170
rect 30268 7310 30270 7362
rect 30322 7310 30324 7362
rect 30268 7298 30324 7310
rect 30828 8652 31108 8708
rect 30156 3390 30158 3442
rect 30210 3390 30212 3442
rect 30156 3378 30212 3390
rect 30268 3444 30324 3454
rect 30492 3442 30548 3454
rect 30492 3390 30494 3442
rect 30546 3390 30548 3442
rect 30492 3388 30548 3390
rect 29596 2268 29876 2324
rect 30268 3332 30548 3388
rect 30828 3442 30884 8652
rect 31500 8484 31556 10444
rect 31836 9716 31892 9726
rect 31836 9622 31892 9660
rect 31500 8428 31668 8484
rect 31500 8260 31556 8270
rect 31500 8166 31556 8204
rect 30828 3390 30830 3442
rect 30882 3390 30884 3442
rect 30828 3378 30884 3390
rect 30940 4226 30996 4238
rect 30940 4174 30942 4226
rect 30994 4174 30996 4226
rect 30940 3556 30996 4174
rect 31164 3556 31220 3566
rect 30940 3554 31220 3556
rect 30940 3502 31166 3554
rect 31218 3502 31220 3554
rect 30940 3500 31220 3502
rect 29596 800 29652 2268
rect 30268 800 30324 3332
rect 30940 800 30996 3500
rect 31164 3490 31220 3500
rect 31500 3444 31556 3454
rect 31612 3444 31668 8428
rect 32172 8372 32228 8382
rect 32284 8372 32340 11118
rect 32396 11170 32452 11182
rect 32396 11118 32398 11170
rect 32450 11118 32452 11170
rect 32396 10612 32452 11118
rect 32396 10546 32452 10556
rect 32732 10052 32788 15484
rect 33068 15428 33124 15438
rect 33068 15334 33124 15372
rect 33292 15314 33348 15326
rect 33292 15262 33294 15314
rect 33346 15262 33348 15314
rect 33292 15092 33348 15262
rect 33292 15026 33348 15036
rect 33180 14642 33236 14654
rect 33180 14590 33182 14642
rect 33234 14590 33236 14642
rect 32844 14418 32900 14430
rect 32844 14366 32846 14418
rect 32898 14366 32900 14418
rect 32844 12852 32900 14366
rect 33180 13524 33236 14590
rect 33292 14532 33348 14542
rect 33292 14438 33348 14476
rect 33404 14308 33460 15820
rect 33516 15314 33572 16044
rect 33740 15540 33796 21420
rect 33964 21410 34020 21420
rect 33964 20804 34020 20814
rect 33964 20710 34020 20748
rect 33964 17444 34020 17454
rect 33964 17350 34020 17388
rect 34188 17220 34244 23324
rect 34300 22484 34356 23884
rect 34524 23548 34580 29484
rect 34636 28756 34692 30156
rect 34860 30146 34916 30156
rect 34860 29988 34916 29998
rect 34860 29894 34916 29932
rect 35084 29538 35140 30268
rect 35532 30212 35588 30222
rect 35420 30100 35476 30110
rect 35532 30100 35588 30156
rect 35868 30212 35924 30222
rect 36316 30212 36372 30604
rect 36428 30548 36484 32956
rect 36652 31892 36708 33964
rect 36764 33908 36820 33918
rect 36764 33814 36820 33852
rect 37436 33684 37492 34636
rect 37660 34626 37716 34636
rect 37436 33618 37492 33628
rect 37548 34132 37604 34142
rect 38108 34132 38164 35532
rect 39116 35140 39172 36430
rect 39228 36260 39284 38444
rect 39564 38500 39620 40462
rect 39564 38434 39620 38444
rect 39676 38276 39732 38286
rect 39452 38274 39732 38276
rect 39452 38222 39678 38274
rect 39730 38222 39732 38274
rect 39452 38220 39732 38222
rect 39452 37490 39508 38220
rect 39676 38210 39732 38220
rect 39788 37492 39844 40572
rect 39900 40404 39956 40414
rect 40012 40404 40068 42140
rect 40124 42130 40180 42140
rect 40236 40628 40292 42588
rect 40348 42578 40404 42588
rect 40348 41858 40404 41870
rect 40348 41806 40350 41858
rect 40402 41806 40404 41858
rect 40348 40740 40404 41806
rect 41020 41412 41076 43374
rect 41580 42980 41636 44046
rect 41580 42914 41636 42924
rect 41692 42308 41748 45726
rect 42140 45108 42196 45118
rect 41804 44994 41860 45006
rect 41804 44942 41806 44994
rect 41858 44942 41860 44994
rect 41804 44322 41860 44942
rect 41804 44270 41806 44322
rect 41858 44270 41860 44322
rect 41804 44258 41860 44270
rect 42140 44324 42196 45052
rect 42252 44996 42308 45006
rect 42252 44994 42420 44996
rect 42252 44942 42254 44994
rect 42306 44942 42420 44994
rect 42252 44940 42420 44942
rect 42252 44930 42308 44940
rect 42140 43764 42196 44268
rect 42140 43538 42196 43708
rect 42140 43486 42142 43538
rect 42194 43486 42196 43538
rect 42140 43474 42196 43486
rect 42028 43316 42084 43326
rect 41692 42252 41860 42308
rect 41580 42196 41636 42206
rect 41580 42102 41636 42140
rect 41020 41346 41076 41356
rect 41244 41970 41300 41982
rect 41244 41918 41246 41970
rect 41298 41918 41300 41970
rect 41244 40740 41300 41918
rect 41580 41860 41636 41870
rect 40348 40684 41300 40740
rect 41468 41412 41524 41422
rect 41468 40852 41524 41356
rect 40236 40572 40740 40628
rect 39900 40402 40068 40404
rect 39900 40350 39902 40402
rect 39954 40350 40068 40402
rect 39900 40348 40068 40350
rect 39900 40338 39956 40348
rect 40348 39956 40404 39966
rect 40348 38722 40404 39900
rect 40348 38670 40350 38722
rect 40402 38670 40404 38722
rect 40348 38658 40404 38670
rect 40012 38274 40068 38286
rect 40012 38222 40014 38274
rect 40066 38222 40068 38274
rect 40012 38052 40068 38222
rect 40348 38164 40404 38174
rect 40236 38052 40292 38062
rect 40012 38050 40292 38052
rect 40012 37998 40238 38050
rect 40290 37998 40292 38050
rect 40012 37996 40292 37998
rect 40236 37986 40292 37996
rect 40012 37828 40068 37838
rect 40348 37828 40404 38108
rect 40684 38050 40740 40572
rect 40908 39844 40964 40684
rect 41468 40626 41524 40796
rect 41468 40574 41470 40626
rect 41522 40574 41524 40626
rect 41468 40562 41524 40574
rect 41020 40516 41076 40526
rect 41356 40516 41412 40526
rect 41020 40514 41356 40516
rect 41020 40462 41022 40514
rect 41074 40462 41356 40514
rect 41020 40460 41356 40462
rect 41020 40450 41076 40460
rect 41356 40422 41412 40460
rect 41580 40404 41636 41804
rect 41692 41524 41748 41534
rect 41692 41298 41748 41468
rect 41692 41246 41694 41298
rect 41746 41246 41748 41298
rect 41692 41234 41748 41246
rect 41692 40628 41748 40638
rect 41692 40534 41748 40572
rect 41020 39844 41076 39854
rect 40908 39788 41020 39844
rect 41020 39778 41076 39788
rect 41468 39620 41524 39630
rect 41580 39620 41636 40348
rect 41468 39618 41636 39620
rect 41468 39566 41470 39618
rect 41522 39566 41636 39618
rect 41468 39564 41636 39566
rect 41244 39508 41300 39518
rect 40684 37998 40686 38050
rect 40738 37998 40740 38050
rect 40684 37986 40740 37998
rect 40908 38164 40964 38174
rect 40908 38050 40964 38108
rect 40908 37998 40910 38050
rect 40962 37998 40964 38050
rect 40908 37986 40964 37998
rect 40572 37940 40628 37950
rect 40572 37846 40628 37884
rect 40012 37826 40404 37828
rect 40012 37774 40014 37826
rect 40066 37774 40404 37826
rect 40012 37772 40404 37774
rect 40460 37826 40516 37838
rect 40460 37774 40462 37826
rect 40514 37774 40516 37826
rect 40012 37604 40068 37772
rect 40460 37604 40516 37774
rect 40012 37538 40068 37548
rect 40124 37548 40516 37604
rect 39452 37438 39454 37490
rect 39506 37438 39508 37490
rect 39452 37426 39508 37438
rect 39676 37436 39844 37492
rect 40124 37490 40180 37548
rect 40124 37438 40126 37490
rect 40178 37438 40180 37490
rect 39340 37156 39396 37166
rect 39340 37062 39396 37100
rect 39676 36596 39732 37436
rect 40124 37426 40180 37438
rect 39900 37378 39956 37390
rect 39900 37326 39902 37378
rect 39954 37326 39956 37378
rect 39788 37268 39844 37278
rect 39788 36820 39844 37212
rect 39900 37156 39956 37326
rect 40348 37380 40404 37390
rect 40348 37156 40404 37324
rect 41132 37380 41188 37390
rect 41132 37286 41188 37324
rect 40908 37268 40964 37278
rect 40908 37174 40964 37212
rect 39900 37100 40404 37156
rect 39788 36764 39956 36820
rect 39788 36596 39844 36606
rect 39676 36594 39844 36596
rect 39676 36542 39790 36594
rect 39842 36542 39844 36594
rect 39676 36540 39844 36542
rect 39788 36530 39844 36540
rect 39564 36484 39620 36494
rect 39564 36390 39620 36428
rect 39228 36204 39732 36260
rect 39676 36036 39732 36204
rect 39676 35922 39732 35980
rect 39676 35870 39678 35922
rect 39730 35870 39732 35922
rect 39676 35858 39732 35870
rect 39900 35922 39956 36764
rect 40236 36484 40292 36494
rect 40236 36390 40292 36428
rect 39900 35870 39902 35922
rect 39954 35870 39956 35922
rect 39900 35858 39956 35870
rect 40124 36258 40180 36270
rect 40124 36206 40126 36258
rect 40178 36206 40180 36258
rect 39564 35698 39620 35710
rect 39564 35646 39566 35698
rect 39618 35646 39620 35698
rect 39564 35252 39620 35646
rect 40124 35588 40180 36206
rect 40348 36258 40404 37100
rect 41020 37156 41076 37166
rect 41020 37062 41076 37100
rect 40908 36932 40964 36942
rect 40348 36206 40350 36258
rect 40402 36206 40404 36258
rect 40236 36036 40292 36046
rect 40236 35922 40292 35980
rect 40236 35870 40238 35922
rect 40290 35870 40292 35922
rect 40236 35858 40292 35870
rect 39788 35532 40180 35588
rect 39788 35252 39844 35532
rect 39564 35196 39844 35252
rect 39116 35084 39732 35140
rect 39228 34914 39284 34926
rect 39228 34862 39230 34914
rect 39282 34862 39284 34914
rect 38556 34802 38612 34814
rect 38556 34750 38558 34802
rect 38610 34750 38612 34802
rect 38220 34690 38276 34702
rect 38220 34638 38222 34690
rect 38274 34638 38276 34690
rect 38220 34242 38276 34638
rect 38220 34190 38222 34242
rect 38274 34190 38276 34242
rect 38220 34178 38276 34190
rect 37548 34130 38164 34132
rect 37548 34078 37550 34130
rect 37602 34078 38164 34130
rect 37548 34076 38164 34078
rect 37548 33460 37604 34076
rect 37772 33908 37828 33918
rect 37660 33460 37716 33470
rect 37548 33458 37716 33460
rect 37548 33406 37662 33458
rect 37714 33406 37716 33458
rect 37548 33404 37716 33406
rect 37660 33394 37716 33404
rect 37100 33124 37156 33134
rect 36764 32452 36820 32462
rect 37100 32452 37156 33068
rect 37772 33124 37828 33852
rect 38556 33570 38612 34750
rect 39228 34804 39284 34862
rect 39452 34916 39508 34926
rect 39452 34822 39508 34860
rect 39228 34738 39284 34748
rect 38780 34692 38836 34702
rect 38780 34598 38836 34636
rect 38556 33518 38558 33570
rect 38610 33518 38612 33570
rect 38556 33506 38612 33518
rect 39004 33684 39060 33694
rect 38892 33348 38948 33358
rect 38668 33346 38948 33348
rect 38668 33294 38894 33346
rect 38946 33294 38948 33346
rect 38668 33292 38948 33294
rect 37996 33124 38052 33134
rect 37772 33122 38052 33124
rect 37772 33070 37998 33122
rect 38050 33070 38052 33122
rect 37772 33068 38052 33070
rect 36764 32450 37156 32452
rect 36764 32398 36766 32450
rect 36818 32398 37156 32450
rect 36764 32396 37156 32398
rect 37212 32452 37268 32462
rect 36764 32116 36820 32396
rect 37212 32358 37268 32396
rect 36764 32050 36820 32060
rect 36652 31836 36820 31892
rect 36652 31220 36708 31230
rect 36652 31106 36708 31164
rect 36652 31054 36654 31106
rect 36706 31054 36708 31106
rect 36652 31042 36708 31054
rect 36764 30996 36820 31836
rect 36764 30930 36820 30940
rect 36876 31780 36932 31790
rect 36540 30772 36596 30782
rect 36540 30678 36596 30716
rect 36428 30492 36708 30548
rect 35868 30210 36260 30212
rect 35868 30158 35870 30210
rect 35922 30158 36260 30210
rect 35868 30156 36260 30158
rect 35868 30146 35924 30156
rect 35420 30098 35588 30100
rect 35420 30046 35422 30098
rect 35474 30046 35588 30098
rect 35420 30044 35588 30046
rect 35420 30034 35476 30044
rect 36092 29986 36148 29998
rect 36092 29934 36094 29986
rect 36146 29934 36148 29986
rect 35084 29486 35086 29538
rect 35138 29486 35140 29538
rect 35084 28868 35140 29486
rect 35420 29876 35476 29886
rect 35420 29540 35476 29820
rect 36092 29876 36148 29934
rect 36204 29876 36260 30156
rect 36316 30098 36372 30156
rect 36316 30046 36318 30098
rect 36370 30046 36372 30098
rect 36316 30034 36372 30046
rect 36428 30098 36484 30110
rect 36428 30046 36430 30098
rect 36482 30046 36484 30098
rect 36428 29876 36484 30046
rect 36204 29820 36428 29876
rect 36092 29810 36148 29820
rect 36428 29810 36484 29820
rect 35644 29764 35700 29774
rect 35420 29538 35588 29540
rect 35420 29486 35422 29538
rect 35474 29486 35588 29538
rect 35420 29484 35588 29486
rect 35420 29474 35476 29484
rect 35196 29428 35252 29438
rect 35196 29334 35252 29372
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35084 28812 35252 28868
rect 34748 28756 34804 28766
rect 34636 28754 34804 28756
rect 34636 28702 34750 28754
rect 34802 28702 34804 28754
rect 34636 28700 34804 28702
rect 34748 28690 34804 28700
rect 34860 28756 34916 28766
rect 34860 28530 34916 28700
rect 35196 28642 35252 28812
rect 35196 28590 35198 28642
rect 35250 28590 35252 28642
rect 35196 28578 35252 28590
rect 35532 28644 35588 29484
rect 35644 29538 35700 29708
rect 36652 29764 36708 30492
rect 36652 29698 36708 29708
rect 35644 29486 35646 29538
rect 35698 29486 35700 29538
rect 35644 29474 35700 29486
rect 35980 29596 36484 29652
rect 35756 29092 35812 29102
rect 35644 28756 35700 28766
rect 35756 28756 35812 29036
rect 35980 28980 36036 29596
rect 36428 29540 36484 29596
rect 36540 29540 36596 29550
rect 36428 29538 36596 29540
rect 36428 29486 36542 29538
rect 36594 29486 36596 29538
rect 36428 29484 36596 29486
rect 36540 29474 36596 29484
rect 36316 29428 36372 29438
rect 36316 29334 36372 29372
rect 36652 29426 36708 29438
rect 36652 29374 36654 29426
rect 36706 29374 36708 29426
rect 36428 29316 36484 29326
rect 36428 29222 36484 29260
rect 36652 29092 36708 29374
rect 36876 29316 36932 31724
rect 36988 31444 37044 31454
rect 36988 30548 37044 31388
rect 36988 30482 37044 30492
rect 37100 31220 37156 31230
rect 37100 30434 37156 31164
rect 37212 30884 37268 30894
rect 37660 30884 37716 30894
rect 37268 30828 37380 30884
rect 37212 30790 37268 30828
rect 37100 30382 37102 30434
rect 37154 30382 37156 30434
rect 37100 30370 37156 30382
rect 37212 30324 37268 30334
rect 37212 30230 37268 30268
rect 36988 29428 37044 29438
rect 37212 29428 37268 29438
rect 36988 29426 37268 29428
rect 36988 29374 36990 29426
rect 37042 29374 37214 29426
rect 37266 29374 37268 29426
rect 36988 29372 37268 29374
rect 36988 29362 37044 29372
rect 37212 29362 37268 29372
rect 36876 29250 36932 29260
rect 37324 29204 37380 30828
rect 37436 30882 37716 30884
rect 37436 30830 37662 30882
rect 37714 30830 37716 30882
rect 37436 30828 37716 30830
rect 37436 30210 37492 30828
rect 37660 30818 37716 30828
rect 37772 30660 37828 33068
rect 37996 33058 38052 33068
rect 38332 32452 38388 32462
rect 38108 31666 38164 31678
rect 38108 31614 38110 31666
rect 38162 31614 38164 31666
rect 38108 31220 38164 31614
rect 38108 31154 38164 31164
rect 38108 30996 38164 31006
rect 37660 30604 37828 30660
rect 37884 30772 37940 30782
rect 37436 30158 37438 30210
rect 37490 30158 37492 30210
rect 37436 30100 37492 30158
rect 37436 30034 37492 30044
rect 37548 30548 37604 30558
rect 37548 29764 37604 30492
rect 37436 29652 37492 29662
rect 37548 29652 37604 29708
rect 37436 29650 37604 29652
rect 37436 29598 37438 29650
rect 37490 29598 37604 29650
rect 37436 29596 37604 29598
rect 37436 29586 37492 29596
rect 36652 29026 36708 29036
rect 37100 29148 37380 29204
rect 37548 29428 37604 29438
rect 35980 28914 36036 28924
rect 36428 28980 36484 28990
rect 35644 28754 35812 28756
rect 35644 28702 35646 28754
rect 35698 28702 35812 28754
rect 35644 28700 35812 28702
rect 36428 28756 36484 28924
rect 35644 28690 35700 28700
rect 36428 28690 36484 28700
rect 36764 28756 36820 28766
rect 35868 28644 35924 28654
rect 35532 28550 35588 28588
rect 35756 28642 35924 28644
rect 35756 28590 35870 28642
rect 35922 28590 35924 28642
rect 35756 28588 35924 28590
rect 34860 28478 34862 28530
rect 34914 28478 34916 28530
rect 34860 28466 34916 28478
rect 35084 28532 35140 28542
rect 35084 28438 35140 28476
rect 35756 28532 35812 28588
rect 35868 28578 35924 28588
rect 36316 28644 36372 28654
rect 35756 28466 35812 28476
rect 36204 28532 36260 28542
rect 36204 28438 36260 28476
rect 36316 28530 36372 28588
rect 36540 28644 36596 28654
rect 36540 28550 36596 28588
rect 36316 28478 36318 28530
rect 36370 28478 36372 28530
rect 36316 28466 36372 28478
rect 35868 28420 35924 28430
rect 35868 27970 35924 28364
rect 35868 27918 35870 27970
rect 35922 27918 35924 27970
rect 35868 27906 35924 27918
rect 36652 28420 36708 28430
rect 36092 27858 36148 27870
rect 36316 27860 36372 27870
rect 36092 27806 36094 27858
rect 36146 27806 36148 27858
rect 34748 27746 34804 27758
rect 35196 27748 35252 27758
rect 34748 27694 34750 27746
rect 34802 27694 34804 27746
rect 34748 27524 34804 27694
rect 34748 27188 34804 27468
rect 35084 27746 35252 27748
rect 35084 27694 35198 27746
rect 35250 27694 35252 27746
rect 35084 27692 35252 27694
rect 35084 27300 35140 27692
rect 35196 27682 35252 27692
rect 35980 27748 36036 27758
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35308 27300 35364 27310
rect 35084 27244 35308 27300
rect 34748 27122 34804 27132
rect 35308 27186 35364 27244
rect 35308 27134 35310 27186
rect 35362 27134 35364 27186
rect 35308 27122 35364 27134
rect 35756 27076 35812 27086
rect 34748 26964 34804 27002
rect 34748 26898 34804 26908
rect 34636 26850 34692 26862
rect 34636 26798 34638 26850
rect 34690 26798 34692 26850
rect 34636 26516 34692 26798
rect 34636 26450 34692 26460
rect 35532 26516 35588 26526
rect 35532 26290 35588 26460
rect 35532 26238 35534 26290
rect 35586 26238 35588 26290
rect 35084 26178 35140 26190
rect 35084 26126 35086 26178
rect 35138 26126 35140 26178
rect 35084 26068 35140 26126
rect 35084 26002 35140 26012
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35420 25508 35476 25518
rect 35084 25506 35476 25508
rect 35084 25454 35422 25506
rect 35474 25454 35476 25506
rect 35084 25452 35476 25454
rect 34748 25284 34804 25294
rect 35084 25284 35140 25452
rect 35420 25442 35476 25452
rect 34748 25282 35140 25284
rect 34748 25230 34750 25282
rect 34802 25230 35140 25282
rect 34748 25228 35140 25230
rect 34748 25218 34804 25228
rect 34636 25172 34692 25182
rect 34636 24836 34692 25116
rect 35084 24948 35140 25228
rect 35196 25284 35252 25294
rect 35532 25284 35588 26238
rect 35756 26402 35812 27020
rect 35756 26350 35758 26402
rect 35810 26350 35812 26402
rect 35756 25732 35812 26350
rect 35980 26962 36036 27692
rect 35980 26910 35982 26962
rect 36034 26910 36036 26962
rect 35980 26068 36036 26910
rect 36092 26516 36148 27806
rect 36204 27858 36372 27860
rect 36204 27806 36318 27858
rect 36370 27806 36372 27858
rect 36204 27804 36372 27806
rect 36204 27074 36260 27804
rect 36316 27794 36372 27804
rect 36316 27300 36372 27310
rect 36316 27186 36372 27244
rect 36316 27134 36318 27186
rect 36370 27134 36372 27186
rect 36316 27122 36372 27134
rect 36204 27022 36206 27074
rect 36258 27022 36260 27074
rect 36204 26908 36260 27022
rect 36428 27076 36484 27114
rect 36484 27020 36596 27076
rect 36428 27010 36484 27020
rect 36204 26852 36484 26908
rect 36428 26786 36484 26796
rect 36204 26516 36260 26526
rect 36092 26514 36260 26516
rect 36092 26462 36206 26514
rect 36258 26462 36260 26514
rect 36092 26460 36260 26462
rect 36204 26450 36260 26460
rect 36428 26516 36484 26526
rect 36428 26422 36484 26460
rect 36540 26402 36596 27020
rect 36540 26350 36542 26402
rect 36594 26350 36596 26402
rect 36540 26338 36596 26350
rect 35980 26002 36036 26012
rect 35756 25666 35812 25676
rect 35196 25282 35588 25284
rect 35196 25230 35198 25282
rect 35250 25230 35588 25282
rect 35196 25228 35588 25230
rect 35196 25218 35252 25228
rect 34748 24836 34804 24846
rect 34636 24780 34748 24836
rect 34748 24742 34804 24780
rect 35084 23938 35140 24892
rect 36092 24948 36148 24958
rect 36092 24854 36148 24892
rect 35420 24836 35476 24846
rect 35476 24780 35588 24836
rect 35420 24742 35476 24780
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35084 23886 35086 23938
rect 35138 23886 35140 23938
rect 35084 23874 35140 23886
rect 35532 23938 35588 24780
rect 35756 24834 35812 24846
rect 35756 24782 35758 24834
rect 35810 24782 35812 24834
rect 35756 24724 35812 24782
rect 36428 24836 36484 24846
rect 36428 24742 36484 24780
rect 35812 24668 35924 24724
rect 35756 24658 35812 24668
rect 35532 23886 35534 23938
rect 35586 23886 35588 23938
rect 35532 23874 35588 23886
rect 34748 23716 34804 23726
rect 35756 23716 35812 23726
rect 34524 23492 34692 23548
rect 34636 23380 34692 23492
rect 34748 23492 34804 23660
rect 35644 23714 35812 23716
rect 35644 23662 35758 23714
rect 35810 23662 35812 23714
rect 35644 23660 35812 23662
rect 34748 23436 35140 23492
rect 34636 23324 34804 23380
rect 34636 23156 34692 23166
rect 34636 23062 34692 23100
rect 34524 23044 34580 23054
rect 34412 22932 34468 22942
rect 34412 22838 34468 22876
rect 34524 22930 34580 22988
rect 34524 22878 34526 22930
rect 34578 22878 34580 22930
rect 34524 22866 34580 22878
rect 34748 22820 34804 23324
rect 34972 23044 35028 23054
rect 34972 22950 35028 22988
rect 35084 22820 35140 23436
rect 35196 23268 35252 23278
rect 35196 22932 35252 23212
rect 35532 22932 35588 22942
rect 35196 22930 35588 22932
rect 35196 22878 35198 22930
rect 35250 22878 35534 22930
rect 35586 22878 35588 22930
rect 35196 22876 35588 22878
rect 35196 22866 35252 22876
rect 35532 22866 35588 22876
rect 34636 22764 34804 22820
rect 34972 22764 35140 22820
rect 35196 22764 35460 22774
rect 34524 22708 34580 22718
rect 34412 22484 34468 22494
rect 34300 22482 34468 22484
rect 34300 22430 34414 22482
rect 34466 22430 34468 22482
rect 34300 22428 34468 22430
rect 34412 22418 34468 22428
rect 34524 22370 34580 22652
rect 34524 22318 34526 22370
rect 34578 22318 34580 22370
rect 34524 22306 34580 22318
rect 34300 22260 34356 22270
rect 34300 22146 34356 22204
rect 34300 22094 34302 22146
rect 34354 22094 34356 22146
rect 34300 21924 34356 22094
rect 34412 21924 34468 21934
rect 34300 21868 34412 21924
rect 34412 21810 34468 21868
rect 34412 21758 34414 21810
rect 34466 21758 34468 21810
rect 34412 21746 34468 21758
rect 34300 21700 34356 21710
rect 34300 18004 34356 21644
rect 34412 21252 34468 21262
rect 34468 21196 34580 21252
rect 34412 21186 34468 21196
rect 34300 17444 34356 17948
rect 34300 17378 34356 17388
rect 34412 20804 34468 20814
rect 33852 17164 34244 17220
rect 33852 16100 33908 17164
rect 34412 17108 34468 20748
rect 34524 17332 34580 21196
rect 34524 17266 34580 17276
rect 34412 16882 34468 17052
rect 34412 16830 34414 16882
rect 34466 16830 34468 16882
rect 34412 16818 34468 16830
rect 33852 15986 33908 16044
rect 33852 15934 33854 15986
rect 33906 15934 33908 15986
rect 33852 15652 33908 15934
rect 33852 15586 33908 15596
rect 33964 16772 34020 16782
rect 33516 15262 33518 15314
rect 33570 15262 33572 15314
rect 33516 15250 33572 15262
rect 33628 15484 33796 15540
rect 33292 14252 33460 14308
rect 33516 15092 33572 15102
rect 33292 13860 33348 14252
rect 33404 13972 33460 13982
rect 33516 13972 33572 15036
rect 33404 13970 33572 13972
rect 33404 13918 33406 13970
rect 33458 13918 33572 13970
rect 33404 13916 33572 13918
rect 33404 13906 33460 13916
rect 33292 13766 33348 13804
rect 33404 13524 33460 13534
rect 33180 13522 33460 13524
rect 33180 13470 33406 13522
rect 33458 13470 33460 13522
rect 33180 13468 33460 13470
rect 33404 13458 33460 13468
rect 33180 12852 33236 12862
rect 32844 12850 33236 12852
rect 32844 12798 33182 12850
rect 33234 12798 33236 12850
rect 32844 12796 33236 12798
rect 33180 12786 33236 12796
rect 33404 12852 33460 12862
rect 33404 12758 33460 12796
rect 33292 12738 33348 12750
rect 33292 12686 33294 12738
rect 33346 12686 33348 12738
rect 33180 12404 33236 12414
rect 33180 12310 33236 12348
rect 33292 12290 33348 12686
rect 33292 12238 33294 12290
rect 33346 12238 33348 12290
rect 33292 12226 33348 12238
rect 33404 12628 33460 12638
rect 32956 12178 33012 12190
rect 32956 12126 32958 12178
rect 33010 12126 33012 12178
rect 32844 11396 32900 11406
rect 32956 11396 33012 12126
rect 32844 11394 33012 11396
rect 32844 11342 32846 11394
rect 32898 11342 33012 11394
rect 32844 11340 33012 11342
rect 32844 11330 32900 11340
rect 32172 8370 32340 8372
rect 32172 8318 32174 8370
rect 32226 8318 32340 8370
rect 32172 8316 32340 8318
rect 32508 9996 32788 10052
rect 33068 11170 33124 11182
rect 33068 11118 33070 11170
rect 33122 11118 33124 11170
rect 33068 10052 33124 11118
rect 33180 10612 33236 10622
rect 33180 10518 33236 10556
rect 32172 8306 32228 8316
rect 31500 3442 31668 3444
rect 31500 3390 31502 3442
rect 31554 3390 31668 3442
rect 31500 3388 31668 3390
rect 31948 4228 32004 4238
rect 31948 4226 32228 4228
rect 31948 4174 31950 4226
rect 32002 4174 32228 4226
rect 31948 4172 32228 4174
rect 31948 3388 32004 4172
rect 32172 3554 32228 4172
rect 32172 3502 32174 3554
rect 32226 3502 32228 3554
rect 32172 3490 32228 3502
rect 31500 3378 31556 3388
rect 31724 3332 32004 3388
rect 32508 3442 32564 9996
rect 33068 9986 33124 9996
rect 32620 9826 32676 9838
rect 32620 9774 32622 9826
rect 32674 9774 32676 9826
rect 32620 9604 32676 9774
rect 33068 9604 33124 9614
rect 32620 9602 33236 9604
rect 32620 9550 33070 9602
rect 33122 9550 33236 9602
rect 32620 9548 33236 9550
rect 33068 9538 33124 9548
rect 33180 8260 33236 9548
rect 33180 7700 33236 8204
rect 33180 7474 33236 7644
rect 33180 7422 33182 7474
rect 33234 7422 33236 7474
rect 33180 7410 33236 7422
rect 33404 7252 33460 12572
rect 33628 11620 33684 15484
rect 33852 15204 33908 15214
rect 33964 15204 34020 16716
rect 33908 15148 34020 15204
rect 34076 15874 34132 15886
rect 34076 15822 34078 15874
rect 34130 15822 34132 15874
rect 33852 15138 33908 15148
rect 33740 15090 33796 15102
rect 33740 15038 33742 15090
rect 33794 15038 33796 15090
rect 33740 14756 33796 15038
rect 34076 14980 34132 15822
rect 34188 15874 34244 15886
rect 34188 15822 34190 15874
rect 34242 15822 34244 15874
rect 34188 15316 34244 15822
rect 34300 15876 34356 15886
rect 34636 15876 34692 22764
rect 34748 22596 34804 22606
rect 34748 22258 34804 22540
rect 34748 22206 34750 22258
rect 34802 22206 34804 22258
rect 34748 22194 34804 22206
rect 34860 22148 34916 22158
rect 34860 22036 34916 22092
rect 34748 21980 34916 22036
rect 34748 20802 34804 21980
rect 34860 21812 34916 21822
rect 34860 21718 34916 21756
rect 34748 20750 34750 20802
rect 34802 20750 34804 20802
rect 34748 20580 34804 20750
rect 34748 20514 34804 20524
rect 34972 20132 35028 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35532 22148 35588 22158
rect 35644 22148 35700 23660
rect 35756 23650 35812 23660
rect 35756 23044 35812 23054
rect 35756 22260 35812 22988
rect 35868 22596 35924 24668
rect 36316 23714 36372 23726
rect 36316 23662 36318 23714
rect 36370 23662 36372 23714
rect 35868 22530 35924 22540
rect 36204 23042 36260 23054
rect 36204 22990 36206 23042
rect 36258 22990 36260 23042
rect 35756 22194 35812 22204
rect 36204 22372 36260 22990
rect 35588 22092 35700 22148
rect 35868 22146 35924 22158
rect 35868 22094 35870 22146
rect 35922 22094 35924 22146
rect 35532 22054 35588 22092
rect 35868 22036 35924 22094
rect 35868 21970 35924 21980
rect 35308 21474 35364 21486
rect 35868 21476 35924 21486
rect 35308 21422 35310 21474
rect 35362 21422 35364 21474
rect 35308 21364 35364 21422
rect 35308 21298 35364 21308
rect 35756 21420 35868 21476
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35084 20804 35140 20814
rect 35644 20804 35700 20814
rect 35756 20804 35812 21420
rect 35868 21382 35924 21420
rect 36204 21364 36260 22316
rect 36204 21298 36260 21308
rect 36316 22930 36372 23662
rect 36316 22878 36318 22930
rect 36370 22878 36372 22930
rect 36316 22146 36372 22878
rect 36316 22094 36318 22146
rect 36370 22094 36372 22146
rect 36316 21924 36372 22094
rect 35084 20802 35812 20804
rect 35084 20750 35086 20802
rect 35138 20750 35646 20802
rect 35698 20750 35812 20802
rect 35084 20748 35812 20750
rect 35084 20738 35140 20748
rect 35644 20738 35700 20748
rect 35196 20580 35252 20590
rect 35196 20486 35252 20524
rect 35308 20578 35364 20590
rect 35308 20526 35310 20578
rect 35362 20526 35364 20578
rect 35308 20244 35364 20526
rect 35308 20178 35364 20188
rect 34972 20038 35028 20076
rect 34860 20020 34916 20030
rect 34860 19926 34916 19964
rect 34972 19796 35028 19806
rect 34972 19794 35140 19796
rect 34972 19742 34974 19794
rect 35026 19742 35140 19794
rect 34972 19740 35140 19742
rect 34972 19730 35028 19740
rect 35084 19460 35140 19740
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35084 19404 35364 19460
rect 35308 19346 35364 19404
rect 35308 19294 35310 19346
rect 35362 19294 35364 19346
rect 35308 19282 35364 19294
rect 35756 19234 35812 20748
rect 35868 20804 35924 20814
rect 36092 20804 36148 20814
rect 35868 20802 36036 20804
rect 35868 20750 35870 20802
rect 35922 20750 36036 20802
rect 35868 20748 36036 20750
rect 35868 20738 35924 20748
rect 35868 20580 35924 20590
rect 35868 20018 35924 20524
rect 35868 19966 35870 20018
rect 35922 19966 35924 20018
rect 35868 19954 35924 19966
rect 35980 20020 36036 20748
rect 36092 20244 36148 20748
rect 36316 20244 36372 21868
rect 36540 20578 36596 20590
rect 36540 20526 36542 20578
rect 36594 20526 36596 20578
rect 36540 20468 36596 20526
rect 36540 20402 36596 20412
rect 36316 20188 36596 20244
rect 36092 20178 36148 20188
rect 36316 20020 36372 20030
rect 35980 19964 36316 20020
rect 36316 19926 36372 19964
rect 35756 19182 35758 19234
rect 35810 19182 35812 19234
rect 35756 19170 35812 19182
rect 35868 19348 35924 19358
rect 35756 19012 35812 19022
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 34748 17444 34804 17454
rect 34748 17350 34804 17388
rect 35084 17442 35140 17454
rect 35084 17390 35086 17442
rect 35138 17390 35140 17442
rect 34972 17332 35028 17342
rect 34860 16772 34916 16782
rect 34748 16100 34804 16110
rect 34748 16006 34804 16044
rect 34636 15820 34804 15876
rect 34300 15782 34356 15820
rect 34524 15316 34580 15326
rect 34188 15314 34580 15316
rect 34188 15262 34526 15314
rect 34578 15262 34580 15314
rect 34188 15260 34580 15262
rect 34524 15250 34580 15260
rect 34188 15092 34244 15102
rect 34188 14998 34244 15036
rect 34076 14914 34132 14924
rect 34300 14756 34356 14766
rect 34748 14756 34804 15820
rect 33740 14754 34356 14756
rect 33740 14702 34302 14754
rect 34354 14702 34356 14754
rect 33740 14700 34356 14702
rect 34300 14690 34356 14700
rect 34636 14700 34804 14756
rect 34076 14532 34132 14542
rect 34076 13748 34132 14476
rect 34076 13654 34132 13692
rect 34524 13860 34580 13870
rect 34524 13746 34580 13804
rect 34524 13694 34526 13746
rect 34578 13694 34580 13746
rect 34524 13682 34580 13694
rect 34300 13524 34356 13534
rect 34188 13522 34356 13524
rect 34188 13470 34302 13522
rect 34354 13470 34356 13522
rect 34188 13468 34356 13470
rect 33852 12962 33908 12974
rect 33852 12910 33854 12962
rect 33906 12910 33908 12962
rect 33852 12402 33908 12910
rect 33852 12350 33854 12402
rect 33906 12350 33908 12402
rect 33852 12338 33908 12350
rect 33964 12292 34020 12302
rect 33964 12198 34020 12236
rect 33516 11564 33684 11620
rect 33740 12178 33796 12190
rect 33740 12126 33742 12178
rect 33794 12126 33796 12178
rect 33516 11172 33572 11564
rect 33628 11396 33684 11406
rect 33628 11302 33684 11340
rect 33516 11116 33684 11172
rect 33180 7196 33460 7252
rect 32620 4228 32676 4238
rect 32620 4226 32900 4228
rect 32620 4174 32622 4226
rect 32674 4174 32900 4226
rect 32620 4172 32900 4174
rect 32620 4162 32676 4172
rect 32508 3390 32510 3442
rect 32562 3390 32564 3442
rect 32508 3378 32564 3390
rect 32844 3554 32900 4172
rect 32844 3502 32846 3554
rect 32898 3502 32900 3554
rect 31724 1764 31780 3332
rect 32844 2548 32900 3502
rect 31612 1708 31780 1764
rect 32284 2492 32900 2548
rect 32956 3556 33012 3566
rect 31612 800 31668 1708
rect 32284 800 32340 2492
rect 32956 800 33012 3500
rect 33180 3442 33236 7196
rect 33628 7140 33684 11116
rect 33740 10836 33796 12126
rect 34188 12068 34244 13468
rect 34300 13458 34356 13468
rect 34300 12740 34356 12750
rect 34300 12646 34356 12684
rect 34636 12516 34692 14700
rect 34748 14530 34804 14542
rect 34748 14478 34750 14530
rect 34802 14478 34804 14530
rect 34748 13524 34804 14478
rect 34748 13458 34804 13468
rect 34188 12002 34244 12012
rect 34300 12460 34692 12516
rect 34076 11844 34132 11854
rect 34076 11394 34132 11788
rect 34300 11788 34356 12460
rect 34748 12404 34804 12414
rect 34412 12402 34804 12404
rect 34412 12350 34750 12402
rect 34802 12350 34804 12402
rect 34412 12348 34804 12350
rect 34412 12178 34468 12348
rect 34748 12338 34804 12348
rect 34412 12126 34414 12178
rect 34466 12126 34468 12178
rect 34412 12114 34468 12126
rect 34524 12178 34580 12190
rect 34524 12126 34526 12178
rect 34578 12126 34580 12178
rect 34524 11844 34580 12126
rect 34300 11732 34468 11788
rect 34524 11778 34580 11788
rect 34636 12180 34692 12190
rect 34300 11508 34356 11518
rect 34300 11414 34356 11452
rect 34076 11342 34078 11394
rect 34130 11342 34132 11394
rect 34076 10836 34132 11342
rect 33740 10834 34132 10836
rect 33740 10782 33742 10834
rect 33794 10782 34132 10834
rect 33740 10780 34132 10782
rect 33740 10770 33796 10780
rect 34412 10724 34468 11732
rect 34636 11620 34692 12124
rect 34524 11564 34692 11620
rect 34748 12068 34804 12078
rect 34524 11394 34580 11564
rect 34524 11342 34526 11394
rect 34578 11342 34580 11394
rect 34524 11330 34580 11342
rect 34636 11394 34692 11406
rect 34636 11342 34638 11394
rect 34690 11342 34692 11394
rect 34636 10834 34692 11342
rect 34636 10782 34638 10834
rect 34690 10782 34692 10834
rect 34636 10770 34692 10782
rect 34524 10724 34580 10734
rect 34412 10722 34580 10724
rect 34412 10670 34526 10722
rect 34578 10670 34580 10722
rect 34412 10668 34580 10670
rect 34524 10612 34580 10668
rect 33852 10500 33908 10510
rect 33852 10498 34132 10500
rect 33852 10446 33854 10498
rect 33906 10446 34132 10498
rect 33852 10444 34132 10446
rect 33852 10434 33908 10444
rect 34076 10388 34132 10444
rect 33740 9380 33796 9390
rect 33740 9268 33796 9324
rect 33740 9266 34020 9268
rect 33740 9214 33742 9266
rect 33794 9214 34020 9266
rect 33740 9212 34020 9214
rect 33740 9202 33796 9212
rect 33964 9154 34020 9212
rect 33964 9102 33966 9154
rect 34018 9102 34020 9154
rect 33964 8484 34020 9102
rect 33964 8418 34020 8428
rect 34076 8260 34132 10332
rect 34188 9940 34244 9950
rect 34524 9940 34580 10556
rect 34748 10388 34804 12012
rect 34860 11396 34916 16716
rect 34972 15988 35028 17276
rect 35084 16212 35140 17390
rect 35196 16884 35252 16894
rect 35196 16882 35700 16884
rect 35196 16830 35198 16882
rect 35250 16830 35700 16882
rect 35196 16828 35700 16830
rect 35196 16818 35252 16828
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35084 16156 35588 16212
rect 35532 16100 35588 16156
rect 35644 16210 35700 16828
rect 35644 16158 35646 16210
rect 35698 16158 35700 16210
rect 35644 16146 35700 16158
rect 35756 16436 35812 18956
rect 35868 18676 35924 19292
rect 36204 19122 36260 19134
rect 36204 19070 36206 19122
rect 36258 19070 36260 19122
rect 36204 18788 36260 19070
rect 36204 18722 36260 18732
rect 35868 18610 35924 18620
rect 36428 18676 36484 18686
rect 36428 18450 36484 18620
rect 36428 18398 36430 18450
rect 36482 18398 36484 18450
rect 36428 18228 36484 18398
rect 36428 18162 36484 18172
rect 36428 17442 36484 17454
rect 36428 17390 36430 17442
rect 36482 17390 36484 17442
rect 36428 17332 36484 17390
rect 36428 17266 36484 17276
rect 35532 16006 35588 16044
rect 35756 16098 35812 16380
rect 35756 16046 35758 16098
rect 35810 16046 35812 16098
rect 35756 16034 35812 16046
rect 35196 15988 35252 15998
rect 34972 15986 35252 15988
rect 34972 15934 35198 15986
rect 35250 15934 35252 15986
rect 34972 15932 35252 15934
rect 35196 15540 35252 15932
rect 35196 15474 35252 15484
rect 35644 15988 35700 15998
rect 34972 15316 35028 15326
rect 34972 15314 35140 15316
rect 34972 15262 34974 15314
rect 35026 15262 35140 15314
rect 34972 15260 35140 15262
rect 34972 15250 35028 15260
rect 34972 14532 35028 14570
rect 34972 14466 35028 14476
rect 35084 14532 35140 15260
rect 35420 15204 35476 15242
rect 35420 15138 35476 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 14532 35252 14542
rect 35084 14530 35252 14532
rect 35084 14478 35198 14530
rect 35250 14478 35252 14530
rect 35084 14476 35252 14478
rect 34972 14308 35028 14318
rect 34972 13970 35028 14252
rect 34972 13918 34974 13970
rect 35026 13918 35028 13970
rect 34972 13906 35028 13918
rect 34972 12292 35028 12302
rect 34972 12198 35028 12236
rect 34972 12068 35028 12078
rect 35084 12068 35140 14476
rect 35196 14466 35252 14476
rect 35420 14418 35476 14430
rect 35420 14366 35422 14418
rect 35474 14366 35476 14418
rect 35420 13748 35476 14366
rect 35644 14308 35700 15932
rect 35980 15876 36036 15886
rect 35980 15782 36036 15820
rect 35980 15540 36036 15550
rect 35980 15446 36036 15484
rect 35868 15314 35924 15326
rect 35868 15262 35870 15314
rect 35922 15262 35924 15314
rect 35756 15204 35812 15214
rect 35756 14530 35812 15148
rect 35868 14868 35924 15262
rect 35868 14802 35924 14812
rect 36204 15314 36260 15326
rect 36204 15262 36206 15314
rect 36258 15262 36260 15314
rect 35756 14478 35758 14530
rect 35810 14478 35812 14530
rect 35756 14466 35812 14478
rect 36092 14756 36148 14766
rect 35868 14308 35924 14318
rect 35644 14306 35924 14308
rect 35644 14254 35870 14306
rect 35922 14254 35924 14306
rect 35644 14252 35924 14254
rect 35868 14242 35924 14252
rect 35980 14306 36036 14318
rect 35980 14254 35982 14306
rect 36034 14254 36036 14306
rect 35980 14196 36036 14254
rect 35980 14130 36036 14140
rect 35420 13524 35476 13692
rect 35420 13468 35700 13524
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 12740 35252 12750
rect 35196 12290 35252 12684
rect 35196 12238 35198 12290
rect 35250 12238 35252 12290
rect 35196 12226 35252 12238
rect 35028 12012 35140 12068
rect 34972 12002 35028 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 11508 35252 11518
rect 35196 11414 35252 11452
rect 34860 11330 34916 11340
rect 35420 11394 35476 11406
rect 35420 11342 35422 11394
rect 35474 11342 35476 11394
rect 35420 10724 35476 11342
rect 35420 10658 35476 10668
rect 34860 10610 34916 10622
rect 34860 10558 34862 10610
rect 34914 10558 34916 10610
rect 34860 10500 34916 10558
rect 34860 10444 35140 10500
rect 35084 10388 35140 10444
rect 35532 10388 35588 10398
rect 34748 10332 35028 10388
rect 34636 9940 34692 9950
rect 34860 9940 34916 9950
rect 34188 9938 34916 9940
rect 34188 9886 34190 9938
rect 34242 9886 34638 9938
rect 34690 9886 34862 9938
rect 34914 9886 34916 9938
rect 34188 9884 34916 9886
rect 34188 9874 34244 9884
rect 34636 9874 34692 9884
rect 34860 9874 34916 9884
rect 34524 9716 34580 9726
rect 34972 9716 35028 10332
rect 34524 9268 34580 9660
rect 34300 9266 34580 9268
rect 34300 9214 34526 9266
rect 34578 9214 34580 9266
rect 34300 9212 34580 9214
rect 34300 8370 34356 9212
rect 34524 9202 34580 9212
rect 34860 9660 35028 9716
rect 35084 10386 35588 10388
rect 35084 10334 35534 10386
rect 35586 10334 35588 10386
rect 35084 10332 35588 10334
rect 34860 9044 34916 9660
rect 35084 9492 35140 10332
rect 35532 10322 35588 10332
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35644 10052 35700 13468
rect 36092 11506 36148 14700
rect 36204 14418 36260 15262
rect 36204 14366 36206 14418
rect 36258 14366 36260 14418
rect 36204 14354 36260 14366
rect 36316 14868 36372 14878
rect 36204 13746 36260 13758
rect 36204 13694 36206 13746
rect 36258 13694 36260 13746
rect 36204 13524 36260 13694
rect 36204 13458 36260 13468
rect 36316 13300 36372 14812
rect 36092 11454 36094 11506
rect 36146 11454 36148 11506
rect 36092 11442 36148 11454
rect 36204 13244 36372 13300
rect 36204 12178 36260 13244
rect 36204 12126 36206 12178
rect 36258 12126 36260 12178
rect 35868 10948 35924 10958
rect 35756 10612 35812 10622
rect 35756 10518 35812 10556
rect 35868 10052 35924 10892
rect 36204 10836 36260 12126
rect 36540 11788 36596 20188
rect 36652 19012 36708 28364
rect 36764 23156 36820 28700
rect 36876 26964 36932 27002
rect 36876 26898 36932 26908
rect 36988 24388 37044 24398
rect 36988 23826 37044 24332
rect 36988 23774 36990 23826
rect 37042 23774 37044 23826
rect 36988 23604 37044 23774
rect 36988 23538 37044 23548
rect 36876 23156 36932 23166
rect 36764 23154 36932 23156
rect 36764 23102 36878 23154
rect 36930 23102 36932 23154
rect 36764 23100 36932 23102
rect 37100 23156 37156 29148
rect 37324 28980 37380 28990
rect 37380 28924 37492 28980
rect 37324 28914 37380 28924
rect 37212 28866 37268 28878
rect 37212 28814 37214 28866
rect 37266 28814 37268 28866
rect 37212 28754 37268 28814
rect 37212 28702 37214 28754
rect 37266 28702 37268 28754
rect 37212 28690 37268 28702
rect 37436 28756 37492 28924
rect 37436 28420 37492 28700
rect 37548 28644 37604 29372
rect 37548 28578 37604 28588
rect 37548 28420 37604 28430
rect 37436 28418 37604 28420
rect 37436 28366 37550 28418
rect 37602 28366 37604 28418
rect 37436 28364 37604 28366
rect 37548 28354 37604 28364
rect 37660 28196 37716 30604
rect 37772 30212 37828 30222
rect 37772 28866 37828 30156
rect 37884 30210 37940 30716
rect 38108 30436 38164 30940
rect 38108 30370 38164 30380
rect 37884 30158 37886 30210
rect 37938 30158 37940 30210
rect 37884 30146 37940 30158
rect 38220 30212 38276 30222
rect 38220 30118 38276 30156
rect 38108 30100 38164 30110
rect 37996 29988 38052 29998
rect 37996 29894 38052 29932
rect 38108 29876 38164 30044
rect 37884 29764 37940 29774
rect 37940 29708 38052 29764
rect 37884 29698 37940 29708
rect 37772 28814 37774 28866
rect 37826 28814 37828 28866
rect 37772 28802 37828 28814
rect 37996 28754 38052 29708
rect 38108 29538 38164 29820
rect 38108 29486 38110 29538
rect 38162 29486 38164 29538
rect 38108 29474 38164 29486
rect 37996 28702 37998 28754
rect 38050 28702 38052 28754
rect 37996 28690 38052 28702
rect 37436 28140 37716 28196
rect 37324 27746 37380 27758
rect 37324 27694 37326 27746
rect 37378 27694 37380 27746
rect 37212 27636 37268 27646
rect 37212 27076 37268 27580
rect 37324 27300 37380 27694
rect 37324 27234 37380 27244
rect 37324 27076 37380 27086
rect 37268 27074 37380 27076
rect 37268 27022 37326 27074
rect 37378 27022 37380 27074
rect 37268 27020 37380 27022
rect 37212 27010 37268 27020
rect 37324 27010 37380 27020
rect 37212 26852 37268 26862
rect 37212 26514 37268 26796
rect 37212 26462 37214 26514
rect 37266 26462 37268 26514
rect 37212 26450 37268 26462
rect 37324 23714 37380 23726
rect 37324 23662 37326 23714
rect 37378 23662 37380 23714
rect 37324 23492 37380 23662
rect 37324 23426 37380 23436
rect 37100 23100 37268 23156
rect 36876 21924 36932 23100
rect 37100 22932 37156 22942
rect 37100 22594 37156 22876
rect 37100 22542 37102 22594
rect 37154 22542 37156 22594
rect 37100 22530 37156 22542
rect 37100 22146 37156 22158
rect 37100 22094 37102 22146
rect 37154 22094 37156 22146
rect 37100 21924 37156 22094
rect 36876 21868 37156 21924
rect 36764 21476 36820 21486
rect 36764 21362 36820 21420
rect 36764 21310 36766 21362
rect 36818 21310 36820 21362
rect 36764 21298 36820 21310
rect 36764 19906 36820 19918
rect 36764 19854 36766 19906
rect 36818 19854 36820 19906
rect 36764 19236 36820 19854
rect 36764 19170 36820 19180
rect 36652 18946 36708 18956
rect 36652 18788 36708 18798
rect 36652 18674 36708 18732
rect 36652 18622 36654 18674
rect 36706 18622 36708 18674
rect 36652 18610 36708 18622
rect 36876 18676 36932 21868
rect 37212 21700 37268 23100
rect 37324 22932 37380 22942
rect 37436 22932 37492 28140
rect 37660 27858 37716 27870
rect 37660 27806 37662 27858
rect 37714 27806 37716 27858
rect 37548 27188 37604 27198
rect 37660 27188 37716 27806
rect 38220 27748 38276 27758
rect 38220 27654 38276 27692
rect 37548 27186 37716 27188
rect 37548 27134 37550 27186
rect 37602 27134 37716 27186
rect 37548 27132 37716 27134
rect 37548 27122 37604 27132
rect 37660 26852 37716 27132
rect 38108 27300 38164 27310
rect 37772 27076 37828 27086
rect 38108 27076 38164 27244
rect 38220 27076 38276 27086
rect 37828 27074 38276 27076
rect 37828 27022 38222 27074
rect 38274 27022 38276 27074
rect 37828 27020 38276 27022
rect 37772 26982 37828 27020
rect 37772 26852 37828 26862
rect 37660 26796 37772 26852
rect 37772 26786 37828 26796
rect 38108 26514 38164 27020
rect 38220 27010 38276 27020
rect 38332 26908 38388 32396
rect 38668 32116 38724 33292
rect 38892 33282 38948 33292
rect 39004 33124 39060 33628
rect 39452 33346 39508 33358
rect 39452 33294 39454 33346
rect 39506 33294 39508 33346
rect 39452 33236 39508 33294
rect 39452 33170 39508 33180
rect 38780 33068 39060 33124
rect 38780 32564 38836 33068
rect 38892 32788 38948 32798
rect 38892 32694 38948 32732
rect 39340 32788 39396 32798
rect 39340 32694 39396 32732
rect 38780 32562 39060 32564
rect 38780 32510 38782 32562
rect 38834 32510 39060 32562
rect 38780 32508 39060 32510
rect 38780 32498 38836 32508
rect 38892 32340 38948 32350
rect 38444 32060 38724 32116
rect 38780 32338 38948 32340
rect 38780 32286 38894 32338
rect 38946 32286 38948 32338
rect 38780 32284 38948 32286
rect 38444 31780 38500 32060
rect 38444 31714 38500 31724
rect 38556 31892 38612 31902
rect 38556 31778 38612 31836
rect 38556 31726 38558 31778
rect 38610 31726 38612 31778
rect 38556 31714 38612 31726
rect 38556 30884 38612 30894
rect 38556 30790 38612 30828
rect 38780 30436 38836 32284
rect 38892 32274 38948 32284
rect 39004 31890 39060 32508
rect 39004 31838 39006 31890
rect 39058 31838 39060 31890
rect 39004 31826 39060 31838
rect 39452 32450 39508 32462
rect 39452 32398 39454 32450
rect 39506 32398 39508 32450
rect 39452 32228 39508 32398
rect 39452 31892 39508 32172
rect 39452 31826 39508 31836
rect 39564 31668 39620 35084
rect 39676 35026 39732 35084
rect 39676 34974 39678 35026
rect 39730 34974 39732 35026
rect 39676 34962 39732 34974
rect 39788 34804 39844 35196
rect 39788 34738 39844 34748
rect 40012 35140 40068 35150
rect 39676 34692 39732 34702
rect 39676 33234 39732 34636
rect 39676 33182 39678 33234
rect 39730 33182 39732 33234
rect 39676 33170 39732 33182
rect 40012 33124 40068 35084
rect 40124 34916 40180 34926
rect 40124 34020 40180 34860
rect 40348 34692 40404 36206
rect 40572 36258 40628 36270
rect 40572 36206 40574 36258
rect 40626 36206 40628 36258
rect 40572 36148 40628 36206
rect 40572 36082 40628 36092
rect 40908 35700 40964 36876
rect 41244 36484 41300 39452
rect 41468 38668 41524 39564
rect 41580 39172 41636 39182
rect 41580 38836 41636 39116
rect 41804 39058 41860 42252
rect 42028 41076 42084 43260
rect 42364 42868 42420 44940
rect 42252 42812 42420 42868
rect 42140 42754 42196 42766
rect 42140 42702 42142 42754
rect 42194 42702 42196 42754
rect 42140 41298 42196 42702
rect 42252 41636 42308 42812
rect 42476 42756 42532 46956
rect 42812 45108 42868 45118
rect 42812 45014 42868 45052
rect 43036 44548 43092 47964
rect 44268 47570 44324 48188
rect 44268 47518 44270 47570
rect 44322 47518 44324 47570
rect 44268 46898 44324 47518
rect 44268 46846 44270 46898
rect 44322 46846 44324 46898
rect 44268 46834 44324 46846
rect 44380 46562 44436 46574
rect 44380 46510 44382 46562
rect 44434 46510 44436 46562
rect 43708 46452 43764 46462
rect 43708 45892 43764 46396
rect 44380 46340 44436 46510
rect 44380 46274 44436 46284
rect 44492 46450 44548 48860
rect 44492 46398 44494 46450
rect 44546 46398 44548 46450
rect 43708 45798 43764 45836
rect 43372 45668 43428 45678
rect 43148 45108 43204 45118
rect 43148 45014 43204 45052
rect 43260 44996 43316 45006
rect 43260 44902 43316 44940
rect 42588 44492 43316 44548
rect 42588 43538 42644 44492
rect 43260 44436 43316 44492
rect 42924 44324 42980 44334
rect 42588 43486 42590 43538
rect 42642 43486 42644 43538
rect 42588 43474 42644 43486
rect 42700 44322 42980 44324
rect 42700 44270 42926 44322
rect 42978 44270 42980 44322
rect 42700 44268 42980 44270
rect 42476 42690 42532 42700
rect 42588 42756 42644 42766
rect 42700 42756 42756 44268
rect 42924 44258 42980 44268
rect 43036 44324 43092 44334
rect 43036 44230 43092 44268
rect 43260 44210 43316 44380
rect 43260 44158 43262 44210
rect 43314 44158 43316 44210
rect 43260 44146 43316 44158
rect 42812 44100 42868 44110
rect 42812 43538 42868 44044
rect 43372 43876 43428 45612
rect 43484 45666 43540 45678
rect 43484 45614 43486 45666
rect 43538 45614 43540 45666
rect 43484 45220 43540 45614
rect 43484 45106 43540 45164
rect 43932 45220 43988 45230
rect 43484 45054 43486 45106
rect 43538 45054 43540 45106
rect 43484 45042 43540 45054
rect 43708 45108 43764 45118
rect 43708 44546 43764 45052
rect 43820 44996 43876 45006
rect 43820 44902 43876 44940
rect 43708 44494 43710 44546
rect 43762 44494 43764 44546
rect 43708 44482 43764 44494
rect 43820 44436 43876 44446
rect 43820 44342 43876 44380
rect 43932 44100 43988 45164
rect 44268 45108 44324 45118
rect 44492 45108 44548 46398
rect 44268 45106 44548 45108
rect 44268 45054 44270 45106
rect 44322 45054 44548 45106
rect 44268 45052 44548 45054
rect 44268 45042 44324 45052
rect 43932 44034 43988 44044
rect 43372 43820 43540 43876
rect 42924 43762 42980 43774
rect 42924 43710 42926 43762
rect 42978 43710 42980 43762
rect 42924 43652 42980 43710
rect 43484 43764 43540 43820
rect 43484 43708 43652 43764
rect 43372 43652 43428 43662
rect 42924 43650 43428 43652
rect 42924 43598 43374 43650
rect 43426 43598 43428 43650
rect 42924 43596 43428 43598
rect 43372 43586 43428 43596
rect 42812 43486 42814 43538
rect 42866 43486 42868 43538
rect 42812 43474 42868 43486
rect 43260 43316 43316 43326
rect 42924 43314 43316 43316
rect 42924 43262 43262 43314
rect 43314 43262 43316 43314
rect 42924 43260 43316 43262
rect 42588 42754 42756 42756
rect 42588 42702 42590 42754
rect 42642 42702 42756 42754
rect 42588 42700 42756 42702
rect 42812 42756 42868 42766
rect 42924 42756 42980 43260
rect 43260 43250 43316 43260
rect 42812 42754 42980 42756
rect 42812 42702 42814 42754
rect 42866 42702 42980 42754
rect 42812 42700 42980 42702
rect 42588 42690 42644 42700
rect 42812 42690 42868 42700
rect 42364 42644 42420 42654
rect 42364 42550 42420 42588
rect 42476 42530 42532 42542
rect 42476 42478 42478 42530
rect 42530 42478 42532 42530
rect 42476 42196 42532 42478
rect 43484 42530 43540 42542
rect 43484 42478 43486 42530
rect 43538 42478 43540 42530
rect 42476 42140 43204 42196
rect 43148 42082 43204 42140
rect 43148 42030 43150 42082
rect 43202 42030 43204 42082
rect 43148 42018 43204 42030
rect 42364 41970 42420 41982
rect 42364 41918 42366 41970
rect 42418 41918 42420 41970
rect 42364 41860 42420 41918
rect 42364 41794 42420 41804
rect 42252 41580 42756 41636
rect 42140 41246 42142 41298
rect 42194 41246 42196 41298
rect 42140 41234 42196 41246
rect 42252 41186 42308 41198
rect 42252 41134 42254 41186
rect 42306 41134 42308 41186
rect 42028 41020 42196 41076
rect 42028 40852 42084 40862
rect 42028 40626 42084 40796
rect 42028 40574 42030 40626
rect 42082 40574 42084 40626
rect 42028 40562 42084 40574
rect 42140 40404 42196 41020
rect 42252 40628 42308 41134
rect 42252 40562 42308 40572
rect 42588 40516 42644 40526
rect 42588 40422 42644 40460
rect 42140 40348 42532 40404
rect 42140 39508 42196 39518
rect 42028 39506 42196 39508
rect 42028 39454 42142 39506
rect 42194 39454 42196 39506
rect 42028 39452 42196 39454
rect 41804 39006 41806 39058
rect 41858 39006 41860 39058
rect 41804 38994 41860 39006
rect 41916 39060 41972 39070
rect 42028 39060 42084 39452
rect 42140 39442 42196 39452
rect 42364 39396 42420 39406
rect 42252 39340 42364 39396
rect 42252 39060 42308 39340
rect 42364 39330 42420 39340
rect 42476 39172 42532 40348
rect 41916 39058 42084 39060
rect 41916 39006 41918 39058
rect 41970 39006 42084 39058
rect 41916 39004 42084 39006
rect 42140 39004 42308 39060
rect 42364 39116 42532 39172
rect 41916 38994 41972 39004
rect 42028 38836 42084 38846
rect 42140 38836 42196 39004
rect 42364 38836 42420 39116
rect 42588 38946 42644 38958
rect 42588 38894 42590 38946
rect 42642 38894 42644 38946
rect 41580 38834 42196 38836
rect 41580 38782 41582 38834
rect 41634 38782 42030 38834
rect 42082 38782 42196 38834
rect 41580 38780 42196 38782
rect 42252 38780 42420 38836
rect 42476 38836 42532 38846
rect 42588 38836 42644 38894
rect 42476 38834 42644 38836
rect 42476 38782 42478 38834
rect 42530 38782 42644 38834
rect 42476 38780 42644 38782
rect 41580 38770 41636 38780
rect 42028 38770 42084 38780
rect 42252 38668 42308 38780
rect 42476 38770 42532 38780
rect 41356 38612 41524 38668
rect 42140 38612 42308 38668
rect 42364 38612 42420 38622
rect 41356 38050 41412 38612
rect 41356 37998 41358 38050
rect 41410 37998 41412 38050
rect 41356 37986 41412 37998
rect 42028 37940 42084 37950
rect 42028 37846 42084 37884
rect 41356 37492 41412 37502
rect 41356 37398 41412 37436
rect 42140 37380 42196 38612
rect 41916 37378 42196 37380
rect 41916 37326 42142 37378
rect 42194 37326 42196 37378
rect 41916 37324 42196 37326
rect 41804 37266 41860 37278
rect 41804 37214 41806 37266
rect 41858 37214 41860 37266
rect 41804 37044 41860 37214
rect 40908 35634 40964 35644
rect 41020 36428 41300 36484
rect 41692 36988 41804 37044
rect 41692 36482 41748 36988
rect 41804 36978 41860 36988
rect 41916 36932 41972 37324
rect 42140 37314 42196 37324
rect 41916 36866 41972 36876
rect 42252 36484 42308 36494
rect 41692 36430 41694 36482
rect 41746 36430 41748 36482
rect 40908 35252 40964 35262
rect 40908 35026 40964 35196
rect 40908 34974 40910 35026
rect 40962 34974 40964 35026
rect 40908 34962 40964 34974
rect 40348 34598 40404 34636
rect 40348 34020 40404 34030
rect 40124 34018 40404 34020
rect 40124 33966 40350 34018
rect 40402 33966 40404 34018
rect 40124 33964 40404 33966
rect 40348 33684 40404 33964
rect 40348 33618 40404 33628
rect 40012 33058 40068 33068
rect 40684 32340 40740 32350
rect 40348 32116 40404 32126
rect 39900 31780 39956 31790
rect 39788 31778 39956 31780
rect 39788 31726 39902 31778
rect 39954 31726 39956 31778
rect 39788 31724 39956 31726
rect 39676 31668 39732 31678
rect 39340 31666 39732 31668
rect 39340 31614 39678 31666
rect 39730 31614 39732 31666
rect 39340 31612 39732 31614
rect 39340 31106 39396 31612
rect 39676 31602 39732 31612
rect 39340 31054 39342 31106
rect 39394 31054 39396 31106
rect 39340 30772 39396 31054
rect 39676 31444 39732 31454
rect 39676 31106 39732 31388
rect 39676 31054 39678 31106
rect 39730 31054 39732 31106
rect 39676 31042 39732 31054
rect 39340 30706 39396 30716
rect 39676 30884 39732 30894
rect 39788 30884 39844 31724
rect 39900 31714 39956 31724
rect 39732 30828 39844 30884
rect 40124 31108 40180 31118
rect 38556 30380 38836 30436
rect 39676 30434 39732 30828
rect 39676 30382 39678 30434
rect 39730 30382 39732 30434
rect 38556 30212 38612 30380
rect 39676 30370 39732 30382
rect 39900 30770 39956 30782
rect 39900 30718 39902 30770
rect 39954 30718 39956 30770
rect 39340 30322 39396 30334
rect 39340 30270 39342 30322
rect 39394 30270 39396 30322
rect 38444 30156 38612 30212
rect 38668 30212 38724 30222
rect 38444 30098 38500 30156
rect 38668 30118 38724 30156
rect 39004 30212 39060 30222
rect 39340 30212 39396 30270
rect 39004 30210 39396 30212
rect 39004 30158 39006 30210
rect 39058 30158 39396 30210
rect 39004 30156 39396 30158
rect 39004 30146 39060 30156
rect 38444 30046 38446 30098
rect 38498 30046 38500 30098
rect 38444 29764 38500 30046
rect 38444 29426 38500 29708
rect 38556 29986 38612 29998
rect 38556 29934 38558 29986
rect 38610 29934 38612 29986
rect 38556 29652 38612 29934
rect 39452 29988 39508 29998
rect 39452 29894 39508 29932
rect 38556 29586 38612 29596
rect 39004 29876 39060 29886
rect 39004 29650 39060 29820
rect 39004 29598 39006 29650
rect 39058 29598 39060 29650
rect 39004 29586 39060 29598
rect 39228 29764 39284 29774
rect 39228 29650 39284 29708
rect 39228 29598 39230 29650
rect 39282 29598 39284 29650
rect 39228 29586 39284 29598
rect 38444 29374 38446 29426
rect 38498 29374 38500 29426
rect 38444 29362 38500 29374
rect 38780 29428 38836 29438
rect 38780 29334 38836 29372
rect 39452 29428 39508 29438
rect 39452 29334 39508 29372
rect 38556 29316 38612 29326
rect 38556 29222 38612 29260
rect 39004 29316 39060 29326
rect 39060 29260 39172 29316
rect 39004 29250 39060 29260
rect 38892 29202 38948 29214
rect 38892 29150 38894 29202
rect 38946 29150 38948 29202
rect 38108 26462 38110 26514
rect 38162 26462 38164 26514
rect 38108 26450 38164 26462
rect 38220 26852 38388 26908
rect 38444 28420 38500 28430
rect 38444 26852 38500 28364
rect 37996 26404 38052 26414
rect 37884 25508 37940 25518
rect 37660 25506 37940 25508
rect 37660 25454 37886 25506
rect 37938 25454 37940 25506
rect 37660 25452 37940 25454
rect 37660 24836 37716 25452
rect 37884 25442 37940 25452
rect 37772 25284 37828 25294
rect 37996 25284 38052 26348
rect 37772 25190 37828 25228
rect 37884 25228 38052 25284
rect 37884 25060 37940 25228
rect 37660 23938 37716 24780
rect 37660 23886 37662 23938
rect 37714 23886 37716 23938
rect 37324 22930 37492 22932
rect 37324 22878 37326 22930
rect 37378 22878 37492 22930
rect 37324 22876 37492 22878
rect 37548 22932 37604 22942
rect 37324 22148 37380 22876
rect 37548 22838 37604 22876
rect 37548 22594 37604 22606
rect 37548 22542 37550 22594
rect 37602 22542 37604 22594
rect 37548 22482 37604 22542
rect 37548 22430 37550 22482
rect 37602 22430 37604 22482
rect 37548 22418 37604 22430
rect 37324 22082 37380 22092
rect 37660 21700 37716 23886
rect 37212 21644 37380 21700
rect 37212 21474 37268 21486
rect 37212 21422 37214 21474
rect 37266 21422 37268 21474
rect 36988 21362 37044 21374
rect 36988 21310 36990 21362
rect 37042 21310 37044 21362
rect 36988 20692 37044 21310
rect 37212 20802 37268 21422
rect 37212 20750 37214 20802
rect 37266 20750 37268 20802
rect 36988 20690 37156 20692
rect 36988 20638 36990 20690
rect 37042 20638 37156 20690
rect 36988 20636 37156 20638
rect 36988 20626 37044 20636
rect 37100 19908 37156 20636
rect 37100 19010 37156 19852
rect 37212 20020 37268 20750
rect 37212 19906 37268 19964
rect 37212 19854 37214 19906
rect 37266 19854 37268 19906
rect 37212 19794 37268 19854
rect 37212 19742 37214 19794
rect 37266 19742 37268 19794
rect 37212 19730 37268 19742
rect 37100 18958 37102 19010
rect 37154 18958 37156 19010
rect 36876 18620 37044 18676
rect 36764 18564 36820 18574
rect 36764 18470 36820 18508
rect 36876 18450 36932 18462
rect 36876 18398 36878 18450
rect 36930 18398 36932 18450
rect 36876 18340 36932 18398
rect 36652 18284 36932 18340
rect 36652 18116 36708 18284
rect 36988 18228 37044 18620
rect 36652 14196 36708 18060
rect 36876 18172 37044 18228
rect 36876 16772 36932 18172
rect 36876 16706 36932 16716
rect 37100 16324 37156 18958
rect 37324 18676 37380 21644
rect 37548 21644 37716 21700
rect 37772 25004 37940 25060
rect 38220 25060 38276 26852
rect 38444 26514 38500 26796
rect 38444 26462 38446 26514
rect 38498 26462 38500 26514
rect 38444 26450 38500 26462
rect 38556 28418 38612 28430
rect 38556 28366 38558 28418
rect 38610 28366 38612 28418
rect 38556 27858 38612 28366
rect 38556 27806 38558 27858
rect 38610 27806 38612 27858
rect 38556 26404 38612 27806
rect 38668 27860 38724 27870
rect 38668 27298 38724 27804
rect 38780 27748 38836 27758
rect 38780 27654 38836 27692
rect 38668 27246 38670 27298
rect 38722 27246 38724 27298
rect 38668 27234 38724 27246
rect 38780 27076 38836 27086
rect 38892 27076 38948 29150
rect 39004 28420 39060 28430
rect 39004 28326 39060 28364
rect 39004 28084 39060 28094
rect 39116 28084 39172 29260
rect 39004 28082 39172 28084
rect 39004 28030 39006 28082
rect 39058 28030 39172 28082
rect 39004 28028 39172 28030
rect 39004 28018 39060 28028
rect 39228 27860 39284 27870
rect 39228 27766 39284 27804
rect 39116 27746 39172 27758
rect 39116 27694 39118 27746
rect 39170 27694 39172 27746
rect 39116 27636 39172 27694
rect 39900 27636 39956 30718
rect 40124 30210 40180 31052
rect 40124 30158 40126 30210
rect 40178 30158 40180 30210
rect 40124 30146 40180 30158
rect 40236 30770 40292 30782
rect 40236 30718 40238 30770
rect 40290 30718 40292 30770
rect 40236 30212 40292 30718
rect 40236 30146 40292 30156
rect 40012 29988 40068 29998
rect 40012 29894 40068 29932
rect 39116 27580 39956 27636
rect 40012 28028 40292 28084
rect 38780 27074 38948 27076
rect 38780 27022 38782 27074
rect 38834 27022 38948 27074
rect 38780 27020 38948 27022
rect 39900 27188 39956 27198
rect 38780 27010 38836 27020
rect 38668 26962 38724 26974
rect 38668 26910 38670 26962
rect 38722 26910 38724 26962
rect 38668 26908 38724 26910
rect 39340 26962 39396 26974
rect 39340 26910 39342 26962
rect 39394 26910 39396 26962
rect 39340 26908 39396 26910
rect 38668 26852 39508 26908
rect 38556 26338 38612 26348
rect 39228 26290 39284 26302
rect 39228 26238 39230 26290
rect 39282 26238 39284 26290
rect 39004 26180 39060 26190
rect 38556 26178 39060 26180
rect 38556 26126 39006 26178
rect 39058 26126 39060 26178
rect 38556 26124 39060 26126
rect 38444 25620 38500 25630
rect 38556 25620 38612 26124
rect 39004 26114 39060 26124
rect 39228 25956 39284 26238
rect 39116 25844 39172 25854
rect 38780 25732 38836 25742
rect 38836 25676 38948 25732
rect 38780 25666 38836 25676
rect 38444 25618 38612 25620
rect 38444 25566 38446 25618
rect 38498 25566 38612 25618
rect 38444 25564 38612 25566
rect 38444 25554 38500 25564
rect 38556 25396 38612 25406
rect 38612 25340 38836 25396
rect 38556 25302 38612 25340
rect 38332 25284 38388 25294
rect 38332 25190 38388 25228
rect 38220 25004 38388 25060
rect 37772 23380 37828 25004
rect 37436 20804 37492 20814
rect 37436 20710 37492 20748
rect 37100 16258 37156 16268
rect 37212 18620 37380 18676
rect 37436 19234 37492 19246
rect 37436 19182 37438 19234
rect 37490 19182 37492 19234
rect 37212 16772 37268 18620
rect 37324 18450 37380 18462
rect 37324 18398 37326 18450
rect 37378 18398 37380 18450
rect 37324 18116 37380 18398
rect 37324 18050 37380 18060
rect 37436 17890 37492 19182
rect 37548 18676 37604 21644
rect 37660 21476 37716 21486
rect 37660 21382 37716 21420
rect 37660 21028 37716 21038
rect 37660 20934 37716 20972
rect 37660 19906 37716 19918
rect 37660 19854 37662 19906
rect 37714 19854 37716 19906
rect 37660 19794 37716 19854
rect 37660 19742 37662 19794
rect 37714 19742 37716 19794
rect 37660 18788 37716 19742
rect 37772 19348 37828 23324
rect 37884 24724 37940 24734
rect 37884 22036 37940 24668
rect 38220 24610 38276 24622
rect 38220 24558 38222 24610
rect 38274 24558 38276 24610
rect 37996 23940 38052 23950
rect 37996 23846 38052 23884
rect 38108 23714 38164 23726
rect 38108 23662 38110 23714
rect 38162 23662 38164 23714
rect 37884 21970 37940 21980
rect 37996 23604 38052 23614
rect 37996 21028 38052 23548
rect 38108 23380 38164 23662
rect 38220 23714 38276 24558
rect 38332 23940 38388 25004
rect 38780 24946 38836 25340
rect 38780 24894 38782 24946
rect 38834 24894 38836 24946
rect 38780 24882 38836 24894
rect 38444 24500 38500 24510
rect 38444 24406 38500 24444
rect 38332 23884 38500 23940
rect 38220 23662 38222 23714
rect 38274 23662 38276 23714
rect 38220 23492 38276 23662
rect 38220 23426 38276 23436
rect 38108 23314 38164 23324
rect 38108 23042 38164 23054
rect 38108 22990 38110 23042
rect 38162 22990 38164 23042
rect 38108 22596 38164 22990
rect 38108 22530 38164 22540
rect 38332 22258 38388 22270
rect 38332 22206 38334 22258
rect 38386 22206 38388 22258
rect 38220 22148 38276 22158
rect 38332 22148 38388 22206
rect 38276 22092 38388 22148
rect 38220 22082 38276 22092
rect 38108 21588 38164 21598
rect 38108 21494 38164 21532
rect 38332 21362 38388 21374
rect 38332 21310 38334 21362
rect 38386 21310 38388 21362
rect 38108 21028 38164 21038
rect 37996 21026 38164 21028
rect 37996 20974 38110 21026
rect 38162 20974 38164 21026
rect 37996 20972 38164 20974
rect 38108 20962 38164 20972
rect 38332 21028 38388 21310
rect 38332 20962 38388 20972
rect 38108 19908 38164 19918
rect 38108 19814 38164 19852
rect 37772 19236 37828 19292
rect 37884 19236 37940 19246
rect 37772 19234 37940 19236
rect 37772 19182 37886 19234
rect 37938 19182 37940 19234
rect 37772 19180 37940 19182
rect 37884 19170 37940 19180
rect 38108 19236 38164 19246
rect 38108 19142 38164 19180
rect 37996 19010 38052 19022
rect 37996 18958 37998 19010
rect 38050 18958 38052 19010
rect 37772 18788 37828 18798
rect 37660 18732 37772 18788
rect 37772 18722 37828 18732
rect 37548 18620 37716 18676
rect 37548 18450 37604 18462
rect 37548 18398 37550 18450
rect 37602 18398 37604 18450
rect 37548 18228 37604 18398
rect 37548 18162 37604 18172
rect 37436 17838 37438 17890
rect 37490 17838 37492 17890
rect 37436 17826 37492 17838
rect 37548 17554 37604 17566
rect 37548 17502 37550 17554
rect 37602 17502 37604 17554
rect 37436 17442 37492 17454
rect 37436 17390 37438 17442
rect 37490 17390 37492 17442
rect 37436 17332 37492 17390
rect 37436 17266 37492 17276
rect 37324 16772 37380 16782
rect 37212 16770 37380 16772
rect 37212 16718 37326 16770
rect 37378 16718 37380 16770
rect 37212 16716 37380 16718
rect 36988 15988 37044 15998
rect 36988 15894 37044 15932
rect 37100 15874 37156 15886
rect 37100 15822 37102 15874
rect 37154 15822 37156 15874
rect 37100 15540 37156 15822
rect 37100 15474 37156 15484
rect 36988 15314 37044 15326
rect 36988 15262 36990 15314
rect 37042 15262 37044 15314
rect 36988 14532 37044 15262
rect 37212 15148 37268 16716
rect 37324 16706 37380 16716
rect 37548 16548 37604 17502
rect 37548 16482 37604 16492
rect 37436 15988 37492 15998
rect 37324 15876 37380 15886
rect 37324 15782 37380 15820
rect 37436 15540 37492 15932
rect 37324 15484 37492 15540
rect 37548 15986 37604 15998
rect 37548 15934 37550 15986
rect 37602 15934 37604 15986
rect 37324 15314 37380 15484
rect 37324 15262 37326 15314
rect 37378 15262 37380 15314
rect 37324 15250 37380 15262
rect 37436 15202 37492 15214
rect 37436 15150 37438 15202
rect 37490 15150 37492 15202
rect 37212 15092 37380 15148
rect 37212 14532 37268 14542
rect 36988 14476 37212 14532
rect 37212 14438 37268 14476
rect 36988 14308 37044 14318
rect 36988 14214 37044 14252
rect 37100 14306 37156 14318
rect 37100 14254 37102 14306
rect 37154 14254 37156 14306
rect 36652 14130 36708 14140
rect 37100 13972 37156 14254
rect 37324 14084 37380 15092
rect 36652 13916 37156 13972
rect 37212 14028 37380 14084
rect 36652 13746 36708 13916
rect 36652 13694 36654 13746
rect 36706 13694 36708 13746
rect 36652 13682 36708 13694
rect 36764 13748 36820 13758
rect 36764 13654 36820 13692
rect 36204 10742 36260 10780
rect 36316 11732 36596 11788
rect 36652 13524 36708 13534
rect 35308 9996 35700 10052
rect 35756 10050 35924 10052
rect 35756 9998 35870 10050
rect 35922 9998 35924 10050
rect 35756 9996 35924 9998
rect 35308 9604 35364 9996
rect 35756 9940 35812 9996
rect 35868 9986 35924 9996
rect 35980 10610 36036 10622
rect 35980 10558 35982 10610
rect 36034 10558 36036 10610
rect 35980 10500 36036 10558
rect 36092 10612 36148 10622
rect 36092 10518 36148 10556
rect 35420 9884 35812 9940
rect 35420 9826 35476 9884
rect 35420 9774 35422 9826
rect 35474 9774 35476 9826
rect 35420 9762 35476 9774
rect 35756 9716 35812 9726
rect 35756 9622 35812 9660
rect 35308 9548 35476 9604
rect 34972 9268 35028 9278
rect 34972 9174 35028 9212
rect 35084 9268 35140 9436
rect 35196 9268 35252 9278
rect 35084 9266 35196 9268
rect 35084 9214 35086 9266
rect 35138 9214 35196 9266
rect 35084 9212 35196 9214
rect 35084 9202 35140 9212
rect 35196 9202 35252 9212
rect 35308 9156 35364 9166
rect 35308 9062 35364 9100
rect 34860 8988 35028 9044
rect 34300 8318 34302 8370
rect 34354 8318 34356 8370
rect 34300 8306 34356 8318
rect 34076 8204 34244 8260
rect 34188 8148 34244 8204
rect 34748 8148 34804 8158
rect 34188 8146 34804 8148
rect 34188 8094 34750 8146
rect 34802 8094 34804 8146
rect 34188 8092 34804 8094
rect 34748 8082 34804 8092
rect 33852 7364 33908 7374
rect 33852 7362 34692 7364
rect 33852 7310 33854 7362
rect 33906 7310 34692 7362
rect 33852 7308 34692 7310
rect 33852 7298 33908 7308
rect 33628 7084 34020 7140
rect 33292 4228 33348 4238
rect 33292 4226 33572 4228
rect 33292 4174 33294 4226
rect 33346 4174 33572 4226
rect 33292 4172 33572 4174
rect 33292 4162 33348 4172
rect 33516 3556 33572 4172
rect 33964 3666 34020 7084
rect 34636 6914 34692 7308
rect 34636 6862 34638 6914
rect 34690 6862 34692 6914
rect 34636 6850 34692 6862
rect 34860 6690 34916 6702
rect 34860 6638 34862 6690
rect 34914 6638 34916 6690
rect 34748 6580 34804 6590
rect 34860 6580 34916 6638
rect 34748 6578 34916 6580
rect 34748 6526 34750 6578
rect 34802 6526 34916 6578
rect 34748 6524 34916 6526
rect 34748 6514 34804 6524
rect 34972 5012 35028 8988
rect 35084 8930 35140 8942
rect 35084 8878 35086 8930
rect 35138 8878 35140 8930
rect 35084 6690 35140 8878
rect 35420 8932 35476 9548
rect 35980 9492 36036 10444
rect 35532 9436 36036 9492
rect 35532 9154 35588 9436
rect 35868 9268 35924 9278
rect 35868 9174 35924 9212
rect 35532 9102 35534 9154
rect 35586 9102 35588 9154
rect 35532 9090 35588 9102
rect 36092 9044 36148 9054
rect 35980 9042 36148 9044
rect 35980 8990 36094 9042
rect 36146 8990 36148 9042
rect 35980 8988 36148 8990
rect 35420 8876 35924 8932
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35420 8484 35476 8494
rect 35420 8258 35476 8428
rect 35420 8206 35422 8258
rect 35474 8206 35476 8258
rect 35420 8194 35476 8206
rect 35532 7700 35588 7710
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35308 6804 35364 6814
rect 35532 6804 35588 7644
rect 35308 6802 35588 6804
rect 35308 6750 35310 6802
rect 35362 6750 35588 6802
rect 35308 6748 35588 6750
rect 35308 6738 35364 6748
rect 35084 6638 35086 6690
rect 35138 6638 35140 6690
rect 35084 6626 35140 6638
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35084 5012 35140 5022
rect 34972 4956 35084 5012
rect 35084 4946 35140 4956
rect 34188 4228 34244 4238
rect 34188 4226 34468 4228
rect 34188 4174 34190 4226
rect 34242 4174 34468 4226
rect 34188 4172 34468 4174
rect 34188 4162 34244 4172
rect 33964 3614 33966 3666
rect 34018 3614 34020 3666
rect 33964 3602 34020 3614
rect 33516 3462 33572 3500
rect 34412 3554 34468 4172
rect 34860 4226 34916 4238
rect 34860 4174 34862 4226
rect 34914 4174 34916 4226
rect 34412 3502 34414 3554
rect 34466 3502 34468 3554
rect 33180 3390 33182 3442
rect 33234 3390 33236 3442
rect 33180 3378 33236 3390
rect 34412 2548 34468 3502
rect 34748 3780 34804 3790
rect 34748 3442 34804 3724
rect 34748 3390 34750 3442
rect 34802 3390 34804 3442
rect 34748 3378 34804 3390
rect 33628 2492 34468 2548
rect 34860 2996 34916 4174
rect 35756 4226 35812 4238
rect 35756 4174 35758 4226
rect 35810 4174 35812 4226
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35420 3668 35476 3678
rect 35084 3442 35140 3454
rect 35084 3390 35086 3442
rect 35138 3390 35140 3442
rect 35084 2996 35140 3390
rect 34860 2940 35140 2996
rect 35196 3444 35252 3454
rect 33628 800 33684 2492
rect 34860 2436 34916 2940
rect 35196 2884 35252 3388
rect 35420 3442 35476 3612
rect 35420 3390 35422 3442
rect 35474 3390 35476 3442
rect 35420 3378 35476 3390
rect 35756 3444 35812 4174
rect 35868 3444 35924 8876
rect 35980 8258 36036 8988
rect 36092 8978 36148 8988
rect 35980 8206 35982 8258
rect 36034 8206 36036 8258
rect 35980 7362 36036 8206
rect 35980 7310 35982 7362
rect 36034 7310 36036 7362
rect 35980 7298 36036 7310
rect 36316 4340 36372 11732
rect 36540 10836 36596 10846
rect 36540 9938 36596 10780
rect 36540 9886 36542 9938
rect 36594 9886 36596 9938
rect 36540 9874 36596 9886
rect 36652 8820 36708 13468
rect 37212 13188 37268 14028
rect 37436 13972 37492 15150
rect 37548 14308 37604 15934
rect 37660 15874 37716 18620
rect 37884 18564 37940 18574
rect 37772 18562 37940 18564
rect 37772 18510 37886 18562
rect 37938 18510 37940 18562
rect 37772 18508 37940 18510
rect 37996 18564 38052 18958
rect 38444 19012 38500 23884
rect 38892 23938 38948 25676
rect 39116 25284 39172 25788
rect 39116 24836 39172 25228
rect 39228 25172 39284 25900
rect 39340 25844 39396 25854
rect 39340 25506 39396 25788
rect 39340 25454 39342 25506
rect 39394 25454 39396 25506
rect 39340 25442 39396 25454
rect 39228 25116 39396 25172
rect 39116 24834 39284 24836
rect 39116 24782 39118 24834
rect 39170 24782 39284 24834
rect 39116 24780 39284 24782
rect 39116 24770 39172 24780
rect 39228 24162 39284 24780
rect 39340 24722 39396 25116
rect 39340 24670 39342 24722
rect 39394 24670 39396 24722
rect 39340 24658 39396 24670
rect 39228 24110 39230 24162
rect 39282 24110 39284 24162
rect 39228 24098 39284 24110
rect 39116 23940 39172 23950
rect 38892 23886 38894 23938
rect 38946 23886 38948 23938
rect 38556 23826 38612 23838
rect 38556 23774 38558 23826
rect 38610 23774 38612 23826
rect 38556 23492 38612 23774
rect 38780 23716 38836 23726
rect 38780 23622 38836 23660
rect 38556 22370 38612 23436
rect 38892 23380 38948 23886
rect 38556 22318 38558 22370
rect 38610 22318 38612 22370
rect 38556 22306 38612 22318
rect 38780 23324 38948 23380
rect 39004 23884 39116 23940
rect 38556 22036 38612 22046
rect 38556 20242 38612 21980
rect 38668 21476 38724 21486
rect 38668 21382 38724 21420
rect 38780 21140 38836 23324
rect 38892 23156 38948 23166
rect 38892 23062 38948 23100
rect 38892 22260 38948 22270
rect 39004 22260 39060 23884
rect 39116 23846 39172 23884
rect 39340 23156 39396 23166
rect 39340 23062 39396 23100
rect 39116 23044 39172 23054
rect 39116 22596 39172 22988
rect 39116 22530 39172 22540
rect 39228 22932 39284 22942
rect 39228 22594 39284 22876
rect 39228 22542 39230 22594
rect 39282 22542 39284 22594
rect 39228 22530 39284 22542
rect 39452 22596 39508 26852
rect 39900 26402 39956 27132
rect 40012 26516 40068 28028
rect 40236 27970 40292 28028
rect 40236 27918 40238 27970
rect 40290 27918 40292 27970
rect 40236 27906 40292 27918
rect 40012 26450 40068 26460
rect 40124 27860 40180 27870
rect 39900 26350 39902 26402
rect 39954 26350 39956 26402
rect 39900 26338 39956 26350
rect 40012 26292 40068 26302
rect 39900 25620 39956 25630
rect 40012 25620 40068 26236
rect 39900 25618 40068 25620
rect 39900 25566 39902 25618
rect 39954 25566 40068 25618
rect 39900 25564 40068 25566
rect 39900 25554 39956 25564
rect 39788 25508 39844 25518
rect 39788 25414 39844 25452
rect 40124 24948 40180 27804
rect 40236 27524 40292 27534
rect 40236 27186 40292 27468
rect 40236 27134 40238 27186
rect 40290 27134 40292 27186
rect 40236 27122 40292 27134
rect 40348 26908 40404 32060
rect 40684 31890 40740 32284
rect 40684 31838 40686 31890
rect 40738 31838 40740 31890
rect 40684 31826 40740 31838
rect 41020 31892 41076 36428
rect 41692 36418 41748 36430
rect 42028 36482 42308 36484
rect 42028 36430 42254 36482
rect 42306 36430 42308 36482
rect 42028 36428 42308 36430
rect 41916 36372 41972 36382
rect 41132 36258 41188 36270
rect 41132 36206 41134 36258
rect 41186 36206 41188 36258
rect 41132 36148 41188 36206
rect 41132 36082 41188 36092
rect 41804 36260 41860 36270
rect 41244 35924 41300 35934
rect 41244 35830 41300 35868
rect 41468 35810 41524 35822
rect 41468 35758 41470 35810
rect 41522 35758 41524 35810
rect 41132 35698 41188 35710
rect 41132 35646 41134 35698
rect 41186 35646 41188 35698
rect 41132 34914 41188 35646
rect 41468 35700 41524 35758
rect 41580 35700 41636 35710
rect 41468 35698 41636 35700
rect 41468 35646 41582 35698
rect 41634 35646 41636 35698
rect 41468 35644 41636 35646
rect 41580 35634 41636 35644
rect 41132 34862 41134 34914
rect 41186 34862 41188 34914
rect 41132 34356 41188 34862
rect 41468 35252 41524 35262
rect 41468 34914 41524 35196
rect 41804 35138 41860 36204
rect 41916 36148 41972 36316
rect 41916 36082 41972 36092
rect 41916 35924 41972 35934
rect 42028 35924 42084 36428
rect 42252 36418 42308 36428
rect 41916 35922 42084 35924
rect 41916 35870 41918 35922
rect 41970 35870 42084 35922
rect 41916 35868 42084 35870
rect 42252 36148 42308 36158
rect 41916 35858 41972 35868
rect 42252 35810 42308 36092
rect 42252 35758 42254 35810
rect 42306 35758 42308 35810
rect 42252 35746 42308 35758
rect 41804 35086 41806 35138
rect 41858 35086 41860 35138
rect 41804 35074 41860 35086
rect 42028 35700 42084 35710
rect 41468 34862 41470 34914
rect 41522 34862 41524 34914
rect 41468 34850 41524 34862
rect 42028 34916 42084 35644
rect 42252 34916 42308 34926
rect 42084 34914 42308 34916
rect 42084 34862 42254 34914
rect 42306 34862 42308 34914
rect 42084 34860 42308 34862
rect 42028 34850 42084 34860
rect 42252 34850 42308 34860
rect 42364 34916 42420 38556
rect 42588 36708 42644 36718
rect 42588 36594 42644 36652
rect 42588 36542 42590 36594
rect 42642 36542 42644 36594
rect 42588 36530 42644 36542
rect 42700 36482 42756 41580
rect 42812 41186 42868 41198
rect 42812 41134 42814 41186
rect 42866 41134 42868 41186
rect 42812 40740 42868 41134
rect 43484 40740 43540 42478
rect 42812 40684 43540 40740
rect 43596 41298 43652 43708
rect 43820 43426 43876 43438
rect 43820 43374 43822 43426
rect 43874 43374 43876 43426
rect 43820 43316 43876 43374
rect 43820 43250 43876 43260
rect 43596 41246 43598 41298
rect 43650 41246 43652 41298
rect 42812 40402 42868 40414
rect 42812 40350 42814 40402
rect 42866 40350 42868 40402
rect 42812 40180 42868 40350
rect 42812 40114 42868 40124
rect 43260 40402 43316 40684
rect 43260 40350 43262 40402
rect 43314 40350 43316 40402
rect 43148 39844 43204 39854
rect 42812 38946 42868 38958
rect 42812 38894 42814 38946
rect 42866 38894 42868 38946
rect 42812 38052 42868 38894
rect 42924 38834 42980 38846
rect 42924 38782 42926 38834
rect 42978 38782 42980 38834
rect 42924 38668 42980 38782
rect 42924 38612 43092 38668
rect 42812 37986 42868 37996
rect 42700 36430 42702 36482
rect 42754 36430 42756 36482
rect 42700 36418 42756 36430
rect 42812 36484 42868 36494
rect 42812 36390 42868 36428
rect 42476 36260 42532 36270
rect 42476 36166 42532 36204
rect 43036 36148 43092 38612
rect 42700 36092 43092 36148
rect 42700 36036 42756 36092
rect 42364 34850 42420 34860
rect 42588 35980 42756 36036
rect 41132 34290 41188 34300
rect 41692 34692 41748 34702
rect 41692 33124 41748 34636
rect 42028 34690 42084 34702
rect 42028 34638 42030 34690
rect 42082 34638 42084 34690
rect 42028 34356 42084 34638
rect 42028 34290 42084 34300
rect 42140 34690 42196 34702
rect 42140 34638 42142 34690
rect 42194 34638 42196 34690
rect 41356 33068 41748 33124
rect 42028 34130 42084 34142
rect 42028 34078 42030 34130
rect 42082 34078 42084 34130
rect 42028 34020 42084 34078
rect 41244 32340 41300 32350
rect 41020 31836 41188 31892
rect 41020 31666 41076 31678
rect 41020 31614 41022 31666
rect 41074 31614 41076 31666
rect 41020 31108 41076 31614
rect 41020 31042 41076 31052
rect 40796 30884 40852 30894
rect 41020 30884 41076 30894
rect 40852 30855 40964 30884
rect 40852 30828 40910 30855
rect 40796 30818 40852 30828
rect 40908 30803 40910 30828
rect 40962 30803 40964 30855
rect 40908 30791 40964 30803
rect 40684 30212 40740 30222
rect 40684 30118 40740 30156
rect 41020 30098 41076 30828
rect 41020 30046 41022 30098
rect 41074 30046 41076 30098
rect 41020 30034 41076 30046
rect 40684 29428 40740 29438
rect 40684 28754 40740 29372
rect 40684 28702 40686 28754
rect 40738 28702 40740 28754
rect 40684 28690 40740 28702
rect 40796 29092 40852 29102
rect 40796 28642 40852 29036
rect 41132 28868 41188 31836
rect 41244 31778 41300 32284
rect 41244 31726 41246 31778
rect 41298 31726 41300 31778
rect 41244 31714 41300 31726
rect 41132 28812 41300 28868
rect 40796 28590 40798 28642
rect 40850 28590 40852 28642
rect 40796 28578 40852 28590
rect 41132 28642 41188 28654
rect 41132 28590 41134 28642
rect 41186 28590 41188 28642
rect 40572 28418 40628 28430
rect 40572 28366 40574 28418
rect 40626 28366 40628 28418
rect 40460 27860 40516 27870
rect 40572 27860 40628 28366
rect 40460 27858 40628 27860
rect 40460 27806 40462 27858
rect 40514 27806 40628 27858
rect 40460 27804 40628 27806
rect 40460 27412 40516 27804
rect 40908 27636 40964 27646
rect 40908 27542 40964 27580
rect 40460 27356 40964 27412
rect 40796 27076 40852 27086
rect 40796 26908 40852 27020
rect 40908 27074 40964 27356
rect 41132 27186 41188 28590
rect 41244 28308 41300 28812
rect 41244 28242 41300 28252
rect 41356 28084 41412 33068
rect 41692 32564 41748 32574
rect 41692 32470 41748 32508
rect 42028 32340 42084 33964
rect 42140 34018 42196 34638
rect 42588 34242 42644 35980
rect 42700 35700 42756 35710
rect 42700 35698 42868 35700
rect 42700 35646 42702 35698
rect 42754 35646 42868 35698
rect 42700 35644 42868 35646
rect 42700 35634 42756 35644
rect 42812 35588 42868 35644
rect 42700 35364 42756 35374
rect 42700 34914 42756 35308
rect 42700 34862 42702 34914
rect 42754 34862 42756 34914
rect 42700 34850 42756 34862
rect 42588 34190 42590 34242
rect 42642 34190 42644 34242
rect 42588 34178 42644 34190
rect 42140 33966 42142 34018
rect 42194 33966 42196 34018
rect 42140 33954 42196 33966
rect 42700 33570 42756 33582
rect 42700 33518 42702 33570
rect 42754 33518 42756 33570
rect 42700 33458 42756 33518
rect 42700 33406 42702 33458
rect 42754 33406 42756 33458
rect 42700 33394 42756 33406
rect 42812 32564 42868 35532
rect 42924 34916 42980 34926
rect 42924 33348 42980 34860
rect 43036 34132 43092 34142
rect 43148 34132 43204 39788
rect 43260 38724 43316 40350
rect 43484 40516 43540 40526
rect 43596 40516 43652 41246
rect 43932 41186 43988 41198
rect 43932 41134 43934 41186
rect 43986 41134 43988 41186
rect 43932 40740 43988 41134
rect 43932 40674 43988 40684
rect 44380 40964 44436 40974
rect 43596 40460 43876 40516
rect 43484 40404 43540 40460
rect 43484 40402 43764 40404
rect 43484 40350 43486 40402
rect 43538 40350 43764 40402
rect 43484 40348 43764 40350
rect 43484 40338 43540 40348
rect 43372 40292 43428 40302
rect 43372 40198 43428 40236
rect 43260 38658 43316 38668
rect 43260 36708 43316 36718
rect 43316 36652 43428 36708
rect 43260 36642 43316 36652
rect 43372 35810 43428 36652
rect 43372 35758 43374 35810
rect 43426 35758 43428 35810
rect 43372 35746 43428 35758
rect 43484 36258 43540 36270
rect 43484 36206 43486 36258
rect 43538 36206 43540 36258
rect 43484 35700 43540 36206
rect 43708 36260 43764 40348
rect 43820 40180 43876 40460
rect 44380 40402 44436 40908
rect 44380 40350 44382 40402
rect 44434 40350 44436 40402
rect 44380 40338 44436 40350
rect 43932 40292 43988 40302
rect 43932 40198 43988 40236
rect 44268 40292 44324 40302
rect 43820 39058 43876 40124
rect 44268 39730 44324 40236
rect 44604 40180 44660 49980
rect 44828 49026 44884 50092
rect 44940 49812 44996 49822
rect 45164 49812 45220 52108
rect 45276 50036 45332 55412
rect 45500 55410 46564 55412
rect 45500 55358 45502 55410
rect 45554 55358 46564 55410
rect 45500 55356 46564 55358
rect 45500 55346 45556 55356
rect 46508 55300 46564 55356
rect 48412 55300 48468 55310
rect 48748 55300 48804 55310
rect 46508 55244 46676 55300
rect 46396 55188 46452 55198
rect 46284 54740 46340 54750
rect 45948 54738 46340 54740
rect 45948 54686 46286 54738
rect 46338 54686 46340 54738
rect 45948 54684 46340 54686
rect 45500 54404 45556 54414
rect 45948 54404 46004 54684
rect 46284 54674 46340 54684
rect 46396 54738 46452 55132
rect 46396 54686 46398 54738
rect 46450 54686 46452 54738
rect 46396 54674 46452 54686
rect 45500 54402 46004 54404
rect 45500 54350 45502 54402
rect 45554 54350 46004 54402
rect 45500 54348 46004 54350
rect 46060 54514 46116 54526
rect 46060 54462 46062 54514
rect 46114 54462 46116 54514
rect 45500 53844 45556 54348
rect 45388 53508 45444 53518
rect 45388 52946 45444 53452
rect 45388 52894 45390 52946
rect 45442 52894 45444 52946
rect 45388 52882 45444 52894
rect 45388 51490 45444 51502
rect 45388 51438 45390 51490
rect 45442 51438 45444 51490
rect 45388 51380 45444 51438
rect 45388 51314 45444 51324
rect 45500 50148 45556 53788
rect 45612 53844 45668 53854
rect 45724 53844 45780 53854
rect 45612 53842 45724 53844
rect 45612 53790 45614 53842
rect 45666 53790 45724 53842
rect 45612 53788 45724 53790
rect 45612 53778 45668 53788
rect 45612 53508 45668 53518
rect 45612 53170 45668 53452
rect 45612 53118 45614 53170
rect 45666 53118 45668 53170
rect 45612 53106 45668 53118
rect 45724 52948 45780 53788
rect 46060 53620 46116 54462
rect 46508 54514 46564 54526
rect 46508 54462 46510 54514
rect 46562 54462 46564 54514
rect 46396 54404 46452 54414
rect 46396 54180 46452 54348
rect 46060 53554 46116 53564
rect 46284 54124 46452 54180
rect 46172 53508 46228 53518
rect 46172 53170 46228 53452
rect 46172 53118 46174 53170
rect 46226 53118 46228 53170
rect 46172 53106 46228 53118
rect 46284 53170 46340 54124
rect 46508 54068 46564 54462
rect 46508 54002 46564 54012
rect 46620 54514 46676 55244
rect 48412 55298 48916 55300
rect 48412 55246 48414 55298
rect 48466 55246 48750 55298
rect 48802 55246 48916 55298
rect 48412 55244 48916 55246
rect 47628 55188 47684 55198
rect 47628 55186 48132 55188
rect 47628 55134 47630 55186
rect 47682 55134 48132 55186
rect 47628 55132 48132 55134
rect 47628 55122 47684 55132
rect 48076 54738 48132 55132
rect 48076 54686 48078 54738
rect 48130 54686 48132 54738
rect 48076 54674 48132 54686
rect 47068 54516 47124 54526
rect 46620 54462 46622 54514
rect 46674 54462 46676 54514
rect 46620 53844 46676 54462
rect 46284 53118 46286 53170
rect 46338 53118 46340 53170
rect 46284 53106 46340 53118
rect 46396 53788 46676 53844
rect 46956 54514 47124 54516
rect 46956 54462 47070 54514
rect 47122 54462 47124 54514
rect 46956 54460 47124 54462
rect 46060 52948 46116 52958
rect 45724 52946 46116 52948
rect 45724 52894 46062 52946
rect 46114 52894 46116 52946
rect 45724 52892 46116 52894
rect 46060 52052 46116 52892
rect 46396 52946 46452 53788
rect 46508 53620 46564 53630
rect 46508 53172 46564 53564
rect 46956 53172 47012 54460
rect 47068 54450 47124 54460
rect 47292 54514 47348 54526
rect 47292 54462 47294 54514
rect 47346 54462 47348 54514
rect 47292 53844 47348 54462
rect 47516 54514 47572 54526
rect 47516 54462 47518 54514
rect 47570 54462 47572 54514
rect 47292 53778 47348 53788
rect 47404 54402 47460 54414
rect 47404 54350 47406 54402
rect 47458 54350 47460 54402
rect 46508 53170 47012 53172
rect 46508 53118 46510 53170
rect 46562 53118 46958 53170
rect 47010 53118 47012 53170
rect 46508 53116 47012 53118
rect 46508 53106 46564 53116
rect 46956 53106 47012 53116
rect 47404 53060 47460 54350
rect 47516 53620 47572 54462
rect 47740 54516 47796 54526
rect 47740 54422 47796 54460
rect 48188 54404 48244 54414
rect 48188 54310 48244 54348
rect 48412 53732 48468 55244
rect 48748 55234 48804 55244
rect 48860 54738 48916 55244
rect 49532 55188 49588 55198
rect 48860 54686 48862 54738
rect 48914 54686 48916 54738
rect 48860 53844 48916 54686
rect 49420 55186 49588 55188
rect 49420 55134 49534 55186
rect 49586 55134 49588 55186
rect 49420 55132 49588 55134
rect 49420 54738 49476 55132
rect 49532 55122 49588 55132
rect 49420 54686 49422 54738
rect 49474 54686 49476 54738
rect 49420 54674 49476 54686
rect 49644 54516 49700 55356
rect 51660 55412 51716 55422
rect 51660 55318 51716 55356
rect 52108 55074 52164 55086
rect 52108 55022 52110 55074
rect 52162 55022 52164 55074
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 49308 54404 49364 54414
rect 49308 54402 49588 54404
rect 49308 54350 49310 54402
rect 49362 54350 49588 54402
rect 49308 54348 49588 54350
rect 49308 54338 49364 54348
rect 48972 53844 49028 53854
rect 48860 53842 49028 53844
rect 48860 53790 48974 53842
rect 49026 53790 49028 53842
rect 48860 53788 49028 53790
rect 48972 53778 49028 53788
rect 49532 53842 49588 54348
rect 49532 53790 49534 53842
rect 49586 53790 49588 53842
rect 49532 53778 49588 53790
rect 48412 53638 48468 53676
rect 49644 53730 49700 54460
rect 52108 54628 52164 55022
rect 52108 54572 53060 54628
rect 49868 54402 49924 54414
rect 50204 54404 50260 54414
rect 49868 54350 49870 54402
rect 49922 54350 49924 54402
rect 49868 53732 49924 54350
rect 49644 53678 49646 53730
rect 49698 53678 49700 53730
rect 47516 53554 47572 53564
rect 47740 53618 47796 53630
rect 47740 53566 47742 53618
rect 47794 53566 47796 53618
rect 47740 53170 47796 53566
rect 49532 53508 49588 53518
rect 47740 53118 47742 53170
rect 47794 53118 47796 53170
rect 47740 53106 47796 53118
rect 49084 53452 49532 53508
rect 49084 53170 49140 53452
rect 49532 53414 49588 53452
rect 49084 53118 49086 53170
rect 49138 53118 49140 53170
rect 49084 53106 49140 53118
rect 47628 53060 47684 53070
rect 47404 53058 47684 53060
rect 47404 53006 47630 53058
rect 47682 53006 47684 53058
rect 47404 53004 47684 53006
rect 47628 52994 47684 53004
rect 46396 52894 46398 52946
rect 46450 52894 46452 52946
rect 46396 52052 46452 52894
rect 47180 52946 47236 52958
rect 47180 52894 47182 52946
rect 47234 52894 47236 52946
rect 47180 52836 47236 52894
rect 48748 52946 48804 52958
rect 48748 52894 48750 52946
rect 48802 52894 48804 52946
rect 46620 52276 46676 52286
rect 46620 52182 46676 52220
rect 47180 52276 47236 52780
rect 48188 52836 48244 52846
rect 48188 52742 48244 52780
rect 48748 52836 48804 52894
rect 49532 52836 49588 52846
rect 48748 52770 48804 52780
rect 49420 52834 49588 52836
rect 49420 52782 49534 52834
rect 49586 52782 49588 52834
rect 49420 52780 49588 52782
rect 47180 52210 47236 52220
rect 48748 52386 48804 52398
rect 48748 52334 48750 52386
rect 48802 52334 48804 52386
rect 48748 52274 48804 52334
rect 48748 52222 48750 52274
rect 48802 52222 48804 52274
rect 48748 52210 48804 52222
rect 49308 52162 49364 52174
rect 49308 52110 49310 52162
rect 49362 52110 49364 52162
rect 46956 52052 47012 52062
rect 46396 51996 46900 52052
rect 46060 51986 46116 51996
rect 46060 51492 46116 51502
rect 46060 51398 46116 51436
rect 46620 51380 46676 51390
rect 46620 51286 46676 51324
rect 46060 51266 46116 51278
rect 46060 51214 46062 51266
rect 46114 51214 46116 51266
rect 45500 50092 45892 50148
rect 45276 49970 45332 49980
rect 45388 49812 45444 49822
rect 45164 49756 45388 49812
rect 44940 49718 44996 49756
rect 45388 49718 45444 49756
rect 44828 48974 44830 49026
rect 44882 48974 44884 49026
rect 44828 48962 44884 48974
rect 45836 49700 45892 50092
rect 46060 49922 46116 51214
rect 46732 51266 46788 51278
rect 46732 51214 46734 51266
rect 46786 51214 46788 51266
rect 46284 51156 46340 51166
rect 46732 51156 46788 51214
rect 46284 51154 46788 51156
rect 46284 51102 46286 51154
rect 46338 51102 46788 51154
rect 46284 51100 46788 51102
rect 46284 51090 46340 51100
rect 46060 49870 46062 49922
rect 46114 49870 46116 49922
rect 46060 49858 46116 49870
rect 46396 50594 46452 50606
rect 46396 50542 46398 50594
rect 46450 50542 46452 50594
rect 46396 49700 46452 50542
rect 45836 49644 46452 49700
rect 46844 50594 46900 51996
rect 46844 50542 46846 50594
rect 46898 50542 46900 50594
rect 45164 48804 45220 48814
rect 45220 48748 45444 48804
rect 45164 48710 45220 48748
rect 45388 48242 45444 48748
rect 45388 48190 45390 48242
rect 45442 48190 45444 48242
rect 45388 48178 45444 48190
rect 45724 48466 45780 48478
rect 45724 48414 45726 48466
rect 45778 48414 45780 48466
rect 45724 47684 45780 48414
rect 45836 48354 45892 49644
rect 45836 48302 45838 48354
rect 45890 48302 45892 48354
rect 45836 48290 45892 48302
rect 46396 48804 46452 48814
rect 46060 48244 46116 48254
rect 46060 48242 46228 48244
rect 46060 48190 46062 48242
rect 46114 48190 46228 48242
rect 46060 48188 46228 48190
rect 46060 48178 46116 48188
rect 45836 47684 45892 47694
rect 45724 47682 45892 47684
rect 45724 47630 45838 47682
rect 45890 47630 45892 47682
rect 45724 47628 45892 47630
rect 45836 47618 45892 47628
rect 44940 47236 44996 47246
rect 44940 46676 44996 47180
rect 45948 47234 46004 47246
rect 45948 47182 45950 47234
rect 46002 47182 46004 47234
rect 45836 46788 45892 46798
rect 45948 46788 46004 47182
rect 46060 47234 46116 47246
rect 46060 47182 46062 47234
rect 46114 47182 46116 47234
rect 46060 47124 46116 47182
rect 46060 47058 46116 47068
rect 45836 46786 46004 46788
rect 45836 46734 45838 46786
rect 45890 46734 46004 46786
rect 45836 46732 46004 46734
rect 45836 46722 45892 46732
rect 45052 46676 45108 46686
rect 44940 46674 45108 46676
rect 44940 46622 45054 46674
rect 45106 46622 45108 46674
rect 44940 46620 45108 46622
rect 44716 44994 44772 45006
rect 44716 44942 44718 44994
rect 44770 44942 44772 44994
rect 44716 42868 44772 44942
rect 44940 44548 44996 46620
rect 45052 46610 45108 46620
rect 45052 46340 45108 46350
rect 45108 46284 45332 46340
rect 45052 45218 45108 46284
rect 45164 45892 45220 45902
rect 45164 45798 45220 45836
rect 45276 45890 45332 46284
rect 45836 46228 45892 46238
rect 45276 45838 45278 45890
rect 45330 45838 45332 45890
rect 45276 45826 45332 45838
rect 45724 46172 45836 46228
rect 45388 45780 45444 45790
rect 45388 45686 45444 45724
rect 45052 45166 45054 45218
rect 45106 45166 45108 45218
rect 45052 45154 45108 45166
rect 45164 45220 45220 45230
rect 45164 45126 45220 45164
rect 45164 44884 45220 44894
rect 45164 44790 45220 44828
rect 45388 44772 45444 44782
rect 44940 44492 45332 44548
rect 44716 42812 45220 42868
rect 45052 42530 45108 42542
rect 45052 42478 45054 42530
rect 45106 42478 45108 42530
rect 45052 41972 45108 42478
rect 45052 41076 45108 41916
rect 45164 41186 45220 42812
rect 45276 42084 45332 44492
rect 45388 44436 45444 44716
rect 45724 44660 45780 46172
rect 45836 46162 45892 46172
rect 46172 45892 46228 48188
rect 46396 48242 46452 48748
rect 46844 48354 46900 50542
rect 46956 51378 47012 51996
rect 49308 52052 49364 52110
rect 47740 51660 48244 51716
rect 47180 51492 47236 51502
rect 47740 51492 47796 51660
rect 47180 51490 47796 51492
rect 47180 51438 47182 51490
rect 47234 51438 47796 51490
rect 47180 51436 47796 51438
rect 47852 51492 47908 51502
rect 47180 51426 47236 51436
rect 46956 51326 46958 51378
rect 47010 51326 47012 51378
rect 46956 50484 47012 51326
rect 47404 50484 47460 50494
rect 46956 50482 47460 50484
rect 46956 50430 47406 50482
rect 47458 50430 47460 50482
rect 46956 50428 47460 50430
rect 47852 50428 47908 51436
rect 47404 50418 47460 50428
rect 47740 50372 47908 50428
rect 47964 51266 48020 51278
rect 47964 51214 47966 51266
rect 48018 51214 48020 51266
rect 47068 49812 47124 49822
rect 47068 49138 47124 49756
rect 47068 49086 47070 49138
rect 47122 49086 47124 49138
rect 47068 49074 47124 49086
rect 46844 48302 46846 48354
rect 46898 48302 46900 48354
rect 46844 48290 46900 48302
rect 47292 49026 47348 49038
rect 47292 48974 47294 49026
rect 47346 48974 47348 49026
rect 46396 48190 46398 48242
rect 46450 48190 46452 48242
rect 46396 48178 46452 48190
rect 47068 48242 47124 48254
rect 47068 48190 47070 48242
rect 47122 48190 47124 48242
rect 46620 48130 46676 48142
rect 46620 48078 46622 48130
rect 46674 48078 46676 48130
rect 46620 46788 46676 48078
rect 46620 46722 46676 46732
rect 46844 47570 46900 47582
rect 46844 47518 46846 47570
rect 46898 47518 46900 47570
rect 46844 46116 46900 47518
rect 46844 46050 46900 46060
rect 47068 46900 47124 48190
rect 47292 47236 47348 48974
rect 47740 48354 47796 50372
rect 47964 49140 48020 51214
rect 48076 51154 48132 51166
rect 48076 51102 48078 51154
rect 48130 51102 48132 51154
rect 48076 50036 48132 51102
rect 48076 49970 48132 49980
rect 48188 49700 48244 51660
rect 48748 51380 48804 51390
rect 48748 49922 48804 51324
rect 49196 51268 49252 51278
rect 49196 51174 49252 51212
rect 49308 50596 49364 51996
rect 49420 51828 49476 52780
rect 49532 52770 49588 52780
rect 49420 51762 49476 51772
rect 49532 52386 49588 52398
rect 49532 52334 49534 52386
rect 49586 52334 49588 52386
rect 49308 50530 49364 50540
rect 49532 50594 49588 52334
rect 49532 50542 49534 50594
rect 49586 50542 49588 50594
rect 48860 50036 48916 50046
rect 48860 49942 48916 49980
rect 48748 49870 48750 49922
rect 48802 49870 48804 49922
rect 48748 49858 48804 49870
rect 49084 49924 49140 49934
rect 49084 49830 49140 49868
rect 49196 49810 49252 49822
rect 49196 49758 49198 49810
rect 49250 49758 49252 49810
rect 48188 49698 48580 49700
rect 48188 49646 48190 49698
rect 48242 49646 48580 49698
rect 48188 49644 48580 49646
rect 48188 49634 48244 49644
rect 48076 49140 48132 49150
rect 47964 49138 48132 49140
rect 47964 49086 48078 49138
rect 48130 49086 48132 49138
rect 47964 49084 48132 49086
rect 48076 49074 48132 49084
rect 47740 48302 47742 48354
rect 47794 48302 47796 48354
rect 47404 48242 47460 48254
rect 47404 48190 47406 48242
rect 47458 48190 47460 48242
rect 47404 48132 47460 48190
rect 47404 48066 47460 48076
rect 47292 47170 47348 47180
rect 47740 47124 47796 48302
rect 48188 48132 48244 48142
rect 48188 48038 48244 48076
rect 47740 47058 47796 47068
rect 45948 45836 46172 45892
rect 45836 45668 45892 45678
rect 45836 45574 45892 45612
rect 45724 44604 45892 44660
rect 45724 44436 45780 44446
rect 45388 44434 45780 44436
rect 45388 44382 45390 44434
rect 45442 44382 45726 44434
rect 45778 44382 45780 44434
rect 45388 44380 45780 44382
rect 45388 44370 45444 44380
rect 45724 44370 45780 44380
rect 45836 43204 45892 44604
rect 45948 44324 46004 45836
rect 46172 45826 46228 45836
rect 46284 44996 46340 45006
rect 46284 44546 46340 44940
rect 47068 44996 47124 46844
rect 47964 46562 48020 46574
rect 47964 46510 47966 46562
rect 48018 46510 48020 46562
rect 47964 46004 48020 46510
rect 48300 46116 48356 46126
rect 48524 46116 48580 49644
rect 49196 49028 49252 49758
rect 48748 48244 48804 48254
rect 48748 48150 48804 48188
rect 49196 47684 49252 48972
rect 49532 48244 49588 50542
rect 49644 50428 49700 53678
rect 49756 53676 49868 53732
rect 49756 52948 49812 53676
rect 49868 53666 49924 53676
rect 50092 54402 50260 54404
rect 50092 54350 50206 54402
rect 50258 54350 50260 54402
rect 50092 54348 50260 54350
rect 49980 53620 50036 53630
rect 49868 53508 49924 53518
rect 49980 53508 50036 53564
rect 49868 53506 50036 53508
rect 49868 53454 49870 53506
rect 49922 53454 50036 53506
rect 49868 53452 50036 53454
rect 50092 53618 50148 54348
rect 50204 54338 50260 54348
rect 51548 54404 51604 54414
rect 50764 53844 50820 53854
rect 51436 53844 51492 53854
rect 50764 53842 51492 53844
rect 50764 53790 50766 53842
rect 50818 53790 51438 53842
rect 51490 53790 51492 53842
rect 50764 53788 51492 53790
rect 50764 53778 50820 53788
rect 51436 53778 51492 53788
rect 50092 53566 50094 53618
rect 50146 53566 50148 53618
rect 49868 53442 49924 53452
rect 50092 53172 50148 53566
rect 50428 53730 50484 53742
rect 50428 53678 50430 53730
rect 50482 53678 50484 53730
rect 50428 53508 50484 53678
rect 51548 53730 51604 54348
rect 51548 53678 51550 53730
rect 51602 53678 51604 53730
rect 51548 53666 51604 53678
rect 50876 53620 50932 53630
rect 50428 53172 50484 53452
rect 50652 53508 50708 53546
rect 50876 53526 50932 53564
rect 51100 53618 51156 53630
rect 51100 53566 51102 53618
rect 51154 53566 51156 53618
rect 50652 53442 50708 53452
rect 50988 53508 51044 53518
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50988 53172 51044 53452
rect 50428 53116 50708 53172
rect 50092 53106 50148 53116
rect 49756 52882 49812 52892
rect 50540 52948 50596 52958
rect 50428 52834 50484 52846
rect 50428 52782 50430 52834
rect 50482 52782 50484 52834
rect 50428 52388 50484 52782
rect 49980 52332 50484 52388
rect 49756 52162 49812 52174
rect 49756 52110 49758 52162
rect 49810 52110 49812 52162
rect 49756 52052 49812 52110
rect 49756 51986 49812 51996
rect 49980 51938 50036 52332
rect 50316 52164 50372 52174
rect 50316 52070 50372 52108
rect 50540 52052 50596 52892
rect 50652 52164 50708 53116
rect 50876 52948 50932 52958
rect 50876 52854 50932 52892
rect 50988 52500 51044 53116
rect 50876 52444 51044 52500
rect 50652 52098 50708 52108
rect 50764 52162 50820 52174
rect 50764 52110 50766 52162
rect 50818 52110 50820 52162
rect 50428 51996 50596 52052
rect 50764 52052 50820 52110
rect 49980 51886 49982 51938
rect 50034 51886 50036 51938
rect 49980 51828 50036 51886
rect 49980 51762 50036 51772
rect 50092 51938 50148 51950
rect 50092 51886 50094 51938
rect 50146 51886 50148 51938
rect 50092 50708 50148 51886
rect 50092 50642 50148 50652
rect 50204 51938 50260 51950
rect 50204 51886 50206 51938
rect 50258 51886 50260 51938
rect 50204 51828 50260 51886
rect 50204 51268 50260 51772
rect 50204 50484 50260 51212
rect 50428 50706 50484 51996
rect 50764 51986 50820 51996
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50876 51044 50932 52444
rect 51100 52052 51156 53566
rect 51324 52948 51380 52958
rect 51324 52854 51380 52892
rect 51660 52946 51716 52958
rect 51660 52894 51662 52946
rect 51714 52894 51716 52946
rect 51212 52834 51268 52846
rect 51212 52782 51214 52834
rect 51266 52782 51268 52834
rect 51212 52274 51268 52782
rect 51660 52836 51716 52894
rect 52108 52836 52164 54572
rect 53004 54516 53060 54572
rect 53564 54516 53620 54526
rect 53004 54514 53620 54516
rect 53004 54462 53006 54514
rect 53058 54462 53566 54514
rect 53618 54462 53620 54514
rect 53004 54460 53620 54462
rect 53004 54450 53060 54460
rect 53564 54450 53620 54460
rect 52332 54404 52388 54414
rect 52332 54310 52388 54348
rect 52444 52948 52500 52958
rect 52444 52854 52500 52892
rect 51716 52780 52164 52836
rect 54572 52834 54628 52846
rect 54572 52782 54574 52834
rect 54626 52782 54628 52834
rect 51660 52770 51716 52780
rect 51212 52222 51214 52274
rect 51266 52222 51268 52274
rect 51212 52210 51268 52222
rect 51324 52164 51380 52174
rect 51324 52070 51380 52108
rect 51212 52052 51268 52062
rect 51100 52050 51268 52052
rect 51100 51998 51214 52050
rect 51266 51998 51268 52050
rect 51100 51996 51268 51998
rect 50988 51938 51044 51950
rect 50988 51886 50990 51938
rect 51042 51886 51044 51938
rect 50988 51604 51044 51886
rect 50988 51538 51044 51548
rect 50876 50978 50932 50988
rect 50428 50654 50430 50706
rect 50482 50654 50484 50706
rect 50428 50642 50484 50654
rect 50876 50596 50932 50606
rect 51212 50596 51268 51996
rect 51996 51378 52052 52780
rect 53564 52164 53620 52174
rect 52780 51940 52836 51950
rect 53228 51940 53284 51950
rect 52780 51938 53284 51940
rect 52780 51886 52782 51938
rect 52834 51886 53230 51938
rect 53282 51886 53284 51938
rect 52780 51884 53284 51886
rect 52444 51492 52500 51502
rect 52444 51398 52500 51436
rect 52668 51380 52724 51390
rect 51996 51326 51998 51378
rect 52050 51326 52052 51378
rect 51324 51268 51380 51278
rect 51324 51266 51940 51268
rect 51324 51214 51326 51266
rect 51378 51214 51940 51266
rect 51324 51212 51940 51214
rect 51324 51202 51380 51212
rect 50932 50540 51044 50596
rect 50876 50530 50932 50540
rect 50316 50484 50372 50494
rect 50204 50428 50316 50484
rect 49644 50372 49812 50428
rect 50316 50418 50372 50428
rect 49756 49924 49812 50372
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 49756 49830 49812 49868
rect 50764 50034 50820 50046
rect 50764 49982 50766 50034
rect 50818 49982 50820 50034
rect 50204 49138 50260 49150
rect 50204 49086 50206 49138
rect 50258 49086 50260 49138
rect 50204 49028 50260 49086
rect 50764 49140 50820 49982
rect 50764 49074 50820 49084
rect 50204 48962 50260 48972
rect 50876 48916 50932 48926
rect 50876 48822 50932 48860
rect 50540 48804 50596 48814
rect 50428 48802 50596 48804
rect 50428 48750 50542 48802
rect 50594 48750 50596 48802
rect 50428 48748 50596 48750
rect 50428 48468 50484 48748
rect 50540 48738 50596 48748
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 49532 48178 49588 48188
rect 50204 48244 50260 48254
rect 48860 47628 49252 47684
rect 49868 48132 49924 48142
rect 48748 46900 48804 46910
rect 48748 46806 48804 46844
rect 48300 46022 48356 46060
rect 48412 46114 48580 46116
rect 48412 46062 48526 46114
rect 48578 46062 48580 46114
rect 48412 46060 48580 46062
rect 48076 46004 48132 46014
rect 47852 46002 48132 46004
rect 47852 45950 48078 46002
rect 48130 45950 48132 46002
rect 47852 45948 48132 45950
rect 47292 45892 47348 45902
rect 47292 45778 47348 45836
rect 47292 45726 47294 45778
rect 47346 45726 47348 45778
rect 47292 45714 47348 45726
rect 47516 45892 47572 45902
rect 47852 45892 47908 45948
rect 48076 45938 48132 45948
rect 47516 45890 47908 45892
rect 47516 45838 47518 45890
rect 47570 45838 47908 45890
rect 47516 45836 47908 45838
rect 47180 45220 47236 45230
rect 47516 45220 47572 45836
rect 47964 45780 48020 45790
rect 47964 45686 48020 45724
rect 48412 45556 48468 46060
rect 48524 46050 48580 46060
rect 48636 45892 48692 45902
rect 48860 45892 48916 47628
rect 48972 47460 49028 47470
rect 49644 47460 49700 47470
rect 49868 47460 49924 48076
rect 50204 47570 50260 48188
rect 50428 48020 50484 48412
rect 50428 47954 50484 47964
rect 50204 47518 50206 47570
rect 50258 47518 50260 47570
rect 50204 47506 50260 47518
rect 48972 47458 49588 47460
rect 48972 47406 48974 47458
rect 49026 47406 49588 47458
rect 48972 47404 49588 47406
rect 48972 47394 49028 47404
rect 49196 47236 49252 47246
rect 48972 46674 49028 46686
rect 48972 46622 48974 46674
rect 49026 46622 49028 46674
rect 48972 46116 49028 46622
rect 48972 46050 49028 46060
rect 49196 46002 49252 47180
rect 49532 46898 49588 47404
rect 49644 47458 50148 47460
rect 49644 47406 49646 47458
rect 49698 47406 50148 47458
rect 49644 47404 50148 47406
rect 49644 47236 49700 47404
rect 49644 47170 49700 47180
rect 49532 46846 49534 46898
rect 49586 46846 49588 46898
rect 49532 46834 49588 46846
rect 49756 47124 49812 47134
rect 49420 46788 49476 46798
rect 49420 46694 49476 46732
rect 49756 46674 49812 47068
rect 50092 46900 50148 47404
rect 50988 47458 51044 50540
rect 51212 50530 51268 50540
rect 51436 51044 51492 51054
rect 51436 49810 51492 50988
rect 51884 50818 51940 51212
rect 51996 51156 52052 51326
rect 51996 51090 52052 51100
rect 52556 51378 52724 51380
rect 52556 51326 52670 51378
rect 52722 51326 52724 51378
rect 52556 51324 52724 51326
rect 52556 51044 52612 51324
rect 52668 51314 52724 51324
rect 52556 50978 52612 50988
rect 52668 51156 52724 51166
rect 52780 51156 52836 51884
rect 53228 51874 53284 51884
rect 53116 51380 53172 51390
rect 53340 51380 53396 51390
rect 53116 51286 53172 51324
rect 53228 51378 53396 51380
rect 53228 51326 53342 51378
rect 53394 51326 53396 51378
rect 53228 51324 53396 51326
rect 52724 51100 52836 51156
rect 52892 51266 52948 51278
rect 52892 51214 52894 51266
rect 52946 51214 52948 51266
rect 51884 50766 51886 50818
rect 51938 50766 51940 50818
rect 51884 50754 51940 50766
rect 51996 50708 52052 50718
rect 51996 50614 52052 50652
rect 51436 49758 51438 49810
rect 51490 49758 51492 49810
rect 51436 49746 51492 49758
rect 51884 50596 51940 50606
rect 51884 49810 51940 50540
rect 52668 50594 52724 51100
rect 52668 50542 52670 50594
rect 52722 50542 52724 50594
rect 52668 50530 52724 50542
rect 51884 49758 51886 49810
rect 51938 49758 51940 49810
rect 51884 49746 51940 49758
rect 51996 50484 52052 50494
rect 51996 50372 52388 50428
rect 51884 48916 51940 48926
rect 51324 48802 51380 48814
rect 51324 48750 51326 48802
rect 51378 48750 51380 48802
rect 51324 48468 51380 48750
rect 51324 48402 51380 48412
rect 51772 48802 51828 48814
rect 51772 48750 51774 48802
rect 51826 48750 51828 48802
rect 51772 48132 51828 48750
rect 51884 48466 51940 48860
rect 51884 48414 51886 48466
rect 51938 48414 51940 48466
rect 51884 48402 51940 48414
rect 51996 48244 52052 50372
rect 52332 49922 52388 50372
rect 52332 49870 52334 49922
rect 52386 49870 52388 49922
rect 52332 49858 52388 49870
rect 52892 49924 52948 51214
rect 53228 50428 53284 51324
rect 53340 51314 53396 51324
rect 53564 51378 53620 52108
rect 54572 52164 54628 52782
rect 54572 52098 54628 52108
rect 54684 51492 54740 51502
rect 53564 51326 53566 51378
rect 53618 51326 53620 51378
rect 53564 50708 53620 51326
rect 53900 51380 53956 51390
rect 53900 51286 53956 51324
rect 53564 50642 53620 50652
rect 53788 51266 53844 51278
rect 53788 51214 53790 51266
rect 53842 51214 53844 51266
rect 52892 49858 52948 49868
rect 53004 50372 53284 50428
rect 53452 50484 53508 50494
rect 53452 50482 53732 50484
rect 53452 50430 53454 50482
rect 53506 50430 53732 50482
rect 53452 50428 53732 50430
rect 53452 50418 53508 50428
rect 53004 49252 53060 50372
rect 53676 50148 53732 50428
rect 53788 50428 53844 51214
rect 53788 50372 54628 50428
rect 53676 50092 54068 50148
rect 54012 50034 54068 50092
rect 54012 49982 54014 50034
rect 54066 49982 54068 50034
rect 54012 49970 54068 49982
rect 54124 50036 54180 50046
rect 53900 49924 53956 49934
rect 53900 49830 53956 49868
rect 52668 49196 53060 49252
rect 52668 49140 52724 49196
rect 51772 48066 51828 48076
rect 51884 48188 52052 48244
rect 52556 49138 52724 49140
rect 52556 49086 52670 49138
rect 52722 49086 52724 49138
rect 52556 49084 52724 49086
rect 51660 48020 51716 48030
rect 51100 48018 51716 48020
rect 51100 47966 51662 48018
rect 51714 47966 51716 48018
rect 51100 47964 51716 47966
rect 51100 47570 51156 47964
rect 51660 47954 51716 47964
rect 51100 47518 51102 47570
rect 51154 47518 51156 47570
rect 51100 47506 51156 47518
rect 51212 47796 51268 47806
rect 50988 47406 50990 47458
rect 51042 47406 51044 47458
rect 50652 47348 50708 47358
rect 50428 47346 50708 47348
rect 50428 47294 50654 47346
rect 50706 47294 50708 47346
rect 50428 47292 50708 47294
rect 50204 46900 50260 46910
rect 50092 46898 50260 46900
rect 50092 46846 50206 46898
rect 50258 46846 50260 46898
rect 50092 46844 50260 46846
rect 49756 46622 49758 46674
rect 49810 46622 49812 46674
rect 49756 46610 49812 46622
rect 49196 45950 49198 46002
rect 49250 45950 49252 46002
rect 49196 45938 49252 45950
rect 48636 45890 48916 45892
rect 48636 45838 48638 45890
rect 48690 45838 48916 45890
rect 48636 45836 48916 45838
rect 49644 45892 49700 45902
rect 48636 45826 48692 45836
rect 47180 45218 47572 45220
rect 47180 45166 47182 45218
rect 47234 45166 47572 45218
rect 47180 45164 47572 45166
rect 47628 45500 48468 45556
rect 47180 45154 47236 45164
rect 47628 45106 47684 45500
rect 47628 45054 47630 45106
rect 47682 45054 47684 45106
rect 47404 44996 47460 45006
rect 47124 44994 47460 44996
rect 47124 44942 47406 44994
rect 47458 44942 47460 44994
rect 47124 44940 47460 44942
rect 47068 44902 47124 44940
rect 46284 44494 46286 44546
rect 46338 44494 46340 44546
rect 46284 44482 46340 44494
rect 46508 44884 46564 44894
rect 46508 44546 46564 44828
rect 46508 44494 46510 44546
rect 46562 44494 46564 44546
rect 45948 44322 46116 44324
rect 45948 44270 45950 44322
rect 46002 44270 46116 44322
rect 45948 44268 46116 44270
rect 45948 44258 46004 44268
rect 46060 43540 46116 44268
rect 46060 43446 46116 43484
rect 45612 43148 45892 43204
rect 46284 43426 46340 43438
rect 46284 43374 46286 43426
rect 46338 43374 46340 43426
rect 45276 42028 45444 42084
rect 45276 41860 45332 41870
rect 45388 41860 45444 42028
rect 45500 41860 45556 41870
rect 45388 41804 45500 41860
rect 45276 41766 45332 41804
rect 45500 41794 45556 41804
rect 45612 41524 45668 43148
rect 45724 42980 45780 42990
rect 45724 42644 45780 42924
rect 46284 42978 46340 43374
rect 46284 42926 46286 42978
rect 46338 42926 46340 42978
rect 46284 42914 46340 42926
rect 46396 42756 46452 42766
rect 46508 42756 46564 44494
rect 47068 44322 47124 44334
rect 47068 44270 47070 44322
rect 47122 44270 47124 44322
rect 46620 44100 46676 44110
rect 47068 44100 47124 44270
rect 46620 44098 47124 44100
rect 46620 44046 46622 44098
rect 46674 44046 47124 44098
rect 46620 44044 47124 44046
rect 46620 44034 46676 44044
rect 47404 43538 47460 44940
rect 47516 44324 47572 44334
rect 47628 44324 47684 45054
rect 47852 44884 47908 44894
rect 47852 44790 47908 44828
rect 48300 44884 48356 44894
rect 48300 44882 48692 44884
rect 48300 44830 48302 44882
rect 48354 44830 48692 44882
rect 48300 44828 48692 44830
rect 48300 44818 48356 44828
rect 47516 44322 47684 44324
rect 47516 44270 47518 44322
rect 47570 44270 47684 44322
rect 47516 44268 47684 44270
rect 47516 44258 47572 44268
rect 47964 44212 48020 44222
rect 47740 44210 48020 44212
rect 47740 44158 47966 44210
rect 48018 44158 48020 44210
rect 47740 44156 48020 44158
rect 47404 43486 47406 43538
rect 47458 43486 47460 43538
rect 47404 43474 47460 43486
rect 47628 43540 47684 43550
rect 46732 43428 46788 43438
rect 46732 43426 46900 43428
rect 46732 43374 46734 43426
rect 46786 43374 46900 43426
rect 46732 43372 46900 43374
rect 46732 43362 46788 43372
rect 46396 42754 46508 42756
rect 46396 42702 46398 42754
rect 46450 42702 46508 42754
rect 46396 42700 46508 42702
rect 46396 42690 46452 42700
rect 46508 42662 46564 42700
rect 46284 42644 46340 42654
rect 45724 42642 46340 42644
rect 45724 42590 46286 42642
rect 46338 42590 46340 42642
rect 45724 42588 46340 42590
rect 45724 42194 45780 42588
rect 46284 42578 46340 42588
rect 45724 42142 45726 42194
rect 45778 42142 45780 42194
rect 45724 42130 45780 42142
rect 46060 41970 46116 41982
rect 46060 41918 46062 41970
rect 46114 41918 46116 41970
rect 45612 41458 45668 41468
rect 45836 41636 45892 41646
rect 45164 41134 45166 41186
rect 45218 41134 45220 41186
rect 45164 41122 45220 41134
rect 45836 41188 45892 41580
rect 45052 41010 45108 41020
rect 45276 41076 45332 41086
rect 45276 40982 45332 41020
rect 45500 40964 45556 40974
rect 45388 40962 45556 40964
rect 45388 40910 45502 40962
rect 45554 40910 45556 40962
rect 45388 40908 45556 40910
rect 44940 40404 44996 40414
rect 44604 40114 44660 40124
rect 44828 40290 44884 40302
rect 44828 40238 44830 40290
rect 44882 40238 44884 40290
rect 44268 39678 44270 39730
rect 44322 39678 44324 39730
rect 44268 39666 44324 39678
rect 44828 39620 44884 40238
rect 44940 39732 44996 40348
rect 45276 40404 45332 40414
rect 45276 40310 45332 40348
rect 45388 40180 45444 40908
rect 45500 40898 45556 40908
rect 45612 40964 45668 40974
rect 45276 40124 45444 40180
rect 44940 39730 45108 39732
rect 44940 39678 44942 39730
rect 44994 39678 45108 39730
rect 44940 39676 45108 39678
rect 44940 39666 44996 39676
rect 44828 39554 44884 39564
rect 43820 39006 43822 39058
rect 43874 39006 43876 39058
rect 43820 38994 43876 39006
rect 44268 38836 44324 38846
rect 44156 38724 44212 38762
rect 44156 38658 44212 38668
rect 44156 38164 44212 38174
rect 44268 38164 44324 38780
rect 44156 38162 44324 38164
rect 44156 38110 44158 38162
rect 44210 38110 44324 38162
rect 44156 38108 44324 38110
rect 45052 38162 45108 39676
rect 45276 39618 45332 40124
rect 45612 39956 45668 40908
rect 45836 40516 45892 41132
rect 45948 40964 46004 40974
rect 46060 40964 46116 41918
rect 46508 41860 46564 41870
rect 46396 40964 46452 40974
rect 46060 40962 46452 40964
rect 46060 40910 46398 40962
rect 46450 40910 46452 40962
rect 46060 40908 46452 40910
rect 45948 40870 46004 40908
rect 46396 40740 46452 40908
rect 46396 40674 46452 40684
rect 46508 40516 46564 41804
rect 45836 40460 46116 40516
rect 45948 40292 46004 40302
rect 45276 39566 45278 39618
rect 45330 39566 45332 39618
rect 45276 39554 45332 39566
rect 45388 39900 45668 39956
rect 45724 40290 46004 40292
rect 45724 40238 45950 40290
rect 46002 40238 46004 40290
rect 45724 40236 46004 40238
rect 45052 38110 45054 38162
rect 45106 38110 45108 38162
rect 44156 38098 44212 38108
rect 45052 38098 45108 38110
rect 45388 37154 45444 39900
rect 45724 39730 45780 40236
rect 45948 40226 46004 40236
rect 45724 39678 45726 39730
rect 45778 39678 45780 39730
rect 45724 39666 45780 39678
rect 45836 39620 45892 39630
rect 46060 39620 46116 40460
rect 46508 40450 46564 40460
rect 46732 41860 46788 41870
rect 46732 41074 46788 41804
rect 46732 41022 46734 41074
rect 46786 41022 46788 41074
rect 45836 39526 45892 39564
rect 45948 39564 46116 39620
rect 45612 39396 45668 39406
rect 45948 39396 46004 39564
rect 45612 39394 46004 39396
rect 45612 39342 45614 39394
rect 45666 39342 46004 39394
rect 45612 39340 46004 39342
rect 45612 39330 45668 39340
rect 45500 38948 45556 38958
rect 45500 38854 45556 38892
rect 45836 38834 45892 38846
rect 45836 38782 45838 38834
rect 45890 38782 45892 38834
rect 45388 37102 45390 37154
rect 45442 37102 45444 37154
rect 45276 36484 45332 36494
rect 45388 36484 45444 37102
rect 45276 36482 45444 36484
rect 45276 36430 45278 36482
rect 45330 36430 45444 36482
rect 45276 36428 45444 36430
rect 45500 38724 45556 38734
rect 45500 36484 45556 38668
rect 45836 37492 45892 38782
rect 46508 38722 46564 38734
rect 46508 38670 46510 38722
rect 46562 38670 46564 38722
rect 46508 38668 46564 38670
rect 45836 37398 45892 37436
rect 46172 38612 46564 38668
rect 46620 38612 46676 38622
rect 46172 37490 46228 38612
rect 46620 38518 46676 38556
rect 46620 38052 46676 38062
rect 46620 37958 46676 37996
rect 46172 37438 46174 37490
rect 46226 37438 46228 37490
rect 46172 37426 46228 37438
rect 46284 37938 46340 37950
rect 46284 37886 46286 37938
rect 46338 37886 46340 37938
rect 46284 37380 46340 37886
rect 46284 37286 46340 37324
rect 46396 37826 46452 37838
rect 46396 37774 46398 37826
rect 46450 37774 46452 37826
rect 46060 37268 46116 37278
rect 45724 36484 45780 36494
rect 45500 36482 45668 36484
rect 45500 36430 45502 36482
rect 45554 36430 45668 36482
rect 45500 36428 45668 36430
rect 43708 36194 43764 36204
rect 44940 36260 44996 36270
rect 44940 36166 44996 36204
rect 45276 35812 45332 36428
rect 45500 36418 45556 36428
rect 45276 35746 45332 35756
rect 45500 35924 45556 35934
rect 43260 35364 43316 35374
rect 43260 34354 43316 35308
rect 43484 35140 43540 35644
rect 45500 35586 45556 35868
rect 45500 35534 45502 35586
rect 45554 35534 45556 35586
rect 45500 35522 45556 35534
rect 45612 35476 45668 36428
rect 45724 36482 45892 36484
rect 45724 36430 45726 36482
rect 45778 36430 45892 36482
rect 45724 36428 45892 36430
rect 45724 36418 45780 36428
rect 45836 36260 45892 36428
rect 45724 35476 45780 35486
rect 45612 35474 45780 35476
rect 45612 35422 45726 35474
rect 45778 35422 45780 35474
rect 45612 35420 45780 35422
rect 45724 35410 45780 35420
rect 43484 35074 43540 35084
rect 44940 35140 44996 35150
rect 44940 35026 44996 35084
rect 44940 34974 44942 35026
rect 44994 34974 44996 35026
rect 44940 34962 44996 34974
rect 43484 34916 43540 34926
rect 43484 34914 43652 34916
rect 43484 34862 43486 34914
rect 43538 34862 43652 34914
rect 43484 34860 43652 34862
rect 43484 34850 43540 34860
rect 43260 34302 43262 34354
rect 43314 34302 43316 34354
rect 43260 34290 43316 34302
rect 43036 34130 43204 34132
rect 43036 34078 43038 34130
rect 43090 34078 43204 34130
rect 43036 34076 43204 34078
rect 43036 33570 43092 34076
rect 43596 33684 43652 34860
rect 44044 34692 44100 34702
rect 44044 34598 44100 34636
rect 45836 34580 45892 36204
rect 46060 36148 46116 37212
rect 46396 37268 46452 37774
rect 46396 37202 46452 37212
rect 46508 37380 46564 37390
rect 46172 36260 46228 36270
rect 46172 36166 46228 36204
rect 45948 35588 46004 35598
rect 45948 35494 46004 35532
rect 45836 34514 45892 34524
rect 45948 34692 46004 34702
rect 45388 34242 45444 34254
rect 45388 34190 45390 34242
rect 45442 34190 45444 34242
rect 43708 34020 43764 34030
rect 43708 33926 43764 33964
rect 44828 33908 44884 33918
rect 44044 33906 44884 33908
rect 44044 33854 44830 33906
rect 44882 33854 44884 33906
rect 44044 33852 44884 33854
rect 43596 33628 43764 33684
rect 43036 33518 43038 33570
rect 43090 33518 43092 33570
rect 43036 33506 43092 33518
rect 43036 33348 43092 33358
rect 42924 33346 43092 33348
rect 42924 33294 43038 33346
rect 43090 33294 43092 33346
rect 42924 33292 43092 33294
rect 43036 33282 43092 33292
rect 42812 32498 42868 32508
rect 42476 32452 42532 32462
rect 42252 32450 42532 32452
rect 42252 32398 42478 32450
rect 42530 32398 42532 32450
rect 42252 32396 42532 32398
rect 42140 32340 42196 32350
rect 42028 32284 42140 32340
rect 42140 32274 42196 32284
rect 41468 32228 41524 32238
rect 41468 31778 41524 32172
rect 42140 32004 42196 32014
rect 42252 32004 42308 32396
rect 42476 32386 42532 32396
rect 42140 32002 42308 32004
rect 42140 31950 42142 32002
rect 42194 31950 42308 32002
rect 42140 31948 42308 31950
rect 42140 31938 42196 31948
rect 41580 31892 41636 31902
rect 42028 31892 42084 31902
rect 41580 31890 42084 31892
rect 41580 31838 41582 31890
rect 41634 31838 42030 31890
rect 42082 31838 42084 31890
rect 41580 31836 42084 31838
rect 41580 31826 41636 31836
rect 42028 31826 42084 31836
rect 43596 31892 43652 31902
rect 41468 31726 41470 31778
rect 41522 31726 41524 31778
rect 41468 31714 41524 31726
rect 41580 31554 41636 31566
rect 41580 31502 41582 31554
rect 41634 31502 41636 31554
rect 41580 31220 41636 31502
rect 42700 31554 42756 31566
rect 42700 31502 42702 31554
rect 42754 31502 42756 31554
rect 41692 31220 41748 31230
rect 41580 31164 41692 31220
rect 41692 31154 41748 31164
rect 42700 31220 42756 31502
rect 43148 31556 43204 31566
rect 43148 31462 43204 31500
rect 43596 31444 43652 31836
rect 43596 31378 43652 31388
rect 42700 31154 42756 31164
rect 43036 30884 43092 30894
rect 43036 30790 43092 30828
rect 43708 30548 43764 33628
rect 44044 33346 44100 33852
rect 44828 33842 44884 33852
rect 45164 33906 45220 33918
rect 45164 33854 45166 33906
rect 45218 33854 45220 33906
rect 44044 33294 44046 33346
rect 44098 33294 44100 33346
rect 44044 33282 44100 33294
rect 44940 33348 44996 33358
rect 44940 33346 45108 33348
rect 44940 33294 44942 33346
rect 44994 33294 45108 33346
rect 44940 33292 45108 33294
rect 44940 33282 44996 33292
rect 44268 33236 44324 33246
rect 44268 33142 44324 33180
rect 45052 32564 45108 33292
rect 45052 32470 45108 32508
rect 44604 32450 44660 32462
rect 44604 32398 44606 32450
rect 44658 32398 44660 32450
rect 44604 32228 44660 32398
rect 44604 32162 44660 32172
rect 44156 31556 44212 31566
rect 44156 31462 44212 31500
rect 44604 31108 44660 31118
rect 44604 31014 44660 31052
rect 43820 30994 43876 31006
rect 43820 30942 43822 30994
rect 43874 30942 43876 30994
rect 43820 30884 43876 30942
rect 44380 30996 44436 31006
rect 44380 30994 44548 30996
rect 44380 30942 44382 30994
rect 44434 30942 44548 30994
rect 44380 30940 44548 30942
rect 44380 30930 44436 30940
rect 44044 30884 44100 30894
rect 43820 30828 44044 30884
rect 43708 30482 43764 30492
rect 44044 30322 44100 30828
rect 44492 30548 44548 30940
rect 45052 30994 45108 31006
rect 45052 30942 45054 30994
rect 45106 30942 45108 30994
rect 45052 30884 45108 30942
rect 45052 30818 45108 30828
rect 44492 30492 44996 30548
rect 44940 30434 44996 30492
rect 44940 30382 44942 30434
rect 44994 30382 44996 30434
rect 44940 30370 44996 30382
rect 44044 30270 44046 30322
rect 44098 30270 44100 30322
rect 44044 30258 44100 30270
rect 44380 30100 44436 30110
rect 41916 29652 41972 29662
rect 41468 29314 41524 29326
rect 41468 29262 41470 29314
rect 41522 29262 41524 29314
rect 41468 29092 41524 29262
rect 41468 29026 41524 29036
rect 41916 28644 41972 29596
rect 43260 29538 43316 29550
rect 43260 29486 43262 29538
rect 43314 29486 43316 29538
rect 42700 29428 42756 29438
rect 42700 29334 42756 29372
rect 43036 29428 43092 29438
rect 43036 29426 43204 29428
rect 43036 29374 43038 29426
rect 43090 29374 43204 29426
rect 43036 29372 43204 29374
rect 43036 29362 43092 29372
rect 42476 29316 42532 29326
rect 42476 28980 42532 29260
rect 42476 28914 42532 28924
rect 42588 29204 42644 29214
rect 41804 28642 41972 28644
rect 41804 28590 41918 28642
rect 41970 28590 41972 28642
rect 41804 28588 41972 28590
rect 41804 28308 41860 28588
rect 41916 28578 41972 28588
rect 42252 28754 42308 28766
rect 42252 28702 42254 28754
rect 42306 28702 42308 28754
rect 41580 28252 41860 28308
rect 41132 27134 41134 27186
rect 41186 27134 41188 27186
rect 41132 27122 41188 27134
rect 41244 28028 41412 28084
rect 41468 28084 41524 28094
rect 40908 27022 40910 27074
rect 40962 27022 40964 27074
rect 40908 27010 40964 27022
rect 40348 26852 40516 26908
rect 40348 26178 40404 26190
rect 40348 26126 40350 26178
rect 40402 26126 40404 26178
rect 40348 25956 40404 26126
rect 40348 25890 40404 25900
rect 40236 25396 40292 25406
rect 40236 25302 40292 25340
rect 40348 25282 40404 25294
rect 40348 25230 40350 25282
rect 40402 25230 40404 25282
rect 40236 24948 40292 24958
rect 40124 24946 40292 24948
rect 40124 24894 40238 24946
rect 40290 24894 40292 24946
rect 40124 24892 40292 24894
rect 40236 24882 40292 24892
rect 40348 24724 40404 25230
rect 40348 24658 40404 24668
rect 39564 24498 39620 24510
rect 39564 24446 39566 24498
rect 39618 24446 39620 24498
rect 39564 24388 39620 24446
rect 39788 24500 39844 24510
rect 39844 24444 39956 24500
rect 39788 24406 39844 24444
rect 39564 23828 39620 24332
rect 39788 24162 39844 24174
rect 39788 24110 39790 24162
rect 39842 24110 39844 24162
rect 39788 24050 39844 24110
rect 39900 24162 39956 24444
rect 39900 24110 39902 24162
rect 39954 24110 39956 24162
rect 39900 24098 39956 24110
rect 39788 23998 39790 24050
rect 39842 23998 39844 24050
rect 39788 23986 39844 23998
rect 40348 24052 40404 24062
rect 40348 23958 40404 23996
rect 39564 23762 39620 23772
rect 40460 23716 40516 26852
rect 40684 26852 40852 26908
rect 41244 26908 41300 28028
rect 41356 27860 41412 27870
rect 41356 27766 41412 27804
rect 41468 27636 41524 28028
rect 41580 27858 41636 28252
rect 41580 27806 41582 27858
rect 41634 27806 41636 27858
rect 41580 27794 41636 27806
rect 41804 28084 41860 28094
rect 41804 27858 41860 28028
rect 42252 28082 42308 28702
rect 42588 28642 42644 29148
rect 42588 28590 42590 28642
rect 42642 28590 42644 28642
rect 42588 28578 42644 28590
rect 43036 28980 43092 28990
rect 43148 28980 43204 29372
rect 43260 29316 43316 29486
rect 43708 29540 43764 29550
rect 43708 29446 43764 29484
rect 44156 29540 44212 29550
rect 43372 29428 43428 29438
rect 43372 29334 43428 29372
rect 44156 29426 44212 29484
rect 44380 29538 44436 30044
rect 44380 29486 44382 29538
rect 44434 29486 44436 29538
rect 44380 29474 44436 29486
rect 44156 29374 44158 29426
rect 44210 29374 44212 29426
rect 44156 29362 44212 29374
rect 43260 29250 43316 29260
rect 43820 29316 43876 29326
rect 43148 28924 43540 28980
rect 42252 28030 42254 28082
rect 42306 28030 42308 28082
rect 42252 28018 42308 28030
rect 42364 28084 42420 28094
rect 42364 27990 42420 28028
rect 43036 28084 43092 28924
rect 43260 28644 43316 28654
rect 43260 28550 43316 28588
rect 43484 28642 43540 28924
rect 43484 28590 43486 28642
rect 43538 28590 43540 28642
rect 43484 28578 43540 28590
rect 43596 28644 43652 28654
rect 43596 28532 43652 28588
rect 43708 28532 43764 28542
rect 43596 28476 43708 28532
rect 43708 28438 43764 28476
rect 43820 28530 43876 29260
rect 44940 29204 44996 29214
rect 44940 29110 44996 29148
rect 44268 28980 44324 28990
rect 43820 28478 43822 28530
rect 43874 28478 43876 28530
rect 43820 28466 43876 28478
rect 43932 28868 43988 28878
rect 43484 28308 43540 28318
rect 43148 28084 43204 28094
rect 43092 28082 43204 28084
rect 43092 28030 43150 28082
rect 43202 28030 43204 28082
rect 43092 28028 43204 28030
rect 43036 27990 43092 28028
rect 43148 28018 43204 28028
rect 42588 27972 42644 27982
rect 42644 27916 42756 27972
rect 42588 27878 42644 27916
rect 41804 27806 41806 27858
rect 41858 27806 41860 27858
rect 41356 27580 41524 27636
rect 41356 27074 41412 27580
rect 41356 27022 41358 27074
rect 41410 27022 41412 27074
rect 41356 27010 41412 27022
rect 41468 27076 41524 27086
rect 41468 26982 41524 27020
rect 41244 26852 41748 26908
rect 40684 26850 40740 26852
rect 40684 26798 40686 26850
rect 40738 26798 40740 26850
rect 40572 25508 40628 25518
rect 40572 25414 40628 25452
rect 40684 24612 40740 26798
rect 41132 26178 41188 26190
rect 41132 26126 41134 26178
rect 41186 26126 41188 26178
rect 41132 25844 41188 26126
rect 41468 25956 41524 25966
rect 41524 25900 41636 25956
rect 41468 25890 41524 25900
rect 41132 25778 41188 25788
rect 41468 25508 41524 25518
rect 41244 25506 41524 25508
rect 41244 25454 41470 25506
rect 41522 25454 41524 25506
rect 41244 25452 41524 25454
rect 40684 24546 40740 24556
rect 40796 25394 40852 25406
rect 40796 25342 40798 25394
rect 40850 25342 40852 25394
rect 40572 24500 40628 24510
rect 40572 24162 40628 24444
rect 40572 24110 40574 24162
rect 40626 24110 40628 24162
rect 40572 24098 40628 24110
rect 40796 24164 40852 25342
rect 40908 25282 40964 25294
rect 40908 25230 40910 25282
rect 40962 25230 40964 25282
rect 40908 24724 40964 25230
rect 41244 24946 41300 25452
rect 41468 25442 41524 25452
rect 41244 24894 41246 24946
rect 41298 24894 41300 24946
rect 41244 24882 41300 24894
rect 41020 24836 41076 24846
rect 41020 24742 41076 24780
rect 40908 24630 40964 24668
rect 41356 24164 41412 24174
rect 40796 24162 41412 24164
rect 40796 24110 41358 24162
rect 41410 24110 41412 24162
rect 40796 24108 41412 24110
rect 41356 24098 41412 24108
rect 40796 23940 40852 23950
rect 41468 23940 41524 23950
rect 40796 23938 40964 23940
rect 40796 23886 40798 23938
rect 40850 23886 40964 23938
rect 40796 23884 40964 23886
rect 40796 23874 40852 23884
rect 40460 23660 40852 23716
rect 40236 23156 40292 23166
rect 40236 23062 40292 23100
rect 39788 23044 39844 23054
rect 39788 23042 39956 23044
rect 39788 22990 39790 23042
rect 39842 22990 39956 23042
rect 39788 22988 39956 22990
rect 39788 22978 39844 22988
rect 39452 22530 39508 22540
rect 39116 22260 39172 22270
rect 39452 22260 39508 22270
rect 39004 22258 39508 22260
rect 39004 22206 39118 22258
rect 39170 22206 39454 22258
rect 39506 22206 39508 22258
rect 39004 22204 39508 22206
rect 38892 22166 38948 22204
rect 39116 22194 39172 22204
rect 39452 22194 39508 22204
rect 39564 22260 39620 22270
rect 39564 21698 39620 22204
rect 39788 22260 39844 22270
rect 39788 22166 39844 22204
rect 39564 21646 39566 21698
rect 39618 21646 39620 21698
rect 39564 21634 39620 21646
rect 39900 21700 39956 22988
rect 40460 22820 40516 22830
rect 40348 22764 40460 22820
rect 40236 22484 40292 22494
rect 40124 22428 40236 22484
rect 40012 21812 40068 21822
rect 40124 21812 40180 22428
rect 40236 22418 40292 22428
rect 40236 22260 40292 22270
rect 40348 22260 40404 22764
rect 40460 22754 40516 22764
rect 40684 22484 40740 22494
rect 40684 22390 40740 22428
rect 40292 22204 40404 22260
rect 40236 22166 40292 22204
rect 40684 21924 40740 21934
rect 40236 21812 40292 21822
rect 40124 21810 40292 21812
rect 40124 21758 40238 21810
rect 40290 21758 40292 21810
rect 40124 21756 40292 21758
rect 40012 21718 40068 21756
rect 40236 21746 40292 21756
rect 39900 21634 39956 21644
rect 38892 21588 38948 21598
rect 38892 21494 38948 21532
rect 39116 21586 39172 21598
rect 39116 21534 39118 21586
rect 39170 21534 39172 21586
rect 38556 20190 38558 20242
rect 38610 20190 38612 20242
rect 38556 20178 38612 20190
rect 38668 21084 38836 21140
rect 39004 21476 39060 21486
rect 38668 19796 38724 21084
rect 38780 20914 38836 20926
rect 38780 20862 38782 20914
rect 38834 20862 38836 20914
rect 38780 20244 38836 20862
rect 39004 20802 39060 21420
rect 39004 20750 39006 20802
rect 39058 20750 39060 20802
rect 39004 20468 39060 20750
rect 39004 20402 39060 20412
rect 39116 20580 39172 21534
rect 39788 21588 39844 21598
rect 39340 21474 39396 21486
rect 39340 21422 39342 21474
rect 39394 21422 39396 21474
rect 39340 20692 39396 21422
rect 39340 20626 39396 20636
rect 39564 20692 39620 20702
rect 39564 20690 39732 20692
rect 39564 20638 39566 20690
rect 39618 20638 39732 20690
rect 39564 20636 39732 20638
rect 39564 20626 39620 20636
rect 38892 20244 38948 20254
rect 38780 20242 38948 20244
rect 38780 20190 38894 20242
rect 38946 20190 38948 20242
rect 38780 20188 38948 20190
rect 38892 20178 38948 20188
rect 39004 20244 39060 20254
rect 39116 20244 39172 20524
rect 39340 20468 39396 20478
rect 39004 20242 39284 20244
rect 39004 20190 39006 20242
rect 39058 20190 39284 20242
rect 39004 20188 39284 20190
rect 39004 20178 39060 20188
rect 38668 19730 38724 19740
rect 38780 20018 38836 20030
rect 38780 19966 38782 20018
rect 38834 19966 38836 20018
rect 38780 19684 38836 19966
rect 39228 20018 39284 20188
rect 39228 19966 39230 20018
rect 39282 19966 39284 20018
rect 39228 19954 39284 19966
rect 39116 19684 39172 19694
rect 38780 19628 39116 19684
rect 38556 19348 38612 19358
rect 38556 19254 38612 19292
rect 39116 19346 39172 19628
rect 39340 19458 39396 20412
rect 39340 19406 39342 19458
rect 39394 19406 39396 19458
rect 39340 19394 39396 19406
rect 39452 20356 39508 20366
rect 39116 19294 39118 19346
rect 39170 19294 39172 19346
rect 39116 19282 39172 19294
rect 38556 19012 38612 19022
rect 38444 18956 38556 19012
rect 39452 19012 39508 20300
rect 39564 20018 39620 20030
rect 39564 19966 39566 20018
rect 39618 19966 39620 20018
rect 39564 19796 39620 19966
rect 39676 19908 39732 20636
rect 39676 19842 39732 19852
rect 39788 20130 39844 21532
rect 40348 21586 40404 21598
rect 40348 21534 40350 21586
rect 40402 21534 40404 21586
rect 40348 20916 40404 21534
rect 40348 20850 40404 20860
rect 40460 20914 40516 20926
rect 40460 20862 40462 20914
rect 40514 20862 40516 20914
rect 40460 20804 40516 20862
rect 40012 20748 40292 20804
rect 39900 20690 39956 20702
rect 39900 20638 39902 20690
rect 39954 20638 39956 20690
rect 39900 20356 39956 20638
rect 39900 20290 39956 20300
rect 39788 20078 39790 20130
rect 39842 20078 39844 20130
rect 39564 19730 39620 19740
rect 39788 19796 39844 20078
rect 39900 20132 39956 20142
rect 40012 20132 40068 20748
rect 40236 20692 40292 20748
rect 40460 20738 40516 20748
rect 40572 20802 40628 20814
rect 40572 20750 40574 20802
rect 40626 20750 40628 20802
rect 40348 20692 40404 20702
rect 40236 20690 40404 20692
rect 40236 20638 40350 20690
rect 40402 20638 40404 20690
rect 40236 20636 40404 20638
rect 40348 20626 40404 20636
rect 39900 20130 40068 20132
rect 39900 20078 39902 20130
rect 39954 20078 40068 20130
rect 39900 20076 40068 20078
rect 40124 20578 40180 20590
rect 40124 20526 40126 20578
rect 40178 20526 40180 20578
rect 39900 20066 39956 20076
rect 39788 19730 39844 19740
rect 40012 19458 40068 19470
rect 40012 19406 40014 19458
rect 40066 19406 40068 19458
rect 39564 19012 39620 19022
rect 39452 19010 39620 19012
rect 39452 18958 39566 19010
rect 39618 18958 39620 19010
rect 39452 18956 39620 18958
rect 38556 18946 38612 18956
rect 39564 18900 39620 18956
rect 39564 18834 39620 18844
rect 40012 19010 40068 19406
rect 40012 18958 40014 19010
rect 40066 18958 40068 19010
rect 39900 18676 39956 18686
rect 39564 18674 39956 18676
rect 39564 18622 39902 18674
rect 39954 18622 39956 18674
rect 39564 18620 39956 18622
rect 38220 18564 38276 18574
rect 37996 18562 38276 18564
rect 37996 18510 38222 18562
rect 38274 18510 38276 18562
rect 37996 18508 38276 18510
rect 37772 17444 37828 18508
rect 37884 18498 37940 18508
rect 38220 18498 38276 18508
rect 38332 18562 38388 18574
rect 38332 18510 38334 18562
rect 38386 18510 38388 18562
rect 38332 17892 38388 18510
rect 38556 18452 38612 18462
rect 38556 18358 38612 18396
rect 39228 18452 39284 18462
rect 39228 18358 39284 18396
rect 38108 17836 38388 17892
rect 37884 17668 37940 17678
rect 37884 17574 37940 17612
rect 37996 17444 38052 17454
rect 38108 17444 38164 17836
rect 38220 17668 38276 17678
rect 38556 17668 38612 17678
rect 39228 17668 39284 17678
rect 39564 17668 39620 18620
rect 39900 18610 39956 18620
rect 39676 18452 39732 18462
rect 40012 18452 40068 18958
rect 40124 18676 40180 20526
rect 40572 20580 40628 20750
rect 40572 20514 40628 20524
rect 40236 19906 40292 19918
rect 40236 19854 40238 19906
rect 40290 19854 40292 19906
rect 40236 19796 40292 19854
rect 40236 19012 40292 19740
rect 40460 19012 40516 19022
rect 40236 19010 40516 19012
rect 40236 18958 40462 19010
rect 40514 18958 40516 19010
rect 40236 18956 40516 18958
rect 40124 18610 40180 18620
rect 39676 18358 39732 18396
rect 39900 18396 40068 18452
rect 40348 18452 40404 18462
rect 39788 18338 39844 18350
rect 39788 18286 39790 18338
rect 39842 18286 39844 18338
rect 39788 18004 39844 18286
rect 39788 17938 39844 17948
rect 38220 17666 38612 17668
rect 38220 17614 38222 17666
rect 38274 17614 38558 17666
rect 38610 17614 38612 17666
rect 38220 17612 38612 17614
rect 38220 17602 38276 17612
rect 38556 17602 38612 17612
rect 38892 17666 39620 17668
rect 38892 17614 39230 17666
rect 39282 17614 39620 17666
rect 38892 17612 39620 17614
rect 39676 17668 39732 17678
rect 37772 17442 38164 17444
rect 37772 17390 37998 17442
rect 38050 17390 38164 17442
rect 37772 17388 38164 17390
rect 37660 15822 37662 15874
rect 37714 15822 37716 15874
rect 37660 15540 37716 15822
rect 37772 17108 37828 17118
rect 37772 15764 37828 17052
rect 37996 16772 38052 17388
rect 37996 16706 38052 16716
rect 38220 16436 38276 16446
rect 38220 16210 38276 16380
rect 38220 16158 38222 16210
rect 38274 16158 38276 16210
rect 38220 16146 38276 16158
rect 38108 16100 38164 16110
rect 37884 15988 37940 15998
rect 37884 15894 37940 15932
rect 37772 15708 37940 15764
rect 37660 15484 37828 15540
rect 37772 15148 37828 15484
rect 37660 15092 37828 15148
rect 37660 14530 37716 15092
rect 37660 14478 37662 14530
rect 37714 14478 37716 14530
rect 37660 14466 37716 14478
rect 37884 14530 37940 15708
rect 38108 15652 38164 16044
rect 38892 15652 38948 17612
rect 39228 17602 39284 17612
rect 39004 17442 39060 17454
rect 39004 17390 39006 17442
rect 39058 17390 39060 17442
rect 39004 16996 39060 17390
rect 39116 17444 39172 17454
rect 39116 17442 39396 17444
rect 39116 17390 39118 17442
rect 39170 17390 39396 17442
rect 39116 17388 39396 17390
rect 39116 17378 39172 17388
rect 39004 16930 39060 16940
rect 39116 16884 39172 16894
rect 39116 16098 39172 16828
rect 39116 16046 39118 16098
rect 39170 16046 39172 16098
rect 39116 16034 39172 16046
rect 39228 16772 39284 16782
rect 38108 15540 38164 15596
rect 38332 15596 38724 15652
rect 38220 15540 38276 15550
rect 38108 15538 38276 15540
rect 38108 15486 38222 15538
rect 38274 15486 38276 15538
rect 38108 15484 38276 15486
rect 38220 15474 38276 15484
rect 38332 15538 38388 15596
rect 38332 15486 38334 15538
rect 38386 15486 38388 15538
rect 38332 15474 38388 15486
rect 38444 15426 38500 15438
rect 38444 15374 38446 15426
rect 38498 15374 38500 15426
rect 38220 15316 38276 15326
rect 37884 14478 37886 14530
rect 37938 14478 37940 14530
rect 37884 14466 37940 14478
rect 37996 14980 38052 14990
rect 37548 14242 37604 14252
rect 37884 14084 37940 14094
rect 37660 13972 37716 13982
rect 37436 13970 37716 13972
rect 37436 13918 37662 13970
rect 37714 13918 37716 13970
rect 37436 13916 37716 13918
rect 37660 13906 37716 13916
rect 37772 13972 37828 13982
rect 37772 13878 37828 13916
rect 37884 13970 37940 14028
rect 37884 13918 37886 13970
rect 37938 13918 37940 13970
rect 37324 13748 37380 13758
rect 37884 13748 37940 13918
rect 37324 13746 37940 13748
rect 37324 13694 37326 13746
rect 37378 13694 37940 13746
rect 37324 13692 37940 13694
rect 37324 13682 37380 13692
rect 37100 13132 37492 13188
rect 37100 12290 37156 13132
rect 37436 13076 37492 13132
rect 37436 13074 37716 13076
rect 37436 13022 37438 13074
rect 37490 13022 37716 13074
rect 37436 13020 37716 13022
rect 37436 13010 37492 13020
rect 37100 12238 37102 12290
rect 37154 12238 37156 12290
rect 37100 12226 37156 12238
rect 36764 12178 36820 12190
rect 37548 12180 37604 12190
rect 36764 12126 36766 12178
rect 36818 12126 36820 12178
rect 36764 11844 36820 12126
rect 37324 12124 37548 12180
rect 37212 11954 37268 11966
rect 37212 11902 37214 11954
rect 37266 11902 37268 11954
rect 37212 11844 37268 11902
rect 36764 11788 37268 11844
rect 37100 11396 37156 11406
rect 37100 11302 37156 11340
rect 37212 11282 37268 11788
rect 37212 11230 37214 11282
rect 37266 11230 37268 11282
rect 37212 11218 37268 11230
rect 36988 10836 37044 10846
rect 36988 10722 37044 10780
rect 37324 10836 37380 12124
rect 37548 12114 37604 12124
rect 37324 10834 37492 10836
rect 37324 10782 37326 10834
rect 37378 10782 37492 10834
rect 37324 10780 37492 10782
rect 37324 10770 37380 10780
rect 36988 10670 36990 10722
rect 37042 10670 37044 10722
rect 36988 10276 37044 10670
rect 37100 10722 37156 10734
rect 37100 10670 37102 10722
rect 37154 10670 37156 10722
rect 37100 10500 37156 10670
rect 37100 10434 37156 10444
rect 37324 10612 37380 10622
rect 36988 10220 37268 10276
rect 37212 9938 37268 10220
rect 37212 9886 37214 9938
rect 37266 9886 37268 9938
rect 37212 9874 37268 9886
rect 37324 9716 37380 10556
rect 37436 9828 37492 10780
rect 37660 10612 37716 13020
rect 37772 12740 37828 12750
rect 37772 12292 37828 12684
rect 37772 12198 37828 12236
rect 37884 11954 37940 11966
rect 37884 11902 37886 11954
rect 37938 11902 37940 11954
rect 37772 11394 37828 11406
rect 37772 11342 37774 11394
rect 37826 11342 37828 11394
rect 37772 11284 37828 11342
rect 37772 11218 37828 11228
rect 37884 10722 37940 11902
rect 37884 10670 37886 10722
rect 37938 10670 37940 10722
rect 37884 10658 37940 10670
rect 37660 10556 37828 10612
rect 37660 10388 37716 10398
rect 37548 10386 37716 10388
rect 37548 10334 37662 10386
rect 37714 10334 37716 10386
rect 37548 10332 37716 10334
rect 37548 10050 37604 10332
rect 37660 10322 37716 10332
rect 37548 9998 37550 10050
rect 37602 9998 37604 10050
rect 37548 9986 37604 9998
rect 37436 9772 37604 9828
rect 37324 9660 37492 9716
rect 37436 9658 37492 9660
rect 37436 9606 37438 9658
rect 37490 9606 37492 9658
rect 37548 9714 37604 9772
rect 37548 9662 37550 9714
rect 37602 9662 37604 9714
rect 37548 9650 37604 9662
rect 37436 9594 37492 9606
rect 37212 9044 37268 9054
rect 37660 9044 37716 9054
rect 37772 9044 37828 10556
rect 37884 10500 37940 10510
rect 37884 10164 37940 10444
rect 37884 10098 37940 10108
rect 37212 9042 37828 9044
rect 37212 8990 37214 9042
rect 37266 8990 37662 9042
rect 37714 8990 37828 9042
rect 37212 8988 37828 8990
rect 37212 8978 37268 8988
rect 37660 8978 37716 8988
rect 36652 8764 37268 8820
rect 36428 7700 36484 7710
rect 36428 7606 36484 7644
rect 36876 7700 36932 7710
rect 36876 7474 36932 7644
rect 36876 7422 36878 7474
rect 36930 7422 36932 7474
rect 36876 7410 36932 7422
rect 36092 4284 36372 4340
rect 36652 5012 36708 5022
rect 36092 3668 36148 4284
rect 36092 3602 36148 3612
rect 36428 4226 36484 4238
rect 36428 4174 36430 4226
rect 36482 4174 36484 4226
rect 36204 3554 36260 3566
rect 36204 3502 36206 3554
rect 36258 3502 36260 3554
rect 35980 3444 36036 3454
rect 35868 3442 36036 3444
rect 35868 3390 35982 3442
rect 36034 3390 36036 3442
rect 35868 3388 36036 3390
rect 35756 3378 35812 3388
rect 35980 3378 36036 3388
rect 36204 3444 36260 3502
rect 36204 3378 36260 3388
rect 36316 3556 36372 3566
rect 34300 2380 34916 2436
rect 34972 2828 35252 2884
rect 34300 800 34356 2380
rect 34972 800 35028 2828
rect 35644 2546 35700 2558
rect 35644 2494 35646 2546
rect 35698 2494 35700 2546
rect 35644 800 35700 2494
rect 36316 800 36372 3500
rect 36428 2546 36484 4174
rect 36652 3442 36708 4956
rect 37100 4226 37156 4238
rect 37100 4174 37102 4226
rect 37154 4174 37156 4226
rect 36652 3390 36654 3442
rect 36706 3390 36708 3442
rect 36652 3378 36708 3390
rect 36876 3554 36932 3566
rect 36876 3502 36878 3554
rect 36930 3502 36932 3554
rect 36428 2494 36430 2546
rect 36482 2494 36484 2546
rect 36428 2482 36484 2494
rect 36876 2546 36932 3502
rect 37100 3556 37156 4174
rect 37100 3490 37156 3500
rect 37212 3444 37268 8764
rect 37548 8036 37604 8046
rect 37548 7586 37604 7980
rect 37996 7812 38052 14924
rect 38108 13634 38164 13646
rect 38108 13582 38110 13634
rect 38162 13582 38164 13634
rect 38108 12068 38164 13582
rect 38220 13524 38276 15260
rect 38444 15316 38500 15374
rect 38444 15250 38500 15260
rect 38668 14642 38724 15596
rect 38892 15586 38948 15596
rect 39228 15540 39284 16716
rect 39340 16660 39396 17388
rect 39452 16996 39508 17006
rect 39452 16902 39508 16940
rect 39676 16884 39732 17612
rect 39676 16818 39732 16828
rect 39340 16604 39844 16660
rect 39788 16210 39844 16604
rect 39788 16158 39790 16210
rect 39842 16158 39844 16210
rect 39788 16146 39844 16158
rect 39228 15446 39284 15484
rect 39004 15426 39060 15438
rect 39004 15374 39006 15426
rect 39058 15374 39060 15426
rect 38892 15316 38948 15326
rect 39004 15316 39060 15374
rect 38892 15314 39060 15316
rect 38892 15262 38894 15314
rect 38946 15262 39060 15314
rect 38892 15260 39060 15262
rect 39340 15314 39396 15326
rect 39340 15262 39342 15314
rect 39394 15262 39396 15314
rect 38892 15250 38948 15260
rect 38668 14590 38670 14642
rect 38722 14590 38724 14642
rect 38668 14578 38724 14590
rect 38780 15204 38836 15214
rect 38780 13970 38836 15148
rect 38780 13918 38782 13970
rect 38834 13918 38836 13970
rect 38780 13906 38836 13918
rect 39340 13972 39396 15262
rect 39564 14532 39620 14542
rect 39340 13906 39396 13916
rect 39452 14420 39508 14430
rect 39452 13970 39508 14364
rect 39452 13918 39454 13970
rect 39506 13918 39508 13970
rect 39452 13906 39508 13918
rect 39564 13858 39620 14476
rect 39564 13806 39566 13858
rect 39618 13806 39620 13858
rect 38332 13748 38388 13758
rect 38556 13748 38612 13758
rect 38332 13746 38612 13748
rect 38332 13694 38334 13746
rect 38386 13694 38558 13746
rect 38610 13694 38612 13746
rect 38332 13692 38612 13694
rect 38332 13682 38388 13692
rect 38556 13682 38612 13692
rect 38780 13748 38836 13758
rect 38220 13468 38388 13524
rect 38108 12002 38164 12012
rect 38220 12178 38276 12190
rect 38220 12126 38222 12178
rect 38274 12126 38276 12178
rect 38220 11844 38276 12126
rect 38108 11788 38276 11844
rect 38108 10612 38164 11788
rect 38332 11732 38388 13468
rect 38780 12962 38836 13692
rect 38892 13748 38948 13758
rect 39452 13748 39508 13758
rect 38892 13746 39396 13748
rect 38892 13694 38894 13746
rect 38946 13694 39396 13746
rect 38892 13692 39396 13694
rect 38892 13682 38948 13692
rect 38780 12910 38782 12962
rect 38834 12910 38836 12962
rect 38780 12898 38836 12910
rect 38556 12740 38612 12750
rect 38556 12646 38612 12684
rect 38556 12516 38612 12526
rect 38444 12180 38500 12190
rect 38444 12086 38500 12124
rect 38556 11732 38612 12460
rect 38780 12404 38836 12414
rect 38780 12310 38836 12348
rect 38668 12292 38724 12302
rect 39228 12292 39284 12302
rect 38668 12198 38724 12236
rect 38892 12290 39284 12292
rect 38892 12238 39230 12290
rect 39282 12238 39284 12290
rect 38892 12236 39284 12238
rect 38332 11666 38388 11676
rect 38444 11676 38724 11732
rect 38220 11620 38276 11658
rect 38220 11554 38276 11564
rect 38220 11394 38276 11406
rect 38220 11342 38222 11394
rect 38274 11342 38276 11394
rect 38220 10948 38276 11342
rect 38332 11396 38388 11406
rect 38444 11396 38500 11676
rect 38388 11340 38500 11396
rect 38556 11396 38612 11406
rect 38332 11330 38388 11340
rect 38220 10882 38276 10892
rect 38444 11172 38500 11182
rect 38108 10546 38164 10556
rect 38220 10724 38276 10734
rect 38220 10610 38276 10668
rect 38220 10558 38222 10610
rect 38274 10558 38276 10610
rect 38220 10546 38276 10558
rect 38444 10612 38500 11116
rect 38556 10834 38612 11340
rect 38556 10782 38558 10834
rect 38610 10782 38612 10834
rect 38556 10770 38612 10782
rect 38668 10836 38724 11676
rect 38780 11508 38836 11518
rect 38780 11394 38836 11452
rect 38780 11342 38782 11394
rect 38834 11342 38836 11394
rect 38780 11330 38836 11342
rect 38892 11284 38948 12236
rect 39228 12226 39284 12236
rect 39116 12068 39172 12078
rect 39116 11974 39172 12012
rect 39004 11954 39060 11966
rect 39004 11902 39006 11954
rect 39058 11902 39060 11954
rect 39004 11508 39060 11902
rect 39004 11442 39060 11452
rect 39116 11396 39172 11406
rect 39340 11396 39396 13692
rect 39452 13522 39508 13692
rect 39564 13636 39620 13806
rect 39564 13570 39620 13580
rect 39452 13470 39454 13522
rect 39506 13470 39508 13522
rect 39452 13458 39508 13470
rect 39452 12292 39508 12302
rect 39508 12236 39620 12292
rect 39452 12226 39508 12236
rect 39116 11394 39396 11396
rect 39116 11342 39118 11394
rect 39170 11342 39342 11394
rect 39394 11342 39396 11394
rect 39116 11340 39396 11342
rect 39116 11330 39172 11340
rect 39340 11330 39396 11340
rect 38892 11282 39060 11284
rect 38892 11230 38894 11282
rect 38946 11230 39060 11282
rect 38892 11228 39060 11230
rect 38892 11218 38948 11228
rect 38780 10836 38836 10846
rect 38668 10780 38780 10836
rect 38444 10556 38612 10612
rect 38444 10388 38500 10398
rect 38444 10294 38500 10332
rect 38220 9044 38276 9054
rect 38220 8950 38276 8988
rect 38332 8932 38388 8942
rect 38332 8370 38388 8876
rect 38332 8318 38334 8370
rect 38386 8318 38388 8370
rect 38332 8306 38388 8318
rect 38220 8036 38276 8046
rect 38220 7942 38276 7980
rect 37996 7756 38164 7812
rect 37548 7534 37550 7586
rect 37602 7534 37604 7586
rect 37548 7522 37604 7534
rect 37772 4226 37828 4238
rect 37772 4174 37774 4226
rect 37826 4174 37828 4226
rect 37772 4114 37828 4174
rect 37772 4062 37774 4114
rect 37826 4062 37828 4114
rect 37772 4050 37828 4062
rect 37548 3556 37604 3566
rect 37548 3462 37604 3500
rect 37884 3556 37940 3566
rect 37324 3444 37380 3454
rect 37212 3442 37380 3444
rect 37212 3390 37326 3442
rect 37378 3390 37380 3442
rect 37212 3388 37380 3390
rect 37884 3388 37940 3500
rect 37324 3378 37380 3388
rect 36876 2494 36878 2546
rect 36930 2494 36932 2546
rect 36876 2482 36932 2494
rect 37660 3332 37940 3388
rect 37996 3444 38052 3454
rect 38108 3444 38164 7756
rect 38556 4562 38612 10556
rect 38668 10164 38724 10174
rect 38668 8146 38724 10108
rect 38780 9938 38836 10780
rect 39004 10834 39060 11228
rect 39004 10782 39006 10834
rect 39058 10782 39060 10834
rect 39004 10770 39060 10782
rect 39564 10834 39620 12236
rect 39900 11844 39956 18396
rect 40348 18358 40404 18396
rect 40348 18004 40404 18014
rect 40348 17778 40404 17948
rect 40348 17726 40350 17778
rect 40402 17726 40404 17778
rect 40348 17714 40404 17726
rect 40460 17556 40516 18956
rect 40236 17500 40516 17556
rect 40012 15204 40068 15214
rect 40012 13970 40068 15148
rect 40012 13918 40014 13970
rect 40066 13918 40068 13970
rect 40012 13906 40068 13918
rect 39900 11778 39956 11788
rect 39788 11396 39844 11406
rect 39788 11302 39844 11340
rect 39676 11284 39732 11294
rect 39676 11190 39732 11228
rect 39900 11172 39956 11182
rect 39900 11078 39956 11116
rect 39564 10782 39566 10834
rect 39618 10782 39620 10834
rect 39564 10770 39620 10782
rect 38780 9886 38782 9938
rect 38834 9886 38836 9938
rect 38780 9874 38836 9886
rect 39004 10612 39060 10622
rect 39004 9828 39060 10556
rect 39788 10610 39844 10622
rect 39788 10558 39790 10610
rect 39842 10558 39844 10610
rect 39116 10500 39172 10510
rect 39788 10500 39844 10558
rect 39116 10498 39396 10500
rect 39116 10446 39118 10498
rect 39170 10446 39396 10498
rect 39116 10444 39396 10446
rect 39116 10434 39172 10444
rect 39340 10388 39396 10444
rect 39788 10434 39844 10444
rect 39452 10388 39508 10398
rect 39340 10386 39508 10388
rect 39340 10334 39454 10386
rect 39506 10334 39508 10386
rect 39340 10332 39508 10334
rect 39228 10276 39284 10286
rect 39116 9828 39172 9838
rect 39004 9826 39172 9828
rect 39004 9774 39118 9826
rect 39170 9774 39172 9826
rect 39004 9772 39172 9774
rect 39116 9154 39172 9772
rect 39228 9714 39284 10220
rect 39452 9828 39508 10332
rect 39452 9762 39508 9772
rect 40012 10164 40068 10174
rect 39228 9662 39230 9714
rect 39282 9662 39284 9714
rect 39228 9650 39284 9662
rect 40012 9266 40068 10108
rect 40012 9214 40014 9266
rect 40066 9214 40068 9266
rect 40012 9202 40068 9214
rect 40124 9716 40180 9726
rect 40124 9266 40180 9660
rect 40124 9214 40126 9266
rect 40178 9214 40180 9266
rect 40124 9202 40180 9214
rect 39116 9102 39118 9154
rect 39170 9102 39172 9154
rect 39116 9090 39172 9102
rect 39788 9156 39844 9166
rect 39788 9062 39844 9100
rect 38892 9044 38948 9054
rect 38892 8260 38948 8988
rect 39564 9042 39620 9054
rect 39564 8990 39566 9042
rect 39618 8990 39620 9042
rect 39564 8484 39620 8990
rect 39564 8418 39620 8428
rect 39676 9044 39732 9054
rect 39676 8370 39732 8988
rect 39900 8932 39956 8942
rect 39900 8838 39956 8876
rect 39676 8318 39678 8370
rect 39730 8318 39732 8370
rect 39676 8306 39732 8318
rect 38892 8258 39620 8260
rect 38892 8206 38894 8258
rect 38946 8206 39620 8258
rect 38892 8204 39620 8206
rect 38892 8194 38948 8204
rect 38668 8094 38670 8146
rect 38722 8094 38724 8146
rect 38668 8082 38724 8094
rect 39564 7364 39620 8204
rect 40124 7700 40180 7710
rect 40124 7606 40180 7644
rect 39676 7364 39732 7374
rect 39564 7362 39732 7364
rect 39564 7310 39678 7362
rect 39730 7310 39732 7362
rect 39564 7308 39732 7310
rect 39676 7298 39732 7308
rect 38556 4510 38558 4562
rect 38610 4510 38612 4562
rect 38556 4498 38612 4510
rect 38780 4338 38836 4350
rect 38780 4286 38782 4338
rect 38834 4286 38836 4338
rect 38332 4228 38388 4238
rect 38780 4228 38836 4286
rect 39340 4228 39396 4238
rect 38332 4226 38836 4228
rect 38332 4174 38334 4226
rect 38386 4174 38836 4226
rect 38332 4172 38836 4174
rect 39004 4226 39396 4228
rect 39004 4174 39342 4226
rect 39394 4174 39396 4226
rect 39004 4172 39396 4174
rect 38332 4162 38388 4172
rect 37996 3442 38164 3444
rect 37996 3390 37998 3442
rect 38050 3390 38164 3442
rect 37996 3388 38164 3390
rect 38220 4114 38276 4126
rect 38220 4062 38222 4114
rect 38274 4062 38276 4114
rect 38220 3554 38276 4062
rect 38220 3502 38222 3554
rect 38274 3502 38276 3554
rect 37996 3378 38052 3388
rect 36988 2434 37044 2446
rect 36988 2382 36990 2434
rect 37042 2382 37044 2434
rect 36988 800 37044 2382
rect 37660 800 37716 3332
rect 38220 2434 38276 3502
rect 38444 3332 38500 4172
rect 38668 4004 38724 4014
rect 38668 3442 38724 3948
rect 39004 3556 39060 4172
rect 39340 4162 39396 4172
rect 39788 4226 39844 4238
rect 39788 4174 39790 4226
rect 39842 4174 39844 4226
rect 39004 3462 39060 3500
rect 39788 3554 39844 4174
rect 39788 3502 39790 3554
rect 39842 3502 39844 3554
rect 38668 3390 38670 3442
rect 38722 3390 38724 3442
rect 38668 3378 38724 3390
rect 38220 2382 38222 2434
rect 38274 2382 38276 2434
rect 38220 2370 38276 2382
rect 38332 3276 38500 3332
rect 38332 800 38388 3276
rect 39788 2884 39844 3502
rect 39564 2828 39844 2884
rect 39900 3444 39956 3454
rect 39564 2548 39620 2828
rect 39900 2772 39956 3388
rect 40124 3444 40180 3454
rect 40236 3444 40292 17500
rect 40684 15148 40740 21868
rect 40572 15092 40740 15148
rect 40348 12740 40404 12750
rect 40348 12402 40404 12684
rect 40348 12350 40350 12402
rect 40402 12350 40404 12402
rect 40348 12338 40404 12350
rect 40572 11956 40628 15092
rect 40796 14644 40852 23660
rect 40908 23156 40964 23884
rect 41468 23846 41524 23884
rect 41020 23826 41076 23838
rect 41020 23774 41022 23826
rect 41074 23774 41076 23826
rect 41020 23268 41076 23774
rect 41020 23212 41300 23268
rect 40908 22484 40964 23100
rect 41132 23042 41188 23054
rect 41132 22990 41134 23042
rect 41186 22990 41188 23042
rect 41132 22930 41188 22990
rect 41244 23044 41300 23212
rect 41468 23044 41524 23054
rect 41244 23042 41524 23044
rect 41244 22990 41470 23042
rect 41522 22990 41524 23042
rect 41244 22988 41524 22990
rect 41132 22878 41134 22930
rect 41186 22878 41188 22930
rect 41132 22866 41188 22878
rect 41468 22820 41524 22988
rect 41580 22930 41636 25900
rect 41692 24164 41748 26852
rect 41804 26516 41860 27806
rect 42140 27860 42196 27870
rect 42140 27766 42196 27804
rect 42588 27524 42644 27534
rect 42588 27074 42644 27468
rect 42588 27022 42590 27074
rect 42642 27022 42644 27074
rect 42588 27010 42644 27022
rect 42028 26850 42084 26862
rect 42028 26798 42030 26850
rect 42082 26798 42084 26850
rect 42028 26740 42084 26798
rect 42028 26674 42084 26684
rect 42700 26740 42756 27916
rect 42700 26674 42756 26684
rect 42812 27860 42868 27870
rect 41916 26516 41972 26526
rect 41804 26514 41972 26516
rect 41804 26462 41918 26514
rect 41970 26462 41972 26514
rect 41804 26460 41972 26462
rect 41916 26450 41972 26460
rect 42028 26516 42084 26526
rect 41916 25506 41972 25518
rect 41916 25454 41918 25506
rect 41970 25454 41972 25506
rect 41916 24500 41972 25454
rect 41916 24434 41972 24444
rect 41692 24108 41972 24164
rect 41692 23938 41748 23950
rect 41692 23886 41694 23938
rect 41746 23886 41748 23938
rect 41692 23042 41748 23886
rect 41804 23938 41860 23950
rect 41804 23886 41806 23938
rect 41858 23886 41860 23938
rect 41804 23828 41860 23886
rect 41804 23762 41860 23772
rect 41916 23268 41972 24108
rect 41692 22990 41694 23042
rect 41746 22990 41748 23042
rect 41692 22978 41748 22990
rect 41804 23212 41972 23268
rect 41580 22878 41582 22930
rect 41634 22878 41636 22930
rect 41580 22866 41636 22878
rect 41468 22754 41524 22764
rect 41692 22596 41748 22606
rect 41692 22502 41748 22540
rect 41244 22484 41300 22494
rect 40908 22428 41244 22484
rect 41244 22390 41300 22428
rect 41804 22372 41860 23212
rect 41916 23042 41972 23054
rect 41916 22990 41918 23042
rect 41970 22990 41972 23042
rect 41916 22930 41972 22990
rect 41916 22878 41918 22930
rect 41970 22878 41972 22930
rect 41916 22484 41972 22878
rect 41916 22418 41972 22428
rect 41580 22370 41860 22372
rect 41580 22318 41806 22370
rect 41858 22318 41860 22370
rect 41580 22316 41860 22318
rect 41020 21812 41076 21822
rect 41020 21718 41076 21756
rect 41468 21700 41524 21710
rect 41468 21606 41524 21644
rect 41244 21586 41300 21598
rect 41244 21534 41246 21586
rect 41298 21534 41300 21586
rect 40908 20692 40964 20702
rect 41244 20692 41300 21534
rect 41356 21474 41412 21486
rect 41356 21422 41358 21474
rect 41410 21422 41412 21474
rect 41356 21028 41412 21422
rect 41356 20962 41412 20972
rect 41244 20636 41524 20692
rect 40908 20598 40964 20636
rect 41020 20580 41076 20618
rect 41020 20514 41076 20524
rect 41132 20578 41188 20590
rect 41132 20526 41134 20578
rect 41186 20526 41188 20578
rect 41020 20356 41076 20366
rect 41020 20242 41076 20300
rect 41020 20190 41022 20242
rect 41074 20190 41076 20242
rect 41020 20178 41076 20190
rect 41132 19908 41188 20526
rect 41468 20356 41524 20636
rect 41468 20290 41524 20300
rect 41468 19908 41524 19918
rect 41132 19906 41524 19908
rect 41132 19854 41470 19906
rect 41522 19854 41524 19906
rect 41132 19852 41524 19854
rect 41020 19460 41076 19470
rect 41020 19346 41076 19404
rect 41020 19294 41022 19346
rect 41074 19294 41076 19346
rect 41020 19282 41076 19294
rect 41356 18564 41412 19852
rect 41468 19842 41524 19852
rect 41244 17780 41300 17790
rect 41356 17780 41412 18508
rect 41300 17724 41412 17780
rect 41244 17714 41300 17724
rect 41244 17556 41300 17566
rect 41244 15538 41300 17500
rect 41244 15486 41246 15538
rect 41298 15486 41300 15538
rect 40796 14642 40964 14644
rect 40796 14590 40798 14642
rect 40850 14590 40964 14642
rect 40796 14588 40964 14590
rect 40796 14578 40852 14588
rect 40684 13076 40740 13086
rect 40684 12982 40740 13020
rect 40572 11890 40628 11900
rect 40908 12290 40964 14588
rect 41132 13860 41188 13870
rect 41132 13766 41188 13804
rect 41132 13636 41188 13646
rect 40908 12238 40910 12290
rect 40962 12238 40964 12290
rect 40908 12180 40964 12238
rect 41020 13524 41076 13534
rect 41020 12850 41076 13468
rect 41132 13186 41188 13580
rect 41132 13134 41134 13186
rect 41186 13134 41188 13186
rect 41132 13122 41188 13134
rect 41020 12798 41022 12850
rect 41074 12798 41076 12850
rect 41020 12180 41076 12798
rect 41132 12852 41188 12862
rect 41132 12758 41188 12796
rect 41244 12292 41300 15486
rect 41356 14980 41412 17724
rect 41468 19458 41524 19470
rect 41468 19406 41470 19458
rect 41522 19406 41524 19458
rect 41468 19346 41524 19406
rect 41468 19294 41470 19346
rect 41522 19294 41524 19346
rect 41468 18116 41524 19294
rect 41468 15148 41524 18060
rect 41580 16996 41636 22316
rect 41804 22260 41860 22316
rect 42028 22372 42084 26460
rect 42812 26514 42868 27804
rect 43484 27858 43540 28252
rect 43484 27806 43486 27858
rect 43538 27806 43540 27858
rect 43036 27186 43092 27198
rect 43036 27134 43038 27186
rect 43090 27134 43092 27186
rect 43036 26964 43092 27134
rect 43484 27074 43540 27806
rect 43820 27860 43876 27870
rect 43820 27766 43876 27804
rect 43932 27186 43988 28812
rect 44268 28754 44324 28924
rect 44268 28702 44270 28754
rect 44322 28702 44324 28754
rect 44268 28690 44324 28702
rect 44380 28756 44436 28766
rect 44156 28644 44212 28654
rect 44156 28082 44212 28588
rect 44156 28030 44158 28082
rect 44210 28030 44212 28082
rect 44156 28018 44212 28030
rect 44268 28084 44324 28094
rect 44380 28084 44436 28700
rect 44268 28082 44436 28084
rect 44268 28030 44270 28082
rect 44322 28030 44436 28082
rect 44268 28028 44436 28030
rect 44604 28532 44660 28542
rect 44268 28018 44324 28028
rect 43932 27134 43934 27186
rect 43986 27134 43988 27186
rect 43932 27122 43988 27134
rect 44044 27970 44100 27982
rect 44044 27918 44046 27970
rect 44098 27918 44100 27970
rect 44044 27748 44100 27918
rect 43484 27022 43486 27074
rect 43538 27022 43540 27074
rect 43036 26898 43092 26908
rect 43260 26964 43316 26974
rect 42812 26462 42814 26514
rect 42866 26462 42868 26514
rect 42812 26450 42868 26462
rect 42588 26404 42644 26414
rect 42476 26292 42532 26302
rect 42476 26198 42532 26236
rect 42588 26068 42644 26348
rect 43148 26404 43204 26414
rect 43148 26310 43204 26348
rect 43036 26292 43092 26302
rect 42252 26012 42644 26068
rect 42700 26290 43092 26292
rect 42700 26238 43038 26290
rect 43090 26238 43092 26290
rect 42700 26236 43092 26238
rect 42252 25620 42308 26012
rect 42700 25844 42756 26236
rect 43036 26226 43092 26236
rect 42252 25554 42308 25564
rect 42364 25788 42756 25844
rect 42364 25618 42420 25788
rect 42364 25566 42366 25618
rect 42418 25566 42420 25618
rect 42364 25554 42420 25566
rect 42924 25282 42980 25294
rect 42924 25230 42926 25282
rect 42978 25230 42980 25282
rect 42924 25172 42980 25230
rect 43260 25172 43316 26908
rect 43484 26740 43540 27022
rect 43932 26962 43988 26974
rect 43932 26910 43934 26962
rect 43986 26910 43988 26962
rect 43820 26740 43876 26750
rect 43484 26684 43764 26740
rect 43372 26516 43428 26526
rect 43372 26422 43428 26460
rect 43484 25618 43540 26684
rect 43708 26514 43764 26684
rect 43708 26462 43710 26514
rect 43762 26462 43764 26514
rect 43708 26450 43764 26462
rect 43820 25620 43876 26684
rect 43932 26516 43988 26910
rect 44044 26964 44100 27692
rect 44044 26898 44100 26908
rect 44156 27076 44212 27086
rect 43932 26450 43988 26460
rect 44044 26404 44100 26414
rect 44156 26404 44212 27020
rect 44268 26852 44324 26862
rect 44268 26850 44436 26852
rect 44268 26798 44270 26850
rect 44322 26798 44436 26850
rect 44268 26796 44436 26798
rect 44268 26786 44324 26796
rect 44156 26348 44324 26404
rect 44044 26180 44100 26348
rect 44156 26180 44212 26190
rect 44044 26178 44212 26180
rect 44044 26126 44158 26178
rect 44210 26126 44212 26178
rect 44044 26124 44212 26126
rect 44156 26114 44212 26124
rect 43484 25566 43486 25618
rect 43538 25566 43540 25618
rect 43484 25554 43540 25566
rect 43596 25618 43876 25620
rect 43596 25566 43822 25618
rect 43874 25566 43876 25618
rect 43596 25564 43876 25566
rect 42924 25116 43316 25172
rect 43036 24948 43092 24958
rect 42812 24946 43092 24948
rect 42812 24894 43038 24946
rect 43090 24894 43092 24946
rect 42812 24892 43092 24894
rect 42140 24722 42196 24734
rect 42140 24670 42142 24722
rect 42194 24670 42196 24722
rect 42140 24052 42196 24670
rect 42364 24724 42420 24734
rect 42812 24724 42868 24892
rect 43036 24882 43092 24892
rect 42364 24722 42868 24724
rect 42364 24670 42366 24722
rect 42418 24670 42868 24722
rect 42364 24668 42868 24670
rect 42924 24724 42980 24734
rect 42364 24658 42420 24668
rect 42924 24630 42980 24668
rect 43148 24722 43204 24734
rect 43148 24670 43150 24722
rect 43202 24670 43204 24722
rect 42476 24500 42532 24510
rect 43148 24500 43204 24670
rect 42476 24498 42756 24500
rect 42476 24446 42478 24498
rect 42530 24446 42756 24498
rect 42476 24444 42756 24446
rect 42476 24434 42532 24444
rect 42140 23380 42196 23996
rect 42476 23826 42532 23838
rect 42476 23774 42478 23826
rect 42530 23774 42532 23826
rect 42364 23380 42420 23390
rect 42140 23324 42364 23380
rect 42364 23286 42420 23324
rect 42476 22932 42532 23774
rect 42588 23714 42644 23726
rect 42588 23662 42590 23714
rect 42642 23662 42644 23714
rect 42588 23044 42644 23662
rect 42700 23268 42756 24444
rect 43260 24500 43316 25116
rect 43596 24722 43652 25564
rect 43820 25554 43876 25564
rect 44268 25282 44324 26348
rect 44380 26180 44436 26796
rect 44604 26740 44660 28476
rect 44716 27748 44772 27758
rect 44716 27654 44772 27692
rect 44828 27188 44884 27198
rect 44828 26962 44884 27132
rect 44940 27188 44996 27198
rect 45164 27188 45220 33854
rect 45388 31892 45444 34190
rect 45836 34242 45892 34254
rect 45836 34190 45838 34242
rect 45890 34190 45892 34242
rect 45836 33572 45892 34190
rect 45836 33506 45892 33516
rect 45612 33236 45668 33246
rect 45612 33142 45668 33180
rect 45276 30210 45332 30222
rect 45276 30158 45278 30210
rect 45330 30158 45332 30210
rect 45276 29650 45332 30158
rect 45388 30100 45444 31836
rect 45836 32004 45892 32014
rect 45724 31108 45780 31118
rect 45724 31014 45780 31052
rect 45500 30100 45556 30110
rect 45388 30098 45556 30100
rect 45388 30046 45502 30098
rect 45554 30046 45556 30098
rect 45388 30044 45556 30046
rect 45500 30034 45556 30044
rect 45276 29598 45278 29650
rect 45330 29598 45332 29650
rect 45276 29586 45332 29598
rect 45836 29652 45892 31948
rect 45948 31668 46004 34636
rect 45948 31602 46004 31612
rect 46060 34692 46116 36092
rect 46396 35586 46452 35598
rect 46396 35534 46398 35586
rect 46450 35534 46452 35586
rect 46396 35474 46452 35534
rect 46396 35422 46398 35474
rect 46450 35422 46452 35474
rect 46284 34692 46340 34702
rect 46060 34690 46340 34692
rect 46060 34638 46286 34690
rect 46338 34638 46340 34690
rect 46060 34636 46340 34638
rect 46060 31108 46116 34636
rect 46284 34626 46340 34636
rect 46060 31042 46116 31052
rect 46060 30436 46116 30446
rect 46060 30098 46116 30380
rect 46060 30046 46062 30098
rect 46114 30046 46116 30098
rect 46060 30034 46116 30046
rect 45948 29652 46004 29662
rect 45836 29650 46004 29652
rect 45836 29598 45950 29650
rect 46002 29598 46004 29650
rect 45836 29596 46004 29598
rect 45948 29540 46004 29596
rect 45948 29474 46004 29484
rect 46172 28868 46228 28878
rect 45948 28642 46004 28654
rect 45948 28590 45950 28642
rect 46002 28590 46004 28642
rect 45276 28420 45332 28430
rect 45276 28326 45332 28364
rect 45388 28418 45444 28430
rect 45388 28366 45390 28418
rect 45442 28366 45444 28418
rect 45388 28196 45444 28366
rect 45500 28420 45556 28430
rect 45500 28418 45892 28420
rect 45500 28366 45502 28418
rect 45554 28366 45892 28418
rect 45500 28364 45892 28366
rect 45500 28354 45556 28364
rect 45388 28140 45556 28196
rect 45388 27972 45444 27982
rect 45388 27858 45444 27916
rect 45388 27806 45390 27858
rect 45442 27806 45444 27858
rect 45388 27794 45444 27806
rect 44940 27186 45220 27188
rect 44940 27134 44942 27186
rect 44994 27134 45220 27186
rect 44940 27132 45220 27134
rect 45388 27524 45444 27534
rect 44940 27122 44996 27132
rect 44828 26910 44830 26962
rect 44882 26910 44884 26962
rect 44828 26898 44884 26910
rect 45388 26908 45444 27468
rect 45500 27074 45556 28140
rect 45500 27022 45502 27074
rect 45554 27022 45556 27074
rect 45500 27010 45556 27022
rect 45836 27188 45892 28364
rect 45948 27636 46004 28590
rect 46172 28642 46228 28812
rect 46172 28590 46174 28642
rect 46226 28590 46228 28642
rect 46172 28578 46228 28590
rect 46172 28196 46228 28206
rect 46060 28140 46172 28196
rect 46060 27970 46116 28140
rect 46172 28130 46228 28140
rect 46060 27918 46062 27970
rect 46114 27918 46116 27970
rect 46060 27906 46116 27918
rect 46396 27860 46452 35422
rect 46508 35476 46564 37324
rect 46620 37268 46676 37278
rect 46620 35588 46676 37212
rect 46732 36708 46788 41022
rect 46844 38276 46900 43372
rect 47516 43426 47572 43438
rect 47516 43374 47518 43426
rect 47570 43374 47572 43426
rect 47516 42866 47572 43374
rect 47516 42814 47518 42866
rect 47570 42814 47572 42866
rect 47516 42802 47572 42814
rect 47404 42756 47460 42766
rect 47404 42662 47460 42700
rect 47628 42754 47684 43484
rect 47628 42702 47630 42754
rect 47682 42702 47684 42754
rect 47628 42690 47684 42702
rect 47516 41972 47572 41982
rect 47516 41878 47572 41916
rect 47628 41636 47684 41646
rect 47068 41412 47124 41422
rect 47068 40292 47124 41356
rect 47628 41188 47684 41580
rect 47628 41094 47684 41132
rect 47516 41076 47572 41086
rect 47516 40982 47572 41020
rect 47068 40226 47124 40236
rect 47404 40962 47460 40974
rect 47404 40910 47406 40962
rect 47458 40910 47460 40962
rect 47180 38724 47236 38734
rect 46844 38210 46900 38220
rect 46956 38612 47012 38622
rect 46956 38050 47012 38556
rect 47180 38162 47236 38668
rect 47404 38668 47460 40910
rect 47404 38612 47684 38668
rect 47180 38110 47182 38162
rect 47234 38110 47236 38162
rect 47180 38098 47236 38110
rect 47292 38276 47348 38286
rect 46956 37998 46958 38050
rect 47010 37998 47012 38050
rect 46956 37986 47012 37998
rect 47068 38052 47124 38062
rect 47068 37958 47124 37996
rect 47292 38050 47348 38220
rect 47292 37998 47294 38050
rect 47346 37998 47348 38050
rect 47292 37986 47348 37998
rect 47516 37938 47572 37950
rect 47516 37886 47518 37938
rect 47570 37886 47572 37938
rect 47068 37268 47124 37278
rect 47068 37174 47124 37212
rect 46844 37156 46900 37166
rect 46844 37154 47012 37156
rect 46844 37102 46846 37154
rect 46898 37102 47012 37154
rect 46844 37100 47012 37102
rect 46844 37090 46900 37100
rect 46732 36370 46788 36652
rect 46956 36596 47012 37100
rect 47068 36596 47124 36606
rect 46956 36594 47124 36596
rect 46956 36542 47070 36594
rect 47122 36542 47124 36594
rect 46956 36540 47124 36542
rect 47068 36530 47124 36540
rect 47516 36484 47572 37886
rect 47628 37378 47684 38612
rect 47628 37326 47630 37378
rect 47682 37326 47684 37378
rect 47628 37314 47684 37326
rect 47516 36390 47572 36428
rect 47740 36482 47796 44156
rect 47964 44146 48020 44156
rect 47852 43652 47908 43662
rect 48636 43652 48692 44828
rect 48748 44324 48804 45836
rect 49420 44546 49476 44558
rect 49420 44494 49422 44546
rect 49474 44494 49476 44546
rect 49084 44434 49140 44446
rect 49084 44382 49086 44434
rect 49138 44382 49140 44434
rect 48972 44324 49028 44334
rect 48748 44322 49028 44324
rect 48748 44270 48974 44322
rect 49026 44270 49028 44322
rect 48748 44268 49028 44270
rect 48972 44258 49028 44268
rect 49084 43762 49140 44382
rect 49084 43710 49086 43762
rect 49138 43710 49140 43762
rect 49084 43698 49140 43710
rect 48748 43652 48804 43662
rect 48636 43650 48804 43652
rect 48636 43598 48750 43650
rect 48802 43598 48804 43650
rect 48636 43596 48804 43598
rect 47852 42642 47908 43596
rect 48748 43586 48804 43596
rect 48860 43652 48916 43662
rect 48860 43558 48916 43596
rect 47852 42590 47854 42642
rect 47906 42590 47908 42642
rect 47852 42196 47908 42590
rect 47852 42130 47908 42140
rect 48076 43314 48132 43326
rect 48076 43262 48078 43314
rect 48130 43262 48132 43314
rect 47964 42082 48020 42094
rect 47964 42030 47966 42082
rect 48018 42030 48020 42082
rect 47964 41972 48020 42030
rect 48076 42082 48132 43262
rect 49420 42754 49476 44494
rect 49420 42702 49422 42754
rect 49474 42702 49476 42754
rect 49420 42690 49476 42702
rect 48860 42532 48916 42542
rect 48860 42438 48916 42476
rect 49084 42532 49140 42542
rect 49308 42532 49364 42542
rect 49084 42530 49252 42532
rect 49084 42478 49086 42530
rect 49138 42478 49252 42530
rect 49084 42476 49252 42478
rect 49084 42466 49140 42476
rect 49196 42308 49252 42476
rect 49308 42438 49364 42476
rect 49196 42252 49588 42308
rect 49532 42194 49588 42252
rect 49532 42142 49534 42194
rect 49586 42142 49588 42194
rect 49532 42130 49588 42142
rect 48076 42030 48078 42082
rect 48130 42030 48132 42082
rect 48076 42018 48132 42030
rect 49308 42082 49364 42094
rect 49308 42030 49310 42082
rect 49362 42030 49364 42082
rect 47964 41906 48020 41916
rect 49084 41970 49140 41982
rect 49084 41918 49086 41970
rect 49138 41918 49140 41970
rect 47964 41746 48020 41758
rect 47964 41694 47966 41746
rect 48018 41694 48020 41746
rect 47964 41186 48020 41694
rect 49084 41300 49140 41918
rect 49196 41858 49252 41870
rect 49196 41806 49198 41858
rect 49250 41806 49252 41858
rect 49196 41412 49252 41806
rect 49308 41636 49364 42030
rect 49644 41748 49700 45836
rect 50204 45780 50260 46844
rect 50428 46564 50484 47292
rect 50652 47282 50708 47292
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50540 46564 50596 46574
rect 50428 46508 50540 46564
rect 50540 46470 50596 46508
rect 50428 46004 50484 46042
rect 50428 45938 50484 45948
rect 50988 46004 51044 47406
rect 51212 47460 51268 47740
rect 51772 47572 51828 47582
rect 51436 47460 51492 47470
rect 51212 47458 51492 47460
rect 51212 47406 51214 47458
rect 51266 47406 51438 47458
rect 51490 47406 51492 47458
rect 51212 47404 51492 47406
rect 51212 47394 51268 47404
rect 51436 47394 51492 47404
rect 51772 47234 51828 47516
rect 51884 47458 51940 48188
rect 51884 47406 51886 47458
rect 51938 47406 51940 47458
rect 51884 47394 51940 47406
rect 51996 48018 52052 48030
rect 51996 47966 51998 48018
rect 52050 47966 52052 48018
rect 51772 47182 51774 47234
rect 51826 47182 51828 47234
rect 51772 47170 51828 47182
rect 51996 46788 52052 47966
rect 52332 48018 52388 48030
rect 52332 47966 52334 48018
rect 52386 47966 52388 48018
rect 52332 47572 52388 47966
rect 52332 47506 52388 47516
rect 51996 46722 52052 46732
rect 52108 47346 52164 47358
rect 52108 47294 52110 47346
rect 52162 47294 52164 47346
rect 50988 45938 51044 45948
rect 51884 45780 51940 45790
rect 50204 45724 50932 45780
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50764 45332 50820 45342
rect 50764 44210 50820 45276
rect 50876 45330 50932 45724
rect 50876 45278 50878 45330
rect 50930 45278 50932 45330
rect 50876 45266 50932 45278
rect 50988 45778 51940 45780
rect 50988 45726 51886 45778
rect 51938 45726 51940 45778
rect 50988 45724 51940 45726
rect 50876 44436 50932 44446
rect 50988 44436 51044 45724
rect 51884 45714 51940 45724
rect 51996 45668 52052 45678
rect 51996 45574 52052 45612
rect 51660 45444 51716 45454
rect 51212 44996 51268 45006
rect 51212 44902 51268 44940
rect 50876 44434 51044 44436
rect 50876 44382 50878 44434
rect 50930 44382 51044 44434
rect 50876 44380 51044 44382
rect 51100 44548 51156 44558
rect 50876 44370 50932 44380
rect 50764 44158 50766 44210
rect 50818 44158 50820 44210
rect 50764 44100 50820 44158
rect 50988 44212 51044 44222
rect 51100 44212 51156 44492
rect 51660 44546 51716 45388
rect 51660 44494 51662 44546
rect 51714 44494 51716 44546
rect 50988 44210 51156 44212
rect 50988 44158 50990 44210
rect 51042 44158 51156 44210
rect 50988 44156 51156 44158
rect 51212 44212 51268 44222
rect 50988 44146 51044 44156
rect 51212 44118 51268 44156
rect 50764 44034 50820 44044
rect 50988 43988 51044 43998
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50876 43932 50988 43988
rect 49868 43652 49924 43662
rect 49756 43650 49924 43652
rect 49756 43598 49870 43650
rect 49922 43598 49924 43650
rect 49756 43596 49924 43598
rect 49756 42980 49812 43596
rect 49868 43586 49924 43596
rect 49980 43652 50036 43662
rect 49980 43558 50036 43596
rect 50876 43538 50932 43932
rect 50988 43922 51044 43932
rect 51660 43988 51716 44494
rect 52108 44996 52164 47294
rect 52220 45666 52276 45678
rect 52220 45614 52222 45666
rect 52274 45614 52276 45666
rect 52220 45444 52276 45614
rect 52220 45378 52276 45388
rect 51884 44436 51940 44446
rect 51884 44342 51940 44380
rect 52108 44434 52164 44940
rect 52108 44382 52110 44434
rect 52162 44382 52164 44434
rect 51660 43922 51716 43932
rect 50876 43486 50878 43538
rect 50930 43486 50932 43538
rect 50876 43474 50932 43486
rect 51212 43538 51268 43550
rect 51212 43486 51214 43538
rect 51266 43486 51268 43538
rect 49868 43316 49924 43326
rect 49868 43222 49924 43260
rect 51212 43204 51268 43486
rect 51772 43540 51828 43550
rect 52108 43540 52164 44382
rect 51772 43446 51828 43484
rect 51884 43538 52164 43540
rect 51884 43486 52110 43538
rect 52162 43486 52164 43538
rect 51884 43484 52164 43486
rect 51324 43428 51380 43438
rect 51324 43426 51604 43428
rect 51324 43374 51326 43426
rect 51378 43374 51604 43426
rect 51324 43372 51604 43374
rect 51324 43362 51380 43372
rect 49756 42914 49812 42924
rect 50428 43148 50820 43204
rect 51212 43148 51380 43204
rect 50428 42754 50484 43148
rect 50764 43092 50820 43148
rect 50764 43036 51268 43092
rect 50428 42702 50430 42754
rect 50482 42702 50484 42754
rect 50428 42690 50484 42702
rect 50652 42980 50708 42990
rect 50652 42642 50708 42924
rect 50988 42868 51044 42878
rect 51044 42812 51156 42868
rect 50988 42802 51044 42812
rect 50764 42756 50820 42766
rect 50764 42662 50820 42700
rect 50652 42590 50654 42642
rect 50706 42590 50708 42642
rect 50652 42578 50708 42590
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50988 42308 51044 42318
rect 50876 41860 50932 41870
rect 50876 41766 50932 41804
rect 49644 41682 49700 41692
rect 49308 41570 49364 41580
rect 49196 41356 50148 41412
rect 49084 41244 49252 41300
rect 47964 41134 47966 41186
rect 48018 41134 48020 41186
rect 47964 41122 48020 41134
rect 48412 41186 48468 41198
rect 48412 41134 48414 41186
rect 48466 41134 48468 41186
rect 48412 40404 48468 41134
rect 48412 40338 48468 40348
rect 48748 41188 48804 41198
rect 48076 40290 48132 40302
rect 48076 40238 48078 40290
rect 48130 40238 48132 40290
rect 48076 40180 48132 40238
rect 48076 40114 48132 40124
rect 48748 39956 48804 41132
rect 49084 41076 49140 41086
rect 49084 40982 49140 41020
rect 48748 39890 48804 39900
rect 48860 40404 48916 40414
rect 48860 39732 48916 40348
rect 48972 39732 49028 39742
rect 48860 39730 49028 39732
rect 48860 39678 48974 39730
rect 49026 39678 49028 39730
rect 48860 39676 49028 39678
rect 48860 38836 48916 39676
rect 48972 39666 49028 39676
rect 48748 38834 48916 38836
rect 48748 38782 48862 38834
rect 48914 38782 48916 38834
rect 48748 38780 48916 38782
rect 48748 38052 48804 38780
rect 48860 38770 48916 38780
rect 49196 38668 49252 41244
rect 50092 40514 50148 41356
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50092 40462 50094 40514
rect 50146 40462 50148 40514
rect 50092 40450 50148 40462
rect 49308 40404 49364 40414
rect 49308 40310 49364 40348
rect 50316 39396 50372 39406
rect 50316 39302 50372 39340
rect 50764 39396 50820 39406
rect 50764 39394 50932 39396
rect 50764 39342 50766 39394
rect 50818 39342 50932 39394
rect 50764 39340 50932 39342
rect 50764 39330 50820 39340
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50876 38948 50932 39340
rect 50988 39060 51044 42252
rect 51100 42196 51156 42812
rect 51212 42866 51268 43036
rect 51212 42814 51214 42866
rect 51266 42814 51268 42866
rect 51212 42802 51268 42814
rect 51212 42196 51268 42206
rect 51100 42194 51268 42196
rect 51100 42142 51214 42194
rect 51266 42142 51268 42194
rect 51100 42140 51268 42142
rect 51212 42130 51268 42140
rect 51324 42194 51380 43148
rect 51436 43092 51492 43102
rect 51436 42754 51492 43036
rect 51436 42702 51438 42754
rect 51490 42702 51492 42754
rect 51436 42690 51492 42702
rect 51324 42142 51326 42194
rect 51378 42142 51380 42194
rect 51324 42130 51380 42142
rect 51436 42196 51492 42206
rect 51436 42102 51492 42140
rect 51324 41972 51380 41982
rect 51212 41300 51268 41310
rect 51324 41300 51380 41916
rect 51212 41298 51380 41300
rect 51212 41246 51214 41298
rect 51266 41246 51380 41298
rect 51212 41244 51380 41246
rect 51212 41234 51268 41244
rect 51212 40404 51268 40414
rect 51212 39732 51268 40348
rect 51212 39638 51268 39676
rect 51548 39618 51604 43372
rect 51660 43426 51716 43438
rect 51660 43374 51662 43426
rect 51714 43374 51716 43426
rect 51660 41188 51716 43374
rect 51884 42196 51940 43484
rect 52108 43474 52164 43484
rect 52556 44548 52612 49084
rect 52668 49074 52724 49084
rect 52668 48916 52724 48926
rect 52668 48242 52724 48860
rect 54124 48916 54180 49980
rect 54572 49922 54628 50372
rect 54572 49870 54574 49922
rect 54626 49870 54628 49922
rect 54572 49858 54628 49870
rect 54124 48850 54180 48860
rect 52668 48190 52670 48242
rect 52722 48190 52724 48242
rect 52668 48178 52724 48190
rect 53340 48804 53396 48814
rect 53116 48132 53172 48142
rect 53340 48132 53396 48748
rect 53172 48076 53396 48132
rect 53116 48038 53172 48076
rect 52668 48020 52724 48030
rect 52668 48018 53060 48020
rect 52668 47966 52670 48018
rect 52722 47966 53060 48018
rect 52668 47964 53060 47966
rect 52668 47954 52724 47964
rect 52668 46788 52724 46798
rect 52668 46694 52724 46732
rect 53004 46452 53060 47964
rect 53340 46900 53396 48076
rect 53900 46900 53956 46910
rect 53340 46898 54068 46900
rect 53340 46846 53902 46898
rect 53954 46846 54068 46898
rect 53340 46844 54068 46846
rect 53340 46674 53396 46844
rect 53900 46834 53956 46844
rect 53340 46622 53342 46674
rect 53394 46622 53396 46674
rect 53340 46610 53396 46622
rect 53004 46396 53396 46452
rect 52668 45892 52724 45902
rect 52668 45798 52724 45836
rect 52108 42644 52164 42654
rect 51884 42130 51940 42140
rect 51996 42642 52164 42644
rect 51996 42590 52110 42642
rect 52162 42590 52164 42642
rect 51996 42588 52164 42590
rect 51884 41972 51940 41982
rect 51884 41878 51940 41916
rect 51660 41132 51940 41188
rect 51660 40964 51716 40974
rect 51660 40870 51716 40908
rect 51660 40404 51716 40414
rect 51660 39730 51716 40348
rect 51660 39678 51662 39730
rect 51714 39678 51716 39730
rect 51660 39666 51716 39678
rect 51548 39566 51550 39618
rect 51602 39566 51604 39618
rect 51548 39554 51604 39566
rect 51772 39396 51828 39406
rect 51772 39302 51828 39340
rect 50988 39004 51716 39060
rect 50876 38882 50932 38892
rect 48412 38050 48804 38052
rect 48412 37998 48750 38050
rect 48802 37998 48804 38050
rect 48412 37996 48804 37998
rect 47852 37940 47908 37950
rect 47852 36594 47908 37884
rect 48412 37492 48468 37996
rect 48748 37986 48804 37996
rect 48972 38612 49252 38668
rect 49532 38724 49588 38762
rect 49532 38658 49588 38668
rect 51660 38722 51716 39004
rect 51660 38670 51662 38722
rect 51714 38670 51716 38722
rect 51660 38658 51716 38670
rect 51884 38668 51940 41132
rect 51996 40404 52052 42588
rect 52108 42578 52164 42588
rect 52556 41970 52612 44492
rect 53004 45668 53060 45678
rect 52668 44322 52724 44334
rect 52668 44270 52670 44322
rect 52722 44270 52724 44322
rect 52668 42084 52724 44270
rect 53004 43650 53060 45612
rect 53340 45218 53396 46396
rect 53340 45166 53342 45218
rect 53394 45166 53396 45218
rect 53340 45154 53396 45166
rect 54012 45106 54068 46844
rect 54684 45332 54740 51436
rect 55580 51492 55636 51502
rect 55580 50706 55636 51436
rect 55580 50654 55582 50706
rect 55634 50654 55636 50706
rect 55580 50642 55636 50654
rect 54796 50036 54852 50046
rect 54796 49942 54852 49980
rect 54796 49698 54852 49710
rect 54796 49646 54798 49698
rect 54850 49646 54852 49698
rect 54796 49138 54852 49646
rect 54796 49086 54798 49138
rect 54850 49086 54852 49138
rect 54796 49074 54852 49086
rect 55468 49026 55524 49038
rect 55468 48974 55470 49026
rect 55522 48974 55524 49026
rect 55468 48804 55524 48974
rect 55468 48738 55524 48748
rect 57932 47570 57988 47582
rect 57932 47518 57934 47570
rect 57986 47518 57988 47570
rect 55580 47458 55636 47470
rect 55580 47406 55582 47458
rect 55634 47406 55636 47458
rect 55244 47236 55300 47246
rect 55580 47236 55636 47406
rect 55244 47234 55636 47236
rect 55244 47182 55246 47234
rect 55298 47182 55636 47234
rect 55244 47180 55636 47182
rect 55244 46228 55300 47180
rect 55244 46162 55300 46172
rect 54684 45238 54740 45276
rect 54908 46002 54964 46014
rect 54908 45950 54910 46002
rect 54962 45950 54964 46002
rect 54012 45054 54014 45106
rect 54066 45054 54068 45106
rect 54012 45042 54068 45054
rect 54460 45106 54516 45118
rect 54460 45054 54462 45106
rect 54514 45054 54516 45106
rect 53004 43598 53006 43650
rect 53058 43598 53060 43650
rect 53004 43586 53060 43598
rect 53116 43652 53172 43662
rect 52668 42018 52724 42028
rect 53004 43204 53060 43214
rect 52556 41918 52558 41970
rect 52610 41918 52612 41970
rect 52556 41906 52612 41918
rect 53004 41970 53060 43148
rect 53116 42756 53172 43596
rect 54460 43652 54516 45054
rect 54460 43586 54516 43596
rect 54572 44994 54628 45006
rect 54572 44942 54574 44994
rect 54626 44942 54628 44994
rect 53452 43540 53508 43550
rect 53452 43538 53620 43540
rect 53452 43486 53454 43538
rect 53506 43486 53620 43538
rect 53452 43484 53620 43486
rect 53452 43474 53508 43484
rect 53116 42690 53172 42700
rect 53004 41918 53006 41970
rect 53058 41918 53060 41970
rect 53004 41906 53060 41918
rect 53452 41970 53508 41982
rect 53452 41918 53454 41970
rect 53506 41918 53508 41970
rect 53116 41858 53172 41870
rect 53116 41806 53118 41858
rect 53170 41806 53172 41858
rect 52668 41188 52724 41198
rect 52668 41094 52724 41132
rect 52108 40964 52164 40974
rect 52108 40516 52164 40908
rect 53116 40628 53172 41806
rect 53452 41412 53508 41918
rect 53452 41346 53508 41356
rect 53116 40562 53172 40572
rect 53228 41188 53284 41198
rect 52108 40460 52388 40516
rect 52332 40404 52388 40460
rect 52780 40404 52836 40414
rect 51996 40348 52164 40404
rect 52332 40402 52836 40404
rect 52332 40350 52782 40402
rect 52834 40350 52836 40402
rect 52332 40348 52836 40350
rect 51772 38612 51940 38668
rect 52108 38668 52164 40348
rect 52220 40292 52276 40302
rect 52220 40198 52276 40236
rect 52780 39732 52836 40348
rect 52220 39618 52276 39630
rect 52220 39566 52222 39618
rect 52274 39566 52276 39618
rect 52220 39058 52276 39566
rect 52220 39006 52222 39058
rect 52274 39006 52276 39058
rect 52220 38994 52276 39006
rect 52444 38948 52500 38958
rect 52444 38854 52500 38892
rect 52556 38834 52612 38846
rect 52556 38782 52558 38834
rect 52610 38782 52612 38834
rect 52108 38612 52500 38668
rect 48076 37268 48132 37278
rect 48076 37174 48132 37212
rect 47852 36542 47854 36594
rect 47906 36542 47908 36594
rect 47852 36530 47908 36542
rect 48412 36484 48468 37436
rect 48860 37268 48916 37278
rect 48860 37174 48916 37212
rect 48972 36932 49028 38612
rect 51772 38388 51828 38612
rect 51436 38332 51828 38388
rect 50876 38164 50932 38174
rect 49532 37940 49588 37950
rect 49532 37846 49588 37884
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50428 37492 50484 37502
rect 50428 37398 50484 37436
rect 50876 37492 50932 38108
rect 50876 37490 51268 37492
rect 50876 37438 50878 37490
rect 50930 37438 51268 37490
rect 50876 37436 51268 37438
rect 50876 37426 50932 37436
rect 51212 37380 51268 37436
rect 51436 37490 51492 38332
rect 51660 38162 51716 38174
rect 51660 38110 51662 38162
rect 51714 38110 51716 38162
rect 51660 37604 51716 38110
rect 52220 37826 52276 37838
rect 52220 37774 52222 37826
rect 52274 37774 52276 37826
rect 51660 37548 52052 37604
rect 51436 37438 51438 37490
rect 51490 37438 51492 37490
rect 51436 37426 51492 37438
rect 51212 37286 51268 37324
rect 51548 37268 51604 37278
rect 51548 37174 51604 37212
rect 51660 37266 51716 37278
rect 51660 37214 51662 37266
rect 51714 37214 51716 37266
rect 47740 36430 47742 36482
rect 47794 36430 47796 36482
rect 47740 36418 47796 36430
rect 48188 36428 48468 36484
rect 48748 36876 49028 36932
rect 51324 37044 51380 37054
rect 46732 36318 46734 36370
rect 46786 36318 46788 36370
rect 46732 36306 46788 36318
rect 46956 36258 47012 36270
rect 46956 36206 46958 36258
rect 47010 36206 47012 36258
rect 46956 36148 47012 36206
rect 46956 36082 47012 36092
rect 47180 36260 47236 36270
rect 47964 36260 48020 36270
rect 47180 35812 47236 36204
rect 47180 35698 47236 35756
rect 47628 36258 48020 36260
rect 47628 36206 47966 36258
rect 48018 36206 48020 36258
rect 47628 36204 48020 36206
rect 47628 35700 47684 36204
rect 47964 36194 48020 36204
rect 48076 36260 48132 36270
rect 48076 36166 48132 36204
rect 47852 35812 47908 35822
rect 47852 35718 47908 35756
rect 47964 35812 48020 35822
rect 48076 35812 48132 35822
rect 47964 35810 48076 35812
rect 47964 35758 47966 35810
rect 48018 35758 48076 35810
rect 47964 35756 48076 35758
rect 47964 35746 48020 35756
rect 47180 35646 47182 35698
rect 47234 35646 47236 35698
rect 47180 35634 47236 35646
rect 47516 35644 47684 35700
rect 46732 35588 46788 35598
rect 46620 35586 46788 35588
rect 46620 35534 46734 35586
rect 46786 35534 46788 35586
rect 46620 35532 46788 35534
rect 46508 35410 46564 35420
rect 46620 35140 46676 35150
rect 46620 34690 46676 35084
rect 46620 34638 46622 34690
rect 46674 34638 46676 34690
rect 46620 33684 46676 34638
rect 46620 33618 46676 33628
rect 46396 27794 46452 27804
rect 46508 31668 46564 31678
rect 46396 27636 46452 27646
rect 45948 27580 46228 27636
rect 45836 27076 45892 27132
rect 46172 27186 46228 27580
rect 46172 27134 46174 27186
rect 46226 27134 46228 27186
rect 46172 27122 46228 27134
rect 45948 27076 46004 27086
rect 45836 27074 46004 27076
rect 45836 27022 45950 27074
rect 46002 27022 46004 27074
rect 45836 27020 46004 27022
rect 45948 27010 46004 27020
rect 46396 27074 46452 27580
rect 46396 27022 46398 27074
rect 46450 27022 46452 27074
rect 46396 27010 46452 27022
rect 45724 26962 45780 26974
rect 45724 26910 45726 26962
rect 45778 26910 45780 26962
rect 45724 26908 45780 26910
rect 45052 26850 45108 26862
rect 45388 26852 45780 26908
rect 45052 26798 45054 26850
rect 45106 26798 45108 26850
rect 45052 26740 45108 26798
rect 44604 26684 45108 26740
rect 45052 26514 45108 26684
rect 45052 26462 45054 26514
rect 45106 26462 45108 26514
rect 45052 26450 45108 26462
rect 45500 26514 45556 26852
rect 45500 26462 45502 26514
rect 45554 26462 45556 26514
rect 45500 26450 45556 26462
rect 46060 26740 46116 26750
rect 44604 26404 44660 26414
rect 44604 26310 44660 26348
rect 44380 26124 44660 26180
rect 44268 25230 44270 25282
rect 44322 25230 44324 25282
rect 43596 24670 43598 24722
rect 43650 24670 43652 24722
rect 43596 24658 43652 24670
rect 43820 24722 43876 24734
rect 43820 24670 43822 24722
rect 43874 24670 43876 24722
rect 43260 24444 43652 24500
rect 43148 24434 43204 24444
rect 42812 23716 42868 23726
rect 43260 23716 43316 23726
rect 42812 23714 43316 23716
rect 42812 23662 42814 23714
rect 42866 23662 43262 23714
rect 43314 23662 43316 23714
rect 42812 23660 43316 23662
rect 42812 23650 42868 23660
rect 43260 23650 43316 23660
rect 43372 23714 43428 23726
rect 43372 23662 43374 23714
rect 43426 23662 43428 23714
rect 42812 23492 42868 23502
rect 43148 23492 43204 23502
rect 42868 23436 43092 23492
rect 42812 23426 42868 23436
rect 42812 23268 42868 23278
rect 42700 23266 42868 23268
rect 42700 23214 42814 23266
rect 42866 23214 42868 23266
rect 42700 23212 42868 23214
rect 42812 23202 42868 23212
rect 42924 23266 42980 23278
rect 42924 23214 42926 23266
rect 42978 23214 42980 23266
rect 42924 23044 42980 23214
rect 42588 22988 42924 23044
rect 42476 22866 42532 22876
rect 42028 22306 42084 22316
rect 41804 22194 41860 22204
rect 42364 22258 42420 22270
rect 42364 22206 42366 22258
rect 42418 22206 42420 22258
rect 41692 22146 41748 22158
rect 41692 22094 41694 22146
rect 41746 22094 41748 22146
rect 41692 21924 41748 22094
rect 42364 22148 42420 22206
rect 42364 22082 42420 22092
rect 42476 22146 42532 22158
rect 42476 22094 42478 22146
rect 42530 22094 42532 22146
rect 41692 21868 42308 21924
rect 42028 21588 42084 21598
rect 42028 21586 42196 21588
rect 42028 21534 42030 21586
rect 42082 21534 42196 21586
rect 42028 21532 42196 21534
rect 42028 21522 42084 21532
rect 41916 21476 41972 21486
rect 41916 20914 41972 21420
rect 41916 20862 41918 20914
rect 41970 20862 41972 20914
rect 41916 20850 41972 20862
rect 41804 20804 41860 20814
rect 41804 20710 41860 20748
rect 42028 20802 42084 20814
rect 42028 20750 42030 20802
rect 42082 20750 42084 20802
rect 42028 20132 42084 20750
rect 42140 20356 42196 21532
rect 42252 20580 42308 21868
rect 42364 20804 42420 20814
rect 42476 20804 42532 22094
rect 42588 22146 42644 22158
rect 42588 22094 42590 22146
rect 42642 22094 42644 22146
rect 42588 22036 42644 22094
rect 42588 21970 42644 21980
rect 42924 21924 42980 22988
rect 43036 22596 43092 23436
rect 43148 23378 43204 23436
rect 43148 23326 43150 23378
rect 43202 23326 43204 23378
rect 43148 23314 43204 23326
rect 43372 23156 43428 23662
rect 43484 23716 43540 23726
rect 43484 23622 43540 23660
rect 43484 23380 43540 23390
rect 43484 23286 43540 23324
rect 43372 23090 43428 23100
rect 43596 22596 43652 24444
rect 43708 23938 43764 23950
rect 43708 23886 43710 23938
rect 43762 23886 43764 23938
rect 43708 23268 43764 23886
rect 43820 23604 43876 24670
rect 44268 24722 44324 25230
rect 44268 24670 44270 24722
rect 44322 24670 44324 24722
rect 43932 23940 43988 23950
rect 44268 23940 44324 24670
rect 44492 24724 44548 24734
rect 44492 24630 44548 24668
rect 44380 24610 44436 24622
rect 44380 24558 44382 24610
rect 44434 24558 44436 24610
rect 44380 24164 44436 24558
rect 44604 24612 44660 26124
rect 45164 25394 45220 25406
rect 45164 25342 45166 25394
rect 45218 25342 45220 25394
rect 45164 25060 45220 25342
rect 45500 25284 45556 25294
rect 45500 25282 45892 25284
rect 45500 25230 45502 25282
rect 45554 25230 45892 25282
rect 45500 25228 45892 25230
rect 45500 25218 45556 25228
rect 44604 24546 44660 24556
rect 44940 25004 45220 25060
rect 44380 24098 44436 24108
rect 44940 24162 44996 25004
rect 45836 24834 45892 25228
rect 45836 24782 45838 24834
rect 45890 24782 45892 24834
rect 45836 24770 45892 24782
rect 45948 25172 46004 25182
rect 44940 24110 44942 24162
rect 44994 24110 44996 24162
rect 44940 24098 44996 24110
rect 45164 24722 45220 24734
rect 45164 24670 45166 24722
rect 45218 24670 45220 24722
rect 43932 23938 44324 23940
rect 43932 23886 43934 23938
rect 43986 23886 44324 23938
rect 43932 23884 44324 23886
rect 43932 23874 43988 23884
rect 43820 23538 43876 23548
rect 43708 23202 43764 23212
rect 43932 23044 43988 23054
rect 43932 22950 43988 22988
rect 44044 22930 44100 23884
rect 45052 23492 45108 23502
rect 44380 23044 44436 23054
rect 44380 22950 44436 22988
rect 44044 22878 44046 22930
rect 44098 22878 44100 22930
rect 44044 22866 44100 22878
rect 44604 22930 44660 22942
rect 44604 22878 44606 22930
rect 44658 22878 44660 22930
rect 43036 22540 43316 22596
rect 42924 21858 42980 21868
rect 43036 22372 43092 22382
rect 42700 21476 42756 21486
rect 42700 21382 42756 21420
rect 42364 20802 42532 20804
rect 42364 20750 42366 20802
rect 42418 20750 42532 20802
rect 42364 20748 42532 20750
rect 42364 20738 42420 20748
rect 42700 20580 42756 20590
rect 42252 20578 42756 20580
rect 42252 20526 42702 20578
rect 42754 20526 42756 20578
rect 42252 20524 42756 20526
rect 42140 20290 42196 20300
rect 41916 20076 42084 20132
rect 41916 19458 41972 20076
rect 42252 19906 42308 19918
rect 42252 19854 42254 19906
rect 42306 19854 42308 19906
rect 42140 19796 42196 19806
rect 42140 19702 42196 19740
rect 41916 19406 41918 19458
rect 41970 19406 41972 19458
rect 41916 19394 41972 19406
rect 42140 19460 42196 19470
rect 42140 19234 42196 19404
rect 42140 19182 42142 19234
rect 42194 19182 42196 19234
rect 42140 19170 42196 19182
rect 41692 17780 41748 17790
rect 41692 17106 41748 17724
rect 42252 17668 42308 19854
rect 42476 19796 42532 20524
rect 42700 20514 42756 20524
rect 43036 19796 43092 22316
rect 43148 22260 43204 22270
rect 43148 22166 43204 22204
rect 43260 20914 43316 22540
rect 43260 20862 43262 20914
rect 43314 20862 43316 20914
rect 42476 19730 42532 19740
rect 42812 19740 43092 19796
rect 43148 20018 43204 20030
rect 43148 19966 43150 20018
rect 43202 19966 43204 20018
rect 42700 19124 42756 19134
rect 42700 19030 42756 19068
rect 42812 18900 42868 19740
rect 42700 18844 42868 18900
rect 42924 19460 42980 19470
rect 42364 18676 42420 18686
rect 42364 18674 42644 18676
rect 42364 18622 42366 18674
rect 42418 18622 42644 18674
rect 42364 18620 42644 18622
rect 42364 18610 42420 18620
rect 42476 18450 42532 18462
rect 42476 18398 42478 18450
rect 42530 18398 42532 18450
rect 42364 18228 42420 18238
rect 42364 18134 42420 18172
rect 42476 18004 42532 18398
rect 42476 17938 42532 17948
rect 42476 17778 42532 17790
rect 42476 17726 42478 17778
rect 42530 17726 42532 17778
rect 42476 17668 42532 17726
rect 42252 17612 42532 17668
rect 41692 17054 41694 17106
rect 41746 17054 41748 17106
rect 41692 17042 41748 17054
rect 42364 17108 42420 17118
rect 42364 17014 42420 17052
rect 41580 16930 41636 16940
rect 42140 16994 42196 17006
rect 42140 16942 42142 16994
rect 42194 16942 42196 16994
rect 42028 16884 42084 16894
rect 42028 16790 42084 16828
rect 42140 16772 42196 16942
rect 42140 16706 42196 16716
rect 42252 16548 42308 16558
rect 41916 16436 41972 16446
rect 41916 16212 41972 16380
rect 41916 16210 42084 16212
rect 41916 16158 41918 16210
rect 41970 16158 42084 16210
rect 41916 16156 42084 16158
rect 41916 16146 41972 16156
rect 42028 15538 42084 16156
rect 42028 15486 42030 15538
rect 42082 15486 42084 15538
rect 42028 15474 42084 15486
rect 42252 15426 42308 16492
rect 42252 15374 42254 15426
rect 42306 15374 42308 15426
rect 42252 15362 42308 15374
rect 41468 15092 41972 15148
rect 41356 14924 41636 14980
rect 41356 14532 41412 14542
rect 41356 14438 41412 14476
rect 41468 14420 41524 14430
rect 41468 14326 41524 14364
rect 41580 13860 41636 14924
rect 41468 13858 41636 13860
rect 41468 13806 41582 13858
rect 41634 13806 41636 13858
rect 41468 13804 41636 13806
rect 41468 13076 41524 13804
rect 41580 13794 41636 13804
rect 41804 13524 41860 13534
rect 41468 13010 41524 13020
rect 41580 13522 41860 13524
rect 41580 13470 41806 13522
rect 41858 13470 41860 13522
rect 41580 13468 41860 13470
rect 41244 12226 41300 12236
rect 41468 12180 41524 12190
rect 41020 12124 41188 12180
rect 40460 11844 40516 11854
rect 40348 11396 40404 11406
rect 40348 11302 40404 11340
rect 40124 3442 40292 3444
rect 40124 3390 40126 3442
rect 40178 3390 40292 3442
rect 40124 3388 40292 3390
rect 40348 4226 40404 4238
rect 40348 4174 40350 4226
rect 40402 4174 40404 4226
rect 40348 3444 40404 4174
rect 40124 3378 40180 3388
rect 40348 3378 40404 3388
rect 40460 3442 40516 11788
rect 40796 11394 40852 11406
rect 40796 11342 40798 11394
rect 40850 11342 40852 11394
rect 40796 10500 40852 11342
rect 40908 10948 40964 12124
rect 41020 11954 41076 11966
rect 41020 11902 41022 11954
rect 41074 11902 41076 11954
rect 41020 11172 41076 11902
rect 41020 11106 41076 11116
rect 40908 10892 41076 10948
rect 40796 10434 40852 10444
rect 40908 9828 40964 9838
rect 40908 9154 40964 9772
rect 40908 9102 40910 9154
rect 40962 9102 40964 9154
rect 40908 9090 40964 9102
rect 41020 9268 41076 10892
rect 41132 10388 41188 12124
rect 41468 12086 41524 12124
rect 41580 11844 41636 13468
rect 41804 13458 41860 13468
rect 41804 13076 41860 13086
rect 41916 13076 41972 15092
rect 42028 14644 42084 14654
rect 42476 14644 42532 17612
rect 42588 17108 42644 18620
rect 42588 17042 42644 17052
rect 42588 16660 42644 16670
rect 42588 15652 42644 16604
rect 42700 16436 42756 18844
rect 42812 18004 42868 18014
rect 42812 17890 42868 17948
rect 42812 17838 42814 17890
rect 42866 17838 42868 17890
rect 42812 17826 42868 17838
rect 42924 17780 42980 19404
rect 43148 19348 43204 19966
rect 43148 19254 43204 19292
rect 43036 19236 43092 19246
rect 43036 18674 43092 19180
rect 43036 18622 43038 18674
rect 43090 18622 43092 18674
rect 43036 18610 43092 18622
rect 43260 18452 43316 20862
rect 43372 22540 43652 22596
rect 43372 19124 43428 22540
rect 44604 22484 44660 22878
rect 44940 22932 44996 22942
rect 44940 22838 44996 22876
rect 44940 22484 44996 22494
rect 44604 22482 44996 22484
rect 44604 22430 44942 22482
rect 44994 22430 44996 22482
rect 44604 22428 44996 22430
rect 44940 22418 44996 22428
rect 43596 22260 43652 22270
rect 43596 22166 43652 22204
rect 44044 22148 44100 22158
rect 44044 22054 44100 22092
rect 45052 22036 45108 23436
rect 44828 21474 44884 21486
rect 44828 21422 44830 21474
rect 44882 21422 44884 21474
rect 44268 20804 44324 20814
rect 44268 20710 44324 20748
rect 43708 20578 43764 20590
rect 43708 20526 43710 20578
rect 43762 20526 43764 20578
rect 43708 20132 43764 20526
rect 44828 20356 44884 21422
rect 45052 20914 45108 21980
rect 45164 21588 45220 24670
rect 45276 24164 45332 24174
rect 45276 24070 45332 24108
rect 45612 23826 45668 23838
rect 45612 23774 45614 23826
rect 45666 23774 45668 23826
rect 45612 23266 45668 23774
rect 45948 23826 46004 25116
rect 45948 23774 45950 23826
rect 46002 23774 46004 23826
rect 45948 23762 46004 23774
rect 45612 23214 45614 23266
rect 45666 23214 45668 23266
rect 45276 23156 45332 23166
rect 45276 23062 45332 23100
rect 45500 22932 45556 22942
rect 45500 22370 45556 22876
rect 45500 22318 45502 22370
rect 45554 22318 45556 22370
rect 45500 22306 45556 22318
rect 45388 21588 45444 21598
rect 45164 21586 45444 21588
rect 45164 21534 45390 21586
rect 45442 21534 45444 21586
rect 45164 21532 45444 21534
rect 45052 20862 45054 20914
rect 45106 20862 45108 20914
rect 45052 20850 45108 20862
rect 44828 20290 44884 20300
rect 43596 20076 43764 20132
rect 44940 20244 44996 20254
rect 43484 19236 43540 19246
rect 43484 19142 43540 19180
rect 43372 19058 43428 19068
rect 43260 18386 43316 18396
rect 43484 18340 43540 18350
rect 43596 18340 43652 20076
rect 43708 19908 43764 19918
rect 43708 19346 43764 19852
rect 44940 19906 44996 20188
rect 44940 19854 44942 19906
rect 44994 19854 44996 19906
rect 43708 19294 43710 19346
rect 43762 19294 43764 19346
rect 43708 19282 43764 19294
rect 44044 19460 44100 19470
rect 44044 19346 44100 19404
rect 44044 19294 44046 19346
rect 44098 19294 44100 19346
rect 44044 19282 44100 19294
rect 43932 19012 43988 19022
rect 44156 19012 44212 19022
rect 43540 18284 43652 18340
rect 43820 19010 43988 19012
rect 43820 18958 43934 19010
rect 43986 18958 43988 19010
rect 43820 18956 43988 18958
rect 43484 18246 43540 18284
rect 43596 17780 43652 17790
rect 42924 17778 43652 17780
rect 42924 17726 43598 17778
rect 43650 17726 43652 17778
rect 42924 17724 43652 17726
rect 42924 17554 42980 17724
rect 43596 17714 43652 17724
rect 43148 17556 43204 17566
rect 42924 17502 42926 17554
rect 42978 17502 42980 17554
rect 42924 17490 42980 17502
rect 43036 17554 43204 17556
rect 43036 17502 43150 17554
rect 43202 17502 43204 17554
rect 43036 17500 43204 17502
rect 42812 16994 42868 17006
rect 42812 16942 42814 16994
rect 42866 16942 42868 16994
rect 42812 16772 42868 16942
rect 42812 16548 42868 16716
rect 42924 16772 42980 16782
rect 43036 16772 43092 17500
rect 43148 17490 43204 17500
rect 43820 17444 43876 18956
rect 43932 18946 43988 18956
rect 44044 19010 44212 19012
rect 44044 18958 44158 19010
rect 44210 18958 44212 19010
rect 44044 18956 44212 18958
rect 43932 18676 43988 18686
rect 44044 18676 44100 18956
rect 44156 18946 44212 18956
rect 43932 18674 44100 18676
rect 43932 18622 43934 18674
rect 43986 18622 44100 18674
rect 43932 18620 44100 18622
rect 44604 18676 44660 18686
rect 43932 18610 43988 18620
rect 44156 18564 44212 18574
rect 44156 18470 44212 18508
rect 44268 18562 44324 18574
rect 44268 18510 44270 18562
rect 44322 18510 44324 18562
rect 44044 17780 44100 17790
rect 44044 17686 44100 17724
rect 44268 17668 44324 18510
rect 44268 17602 44324 17612
rect 43820 17378 43876 17388
rect 42924 16770 43036 16772
rect 42924 16718 42926 16770
rect 42978 16718 43036 16770
rect 42924 16716 43036 16718
rect 42924 16706 42980 16716
rect 43036 16678 43092 16716
rect 43148 17164 43540 17220
rect 42924 16548 42980 16558
rect 42812 16492 42924 16548
rect 42924 16482 42980 16492
rect 42700 16370 42756 16380
rect 43148 16212 43204 17164
rect 43484 17106 43540 17164
rect 43484 17054 43486 17106
rect 43538 17054 43540 17106
rect 43484 17042 43540 17054
rect 43260 16996 43316 17006
rect 43260 16770 43316 16940
rect 44044 16996 44100 17006
rect 44044 16902 44100 16940
rect 44604 16994 44660 18620
rect 44716 18564 44772 18574
rect 44716 18470 44772 18508
rect 44940 17780 44996 19854
rect 45164 19796 45220 19806
rect 45164 19234 45220 19740
rect 45164 19182 45166 19234
rect 45218 19182 45220 19234
rect 45164 19170 45220 19182
rect 44940 17714 44996 17724
rect 45052 18452 45108 18462
rect 45276 18452 45332 21532
rect 45388 21522 45444 21532
rect 45612 20804 45668 23214
rect 46060 23266 46116 26684
rect 46060 23214 46062 23266
rect 46114 23214 46116 23266
rect 46060 23202 46116 23214
rect 46396 26740 46452 26750
rect 46284 22372 46340 22382
rect 46284 22278 46340 22316
rect 45836 22148 45892 22158
rect 45836 22146 46116 22148
rect 45836 22094 45838 22146
rect 45890 22094 46116 22146
rect 45836 22092 46116 22094
rect 45836 22082 45892 22092
rect 46060 21698 46116 22092
rect 46060 21646 46062 21698
rect 46114 21646 46116 21698
rect 46060 21634 46116 21646
rect 45836 21028 45892 21038
rect 45836 20934 45892 20972
rect 45612 20738 45668 20748
rect 46284 20804 46340 20814
rect 45500 20692 45556 20702
rect 45500 20598 45556 20636
rect 46284 20130 46340 20748
rect 46396 20690 46452 26684
rect 46396 20638 46398 20690
rect 46450 20638 46452 20690
rect 46396 20580 46452 20638
rect 46396 20514 46452 20524
rect 46284 20078 46286 20130
rect 46338 20078 46340 20130
rect 46284 20066 46340 20078
rect 46508 19908 46564 31612
rect 46732 29204 46788 35532
rect 46956 35474 47012 35486
rect 46956 35422 46958 35474
rect 47010 35422 47012 35474
rect 46844 35252 46900 35262
rect 46844 34356 46900 35196
rect 46956 35140 47012 35422
rect 46956 35074 47012 35084
rect 46956 34914 47012 34926
rect 46956 34862 46958 34914
rect 47010 34862 47012 34914
rect 46956 34692 47012 34862
rect 46956 34626 47012 34636
rect 47180 34692 47236 34702
rect 46956 34356 47012 34366
rect 46844 34354 47012 34356
rect 46844 34302 46958 34354
rect 47010 34302 47012 34354
rect 46844 34300 47012 34302
rect 46956 34132 47012 34300
rect 47180 34244 47236 34636
rect 46956 34066 47012 34076
rect 47068 34242 47236 34244
rect 47068 34190 47182 34242
rect 47234 34190 47236 34242
rect 47068 34188 47236 34190
rect 46732 29138 46788 29148
rect 47068 28644 47124 34188
rect 47180 34178 47236 34188
rect 47292 34580 47348 34590
rect 46620 28588 47124 28644
rect 47180 29540 47236 29550
rect 46620 28530 46676 28588
rect 46620 28478 46622 28530
rect 46674 28478 46676 28530
rect 46620 28466 46676 28478
rect 46732 28418 46788 28430
rect 46732 28366 46734 28418
rect 46786 28366 46788 28418
rect 46732 28196 46788 28366
rect 46844 28418 46900 28430
rect 46844 28366 46846 28418
rect 46898 28366 46900 28418
rect 46844 28308 46900 28366
rect 46844 28242 46900 28252
rect 47180 28308 47236 29484
rect 47180 28242 47236 28252
rect 46732 28130 46788 28140
rect 46844 27860 46900 27870
rect 46844 26964 46900 27804
rect 46620 26908 46900 26964
rect 46956 26962 47012 26974
rect 46956 26910 46958 26962
rect 47010 26910 47012 26962
rect 46956 26908 47012 26910
rect 47292 26908 47348 34524
rect 47404 34132 47460 34142
rect 47404 34038 47460 34076
rect 47516 34018 47572 35644
rect 47628 35474 47684 35486
rect 47628 35422 47630 35474
rect 47682 35422 47684 35474
rect 47628 34244 47684 35422
rect 47964 35476 48020 35486
rect 47964 35382 48020 35420
rect 48076 34354 48132 35756
rect 48076 34302 48078 34354
rect 48130 34302 48132 34354
rect 48076 34290 48132 34302
rect 48188 35026 48244 36428
rect 48524 36372 48580 36382
rect 48188 34974 48190 35026
rect 48242 34974 48244 35026
rect 47964 34244 48020 34254
rect 47628 34242 47964 34244
rect 47628 34190 47630 34242
rect 47682 34190 47964 34242
rect 47628 34188 47964 34190
rect 47628 34178 47684 34188
rect 47964 34150 48020 34188
rect 48188 34132 48244 34974
rect 48300 36370 48580 36372
rect 48300 36318 48526 36370
rect 48578 36318 48580 36370
rect 48300 36316 48580 36318
rect 48300 34354 48356 36316
rect 48524 36306 48580 36316
rect 48636 36260 48692 36270
rect 48636 36166 48692 36204
rect 48748 35810 48804 36876
rect 49532 36708 49588 36718
rect 49532 36596 49588 36652
rect 51324 36706 51380 36988
rect 51324 36654 51326 36706
rect 51378 36654 51380 36706
rect 51324 36642 51380 36654
rect 49420 36594 49588 36596
rect 49420 36542 49534 36594
rect 49586 36542 49588 36594
rect 49420 36540 49588 36542
rect 48860 36372 48916 36382
rect 49084 36372 49140 36382
rect 48860 36370 49028 36372
rect 48860 36318 48862 36370
rect 48914 36318 49028 36370
rect 48860 36316 49028 36318
rect 48860 36306 48916 36316
rect 48748 35758 48750 35810
rect 48802 35758 48804 35810
rect 48748 35746 48804 35758
rect 48300 34302 48302 34354
rect 48354 34302 48356 34354
rect 48300 34290 48356 34302
rect 48860 35698 48916 35710
rect 48860 35646 48862 35698
rect 48914 35646 48916 35698
rect 48860 34354 48916 35646
rect 48860 34302 48862 34354
rect 48914 34302 48916 34354
rect 48860 34290 48916 34302
rect 48748 34244 48804 34254
rect 48748 34150 48804 34188
rect 47516 33966 47518 34018
rect 47570 33966 47572 34018
rect 47516 33954 47572 33966
rect 48076 34076 48244 34132
rect 48972 34132 49028 36316
rect 49084 36278 49140 36316
rect 47740 33572 47796 33582
rect 47740 33458 47796 33516
rect 47740 33406 47742 33458
rect 47794 33406 47796 33458
rect 47740 33394 47796 33406
rect 47964 32564 48020 32574
rect 48076 32564 48132 34076
rect 48020 32508 48132 32564
rect 48188 33346 48244 33358
rect 48188 33294 48190 33346
rect 48242 33294 48244 33346
rect 47964 32470 48020 32508
rect 47516 31892 47572 31902
rect 47516 31778 47572 31836
rect 48188 31892 48244 33294
rect 48188 31826 48244 31836
rect 48860 33234 48916 33246
rect 48860 33182 48862 33234
rect 48914 33182 48916 33234
rect 47516 31726 47518 31778
rect 47570 31726 47572 31778
rect 47516 30884 47572 31726
rect 48188 31668 48244 31678
rect 47964 31666 48244 31668
rect 47964 31614 48190 31666
rect 48242 31614 48244 31666
rect 47964 31612 48244 31614
rect 47852 31108 47908 31118
rect 47516 30818 47572 30828
rect 47740 31052 47852 31108
rect 47404 29428 47460 29438
rect 47404 29334 47460 29372
rect 47740 29316 47796 31052
rect 47852 31042 47908 31052
rect 47852 30882 47908 30894
rect 47852 30830 47854 30882
rect 47906 30830 47908 30882
rect 47852 30436 47908 30830
rect 47852 30370 47908 30380
rect 47964 29650 48020 31612
rect 48188 31602 48244 31612
rect 48860 31108 48916 33182
rect 48860 31042 48916 31052
rect 48860 30884 48916 30894
rect 48748 30210 48804 30222
rect 48748 30158 48750 30210
rect 48802 30158 48804 30210
rect 48188 30100 48244 30110
rect 48188 30006 48244 30044
rect 48748 30100 48804 30158
rect 48748 30034 48804 30044
rect 47964 29598 47966 29650
rect 48018 29598 48020 29650
rect 47964 29586 48020 29598
rect 47852 29540 47908 29550
rect 47852 29446 47908 29484
rect 48076 29426 48132 29438
rect 48076 29374 48078 29426
rect 48130 29374 48132 29426
rect 47740 29260 48020 29316
rect 47964 28754 48020 29260
rect 47964 28702 47966 28754
rect 48018 28702 48020 28754
rect 47964 28690 48020 28702
rect 48076 28756 48132 29374
rect 48524 28756 48580 28766
rect 48076 28754 48580 28756
rect 48076 28702 48526 28754
rect 48578 28702 48580 28754
rect 48076 28700 48580 28702
rect 47404 28644 47460 28654
rect 47404 28550 47460 28588
rect 47852 28418 47908 28430
rect 47852 28366 47854 28418
rect 47906 28366 47908 28418
rect 47852 27972 47908 28366
rect 48076 28418 48132 28700
rect 48524 28690 48580 28700
rect 48076 28366 48078 28418
rect 48130 28366 48132 28418
rect 48076 28308 48132 28366
rect 48076 28242 48132 28252
rect 48860 28084 48916 30828
rect 48860 27990 48916 28028
rect 47852 27906 47908 27916
rect 48636 27972 48692 27982
rect 48188 27746 48244 27758
rect 48188 27694 48190 27746
rect 48242 27694 48244 27746
rect 47740 27186 47796 27198
rect 47740 27134 47742 27186
rect 47794 27134 47796 27186
rect 46620 24050 46676 26908
rect 46956 26852 47124 26908
rect 47068 26066 47124 26852
rect 47068 26014 47070 26066
rect 47122 26014 47124 26066
rect 47068 26002 47124 26014
rect 47180 26852 47348 26908
rect 47516 26962 47572 26974
rect 47516 26910 47518 26962
rect 47570 26910 47572 26962
rect 46620 23998 46622 24050
rect 46674 23998 46676 24050
rect 46620 23492 46676 23998
rect 46620 23426 46676 23436
rect 46956 23938 47012 23950
rect 46956 23886 46958 23938
rect 47010 23886 47012 23938
rect 46956 23828 47012 23886
rect 46620 23156 46676 23166
rect 46620 23042 46676 23100
rect 46620 22990 46622 23042
rect 46674 22990 46676 23042
rect 46620 20804 46676 22990
rect 46620 20738 46676 20748
rect 46732 22146 46788 22158
rect 46732 22094 46734 22146
rect 46786 22094 46788 22146
rect 46732 20244 46788 22094
rect 46956 20356 47012 23772
rect 47068 23044 47124 23054
rect 47180 23044 47236 26852
rect 47292 26292 47348 26302
rect 47292 26178 47348 26236
rect 47292 26126 47294 26178
rect 47346 26126 47348 26178
rect 47292 26066 47348 26126
rect 47292 26014 47294 26066
rect 47346 26014 47348 26066
rect 47292 23156 47348 26014
rect 47516 25060 47572 26910
rect 47516 24994 47572 25004
rect 47628 26068 47684 26078
rect 47740 26068 47796 27134
rect 47852 27074 47908 27086
rect 47852 27022 47854 27074
rect 47906 27022 47908 27074
rect 47852 26402 47908 27022
rect 48188 26908 48244 27694
rect 48636 27074 48692 27916
rect 48636 27022 48638 27074
rect 48690 27022 48692 27074
rect 48636 27010 48692 27022
rect 48972 26908 49028 34076
rect 49196 35698 49252 35710
rect 49196 35646 49198 35698
rect 49250 35646 49252 35698
rect 49084 30322 49140 30334
rect 49084 30270 49086 30322
rect 49138 30270 49140 30322
rect 49084 30212 49140 30270
rect 49084 30146 49140 30156
rect 49084 29316 49140 29326
rect 49084 29222 49140 29260
rect 49196 26908 49252 35646
rect 49420 34130 49476 36540
rect 49532 36530 49588 36540
rect 49980 36596 50036 36606
rect 49980 36502 50036 36540
rect 50428 36596 50484 36606
rect 50428 36502 50484 36540
rect 50988 36596 51044 36606
rect 50652 36482 50708 36494
rect 50652 36430 50654 36482
rect 50706 36430 50708 36482
rect 50652 36260 50708 36430
rect 50988 36484 51044 36540
rect 50988 36482 51380 36484
rect 50988 36430 50990 36482
rect 51042 36430 51380 36482
rect 50988 36428 51380 36430
rect 50988 36418 51044 36428
rect 51212 36260 51268 36270
rect 50428 36204 50708 36260
rect 50988 36258 51268 36260
rect 50988 36206 51214 36258
rect 51266 36206 51268 36258
rect 50988 36204 51268 36206
rect 50092 35812 50148 35822
rect 50092 35718 50148 35756
rect 50316 35698 50372 35710
rect 50316 35646 50318 35698
rect 50370 35646 50372 35698
rect 50316 35476 50372 35646
rect 50316 35410 50372 35420
rect 50428 35588 50484 36204
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50988 35924 51044 36204
rect 51212 36194 51268 36204
rect 50428 35308 50484 35532
rect 50316 35252 50484 35308
rect 50540 35868 51044 35924
rect 51324 35922 51380 36428
rect 51324 35870 51326 35922
rect 51378 35870 51380 35922
rect 49980 34802 50036 34814
rect 49980 34750 49982 34802
rect 50034 34750 50036 34802
rect 49868 34692 49924 34702
rect 49868 34598 49924 34636
rect 49980 34244 50036 34750
rect 50204 34804 50260 34814
rect 50204 34354 50260 34748
rect 50204 34302 50206 34354
rect 50258 34302 50260 34354
rect 50204 34290 50260 34302
rect 49420 34078 49422 34130
rect 49474 34078 49476 34130
rect 49420 33908 49476 34078
rect 49756 34188 50036 34244
rect 49756 34132 49812 34188
rect 49756 34066 49812 34076
rect 49868 34018 49924 34030
rect 49868 33966 49870 34018
rect 49922 33966 49924 34018
rect 49868 33908 49924 33966
rect 49420 33852 49924 33908
rect 50204 33684 50260 33694
rect 50316 33684 50372 35252
rect 50540 34692 50596 35868
rect 51324 35858 51380 35870
rect 51436 36482 51492 36494
rect 51436 36430 51438 36482
rect 51490 36430 51492 36482
rect 50988 35698 51044 35710
rect 50988 35646 50990 35698
rect 51042 35646 51044 35698
rect 50652 35364 50708 35374
rect 50652 34914 50708 35308
rect 50652 34862 50654 34914
rect 50706 34862 50708 34914
rect 50652 34850 50708 34862
rect 50988 34914 51044 35646
rect 50988 34862 50990 34914
rect 51042 34862 51044 34914
rect 50260 33628 50372 33684
rect 50428 34690 50596 34692
rect 50428 34638 50542 34690
rect 50594 34638 50596 34690
rect 50428 34636 50596 34638
rect 49420 31668 49476 31678
rect 49420 31220 49476 31612
rect 50092 31556 50148 31566
rect 49420 31218 49812 31220
rect 49420 31166 49422 31218
rect 49474 31166 49812 31218
rect 49420 31164 49812 31166
rect 49420 31154 49476 31164
rect 49756 30994 49812 31164
rect 49756 30942 49758 30994
rect 49810 30942 49812 30994
rect 49756 30930 49812 30942
rect 49644 30436 49700 30446
rect 49644 30322 49700 30380
rect 49644 30270 49646 30322
rect 49698 30270 49700 30322
rect 49644 30258 49700 30270
rect 50092 30210 50148 31500
rect 50092 30158 50094 30210
rect 50146 30158 50148 30210
rect 50092 30146 50148 30158
rect 49756 29988 49812 29998
rect 49756 29426 49812 29932
rect 49756 29374 49758 29426
rect 49810 29374 49812 29426
rect 49756 29362 49812 29374
rect 49980 29428 50036 29438
rect 49980 29334 50036 29372
rect 49868 28756 49924 28766
rect 49868 28662 49924 28700
rect 49980 28082 50036 28094
rect 49980 28030 49982 28082
rect 50034 28030 50036 28082
rect 49980 27972 50036 28030
rect 49980 27906 50036 27916
rect 50204 26908 50260 33628
rect 50316 32452 50372 32462
rect 50316 31890 50372 32396
rect 50316 31838 50318 31890
rect 50370 31838 50372 31890
rect 50316 31826 50372 31838
rect 50428 30212 50484 34636
rect 50540 34626 50596 34636
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50988 34356 51044 34862
rect 51100 35700 51156 35710
rect 51100 34690 51156 35644
rect 51324 34916 51380 34926
rect 51436 34916 51492 36430
rect 51660 35922 51716 37214
rect 51772 37266 51828 37278
rect 51772 37214 51774 37266
rect 51826 37214 51828 37266
rect 51772 36258 51828 37214
rect 51772 36206 51774 36258
rect 51826 36206 51828 36258
rect 51772 36194 51828 36206
rect 51884 36370 51940 36382
rect 51884 36318 51886 36370
rect 51938 36318 51940 36370
rect 51660 35870 51662 35922
rect 51714 35870 51716 35922
rect 51660 35858 51716 35870
rect 51548 35810 51604 35822
rect 51548 35758 51550 35810
rect 51602 35758 51604 35810
rect 51548 35028 51604 35758
rect 51772 35698 51828 35710
rect 51772 35646 51774 35698
rect 51826 35646 51828 35698
rect 51772 35476 51828 35646
rect 51772 35410 51828 35420
rect 51548 34962 51604 34972
rect 51324 34914 51492 34916
rect 51324 34862 51326 34914
rect 51378 34862 51492 34914
rect 51324 34860 51492 34862
rect 51660 34916 51716 34926
rect 51324 34850 51380 34860
rect 51660 34822 51716 34860
rect 51772 34916 51828 34926
rect 51884 34916 51940 36318
rect 51996 35700 52052 37548
rect 52220 37380 52276 37774
rect 52444 37490 52500 38612
rect 52444 37438 52446 37490
rect 52498 37438 52500 37490
rect 52444 37426 52500 37438
rect 52556 37492 52612 38782
rect 52780 38052 52836 39676
rect 53228 39730 53284 41132
rect 53228 39678 53230 39730
rect 53282 39678 53284 39730
rect 53228 39666 53284 39678
rect 53340 40516 53396 40526
rect 53228 39060 53284 39070
rect 53340 39060 53396 40460
rect 53452 40404 53508 40414
rect 53452 40310 53508 40348
rect 53564 40180 53620 43484
rect 54572 43204 54628 44942
rect 54908 44436 54964 45950
rect 57708 46002 57764 46014
rect 57708 45950 57710 46002
rect 57762 45950 57764 46002
rect 55804 45890 55860 45902
rect 55804 45838 55806 45890
rect 55858 45838 55860 45890
rect 55132 45108 55188 45118
rect 55468 45108 55524 45118
rect 55132 45106 55524 45108
rect 55132 45054 55134 45106
rect 55186 45054 55470 45106
rect 55522 45054 55524 45106
rect 55132 45052 55524 45054
rect 54908 44370 54964 44380
rect 55020 44434 55076 44446
rect 55020 44382 55022 44434
rect 55074 44382 55076 44434
rect 54572 43138 54628 43148
rect 55020 43092 55076 44382
rect 55020 43026 55076 43036
rect 54796 42754 54852 42766
rect 54796 42702 54798 42754
rect 54850 42702 54852 42754
rect 53676 42642 53732 42654
rect 53676 42590 53678 42642
rect 53730 42590 53732 42642
rect 53676 41300 53732 42590
rect 53676 41234 53732 41244
rect 54796 41188 54852 42702
rect 55132 41972 55188 45052
rect 55468 45042 55524 45052
rect 55692 44322 55748 44334
rect 55692 44270 55694 44322
rect 55746 44270 55748 44322
rect 55132 41906 55188 41916
rect 55356 43314 55412 43326
rect 55356 43262 55358 43314
rect 55410 43262 55412 43314
rect 55244 41858 55300 41870
rect 55244 41806 55246 41858
rect 55298 41806 55300 41858
rect 54796 41122 54852 41132
rect 55020 41298 55076 41310
rect 55020 41246 55022 41298
rect 55074 41246 55076 41298
rect 53564 40114 53620 40124
rect 53228 39058 53396 39060
rect 53228 39006 53230 39058
rect 53282 39006 53396 39058
rect 53228 39004 53396 39006
rect 55020 39060 55076 41246
rect 55244 39844 55300 41806
rect 55356 41748 55412 43262
rect 55580 42754 55636 42766
rect 55580 42702 55582 42754
rect 55634 42702 55636 42754
rect 55580 42308 55636 42702
rect 55580 42242 55636 42252
rect 55356 41682 55412 41692
rect 55244 39778 55300 39788
rect 55356 40292 55412 40302
rect 55356 39730 55412 40236
rect 55580 40292 55636 40302
rect 55692 40292 55748 44270
rect 55804 40404 55860 45838
rect 57372 42642 57428 42654
rect 57372 42590 57374 42642
rect 57426 42590 57428 42642
rect 55804 40338 55860 40348
rect 55916 41186 55972 41198
rect 55916 41134 55918 41186
rect 55970 41134 55972 41186
rect 55580 40290 55748 40292
rect 55580 40238 55582 40290
rect 55634 40238 55748 40290
rect 55580 40236 55748 40238
rect 55580 40226 55636 40236
rect 55356 39678 55358 39730
rect 55410 39678 55412 39730
rect 55356 39666 55412 39678
rect 53228 38994 53284 39004
rect 55020 38994 55076 39004
rect 53004 38948 53060 38958
rect 53004 38854 53060 38892
rect 52892 38834 52948 38846
rect 52892 38782 52894 38834
rect 52946 38782 52948 38834
rect 52892 38668 52948 38782
rect 53452 38836 53508 38846
rect 53452 38742 53508 38780
rect 52892 38612 53284 38668
rect 53004 38052 53060 38062
rect 52780 38050 53060 38052
rect 52780 37998 53006 38050
rect 53058 37998 53060 38050
rect 52780 37996 53060 37998
rect 52556 37436 52948 37492
rect 52220 37286 52276 37324
rect 52668 37266 52724 37278
rect 52668 37214 52670 37266
rect 52722 37214 52724 37266
rect 52556 37154 52612 37166
rect 52556 37102 52558 37154
rect 52610 37102 52612 37154
rect 52556 36596 52612 37102
rect 52668 37044 52724 37214
rect 52668 36978 52724 36988
rect 52780 37266 52836 37278
rect 52780 37214 52782 37266
rect 52834 37214 52836 37266
rect 52556 36530 52612 36540
rect 52780 36594 52836 37214
rect 52780 36542 52782 36594
rect 52834 36542 52836 36594
rect 52780 36530 52836 36542
rect 52108 36372 52164 36382
rect 52108 36278 52164 36316
rect 52668 36370 52724 36382
rect 52668 36318 52670 36370
rect 52722 36318 52724 36370
rect 52220 36036 52276 36046
rect 52220 35922 52276 35980
rect 52220 35870 52222 35922
rect 52274 35870 52276 35922
rect 52108 35700 52164 35710
rect 51996 35644 52108 35700
rect 52108 35634 52164 35644
rect 51996 35476 52052 35486
rect 52052 35420 52164 35476
rect 51996 35410 52052 35420
rect 51772 34914 51940 34916
rect 51772 34862 51774 34914
rect 51826 34862 51940 34914
rect 51772 34860 51940 34862
rect 51996 35028 52052 35038
rect 51100 34638 51102 34690
rect 51154 34638 51156 34690
rect 51100 34626 51156 34638
rect 51548 34690 51604 34702
rect 51548 34638 51550 34690
rect 51602 34638 51604 34690
rect 51324 34356 51380 34366
rect 51548 34356 51604 34638
rect 50652 34354 51604 34356
rect 50652 34302 51326 34354
rect 51378 34302 51604 34354
rect 50652 34300 51604 34302
rect 50652 34130 50708 34300
rect 51324 34290 51380 34300
rect 51772 34244 51828 34860
rect 51996 34804 52052 34972
rect 52108 34914 52164 35420
rect 52108 34862 52110 34914
rect 52162 34862 52164 34914
rect 52108 34850 52164 34862
rect 52220 35364 52276 35870
rect 52668 35922 52724 36318
rect 52892 36036 52948 37436
rect 53004 37044 53060 37996
rect 53116 37044 53172 37054
rect 53004 36988 53116 37044
rect 53116 36978 53172 36988
rect 53116 36482 53172 36494
rect 53116 36430 53118 36482
rect 53170 36430 53172 36482
rect 52668 35870 52670 35922
rect 52722 35870 52724 35922
rect 52668 35858 52724 35870
rect 52780 35980 52948 36036
rect 53004 36370 53060 36382
rect 53004 36318 53006 36370
rect 53058 36318 53060 36370
rect 53004 36036 53060 36318
rect 53116 36372 53172 36430
rect 53116 36306 53172 36316
rect 52444 35698 52500 35710
rect 52780 35700 52836 35980
rect 53004 35970 53060 35980
rect 52892 35812 52948 35822
rect 52892 35718 52948 35756
rect 52444 35646 52446 35698
rect 52498 35646 52500 35698
rect 50652 34078 50654 34130
rect 50706 34078 50708 34130
rect 50652 34066 50708 34078
rect 50876 34188 51268 34244
rect 50876 34130 50932 34188
rect 50876 34078 50878 34130
rect 50930 34078 50932 34130
rect 50876 34066 50932 34078
rect 51212 34132 51268 34188
rect 51436 34188 51828 34244
rect 51884 34748 52052 34804
rect 51436 34132 51492 34188
rect 51212 34076 51492 34132
rect 50988 34020 51044 34030
rect 50988 33458 51044 33964
rect 50988 33406 50990 33458
rect 51042 33406 51044 33458
rect 50988 33394 51044 33406
rect 51100 34018 51156 34030
rect 51100 33966 51102 34018
rect 51154 33966 51156 34018
rect 51100 33236 51156 33966
rect 51436 33460 51492 33470
rect 51436 33366 51492 33404
rect 51324 33236 51380 33246
rect 51100 33234 51380 33236
rect 51100 33182 51326 33234
rect 51378 33182 51380 33234
rect 51100 33180 51380 33182
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50540 32788 50596 32798
rect 50540 32694 50596 32732
rect 51324 32564 51380 33180
rect 51660 32676 51716 34188
rect 51772 33908 51828 33918
rect 51772 33814 51828 33852
rect 51884 33684 51940 34748
rect 52220 34692 52276 35308
rect 51996 34636 52276 34692
rect 52332 35586 52388 35598
rect 52332 35534 52334 35586
rect 52386 35534 52388 35586
rect 51996 34130 52052 34636
rect 51996 34078 51998 34130
rect 52050 34078 52052 34130
rect 51996 34020 52052 34078
rect 52332 34132 52388 35534
rect 52444 35588 52500 35646
rect 52444 35522 52500 35532
rect 52668 35644 52836 35700
rect 53004 35698 53060 35710
rect 53004 35646 53006 35698
rect 53058 35646 53060 35698
rect 52668 35026 52724 35644
rect 53004 35588 53060 35646
rect 53004 35522 53060 35532
rect 52668 34974 52670 35026
rect 52722 34974 52724 35026
rect 52668 34962 52724 34974
rect 52780 34916 52836 34926
rect 52780 34822 52836 34860
rect 53228 34692 53284 38612
rect 55356 38610 55412 38622
rect 55356 38558 55358 38610
rect 55410 38558 55412 38610
rect 53788 37938 53844 37950
rect 53788 37886 53790 37938
rect 53842 37886 53844 37938
rect 53788 37268 53844 37886
rect 53788 37202 53844 37212
rect 53788 37044 53844 37054
rect 53788 36482 53844 36988
rect 55020 37042 55076 37054
rect 55020 36990 55022 37042
rect 55074 36990 55076 37042
rect 54460 36596 54516 36606
rect 54460 36502 54516 36540
rect 53788 36430 53790 36482
rect 53842 36430 53844 36482
rect 53452 35700 53508 35710
rect 53452 35606 53508 35644
rect 53788 35028 53844 36430
rect 55020 35700 55076 36990
rect 55356 37044 55412 38558
rect 55916 38162 55972 41134
rect 56588 40628 56644 40638
rect 56588 40534 56644 40572
rect 57148 40516 57204 40526
rect 56812 40402 56868 40414
rect 56812 40350 56814 40402
rect 56866 40350 56868 40402
rect 56028 40290 56084 40302
rect 56028 40238 56030 40290
rect 56082 40238 56084 40290
rect 56028 39732 56084 40238
rect 56700 40292 56756 40302
rect 56700 40198 56756 40236
rect 56028 39618 56084 39676
rect 56028 39566 56030 39618
rect 56082 39566 56084 39618
rect 56028 39554 56084 39566
rect 56588 39396 56644 39406
rect 56812 39396 56868 40350
rect 57148 40402 57204 40460
rect 57148 40350 57150 40402
rect 57202 40350 57204 40402
rect 57148 40338 57204 40350
rect 56644 39340 56868 39396
rect 56588 39302 56644 39340
rect 56700 38948 56756 38958
rect 56700 38854 56756 38892
rect 57372 38388 57428 42590
rect 57708 42420 57764 45950
rect 57708 42354 57764 42364
rect 57820 44434 57876 44446
rect 57820 44382 57822 44434
rect 57874 44382 57876 44434
rect 57820 40404 57876 44382
rect 57932 43764 57988 47518
rect 57932 43698 57988 43708
rect 57820 40338 57876 40348
rect 57932 41298 57988 41310
rect 57932 41246 57934 41298
rect 57986 41246 57988 41298
rect 57372 38322 57428 38332
rect 55916 38110 55918 38162
rect 55970 38110 55972 38162
rect 55916 38098 55972 38110
rect 57932 37716 57988 41246
rect 57932 37650 57988 37660
rect 56028 37268 56084 37278
rect 56028 37266 56644 37268
rect 56028 37214 56030 37266
rect 56082 37214 56644 37266
rect 56028 37212 56644 37214
rect 56028 37202 56084 37212
rect 55356 36978 55412 36988
rect 56588 36594 56644 37212
rect 56588 36542 56590 36594
rect 56642 36542 56644 36594
rect 56588 36530 56644 36542
rect 58044 36372 58100 36382
rect 55020 35634 55076 35644
rect 55580 35924 55636 35934
rect 55356 35474 55412 35486
rect 55356 35422 55358 35474
rect 55410 35422 55412 35474
rect 54124 35028 54180 35038
rect 53788 35026 54180 35028
rect 53788 34974 54126 35026
rect 54178 34974 54180 35026
rect 53788 34972 54180 34974
rect 54124 34962 54180 34972
rect 55356 35028 55412 35422
rect 55356 34962 55412 34972
rect 53340 34916 53396 34926
rect 53340 34914 53620 34916
rect 53340 34862 53342 34914
rect 53394 34862 53620 34914
rect 53340 34860 53620 34862
rect 53340 34850 53396 34860
rect 52780 34636 53284 34692
rect 52780 34242 52836 34636
rect 52780 34190 52782 34242
rect 52834 34190 52836 34242
rect 52780 34178 52836 34190
rect 52332 34076 52724 34132
rect 51996 33954 52052 33964
rect 52220 34018 52276 34030
rect 52220 33966 52222 34018
rect 52274 33966 52276 34018
rect 51884 33618 51940 33628
rect 52220 33572 52276 33966
rect 52668 34020 52724 34076
rect 52892 34130 52948 34142
rect 53228 34132 53284 34142
rect 52892 34078 52894 34130
rect 52946 34078 52948 34130
rect 52892 34020 52948 34078
rect 52668 33964 52948 34020
rect 53004 34130 53284 34132
rect 53004 34078 53230 34130
rect 53282 34078 53284 34130
rect 53004 34076 53284 34078
rect 52220 33506 52276 33516
rect 52556 33684 52612 33694
rect 51884 33122 51940 33134
rect 51884 33070 51886 33122
rect 51938 33070 51940 33122
rect 51884 32788 51940 33070
rect 52556 32788 52612 33628
rect 52668 33572 52724 33582
rect 52668 33346 52724 33516
rect 52668 33294 52670 33346
rect 52722 33294 52724 33346
rect 52668 33282 52724 33294
rect 52780 33572 52836 33582
rect 53004 33572 53060 34076
rect 53228 34066 53284 34076
rect 52780 33570 53060 33572
rect 52780 33518 52782 33570
rect 52834 33518 53060 33570
rect 52780 33516 53060 33518
rect 51940 32732 52052 32788
rect 51884 32722 51940 32732
rect 51772 32676 51828 32686
rect 51716 32674 51828 32676
rect 51716 32622 51774 32674
rect 51826 32622 51828 32674
rect 51716 32620 51828 32622
rect 51660 32582 51716 32620
rect 51772 32610 51828 32620
rect 51884 32564 51940 32574
rect 51324 32508 51492 32564
rect 50876 31780 50932 31790
rect 50876 31686 50932 31724
rect 50988 31556 51044 31566
rect 50988 31554 51380 31556
rect 50988 31502 50990 31554
rect 51042 31502 51380 31554
rect 50988 31500 51380 31502
rect 50988 31490 51044 31500
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50316 30156 50484 30212
rect 50988 30212 51044 30222
rect 50316 27972 50372 30156
rect 50540 30100 50596 30110
rect 50428 30044 50540 30100
rect 50428 29652 50484 30044
rect 50540 30006 50596 30044
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50428 29596 50596 29652
rect 50428 28644 50484 28654
rect 50428 28550 50484 28588
rect 50540 28420 50596 29596
rect 50988 29650 51044 30156
rect 50988 29598 50990 29650
rect 51042 29598 51044 29650
rect 50988 29586 51044 29598
rect 51212 30100 51268 30110
rect 51212 29538 51268 30044
rect 51212 29486 51214 29538
rect 51266 29486 51268 29538
rect 51212 29474 51268 29486
rect 50876 29428 50932 29438
rect 50876 28756 50932 29372
rect 51324 29426 51380 31500
rect 51436 30436 51492 32508
rect 51884 32002 51940 32508
rect 51884 31950 51886 32002
rect 51938 31950 51940 32002
rect 51884 31938 51940 31950
rect 51436 30370 51492 30380
rect 51548 31890 51604 31902
rect 51548 31838 51550 31890
rect 51602 31838 51604 31890
rect 51548 31780 51604 31838
rect 51548 30210 51604 31724
rect 51996 30884 52052 32732
rect 52556 32786 52724 32788
rect 52556 32734 52558 32786
rect 52610 32734 52724 32786
rect 52556 32732 52724 32734
rect 52556 32722 52612 32732
rect 52220 32564 52276 32574
rect 52220 32470 52276 32508
rect 52556 31780 52612 31790
rect 52556 31686 52612 31724
rect 51996 30790 52052 30828
rect 52108 31666 52164 31678
rect 52108 31614 52110 31666
rect 52162 31614 52164 31666
rect 52108 30324 52164 31614
rect 52108 30258 52164 30268
rect 52220 30548 52276 30558
rect 51548 30158 51550 30210
rect 51602 30158 51604 30210
rect 51548 30146 51604 30158
rect 51996 30100 52052 30110
rect 52220 30100 52276 30492
rect 52668 30212 52724 32732
rect 51996 30006 52052 30044
rect 52108 30044 52276 30100
rect 52556 30210 52724 30212
rect 52556 30158 52670 30210
rect 52722 30158 52724 30210
rect 52556 30156 52724 30158
rect 51436 29988 51492 29998
rect 51492 29932 51604 29988
rect 51436 29894 51492 29932
rect 51324 29374 51326 29426
rect 51378 29374 51380 29426
rect 51324 29362 51380 29374
rect 51324 28756 51380 28766
rect 50876 28754 51380 28756
rect 50876 28702 51326 28754
rect 51378 28702 51380 28754
rect 50876 28700 51380 28702
rect 51324 28690 51380 28700
rect 50316 27906 50372 27916
rect 50428 28364 50596 28420
rect 50764 28642 50820 28654
rect 50764 28590 50766 28642
rect 50818 28590 50820 28642
rect 50764 28420 50820 28590
rect 51436 28532 51492 28542
rect 51436 28438 51492 28476
rect 51212 28420 51268 28430
rect 50764 28418 51268 28420
rect 50764 28366 51214 28418
rect 51266 28366 51268 28418
rect 50764 28364 51268 28366
rect 50428 27970 50484 28364
rect 51212 28308 51268 28364
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50428 27918 50430 27970
rect 50482 27918 50484 27970
rect 50428 27906 50484 27918
rect 51212 27298 51268 28252
rect 51548 27858 51604 29932
rect 51996 29426 52052 29438
rect 51996 29374 51998 29426
rect 52050 29374 52052 29426
rect 51996 29316 52052 29374
rect 51884 29260 51996 29316
rect 51884 28642 51940 29260
rect 51996 29250 52052 29260
rect 51884 28590 51886 28642
rect 51938 28590 51940 28642
rect 51884 28578 51940 28590
rect 52108 27972 52164 30044
rect 52444 29988 52500 29998
rect 52444 29650 52500 29932
rect 52444 29598 52446 29650
rect 52498 29598 52500 29650
rect 52444 29586 52500 29598
rect 52556 29650 52612 30156
rect 52668 30146 52724 30156
rect 52780 30212 52836 33516
rect 53228 33460 53284 33470
rect 53564 33460 53620 34860
rect 55580 34914 55636 35868
rect 55580 34862 55582 34914
rect 55634 34862 55636 34914
rect 55580 34850 55636 34862
rect 57932 35026 57988 35038
rect 57932 34974 57934 35026
rect 57986 34974 57988 35026
rect 57932 34356 57988 34974
rect 57932 34290 57988 34300
rect 57932 33572 57988 33582
rect 58044 33572 58100 36316
rect 57932 33570 58100 33572
rect 57932 33518 57934 33570
rect 57986 33518 58100 33570
rect 57932 33516 58100 33518
rect 57932 33506 57988 33516
rect 53284 33404 53396 33460
rect 53228 33394 53284 33404
rect 53228 33122 53284 33134
rect 53228 33070 53230 33122
rect 53282 33070 53284 33122
rect 53228 32788 53284 33070
rect 53228 32722 53284 32732
rect 53116 32452 53172 32462
rect 52892 32450 53172 32452
rect 52892 32398 53118 32450
rect 53170 32398 53172 32450
rect 52892 32396 53172 32398
rect 52892 31556 52948 32396
rect 53116 32386 53172 32396
rect 53228 31780 53284 31790
rect 53340 31780 53396 33404
rect 53564 33394 53620 33404
rect 55580 33346 55636 33358
rect 55580 33294 55582 33346
rect 55634 33294 55636 33346
rect 54460 33234 54516 33246
rect 54460 33182 54462 33234
rect 54514 33182 54516 33234
rect 53228 31778 53396 31780
rect 53228 31726 53230 31778
rect 53282 31726 53396 31778
rect 53228 31724 53396 31726
rect 53788 32228 53844 32238
rect 53788 31778 53844 32172
rect 54348 31892 54404 31902
rect 54460 31892 54516 33182
rect 54572 33124 54628 33134
rect 55356 33124 55412 33134
rect 55580 33124 55636 33294
rect 54572 33122 55300 33124
rect 54572 33070 54574 33122
rect 54626 33070 55300 33122
rect 54572 33068 55300 33070
rect 54572 33058 54628 33068
rect 55244 32674 55300 33068
rect 55412 33068 55636 33124
rect 55356 33030 55412 33068
rect 55244 32622 55246 32674
rect 55298 32622 55300 32674
rect 55244 32610 55300 32622
rect 55916 32788 55972 32798
rect 55916 32562 55972 32732
rect 55916 32510 55918 32562
rect 55970 32510 55972 32562
rect 55916 32498 55972 32510
rect 54348 31890 54516 31892
rect 54348 31838 54350 31890
rect 54402 31838 54516 31890
rect 54348 31836 54516 31838
rect 54348 31826 54404 31836
rect 53788 31726 53790 31778
rect 53842 31726 53844 31778
rect 52892 31490 52948 31500
rect 53004 31554 53060 31566
rect 53004 31502 53006 31554
rect 53058 31502 53060 31554
rect 53004 31332 53060 31502
rect 53004 31266 53060 31276
rect 53116 31554 53172 31566
rect 53116 31502 53118 31554
rect 53170 31502 53172 31554
rect 53004 30996 53060 31006
rect 52780 30146 52836 30156
rect 52892 30994 53060 30996
rect 52892 30942 53006 30994
rect 53058 30942 53060 30994
rect 52892 30940 53060 30942
rect 52780 29988 52836 29998
rect 52780 29894 52836 29932
rect 52556 29598 52558 29650
rect 52610 29598 52612 29650
rect 52556 29540 52612 29598
rect 52892 29540 52948 30940
rect 53004 30930 53060 30940
rect 53116 30882 53172 31502
rect 53116 30830 53118 30882
rect 53170 30830 53172 30882
rect 53116 30818 53172 30830
rect 53004 30772 53060 30782
rect 53004 30678 53060 30716
rect 53228 30210 53284 31724
rect 53788 31714 53844 31726
rect 55020 31778 55076 31790
rect 55020 31726 55022 31778
rect 55074 31726 55076 31778
rect 55020 31668 55076 31726
rect 55020 31602 55076 31612
rect 54012 31554 54068 31566
rect 54012 31502 54014 31554
rect 54066 31502 54068 31554
rect 53228 30158 53230 30210
rect 53282 30158 53284 30210
rect 53228 30146 53284 30158
rect 53340 31332 53396 31342
rect 53004 30100 53060 30110
rect 53004 30006 53060 30044
rect 53340 30098 53396 31276
rect 53676 30996 53732 31006
rect 53564 30994 53732 30996
rect 53564 30942 53678 30994
rect 53730 30942 53732 30994
rect 53564 30940 53732 30942
rect 53564 30210 53620 30940
rect 53676 30930 53732 30940
rect 54012 30548 54068 31502
rect 54236 31554 54292 31566
rect 54236 31502 54238 31554
rect 54290 31502 54292 31554
rect 54236 31332 54292 31502
rect 54348 31556 54404 31566
rect 54348 31554 54516 31556
rect 54348 31502 54350 31554
rect 54402 31502 54516 31554
rect 54348 31500 54516 31502
rect 54348 31490 54404 31500
rect 54292 31276 54404 31332
rect 54236 31266 54292 31276
rect 54348 31106 54404 31276
rect 54460 31220 54516 31500
rect 54796 31554 54852 31566
rect 54796 31502 54798 31554
rect 54850 31502 54852 31554
rect 54796 31332 54852 31502
rect 54796 31266 54852 31276
rect 55692 31554 55748 31566
rect 55692 31502 55694 31554
rect 55746 31502 55748 31554
rect 54460 31154 54516 31164
rect 54908 31220 54964 31230
rect 54908 31126 54964 31164
rect 55692 31220 55748 31502
rect 55692 31154 55748 31164
rect 56364 31220 56420 31230
rect 54348 31054 54350 31106
rect 54402 31054 54404 31106
rect 54348 31042 54404 31054
rect 54572 30994 54628 31006
rect 54572 30942 54574 30994
rect 54626 30942 54628 30994
rect 54572 30548 54628 30942
rect 54684 30996 54740 31006
rect 54684 30902 54740 30940
rect 54796 30994 54852 31006
rect 54796 30942 54798 30994
rect 54850 30942 54852 30994
rect 54012 30492 54628 30548
rect 53564 30158 53566 30210
rect 53618 30158 53620 30210
rect 53564 30146 53620 30158
rect 54236 30212 54292 30222
rect 53340 30046 53342 30098
rect 53394 30046 53396 30098
rect 53340 30034 53396 30046
rect 54124 30100 54180 30110
rect 54124 30006 54180 30044
rect 54012 29764 54068 29774
rect 53116 29652 53172 29662
rect 53116 29650 53732 29652
rect 53116 29598 53118 29650
rect 53170 29598 53732 29650
rect 53116 29596 53732 29598
rect 53116 29586 53172 29596
rect 52556 29474 52612 29484
rect 52780 29484 52948 29540
rect 52220 29426 52276 29438
rect 52220 29374 52222 29426
rect 52274 29374 52276 29426
rect 52220 28084 52276 29374
rect 52556 29314 52612 29326
rect 52556 29262 52558 29314
rect 52610 29262 52612 29314
rect 52556 29204 52612 29262
rect 52780 29204 52836 29484
rect 53228 29426 53284 29438
rect 53228 29374 53230 29426
rect 53282 29374 53284 29426
rect 52556 29148 52836 29204
rect 52892 29204 52948 29214
rect 53116 29204 53172 29214
rect 52892 28644 52948 29148
rect 52892 28530 52948 28588
rect 52892 28478 52894 28530
rect 52946 28478 52948 28530
rect 52892 28466 52948 28478
rect 53004 29202 53172 29204
rect 53004 29150 53118 29202
rect 53170 29150 53172 29202
rect 53004 29148 53172 29150
rect 53004 28532 53060 29148
rect 53116 29138 53172 29148
rect 52668 28418 52724 28430
rect 52668 28366 52670 28418
rect 52722 28366 52724 28418
rect 52668 28308 52724 28366
rect 52780 28420 52836 28430
rect 52780 28326 52836 28364
rect 52668 28242 52724 28252
rect 52220 28028 52836 28084
rect 52108 27916 52388 27972
rect 51548 27806 51550 27858
rect 51602 27806 51604 27858
rect 51548 27794 51604 27806
rect 51996 27860 52052 27870
rect 51996 27858 52164 27860
rect 51996 27806 51998 27858
rect 52050 27806 52164 27858
rect 51996 27804 52164 27806
rect 51996 27794 52052 27804
rect 51212 27246 51214 27298
rect 51266 27246 51268 27298
rect 51212 27234 51268 27246
rect 51100 27186 51156 27198
rect 51100 27134 51102 27186
rect 51154 27134 51156 27186
rect 51100 26908 51156 27134
rect 51548 27076 51604 27114
rect 51548 27010 51604 27020
rect 51772 27076 51828 27086
rect 51772 26908 51828 27020
rect 48188 26852 48916 26908
rect 48972 26852 49140 26908
rect 49196 26852 49700 26908
rect 47852 26350 47854 26402
rect 47906 26350 47908 26402
rect 47852 26292 47908 26350
rect 47852 26226 47908 26236
rect 48748 26740 48804 26750
rect 47964 26180 48020 26190
rect 47964 26086 48020 26124
rect 47628 26066 47796 26068
rect 47628 26014 47630 26066
rect 47682 26014 47796 26066
rect 47628 26012 47796 26014
rect 47628 24164 47684 26012
rect 48748 25732 48804 26684
rect 48860 26290 48916 26852
rect 48860 26238 48862 26290
rect 48914 26238 48916 26290
rect 48860 26180 48916 26238
rect 49084 26402 49140 26852
rect 49084 26350 49086 26402
rect 49138 26350 49140 26402
rect 49084 26292 49140 26350
rect 49084 26236 49588 26292
rect 48860 26124 49252 26180
rect 48748 25730 49140 25732
rect 48748 25678 48750 25730
rect 48802 25678 49140 25730
rect 48748 25676 49140 25678
rect 48748 25666 48804 25676
rect 47740 25620 47796 25630
rect 47740 25282 47796 25564
rect 48972 25508 49028 25518
rect 48860 25506 49028 25508
rect 48860 25454 48974 25506
rect 49026 25454 49028 25506
rect 48860 25452 49028 25454
rect 48076 25284 48132 25294
rect 48300 25284 48356 25294
rect 47740 25230 47742 25282
rect 47794 25230 47796 25282
rect 47740 25172 47796 25230
rect 47740 25106 47796 25116
rect 47964 25228 48076 25284
rect 47964 24610 48020 25228
rect 48076 25190 48132 25228
rect 48188 25282 48356 25284
rect 48188 25230 48302 25282
rect 48354 25230 48356 25282
rect 48188 25228 48356 25230
rect 47964 24558 47966 24610
rect 48018 24558 48020 24610
rect 47964 24546 48020 24558
rect 48076 24164 48132 24174
rect 48188 24164 48244 25228
rect 48300 25218 48356 25228
rect 47628 24108 47796 24164
rect 47404 23940 47460 23950
rect 47404 23846 47460 23884
rect 47628 23938 47684 23950
rect 47628 23886 47630 23938
rect 47682 23886 47684 23938
rect 47628 23828 47684 23886
rect 47628 23762 47684 23772
rect 47516 23156 47572 23166
rect 47292 23100 47516 23156
rect 47516 23062 47572 23100
rect 47124 22988 47236 23044
rect 47068 22950 47124 22988
rect 47740 22930 47796 24108
rect 48076 24162 48244 24164
rect 48076 24110 48078 24162
rect 48130 24110 48244 24162
rect 48076 24108 48244 24110
rect 48636 24164 48692 24174
rect 48076 24098 48132 24108
rect 48636 24050 48692 24108
rect 48636 23998 48638 24050
rect 48690 23998 48692 24050
rect 48636 23986 48692 23998
rect 47852 23938 47908 23950
rect 47852 23886 47854 23938
rect 47906 23886 47908 23938
rect 47852 23044 47908 23886
rect 48524 23940 48580 23950
rect 47852 22978 47908 22988
rect 48076 23156 48132 23166
rect 48076 23042 48132 23100
rect 48076 22990 48078 23042
rect 48130 22990 48132 23042
rect 48076 22978 48132 22990
rect 47740 22878 47742 22930
rect 47794 22878 47796 22930
rect 47740 22820 47796 22878
rect 47292 22764 47796 22820
rect 47068 20692 47124 20702
rect 47068 20598 47124 20636
rect 47292 20356 47348 22764
rect 48188 21812 48244 21822
rect 48188 21474 48244 21756
rect 48188 21422 48190 21474
rect 48242 21422 48244 21474
rect 48188 21410 48244 21422
rect 47404 20580 47460 20590
rect 47852 20580 47908 20590
rect 47404 20578 47796 20580
rect 47404 20526 47406 20578
rect 47458 20526 47796 20578
rect 47404 20524 47796 20526
rect 47404 20514 47460 20524
rect 47516 20356 47572 20366
rect 47292 20300 47460 20356
rect 46956 20290 47012 20300
rect 46732 20178 46788 20188
rect 46620 20132 46676 20142
rect 46620 20038 46676 20076
rect 47292 20132 47348 20142
rect 47292 20018 47348 20076
rect 47292 19966 47294 20018
rect 47346 19966 47348 20018
rect 47292 19954 47348 19966
rect 46172 19852 46564 19908
rect 45612 19796 45668 19806
rect 45612 19702 45668 19740
rect 45948 19794 46004 19806
rect 45948 19742 45950 19794
rect 46002 19742 46004 19794
rect 45948 19460 46004 19742
rect 45948 19394 46004 19404
rect 46172 19348 46228 19852
rect 46172 19254 46228 19292
rect 45388 19012 45444 19022
rect 45388 19010 46116 19012
rect 45388 18958 45390 19010
rect 45442 18958 46116 19010
rect 45388 18956 46116 18958
rect 45388 18946 45444 18956
rect 46060 18562 46116 18956
rect 46060 18510 46062 18562
rect 46114 18510 46116 18562
rect 46060 18498 46116 18510
rect 46396 18788 46452 18798
rect 45388 18452 45444 18462
rect 45276 18396 45388 18452
rect 44604 16942 44606 16994
rect 44658 16942 44660 16994
rect 44604 16930 44660 16942
rect 44940 16884 44996 16894
rect 43260 16718 43262 16770
rect 43314 16718 43316 16770
rect 43260 16706 43316 16718
rect 43372 16772 43428 16782
rect 43428 16716 43540 16772
rect 43372 16706 43428 16716
rect 43372 16548 43428 16558
rect 42924 16156 43204 16212
rect 43260 16436 43316 16446
rect 42924 16100 42980 16156
rect 42588 15586 42644 15596
rect 42700 16098 42980 16100
rect 42700 16046 42926 16098
rect 42978 16046 42980 16098
rect 42700 16044 42980 16046
rect 42700 14868 42756 16044
rect 42924 16034 42980 16044
rect 43260 16098 43316 16380
rect 43260 16046 43262 16098
rect 43314 16046 43316 16098
rect 43260 16034 43316 16046
rect 43372 15986 43428 16492
rect 43484 16324 43540 16716
rect 44940 16770 44996 16828
rect 44940 16718 44942 16770
rect 44994 16718 44996 16770
rect 43596 16660 43652 16670
rect 43596 16658 43988 16660
rect 43596 16606 43598 16658
rect 43650 16606 43988 16658
rect 43596 16604 43988 16606
rect 43596 16594 43652 16604
rect 43708 16324 43764 16334
rect 43484 16322 43764 16324
rect 43484 16270 43710 16322
rect 43762 16270 43764 16322
rect 43484 16268 43764 16270
rect 43708 16258 43764 16268
rect 43372 15934 43374 15986
rect 43426 15934 43428 15986
rect 43148 15876 43204 15886
rect 43372 15876 43428 15934
rect 43932 15986 43988 16604
rect 43932 15934 43934 15986
rect 43986 15934 43988 15986
rect 43820 15876 43876 15886
rect 43372 15820 43764 15876
rect 42924 15316 42980 15326
rect 42924 15222 42980 15260
rect 43148 15314 43204 15820
rect 43148 15262 43150 15314
rect 43202 15262 43204 15314
rect 43148 15250 43204 15262
rect 43484 15652 43540 15662
rect 42700 14802 42756 14812
rect 43484 15204 43540 15596
rect 42924 14644 42980 14654
rect 42476 14642 42980 14644
rect 42476 14590 42926 14642
rect 42978 14590 42980 14642
rect 42476 14588 42980 14590
rect 42028 14550 42084 14588
rect 42924 14578 42980 14588
rect 42252 14530 42308 14542
rect 42252 14478 42254 14530
rect 42306 14478 42308 14530
rect 42252 13636 42308 14478
rect 43372 14532 43428 14542
rect 43372 14438 43428 14476
rect 43484 13970 43540 15148
rect 43596 15316 43652 15326
rect 43708 15316 43764 15820
rect 43820 15782 43876 15820
rect 43932 15428 43988 15934
rect 44156 15540 44212 15550
rect 44716 15540 44772 15550
rect 44156 15538 44772 15540
rect 44156 15486 44158 15538
rect 44210 15486 44718 15538
rect 44770 15486 44772 15538
rect 44156 15484 44772 15486
rect 44156 15474 44212 15484
rect 43932 15362 43988 15372
rect 43820 15316 43876 15326
rect 43708 15314 43876 15316
rect 43708 15262 43822 15314
rect 43874 15262 43876 15314
rect 43708 15260 43876 15262
rect 43596 15148 43652 15260
rect 43820 15250 43876 15260
rect 43596 15092 43876 15148
rect 43820 14642 43876 15092
rect 43820 14590 43822 14642
rect 43874 14590 43876 14642
rect 43820 14578 43876 14590
rect 43484 13918 43486 13970
rect 43538 13918 43540 13970
rect 43484 13906 43540 13918
rect 42700 13858 42756 13870
rect 42700 13806 42702 13858
rect 42754 13806 42756 13858
rect 42252 13570 42308 13580
rect 42588 13746 42644 13758
rect 42588 13694 42590 13746
rect 42642 13694 42644 13746
rect 41804 13074 41916 13076
rect 41804 13022 41806 13074
rect 41858 13022 41916 13074
rect 41804 13020 41916 13022
rect 41804 13010 41860 13020
rect 41916 12982 41972 13020
rect 42140 13522 42196 13534
rect 42140 13470 42142 13522
rect 42194 13470 42196 13522
rect 42140 12962 42196 13470
rect 42588 13524 42644 13694
rect 42700 13748 42756 13806
rect 42700 13682 42756 13692
rect 43036 13748 43092 13758
rect 42588 13458 42644 13468
rect 42140 12910 42142 12962
rect 42194 12910 42196 12962
rect 42140 12898 42196 12910
rect 42364 13076 42420 13086
rect 42364 12962 42420 13020
rect 42364 12910 42366 12962
rect 42418 12910 42420 12962
rect 42364 12898 42420 12910
rect 42588 12962 42644 12974
rect 42588 12910 42590 12962
rect 42642 12910 42644 12962
rect 42140 12740 42196 12750
rect 42140 12290 42196 12684
rect 42364 12740 42420 12750
rect 42364 12646 42420 12684
rect 42140 12238 42142 12290
rect 42194 12238 42196 12290
rect 42140 12226 42196 12238
rect 42364 12290 42420 12302
rect 42588 12292 42644 12910
rect 43036 12962 43092 13692
rect 43484 13746 43540 13758
rect 43484 13694 43486 13746
rect 43538 13694 43540 13746
rect 43036 12910 43038 12962
rect 43090 12910 43092 12962
rect 42364 12238 42366 12290
rect 42418 12238 42420 12290
rect 41244 11788 41636 11844
rect 41244 11506 41300 11788
rect 41244 11454 41246 11506
rect 41298 11454 41300 11506
rect 41244 11442 41300 11454
rect 41804 11618 41860 11630
rect 41804 11566 41806 11618
rect 41858 11566 41860 11618
rect 41580 11396 41636 11406
rect 41468 11394 41636 11396
rect 41468 11342 41582 11394
rect 41634 11342 41636 11394
rect 41468 11340 41636 11342
rect 41468 11284 41524 11340
rect 41580 11330 41636 11340
rect 41468 10722 41524 11228
rect 41804 11172 41860 11566
rect 42364 11508 42420 12238
rect 42476 12236 42644 12292
rect 42812 12292 42868 12302
rect 42476 12066 42532 12236
rect 42476 12014 42478 12066
rect 42530 12014 42532 12066
rect 42476 12002 42532 12014
rect 42812 12178 42868 12236
rect 42812 12126 42814 12178
rect 42866 12126 42868 12178
rect 42364 11442 42420 11452
rect 41804 11106 41860 11116
rect 42140 11282 42196 11294
rect 42140 11230 42142 11282
rect 42194 11230 42196 11282
rect 41468 10670 41470 10722
rect 41522 10670 41524 10722
rect 41244 10612 41300 10622
rect 41244 10610 41412 10612
rect 41244 10558 41246 10610
rect 41298 10558 41412 10610
rect 41244 10556 41412 10558
rect 41244 10546 41300 10556
rect 41132 10332 41300 10388
rect 41244 9938 41300 10332
rect 41244 9886 41246 9938
rect 41298 9886 41300 9938
rect 41244 9874 41300 9886
rect 41132 9828 41188 9838
rect 41132 9734 41188 9772
rect 41244 9716 41300 9726
rect 41244 9604 41300 9660
rect 41020 9042 41076 9212
rect 41020 8990 41022 9042
rect 41074 8990 41076 9042
rect 41020 8978 41076 8990
rect 41132 9548 41300 9604
rect 41132 7698 41188 9548
rect 41356 9044 41412 10556
rect 41356 8950 41412 8988
rect 41132 7646 41134 7698
rect 41186 7646 41188 7698
rect 41132 7634 41188 7646
rect 41244 8372 41300 8382
rect 41468 8372 41524 10670
rect 42140 10724 42196 11230
rect 42252 11284 42308 11294
rect 42252 11190 42308 11228
rect 42364 11282 42420 11294
rect 42364 11230 42366 11282
rect 42418 11230 42420 11282
rect 42364 11172 42420 11230
rect 42700 11284 42756 11294
rect 42700 11190 42756 11228
rect 42252 10836 42308 10846
rect 42364 10836 42420 11116
rect 42812 10948 42868 12126
rect 43036 11618 43092 12910
rect 43148 13412 43204 13422
rect 43148 12738 43204 13356
rect 43372 12964 43428 12974
rect 43484 12964 43540 13694
rect 44044 13748 44100 13758
rect 44044 13654 44100 13692
rect 44268 13746 44324 13758
rect 44268 13694 44270 13746
rect 44322 13694 44324 13746
rect 44268 13412 44324 13694
rect 44268 13346 44324 13356
rect 44380 13748 44436 15484
rect 44716 15474 44772 15484
rect 44492 15316 44548 15354
rect 44492 15250 44548 15260
rect 44604 15316 44660 15326
rect 44940 15316 44996 16718
rect 44604 15314 44996 15316
rect 44604 15262 44606 15314
rect 44658 15262 44996 15314
rect 44604 15260 44996 15262
rect 45052 16212 45108 18396
rect 45388 18358 45444 18396
rect 45612 17668 45668 17678
rect 45612 17666 45892 17668
rect 45612 17614 45614 17666
rect 45666 17614 45892 17666
rect 45612 17612 45892 17614
rect 45612 17602 45668 17612
rect 45276 17554 45332 17566
rect 45276 17502 45278 17554
rect 45330 17502 45332 17554
rect 45164 17442 45220 17454
rect 45164 17390 45166 17442
rect 45218 17390 45220 17442
rect 45164 17108 45220 17390
rect 45164 16882 45220 17052
rect 45164 16830 45166 16882
rect 45218 16830 45220 16882
rect 45164 16818 45220 16830
rect 45276 16324 45332 17502
rect 45724 17444 45780 17454
rect 45724 17350 45780 17388
rect 45836 16996 45892 17612
rect 45948 17556 46004 17566
rect 45948 17462 46004 17500
rect 46172 17556 46228 17566
rect 46172 17462 46228 17500
rect 46396 17220 46452 18732
rect 46508 17666 46564 19852
rect 47068 19234 47124 19246
rect 47068 19182 47070 19234
rect 47122 19182 47124 19234
rect 47068 18452 47124 19182
rect 47068 18386 47124 18396
rect 46508 17614 46510 17666
rect 46562 17614 46564 17666
rect 46508 17602 46564 17614
rect 47180 17668 47236 17678
rect 46732 17556 46788 17566
rect 46788 17500 46900 17556
rect 46732 17490 46788 17500
rect 46172 17164 46452 17220
rect 46060 17108 46116 17118
rect 46060 17014 46116 17052
rect 45836 16660 45892 16940
rect 45948 16884 46004 16894
rect 46172 16884 46228 17164
rect 46620 16996 46676 17006
rect 46676 16940 46788 16996
rect 46620 16930 46676 16940
rect 46172 16828 46340 16884
rect 45948 16790 46004 16828
rect 46060 16660 46116 16670
rect 45836 16658 46116 16660
rect 45836 16606 46062 16658
rect 46114 16606 46116 16658
rect 45836 16604 46116 16606
rect 46060 16594 46116 16604
rect 45276 16258 45332 16268
rect 46060 16212 46116 16222
rect 45052 16210 45220 16212
rect 45052 16158 45054 16210
rect 45106 16158 45220 16210
rect 45052 16156 45220 16158
rect 44604 15250 44660 15260
rect 44828 15092 44884 15102
rect 44716 15036 44828 15092
rect 44604 13748 44660 13758
rect 44380 13746 44660 13748
rect 44380 13694 44606 13746
rect 44658 13694 44660 13746
rect 44380 13692 44660 13694
rect 44268 13188 44324 13198
rect 44380 13188 44436 13692
rect 44604 13682 44660 13692
rect 44604 13524 44660 13534
rect 44716 13524 44772 15036
rect 44828 15026 44884 15036
rect 45052 14644 45108 16156
rect 45164 16100 45220 16156
rect 45388 16100 45444 16110
rect 45164 16098 45444 16100
rect 45164 16046 45390 16098
rect 45442 16046 45444 16098
rect 45164 16044 45444 16046
rect 45388 16034 45444 16044
rect 45612 16044 46004 16100
rect 45500 15876 45556 15886
rect 45612 15876 45668 16044
rect 45500 15874 45668 15876
rect 45500 15822 45502 15874
rect 45554 15822 45668 15874
rect 45500 15820 45668 15822
rect 45724 15874 45780 15886
rect 45724 15822 45726 15874
rect 45778 15822 45780 15874
rect 45500 15810 45556 15820
rect 45612 15538 45668 15550
rect 45612 15486 45614 15538
rect 45666 15486 45668 15538
rect 45276 15428 45332 15438
rect 45164 15314 45220 15326
rect 45164 15262 45166 15314
rect 45218 15262 45220 15314
rect 45164 15204 45220 15262
rect 45276 15316 45332 15372
rect 45388 15316 45444 15326
rect 45276 15314 45444 15316
rect 45276 15262 45390 15314
rect 45442 15262 45444 15314
rect 45276 15260 45444 15262
rect 45388 15250 45444 15260
rect 45500 15202 45556 15214
rect 45500 15150 45502 15202
rect 45554 15150 45556 15202
rect 45500 15148 45556 15150
rect 45164 15092 45556 15148
rect 45612 14754 45668 15486
rect 45724 15540 45780 15822
rect 45836 15540 45892 15550
rect 45724 15538 45892 15540
rect 45724 15486 45838 15538
rect 45890 15486 45892 15538
rect 45724 15484 45892 15486
rect 45836 15474 45892 15484
rect 45612 14702 45614 14754
rect 45666 14702 45668 14754
rect 45612 14690 45668 14702
rect 45276 14644 45332 14654
rect 45052 14642 45332 14644
rect 45052 14590 45054 14642
rect 45106 14590 45278 14642
rect 45330 14590 45332 14642
rect 45052 14588 45332 14590
rect 45052 14578 45108 14588
rect 45276 14578 45332 14588
rect 45612 14532 45668 14542
rect 45948 14532 46004 16044
rect 45612 14530 46004 14532
rect 45612 14478 45614 14530
rect 45666 14478 46004 14530
rect 45612 14476 46004 14478
rect 45612 14466 45668 14476
rect 45948 14196 46004 14476
rect 45948 14130 46004 14140
rect 46060 15428 46116 16156
rect 44828 13972 44884 13982
rect 44828 13878 44884 13916
rect 45948 13972 46004 13982
rect 46060 13972 46116 15372
rect 46172 15874 46228 15886
rect 46172 15822 46174 15874
rect 46226 15822 46228 15874
rect 46172 15316 46228 15822
rect 46172 15250 46228 15260
rect 46172 13972 46228 13982
rect 45948 13970 46228 13972
rect 45948 13918 45950 13970
rect 46002 13918 46174 13970
rect 46226 13918 46228 13970
rect 45948 13916 46228 13918
rect 45948 13906 46004 13916
rect 46172 13906 46228 13916
rect 44268 13186 44436 13188
rect 44268 13134 44270 13186
rect 44322 13134 44436 13186
rect 44268 13132 44436 13134
rect 44492 13522 44772 13524
rect 44492 13470 44606 13522
rect 44658 13470 44772 13522
rect 44492 13468 44772 13470
rect 44268 13122 44324 13132
rect 43372 12962 43540 12964
rect 43372 12910 43374 12962
rect 43426 12910 43540 12962
rect 43372 12908 43540 12910
rect 43372 12898 43428 12908
rect 44156 12852 44212 12862
rect 44156 12758 44212 12796
rect 43148 12686 43150 12738
rect 43202 12686 43204 12738
rect 43148 12404 43204 12686
rect 43260 12740 43316 12750
rect 43316 12684 43652 12740
rect 43260 12674 43316 12684
rect 43148 12338 43204 12348
rect 43596 12290 43652 12684
rect 44044 12738 44100 12750
rect 44492 12740 44548 13468
rect 44604 13458 44660 13468
rect 44044 12686 44046 12738
rect 44098 12686 44100 12738
rect 44044 12628 44100 12686
rect 44268 12684 44548 12740
rect 44268 12628 44324 12684
rect 44044 12572 44324 12628
rect 43596 12238 43598 12290
rect 43650 12238 43652 12290
rect 43596 12226 43652 12238
rect 46172 12292 46228 12302
rect 46172 12198 46228 12236
rect 45724 12066 45780 12078
rect 45724 12014 45726 12066
rect 45778 12014 45780 12066
rect 43036 11566 43038 11618
rect 43090 11566 43092 11618
rect 43036 11554 43092 11566
rect 44716 11844 44772 11854
rect 43372 11508 43428 11518
rect 43372 11394 43428 11452
rect 43372 11342 43374 11394
rect 43426 11342 43428 11394
rect 43372 11330 43428 11342
rect 44716 11508 44772 11788
rect 45724 11844 45780 12014
rect 45724 11778 45780 11788
rect 42700 10892 42868 10948
rect 42924 11170 42980 11182
rect 42924 11118 42926 11170
rect 42978 11118 42980 11170
rect 42308 10780 42644 10836
rect 42252 10742 42308 10780
rect 41300 8316 41524 8372
rect 41580 9828 41636 9838
rect 41580 9156 41636 9772
rect 41244 7698 41300 8316
rect 41244 7646 41246 7698
rect 41298 7646 41300 7698
rect 41244 7634 41300 7646
rect 41356 7812 41412 7822
rect 41356 7698 41412 7756
rect 41356 7646 41358 7698
rect 41410 7646 41412 7698
rect 41356 7634 41412 7646
rect 41468 7700 41524 7710
rect 41580 7700 41636 9100
rect 41468 7698 41636 7700
rect 41468 7646 41470 7698
rect 41522 7646 41636 7698
rect 41468 7644 41636 7646
rect 41692 9604 41748 9614
rect 41468 7634 41524 7644
rect 41692 7586 41748 9548
rect 42140 9604 42196 10668
rect 42588 10722 42644 10780
rect 42588 10670 42590 10722
rect 42642 10670 42644 10722
rect 42588 10658 42644 10670
rect 42140 9538 42196 9548
rect 42364 9268 42420 9278
rect 42364 9174 42420 9212
rect 42700 9268 42756 10892
rect 42812 10724 42868 10762
rect 42812 10658 42868 10668
rect 42812 10500 42868 10510
rect 42812 9714 42868 10444
rect 42924 10498 42980 11118
rect 43484 11172 43540 11182
rect 43484 11078 43540 11116
rect 44156 11172 44212 11182
rect 44156 11078 44212 11116
rect 43596 10836 43652 10846
rect 43596 10742 43652 10780
rect 43260 10724 43316 10734
rect 43260 10722 43540 10724
rect 43260 10670 43262 10722
rect 43314 10670 43540 10722
rect 43260 10668 43540 10670
rect 43260 10658 43316 10668
rect 42924 10446 42926 10498
rect 42978 10446 42980 10498
rect 42924 10434 42980 10446
rect 43372 10388 43428 10398
rect 43372 9826 43428 10332
rect 43372 9774 43374 9826
rect 43426 9774 43428 9826
rect 43372 9762 43428 9774
rect 43484 9828 43540 10668
rect 44716 10610 44772 11452
rect 44940 11732 44996 11742
rect 44940 11170 44996 11676
rect 44940 11118 44942 11170
rect 44994 11118 44996 11170
rect 44940 10836 44996 11118
rect 44940 10770 44996 10780
rect 45836 11620 45892 11630
rect 45836 11506 45892 11564
rect 45836 11454 45838 11506
rect 45890 11454 45892 11506
rect 44716 10558 44718 10610
rect 44770 10558 44772 10610
rect 44716 10546 44772 10558
rect 45164 10610 45220 10622
rect 45164 10558 45166 10610
rect 45218 10558 45220 10610
rect 44044 10500 44100 10510
rect 44044 10406 44100 10444
rect 43484 9734 43540 9772
rect 43932 9828 43988 9838
rect 43932 9734 43988 9772
rect 42812 9662 42814 9714
rect 42866 9662 42868 9714
rect 42812 9650 42868 9662
rect 42700 9042 42756 9212
rect 42700 8990 42702 9042
rect 42754 8990 42756 9042
rect 42588 8260 42644 8270
rect 42700 8260 42756 8990
rect 43596 9602 43652 9614
rect 43596 9550 43598 9602
rect 43650 9550 43652 9602
rect 43484 8930 43540 8942
rect 43484 8878 43486 8930
rect 43538 8878 43540 8930
rect 43484 8482 43540 8878
rect 43484 8430 43486 8482
rect 43538 8430 43540 8482
rect 43484 8418 43540 8430
rect 43596 8370 43652 9550
rect 43708 9604 43764 9614
rect 43708 9510 43764 9548
rect 44828 9604 44884 9614
rect 44828 9510 44884 9548
rect 45164 9602 45220 10558
rect 45836 10388 45892 11454
rect 45836 10322 45892 10332
rect 45164 9550 45166 9602
rect 45218 9550 45220 9602
rect 45164 8932 45220 9550
rect 46060 9268 46116 9278
rect 46060 9174 46116 9212
rect 45612 8932 45668 8942
rect 45164 8930 45668 8932
rect 45164 8878 45614 8930
rect 45666 8878 45668 8930
rect 45164 8876 45668 8878
rect 45612 8866 45668 8876
rect 43596 8318 43598 8370
rect 43650 8318 43652 8370
rect 43596 8306 43652 8318
rect 42588 8258 42756 8260
rect 42588 8206 42590 8258
rect 42642 8206 42756 8258
rect 42588 8204 42756 8206
rect 42588 8194 42644 8204
rect 41804 8148 41860 8158
rect 41804 8054 41860 8092
rect 42700 7700 42756 8204
rect 42924 8148 42980 8158
rect 42924 8054 42980 8092
rect 43036 8146 43092 8158
rect 43036 8094 43038 8146
rect 43090 8094 43092 8146
rect 43036 7812 43092 8094
rect 43036 7746 43092 7756
rect 42812 7700 42868 7710
rect 42756 7698 42868 7700
rect 42756 7646 42814 7698
rect 42866 7646 42868 7698
rect 42756 7644 42868 7646
rect 42700 7606 42756 7644
rect 42812 7634 42868 7644
rect 41692 7534 41694 7586
rect 41746 7534 41748 7586
rect 41692 7522 41748 7534
rect 46284 4004 46340 16828
rect 46732 16882 46788 16940
rect 46732 16830 46734 16882
rect 46786 16830 46788 16882
rect 46732 16818 46788 16830
rect 46508 16324 46564 16334
rect 46508 16230 46564 16268
rect 46732 16212 46788 16222
rect 46844 16212 46900 17500
rect 47068 17444 47124 17454
rect 47068 17106 47124 17388
rect 47068 17054 47070 17106
rect 47122 17054 47124 17106
rect 47068 16548 47124 17054
rect 47180 16770 47236 17612
rect 47292 17556 47348 17566
rect 47292 17106 47348 17500
rect 47292 17054 47294 17106
rect 47346 17054 47348 17106
rect 47292 17042 47348 17054
rect 47180 16718 47182 16770
rect 47234 16718 47236 16770
rect 47180 16706 47236 16718
rect 47068 16492 47348 16548
rect 46732 16210 46900 16212
rect 46732 16158 46734 16210
rect 46786 16158 46900 16210
rect 46732 16156 46900 16158
rect 47068 16324 47124 16334
rect 47068 16210 47124 16268
rect 47068 16158 47070 16210
rect 47122 16158 47124 16210
rect 46732 16146 46788 16156
rect 47068 16146 47124 16158
rect 47180 16212 47236 16222
rect 47180 16098 47236 16156
rect 47180 16046 47182 16098
rect 47234 16046 47236 16098
rect 47180 16034 47236 16046
rect 47292 15876 47348 16492
rect 47180 15820 47348 15876
rect 46956 15428 47012 15438
rect 46956 15334 47012 15372
rect 47180 15426 47236 15820
rect 47180 15374 47182 15426
rect 47234 15374 47236 15426
rect 47180 15362 47236 15374
rect 46508 15314 46564 15326
rect 46508 15262 46510 15314
rect 46562 15262 46564 15314
rect 46396 15204 46452 15214
rect 46508 15204 46564 15262
rect 46620 15316 46676 15326
rect 46620 15222 46676 15260
rect 46844 15316 46900 15326
rect 46452 15148 46564 15204
rect 46396 15138 46452 15148
rect 46844 14754 46900 15260
rect 47292 15316 47348 15326
rect 47292 15222 47348 15260
rect 47404 15148 47460 20300
rect 47516 16884 47572 20300
rect 47740 19348 47796 20524
rect 47852 20486 47908 20524
rect 48524 20132 48580 23884
rect 48748 23268 48804 23278
rect 48748 23174 48804 23212
rect 48860 21700 48916 25452
rect 48972 25442 49028 25452
rect 48860 21634 48916 21644
rect 48972 24610 49028 24622
rect 48972 24558 48974 24610
rect 49026 24558 49028 24610
rect 48860 21476 48916 21486
rect 48972 21476 49028 24558
rect 49084 23940 49140 25676
rect 49196 25508 49252 26124
rect 49532 25508 49588 26236
rect 49644 25732 49700 26852
rect 49644 25666 49700 25676
rect 50092 26852 50260 26908
rect 50876 26852 51156 26908
rect 51548 26852 51828 26908
rect 49868 25508 49924 25518
rect 49532 25506 49924 25508
rect 49532 25454 49870 25506
rect 49922 25454 49924 25506
rect 49532 25452 49924 25454
rect 49196 25414 49252 25452
rect 49868 25442 49924 25452
rect 49420 25394 49476 25406
rect 49420 25342 49422 25394
rect 49474 25342 49476 25394
rect 49420 25284 49476 25342
rect 49420 24612 49476 25228
rect 49756 24612 49812 24622
rect 49420 24610 49812 24612
rect 49420 24558 49758 24610
rect 49810 24558 49812 24610
rect 49420 24556 49812 24558
rect 49756 24546 49812 24556
rect 50092 24164 50148 26852
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50540 26516 50596 26526
rect 50876 26516 50932 26852
rect 50540 26514 50932 26516
rect 50540 26462 50542 26514
rect 50594 26462 50932 26514
rect 50540 26460 50932 26462
rect 51436 26516 51492 26526
rect 51548 26516 51604 26852
rect 51436 26514 51604 26516
rect 51436 26462 51438 26514
rect 51490 26462 51604 26514
rect 51436 26460 51604 26462
rect 50540 26450 50596 26460
rect 51436 26450 51492 26460
rect 50988 26404 51044 26414
rect 50876 26348 50988 26404
rect 50316 26292 50372 26302
rect 50652 26292 50708 26302
rect 50316 26290 50484 26292
rect 50316 26238 50318 26290
rect 50370 26238 50484 26290
rect 50316 26236 50484 26238
rect 50316 26180 50372 26236
rect 50316 26114 50372 26124
rect 50316 25396 50372 25406
rect 50316 25302 50372 25340
rect 50204 25282 50260 25294
rect 50204 25230 50206 25282
rect 50258 25230 50260 25282
rect 50204 25060 50260 25230
rect 50204 24994 50260 25004
rect 50204 24836 50260 24846
rect 50204 24722 50260 24780
rect 50204 24670 50206 24722
rect 50258 24670 50260 24722
rect 50204 24658 50260 24670
rect 50092 24098 50148 24108
rect 50428 23940 50484 26236
rect 50652 26198 50708 26236
rect 50876 25620 50932 26348
rect 50988 26338 51044 26348
rect 51212 26402 51268 26414
rect 51212 26350 51214 26402
rect 51266 26350 51268 26402
rect 51100 26290 51156 26302
rect 51100 26238 51102 26290
rect 51154 26238 51156 26290
rect 51100 25620 51156 26238
rect 51212 26180 51268 26350
rect 51660 26404 51716 26414
rect 51660 26310 51716 26348
rect 51772 26404 51828 26414
rect 51772 26402 51940 26404
rect 51772 26350 51774 26402
rect 51826 26350 51940 26402
rect 51772 26348 51940 26350
rect 51772 26338 51828 26348
rect 51212 26124 51828 26180
rect 51772 26066 51828 26124
rect 51772 26014 51774 26066
rect 51826 26014 51828 26066
rect 51772 26002 51828 26014
rect 51884 25844 51940 26348
rect 52108 26292 52164 27804
rect 52220 27524 52276 27534
rect 52220 27188 52276 27468
rect 52220 27122 52276 27132
rect 52108 26226 52164 26236
rect 52220 26964 52276 26974
rect 51772 25788 51940 25844
rect 51772 25732 51828 25788
rect 51436 25676 51828 25732
rect 51324 25620 51380 25630
rect 51100 25618 51380 25620
rect 51100 25566 51326 25618
rect 51378 25566 51380 25618
rect 51100 25564 51380 25566
rect 50876 25554 50932 25564
rect 51324 25554 51380 25564
rect 50988 25508 51044 25518
rect 51044 25452 51156 25508
rect 50988 25442 51044 25452
rect 50540 25396 50596 25406
rect 50540 25302 50596 25340
rect 50988 25172 51044 25182
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50876 25116 50988 25172
rect 50876 24836 50932 25116
rect 50988 25106 51044 25116
rect 51100 25060 51156 25452
rect 51212 25394 51268 25406
rect 51212 25342 51214 25394
rect 51266 25342 51268 25394
rect 51212 25284 51268 25342
rect 51212 25218 51268 25228
rect 51324 25394 51380 25406
rect 51324 25342 51326 25394
rect 51378 25342 51380 25394
rect 51324 25060 51380 25342
rect 51436 25394 51492 25676
rect 51772 25620 51828 25676
rect 51996 25620 52052 25630
rect 51772 25618 52052 25620
rect 51772 25566 51998 25618
rect 52050 25566 52052 25618
rect 51772 25564 52052 25566
rect 51996 25554 52052 25564
rect 51660 25508 51716 25518
rect 51660 25414 51716 25452
rect 51436 25342 51438 25394
rect 51490 25342 51492 25394
rect 51436 25330 51492 25342
rect 52108 25394 52164 25406
rect 52108 25342 52110 25394
rect 52162 25342 52164 25394
rect 52108 25284 52164 25342
rect 51884 25228 52164 25284
rect 51884 25172 51940 25228
rect 52220 25172 52276 26908
rect 52332 26180 52388 27916
rect 52556 27860 52612 27870
rect 52556 27188 52612 27804
rect 52556 26908 52612 27132
rect 52780 27186 52836 28028
rect 53004 27970 53060 28476
rect 53228 28420 53284 29374
rect 53340 28644 53396 28654
rect 53340 28550 53396 28588
rect 53564 28420 53620 28430
rect 53228 28418 53620 28420
rect 53228 28366 53566 28418
rect 53618 28366 53620 28418
rect 53228 28364 53620 28366
rect 53004 27918 53006 27970
rect 53058 27918 53060 27970
rect 53004 27906 53060 27918
rect 53116 28308 53172 28318
rect 52780 27134 52782 27186
rect 52834 27134 52836 27186
rect 52780 27122 52836 27134
rect 53004 27524 53060 27534
rect 52668 27076 52724 27086
rect 52668 26982 52724 27020
rect 52892 26964 52948 27002
rect 52556 26852 52836 26908
rect 52892 26898 52948 26908
rect 53004 26962 53060 27468
rect 53004 26910 53006 26962
rect 53058 26910 53060 26962
rect 53004 26898 53060 26910
rect 52780 26402 52836 26852
rect 53116 26514 53172 28252
rect 53452 27076 53508 27086
rect 53564 27076 53620 28364
rect 53676 27748 53732 29596
rect 54012 29650 54068 29708
rect 54012 29598 54014 29650
rect 54066 29598 54068 29650
rect 54012 29586 54068 29598
rect 54236 29650 54292 30156
rect 54236 29598 54238 29650
rect 54290 29598 54292 29650
rect 53788 29540 53844 29550
rect 53788 28644 53844 29484
rect 54124 29428 54180 29438
rect 54124 29334 54180 29372
rect 53788 28578 53844 28588
rect 53900 28980 53956 28990
rect 53900 28642 53956 28924
rect 53900 28590 53902 28642
rect 53954 28590 53956 28642
rect 53900 28308 53956 28590
rect 53900 28242 53956 28252
rect 54124 28644 54180 28654
rect 54012 27748 54068 27758
rect 53676 27746 54068 27748
rect 53676 27694 54014 27746
rect 54066 27694 54068 27746
rect 53676 27692 54068 27694
rect 54012 27524 54068 27692
rect 54012 27458 54068 27468
rect 54124 27300 54180 28588
rect 54236 27858 54292 29598
rect 54348 28084 54404 30492
rect 54460 30324 54516 30334
rect 54460 30210 54516 30268
rect 54460 30158 54462 30210
rect 54514 30158 54516 30210
rect 54460 30146 54516 30158
rect 54796 30100 54852 30942
rect 55580 30996 55636 31006
rect 55580 30902 55636 30940
rect 54572 30044 54796 30100
rect 54572 28756 54628 30044
rect 54796 30034 54852 30044
rect 54908 30772 54964 30782
rect 54908 30212 54964 30716
rect 55692 30772 55748 30782
rect 55692 30770 56084 30772
rect 55692 30718 55694 30770
rect 55746 30718 56084 30770
rect 55692 30716 56084 30718
rect 55692 30706 55748 30716
rect 56028 30322 56084 30716
rect 56028 30270 56030 30322
rect 56082 30270 56084 30322
rect 56028 30258 56084 30270
rect 55244 30212 55300 30222
rect 54908 30210 55300 30212
rect 54908 30158 54910 30210
rect 54962 30158 55246 30210
rect 55298 30158 55300 30210
rect 54908 30156 55300 30158
rect 54684 29540 54740 29550
rect 54684 29446 54740 29484
rect 54796 29426 54852 29438
rect 54796 29374 54798 29426
rect 54850 29374 54852 29426
rect 54684 29204 54740 29214
rect 54684 29110 54740 29148
rect 54684 28980 54740 28990
rect 54796 28980 54852 29374
rect 54740 28924 54852 28980
rect 54684 28914 54740 28924
rect 54572 28700 54740 28756
rect 54684 28642 54740 28700
rect 54908 28644 54964 30156
rect 55244 30146 55300 30156
rect 55916 30212 55972 30222
rect 55804 29764 55860 29774
rect 55804 29652 55860 29708
rect 55692 29650 55860 29652
rect 55692 29598 55806 29650
rect 55858 29598 55860 29650
rect 55692 29596 55860 29598
rect 55132 29538 55188 29550
rect 55132 29486 55134 29538
rect 55186 29486 55188 29538
rect 55020 29428 55076 29438
rect 55132 29428 55188 29486
rect 55244 29540 55300 29550
rect 55580 29540 55636 29550
rect 55244 29538 55636 29540
rect 55244 29486 55246 29538
rect 55298 29486 55582 29538
rect 55634 29486 55636 29538
rect 55244 29484 55636 29486
rect 55244 29474 55300 29484
rect 55580 29474 55636 29484
rect 55076 29372 55188 29428
rect 55020 29362 55076 29372
rect 55244 29316 55300 29326
rect 55244 29202 55300 29260
rect 55244 29150 55246 29202
rect 55298 29150 55300 29202
rect 55244 29138 55300 29150
rect 55692 28980 55748 29596
rect 55804 29586 55860 29596
rect 55916 29538 55972 30156
rect 55916 29486 55918 29538
rect 55970 29486 55972 29538
rect 55916 29474 55972 29486
rect 54684 28590 54686 28642
rect 54738 28590 54740 28642
rect 54684 28578 54740 28590
rect 54796 28588 54964 28644
rect 55132 28924 55748 28980
rect 55132 28642 55188 28924
rect 55244 28756 55300 28766
rect 55804 28756 55860 28766
rect 55244 28754 55860 28756
rect 55244 28702 55246 28754
rect 55298 28702 55806 28754
rect 55858 28702 55860 28754
rect 55244 28700 55860 28702
rect 55244 28690 55300 28700
rect 55804 28690 55860 28700
rect 56140 28756 56196 28766
rect 55132 28590 55134 28642
rect 55186 28590 55188 28642
rect 54684 28308 54740 28318
rect 54684 28084 54740 28252
rect 54796 28196 54852 28588
rect 54908 28420 54964 28430
rect 54908 28418 55076 28420
rect 54908 28366 54910 28418
rect 54962 28366 55076 28418
rect 54908 28364 55076 28366
rect 54908 28354 54964 28364
rect 54796 28140 54964 28196
rect 54348 28028 54516 28084
rect 54684 28028 54852 28084
rect 54236 27806 54238 27858
rect 54290 27806 54292 27858
rect 54236 27794 54292 27806
rect 54348 27300 54404 27310
rect 54124 27298 54404 27300
rect 54124 27246 54350 27298
rect 54402 27246 54404 27298
rect 54124 27244 54404 27246
rect 54348 27234 54404 27244
rect 54460 27300 54516 28028
rect 54684 27860 54740 27870
rect 54684 27766 54740 27804
rect 54572 27300 54628 27310
rect 54460 27298 54628 27300
rect 54460 27246 54574 27298
rect 54626 27246 54628 27298
rect 54460 27244 54628 27246
rect 53452 27074 53620 27076
rect 53452 27022 53454 27074
rect 53506 27022 53620 27074
rect 53452 27020 53620 27022
rect 54012 27188 54068 27198
rect 54012 27074 54068 27132
rect 54012 27022 54014 27074
rect 54066 27022 54068 27074
rect 53452 27010 53508 27020
rect 54012 27010 54068 27022
rect 53116 26462 53118 26514
rect 53170 26462 53172 26514
rect 53116 26450 53172 26462
rect 53788 26962 53844 26974
rect 53788 26910 53790 26962
rect 53842 26910 53844 26962
rect 52780 26350 52782 26402
rect 52834 26350 52836 26402
rect 52780 26338 52836 26350
rect 52892 26404 52948 26414
rect 52892 26310 52948 26348
rect 53788 26404 53844 26910
rect 54460 26516 54516 27244
rect 54572 27234 54628 27244
rect 54796 26908 54852 28028
rect 52332 26114 52388 26124
rect 53676 26180 53732 26190
rect 53004 25506 53060 25518
rect 53004 25454 53006 25506
rect 53058 25454 53060 25506
rect 51884 25106 51940 25116
rect 51996 25116 52276 25172
rect 52668 25394 52724 25406
rect 52668 25342 52670 25394
rect 52722 25342 52724 25394
rect 51436 25060 51492 25070
rect 51100 25004 51436 25060
rect 51436 24994 51492 25004
rect 50876 24770 50932 24780
rect 51100 24836 51156 24846
rect 50652 24722 50708 24734
rect 50652 24670 50654 24722
rect 50706 24670 50708 24722
rect 50652 24500 50708 24670
rect 50988 24724 51044 24734
rect 50988 24630 51044 24668
rect 51100 24722 51156 24780
rect 51100 24670 51102 24722
rect 51154 24670 51156 24722
rect 51100 24658 51156 24670
rect 51436 24722 51492 24734
rect 51436 24670 51438 24722
rect 51490 24670 51492 24722
rect 51436 24500 51492 24670
rect 49084 23884 49252 23940
rect 49084 23716 49140 23726
rect 49084 23622 49140 23660
rect 49196 21924 49252 23884
rect 50204 23884 50484 23940
rect 50540 24444 51492 24500
rect 49420 23156 49476 23166
rect 49420 23062 49476 23100
rect 49644 23044 49700 23054
rect 50204 23044 50260 23884
rect 50540 23826 50596 24444
rect 50652 24164 50708 24174
rect 50652 23938 50708 24108
rect 51100 23996 51380 24052
rect 50652 23886 50654 23938
rect 50706 23886 50708 23938
rect 50652 23874 50708 23886
rect 50876 23940 50932 23950
rect 50876 23846 50932 23884
rect 51100 23938 51156 23996
rect 51100 23886 51102 23938
rect 51154 23886 51156 23938
rect 51100 23874 51156 23886
rect 50540 23774 50542 23826
rect 50594 23774 50596 23826
rect 50540 23762 50596 23774
rect 51212 23828 51268 23838
rect 50316 23716 50372 23726
rect 50316 23714 50484 23716
rect 50316 23662 50318 23714
rect 50370 23662 50484 23714
rect 50316 23660 50484 23662
rect 50316 23650 50372 23660
rect 50428 23268 50484 23660
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 51212 23378 51268 23772
rect 51212 23326 51214 23378
rect 51266 23326 51268 23378
rect 51212 23314 51268 23326
rect 50428 23202 50484 23212
rect 51324 23266 51380 23996
rect 51436 23826 51492 24444
rect 51436 23774 51438 23826
rect 51490 23774 51492 23826
rect 51436 23762 51492 23774
rect 51884 24164 51940 24174
rect 51884 23826 51940 24108
rect 51884 23774 51886 23826
rect 51938 23774 51940 23826
rect 51884 23762 51940 23774
rect 51996 23378 52052 25116
rect 52444 24724 52500 24734
rect 52668 24724 52724 25342
rect 52780 25396 52836 25406
rect 52780 25302 52836 25340
rect 52892 25060 52948 25070
rect 52444 24722 52724 24724
rect 52444 24670 52446 24722
rect 52498 24670 52724 24722
rect 52444 24668 52724 24670
rect 52780 24724 52836 24734
rect 52332 24612 52388 24622
rect 52332 24518 52388 24556
rect 52444 23828 52500 24668
rect 52780 24630 52836 24668
rect 52892 24050 52948 25004
rect 53004 24724 53060 25454
rect 53452 25396 53508 25406
rect 53452 25394 53620 25396
rect 53452 25342 53454 25394
rect 53506 25342 53620 25394
rect 53452 25340 53620 25342
rect 53452 25330 53508 25340
rect 53340 25284 53396 25294
rect 53340 25190 53396 25228
rect 53004 24658 53060 24668
rect 53116 24164 53172 24174
rect 53116 24070 53172 24108
rect 52892 23998 52894 24050
rect 52946 23998 52948 24050
rect 52892 23986 52948 23998
rect 52444 23762 52500 23772
rect 53564 23938 53620 25340
rect 53676 25284 53732 26124
rect 53788 25620 53844 26348
rect 54348 26460 54460 26516
rect 54348 26402 54404 26460
rect 54460 26450 54516 26460
rect 54572 26852 54852 26908
rect 54908 27186 54964 28140
rect 55020 27298 55076 28364
rect 55132 28084 55188 28590
rect 55356 28532 55412 28542
rect 55244 28476 55356 28532
rect 55244 28418 55300 28476
rect 55356 28466 55412 28476
rect 55244 28366 55246 28418
rect 55298 28366 55300 28418
rect 55244 28354 55300 28366
rect 55916 28420 55972 28430
rect 55916 28418 56084 28420
rect 55916 28366 55918 28418
rect 55970 28366 56084 28418
rect 55916 28364 56084 28366
rect 55916 28354 55972 28364
rect 55356 28084 55412 28094
rect 55132 28082 55412 28084
rect 55132 28030 55358 28082
rect 55410 28030 55412 28082
rect 55132 28028 55412 28030
rect 55020 27246 55022 27298
rect 55074 27246 55076 27298
rect 55020 27234 55076 27246
rect 54908 27134 54910 27186
rect 54962 27134 54964 27186
rect 54908 27076 54964 27134
rect 55244 27076 55300 27086
rect 54908 27074 55300 27076
rect 54908 27022 55246 27074
rect 55298 27022 55300 27074
rect 54908 27020 55300 27022
rect 54348 26350 54350 26402
rect 54402 26350 54404 26402
rect 54348 26338 54404 26350
rect 54012 26292 54068 26302
rect 53788 25554 53844 25564
rect 53900 26290 54068 26292
rect 53900 26238 54014 26290
rect 54066 26238 54068 26290
rect 53900 26236 54068 26238
rect 53900 25284 53956 26236
rect 54012 26226 54068 26236
rect 53676 25228 53956 25284
rect 53676 24724 53732 24734
rect 53676 24630 53732 24668
rect 53788 24610 53844 24622
rect 53788 24558 53790 24610
rect 53842 24558 53844 24610
rect 53788 24164 53844 24558
rect 53788 24098 53844 24108
rect 53564 23886 53566 23938
rect 53618 23886 53620 23938
rect 51996 23326 51998 23378
rect 52050 23326 52052 23378
rect 51996 23314 52052 23326
rect 51324 23214 51326 23266
rect 51378 23214 51380 23266
rect 50876 23154 50932 23166
rect 50876 23102 50878 23154
rect 50930 23102 50932 23154
rect 49644 23042 50148 23044
rect 49644 22990 49646 23042
rect 49698 22990 50148 23042
rect 49644 22988 50148 22990
rect 50204 22988 50484 23044
rect 49644 22978 49700 22988
rect 50092 22596 50148 22988
rect 49196 21810 49252 21868
rect 49980 22540 50092 22596
rect 49196 21758 49198 21810
rect 49250 21758 49252 21810
rect 49196 21746 49252 21758
rect 49532 21812 49588 21822
rect 49532 21718 49588 21756
rect 48524 20066 48580 20076
rect 48636 21474 49028 21476
rect 48636 21422 48862 21474
rect 48914 21422 49028 21474
rect 48636 21420 49028 21422
rect 47852 20020 47908 20030
rect 47852 20018 48244 20020
rect 47852 19966 47854 20018
rect 47906 19966 48244 20018
rect 47852 19964 48244 19966
rect 47852 19954 47908 19964
rect 47852 19348 47908 19358
rect 47740 19346 47908 19348
rect 47740 19294 47854 19346
rect 47906 19294 47908 19346
rect 47740 19292 47908 19294
rect 47852 19282 47908 19292
rect 47628 18452 47684 18462
rect 47628 17778 47684 18396
rect 47628 17726 47630 17778
rect 47682 17726 47684 17778
rect 47628 17714 47684 17726
rect 48188 18338 48244 19964
rect 48636 18452 48692 21420
rect 48860 21410 48916 21420
rect 48972 21252 49028 21262
rect 48860 20132 48916 20142
rect 48860 20038 48916 20076
rect 48860 18452 48916 18462
rect 48636 18396 48860 18452
rect 48188 18286 48190 18338
rect 48242 18286 48244 18338
rect 47964 17444 48020 17454
rect 47964 17106 48020 17388
rect 47964 17054 47966 17106
rect 48018 17054 48020 17106
rect 47964 17042 48020 17054
rect 47740 16996 47796 17006
rect 47740 16994 47908 16996
rect 47740 16942 47742 16994
rect 47794 16942 47908 16994
rect 47740 16940 47908 16942
rect 47740 16930 47796 16940
rect 47628 16884 47684 16894
rect 47516 16882 47684 16884
rect 47516 16830 47630 16882
rect 47682 16830 47684 16882
rect 47516 16828 47684 16830
rect 47516 16324 47572 16334
rect 47628 16324 47684 16828
rect 47852 16436 47908 16940
rect 48188 16772 48244 18286
rect 48748 17556 48804 17566
rect 48748 16994 48804 17500
rect 48748 16942 48750 16994
rect 48802 16942 48804 16994
rect 48748 16930 48804 16942
rect 48188 16706 48244 16716
rect 48748 16772 48804 16782
rect 47852 16370 47908 16380
rect 47572 16268 47684 16324
rect 48748 16322 48804 16716
rect 48748 16270 48750 16322
rect 48802 16270 48804 16322
rect 47516 16258 47572 16268
rect 48412 16212 48468 16222
rect 47628 16210 48468 16212
rect 47628 16158 48414 16210
rect 48466 16158 48468 16210
rect 47628 16156 48468 16158
rect 47516 16100 47572 16110
rect 47516 16006 47572 16044
rect 47516 15316 47572 15326
rect 47628 15316 47684 16156
rect 48412 16146 48468 16156
rect 48076 15988 48132 15998
rect 47964 15876 48020 15886
rect 47964 15538 48020 15820
rect 47964 15486 47966 15538
rect 48018 15486 48020 15538
rect 47964 15474 48020 15486
rect 47740 15428 47796 15438
rect 47740 15334 47796 15372
rect 48076 15426 48132 15932
rect 48748 15988 48804 16270
rect 48748 15922 48804 15932
rect 48524 15876 48580 15886
rect 48524 15782 48580 15820
rect 48076 15374 48078 15426
rect 48130 15374 48132 15426
rect 48076 15362 48132 15374
rect 47516 15314 47684 15316
rect 47516 15262 47518 15314
rect 47570 15262 47684 15314
rect 47516 15260 47684 15262
rect 47516 15250 47572 15260
rect 47180 15092 47460 15148
rect 46844 14702 46846 14754
rect 46898 14702 46900 14754
rect 46844 14690 46900 14702
rect 47068 14868 47124 14878
rect 46620 14418 46676 14430
rect 46620 14366 46622 14418
rect 46674 14366 46676 14418
rect 46620 13972 46676 14366
rect 46620 13906 46676 13916
rect 47068 14084 47124 14812
rect 47180 14754 47236 15092
rect 48860 14980 48916 18396
rect 48972 15148 49028 21196
rect 49980 20468 50036 22540
rect 50092 22502 50148 22540
rect 50428 22370 50484 22988
rect 50876 22708 50932 23102
rect 50988 23156 51044 23166
rect 50988 23062 51044 23100
rect 50876 22642 50932 22652
rect 50988 22596 51044 22606
rect 50988 22502 51044 22540
rect 51324 22594 51380 23214
rect 52220 23268 52276 23278
rect 51324 22542 51326 22594
rect 51378 22542 51380 22594
rect 51324 22530 51380 22542
rect 51884 23154 51940 23166
rect 51884 23102 51886 23154
rect 51938 23102 51940 23154
rect 51884 22484 51940 23102
rect 52220 23154 52276 23212
rect 53564 23268 53620 23886
rect 53564 23202 53620 23212
rect 52220 23102 52222 23154
rect 52274 23102 52276 23154
rect 52220 23090 52276 23102
rect 50428 22318 50430 22370
rect 50482 22318 50484 22370
rect 50428 22306 50484 22318
rect 51772 22428 51940 22484
rect 52668 23042 52724 23054
rect 52668 22990 52670 23042
rect 52722 22990 52724 23042
rect 51660 22258 51716 22270
rect 51660 22206 51662 22258
rect 51714 22206 51716 22258
rect 50204 22146 50260 22158
rect 51212 22148 51268 22158
rect 50204 22094 50206 22146
rect 50258 22094 50260 22146
rect 50092 21924 50148 21934
rect 50092 21698 50148 21868
rect 50092 21646 50094 21698
rect 50146 21646 50148 21698
rect 50092 21634 50148 21646
rect 50204 21700 50260 22094
rect 50876 22146 51492 22148
rect 50876 22094 51214 22146
rect 51266 22094 51492 22146
rect 50876 22092 51492 22094
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50204 21634 50260 21644
rect 50316 21810 50372 21822
rect 50316 21758 50318 21810
rect 50370 21758 50372 21810
rect 50204 20916 50260 20926
rect 50204 20822 50260 20860
rect 50316 20802 50372 21758
rect 50540 21700 50596 21710
rect 50428 21588 50484 21598
rect 50428 21494 50484 21532
rect 50540 21586 50596 21644
rect 50540 21534 50542 21586
rect 50594 21534 50596 21586
rect 50540 21522 50596 21534
rect 50316 20750 50318 20802
rect 50370 20750 50372 20802
rect 50316 20738 50372 20750
rect 50876 20802 50932 22092
rect 51212 22082 51268 22092
rect 50876 20750 50878 20802
rect 50930 20750 50932 20802
rect 50876 20738 50932 20750
rect 51100 21812 51156 21822
rect 49980 20412 50260 20468
rect 50204 20130 50260 20412
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50204 20078 50206 20130
rect 50258 20078 50260 20130
rect 50204 20066 50260 20078
rect 50876 20018 50932 20030
rect 50876 19966 50878 20018
rect 50930 19966 50932 20018
rect 49980 19908 50036 19918
rect 49980 19346 50036 19852
rect 49980 19294 49982 19346
rect 50034 19294 50036 19346
rect 49980 19282 50036 19294
rect 50428 19010 50484 19022
rect 50428 18958 50430 19010
rect 50482 18958 50484 19010
rect 49756 18452 49812 18462
rect 49756 17780 49812 18396
rect 50428 18452 50484 18958
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50428 18386 50484 18396
rect 49756 17778 50036 17780
rect 49756 17726 49758 17778
rect 49810 17726 50036 17778
rect 49756 17724 50036 17726
rect 49756 17714 49812 17724
rect 49420 16882 49476 16894
rect 49420 16830 49422 16882
rect 49474 16830 49476 16882
rect 49196 16772 49252 16782
rect 49196 16678 49252 16716
rect 49420 16772 49476 16830
rect 49420 16548 49476 16716
rect 49420 16492 49700 16548
rect 49084 16436 49140 16446
rect 49084 16322 49140 16380
rect 49084 16270 49086 16322
rect 49138 16270 49140 16322
rect 49084 16258 49140 16270
rect 49644 16210 49700 16492
rect 49644 16158 49646 16210
rect 49698 16158 49700 16210
rect 49644 16146 49700 16158
rect 49980 16212 50036 17724
rect 50764 17668 50820 17678
rect 50876 17668 50932 19966
rect 51100 20018 51156 21756
rect 51436 20132 51492 22092
rect 51660 21812 51716 22206
rect 51772 22260 51828 22428
rect 51772 22166 51828 22204
rect 51996 22370 52052 22382
rect 51996 22318 51998 22370
rect 52050 22318 52052 22370
rect 51660 21700 51716 21756
rect 51996 21700 52052 22318
rect 52668 22258 52724 22990
rect 52780 22708 52836 22718
rect 52780 22482 52836 22652
rect 52780 22430 52782 22482
rect 52834 22430 52836 22482
rect 52780 22418 52836 22430
rect 52668 22206 52670 22258
rect 52722 22206 52724 22258
rect 52668 22148 52724 22206
rect 52892 22260 52948 22270
rect 52892 22166 52948 22204
rect 51660 21644 51828 21700
rect 51548 21588 51604 21598
rect 51548 21028 51604 21532
rect 51548 20962 51604 20972
rect 51772 20916 51828 21644
rect 51996 21634 52052 21644
rect 52332 22092 52724 22148
rect 53452 22146 53508 22158
rect 53452 22094 53454 22146
rect 53506 22094 53508 22146
rect 52108 21586 52164 21598
rect 52108 21534 52110 21586
rect 52162 21534 52164 21586
rect 52108 21476 52164 21534
rect 51996 20916 52052 20926
rect 51772 20914 52052 20916
rect 51772 20862 51998 20914
rect 52050 20862 52052 20914
rect 51772 20860 52052 20862
rect 51548 20804 51604 20814
rect 51548 20710 51604 20748
rect 51996 20580 52052 20860
rect 52108 20804 52164 21420
rect 52332 21474 52388 22092
rect 53452 22036 53508 22094
rect 53788 22148 53844 22158
rect 53788 22054 53844 22092
rect 52892 21812 52948 21822
rect 52892 21718 52948 21756
rect 52444 21700 52500 21710
rect 52444 21606 52500 21644
rect 53116 21700 53172 21710
rect 52332 21422 52334 21474
rect 52386 21422 52388 21474
rect 52332 21410 52388 21422
rect 52668 21028 52724 21038
rect 52668 20934 52724 20972
rect 53116 21026 53172 21644
rect 53116 20974 53118 21026
rect 53170 20974 53172 21026
rect 53116 20962 53172 20974
rect 53340 21476 53396 21486
rect 53452 21476 53508 21980
rect 53340 21474 53508 21476
rect 53340 21422 53342 21474
rect 53394 21422 53508 21474
rect 53340 21420 53508 21422
rect 53676 21812 53732 21822
rect 53340 21362 53396 21420
rect 53340 21310 53342 21362
rect 53394 21310 53396 21362
rect 52108 20738 52164 20748
rect 52220 20916 52276 20926
rect 51996 20514 52052 20524
rect 51548 20132 51604 20142
rect 51436 20130 51604 20132
rect 51436 20078 51550 20130
rect 51602 20078 51604 20130
rect 51436 20076 51604 20078
rect 51548 20066 51604 20076
rect 51100 19966 51102 20018
rect 51154 19966 51156 20018
rect 51100 19954 51156 19966
rect 52220 20018 52276 20860
rect 53228 20916 53284 20926
rect 53228 20822 53284 20860
rect 52220 19966 52222 20018
rect 52274 19966 52276 20018
rect 52220 19954 52276 19966
rect 52444 20804 52500 20814
rect 52444 20020 52500 20748
rect 52444 19926 52500 19964
rect 52780 20690 52836 20702
rect 53340 20692 53396 21310
rect 53676 20914 53732 21756
rect 53788 21474 53844 21486
rect 53788 21422 53790 21474
rect 53842 21422 53844 21474
rect 53788 21362 53844 21422
rect 53788 21310 53790 21362
rect 53842 21310 53844 21362
rect 53788 21298 53844 21310
rect 53676 20862 53678 20914
rect 53730 20862 53732 20914
rect 53676 20850 53732 20862
rect 52780 20638 52782 20690
rect 52834 20638 52836 20690
rect 52780 19124 52836 20638
rect 51996 18452 52052 18462
rect 51996 18358 52052 18396
rect 52332 18340 52388 18350
rect 52780 18340 52836 19068
rect 53116 20636 53396 20692
rect 52332 18338 52836 18340
rect 52332 18286 52334 18338
rect 52386 18286 52836 18338
rect 52332 18284 52836 18286
rect 53004 18452 53060 18462
rect 51212 17780 51268 17790
rect 51660 17780 51716 17790
rect 51212 17778 51716 17780
rect 51212 17726 51214 17778
rect 51266 17726 51662 17778
rect 51714 17726 51716 17778
rect 51212 17724 51716 17726
rect 51212 17714 51268 17724
rect 51660 17714 51716 17724
rect 50820 17612 50932 17668
rect 52332 17668 52388 18284
rect 50764 17574 50820 17612
rect 52332 17602 52388 17612
rect 51212 17554 51268 17566
rect 51212 17502 51214 17554
rect 51266 17502 51268 17554
rect 50876 17442 50932 17454
rect 50876 17390 50878 17442
rect 50930 17390 50932 17442
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50092 16772 50148 16782
rect 50092 16678 50148 16716
rect 50652 16772 50708 16782
rect 50092 16212 50148 16222
rect 49980 16210 50148 16212
rect 49980 16158 50094 16210
rect 50146 16158 50148 16210
rect 49980 16156 50148 16158
rect 50092 16146 50148 16156
rect 49196 16100 49252 16110
rect 49252 16044 49476 16100
rect 49196 16006 49252 16044
rect 49420 15428 49476 16044
rect 50652 16098 50708 16716
rect 50652 16046 50654 16098
rect 50706 16046 50708 16098
rect 50652 16034 50708 16046
rect 50764 16100 50820 16110
rect 50876 16100 50932 17390
rect 51100 17442 51156 17454
rect 51100 17390 51102 17442
rect 51154 17390 51156 17442
rect 51100 16772 51156 17390
rect 51212 17444 51268 17502
rect 51324 17444 51380 17454
rect 51212 17388 51324 17444
rect 51324 17378 51380 17388
rect 51772 17444 51828 17454
rect 51772 17442 52276 17444
rect 51772 17390 51774 17442
rect 51826 17390 52276 17442
rect 51772 17388 52276 17390
rect 51772 17378 51828 17388
rect 52220 16994 52276 17388
rect 52220 16942 52222 16994
rect 52274 16942 52276 16994
rect 52220 16930 52276 16942
rect 51100 16706 51156 16716
rect 53004 16882 53060 18396
rect 53004 16830 53006 16882
rect 53058 16830 53060 16882
rect 50820 16044 50932 16100
rect 50764 16006 50820 16044
rect 50540 15988 50596 15998
rect 49532 15876 49588 15886
rect 49868 15876 49924 15886
rect 50540 15876 50596 15932
rect 50988 15988 51044 16026
rect 50988 15922 51044 15932
rect 51548 15986 51604 15998
rect 51548 15934 51550 15986
rect 51602 15934 51604 15986
rect 49532 15782 49588 15820
rect 49644 15820 49868 15876
rect 49420 15334 49476 15372
rect 49644 15426 49700 15820
rect 49868 15810 49924 15820
rect 50428 15820 50596 15876
rect 50876 15874 50932 15886
rect 50876 15822 50878 15874
rect 50930 15822 50932 15874
rect 49644 15374 49646 15426
rect 49698 15374 49700 15426
rect 48972 15092 49588 15148
rect 48860 14924 49140 14980
rect 47180 14702 47182 14754
rect 47234 14702 47236 14754
rect 47180 14690 47236 14702
rect 48524 14644 48580 14654
rect 48524 14550 48580 14588
rect 48860 14642 48916 14654
rect 48860 14590 48862 14642
rect 48914 14590 48916 14642
rect 48860 14532 48916 14590
rect 49084 14644 49140 14924
rect 49140 14588 49364 14644
rect 49084 14578 49140 14588
rect 48860 14466 48916 14476
rect 47068 14028 47460 14084
rect 47068 13970 47124 14028
rect 47068 13918 47070 13970
rect 47122 13918 47124 13970
rect 47068 13906 47124 13918
rect 46508 13858 46564 13870
rect 46508 13806 46510 13858
rect 46562 13806 46564 13858
rect 46508 13748 46564 13806
rect 47292 13860 47348 13870
rect 47292 13766 47348 13804
rect 46844 13748 46900 13758
rect 46508 13746 46900 13748
rect 46508 13694 46846 13746
rect 46898 13694 46900 13746
rect 46508 13692 46900 13694
rect 46508 9828 46564 13692
rect 46844 13682 46900 13692
rect 47180 13634 47236 13646
rect 47180 13582 47182 13634
rect 47234 13582 47236 13634
rect 47180 13524 47236 13582
rect 46956 13468 47236 13524
rect 46956 13074 47012 13468
rect 46956 13022 46958 13074
rect 47010 13022 47012 13074
rect 46956 13010 47012 13022
rect 47068 12740 47124 12750
rect 47068 12738 47348 12740
rect 47068 12686 47070 12738
rect 47122 12686 47348 12738
rect 47068 12684 47348 12686
rect 47068 12674 47124 12684
rect 47292 11396 47348 12684
rect 47404 11620 47460 14028
rect 47516 13972 47572 13982
rect 47516 13858 47572 13916
rect 47516 13806 47518 13858
rect 47570 13806 47572 13858
rect 47516 13794 47572 13806
rect 49084 13636 49140 13646
rect 49084 11732 49140 13580
rect 49084 11666 49140 11676
rect 47404 11554 47460 11564
rect 49308 11508 49364 14588
rect 49420 14532 49476 14542
rect 49420 13970 49476 14476
rect 49420 13918 49422 13970
rect 49474 13918 49476 13970
rect 49420 13906 49476 13918
rect 48748 11506 49364 11508
rect 48748 11454 49310 11506
rect 49362 11454 49364 11506
rect 48748 11452 49364 11454
rect 47964 11396 48020 11406
rect 47292 11394 48020 11396
rect 47292 11342 47966 11394
rect 48018 11342 48020 11394
rect 47292 11340 48020 11342
rect 47964 11330 48020 11340
rect 48748 11394 48804 11452
rect 49308 11442 49364 11452
rect 48748 11342 48750 11394
rect 48802 11342 48804 11394
rect 48748 11330 48804 11342
rect 46508 9762 46564 9772
rect 46284 3938 46340 3948
rect 49532 3780 49588 15092
rect 49644 13860 49700 15374
rect 50092 15540 50148 15550
rect 49868 15314 49924 15326
rect 49868 15262 49870 15314
rect 49922 15262 49924 15314
rect 49756 15202 49812 15214
rect 49756 15150 49758 15202
rect 49810 15150 49812 15202
rect 49756 14196 49812 15150
rect 49756 14130 49812 14140
rect 49756 13972 49812 13982
rect 49868 13972 49924 15262
rect 50092 15314 50148 15484
rect 50092 15262 50094 15314
rect 50146 15262 50148 15314
rect 50092 15250 50148 15262
rect 50428 15428 50484 15820
rect 50876 15764 50932 15822
rect 51100 15876 51156 15886
rect 50988 15764 51044 15774
rect 50556 15708 50820 15718
rect 50876 15708 50988 15764
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50988 15698 51044 15708
rect 50556 15642 50820 15652
rect 51100 15540 51156 15820
rect 51548 15764 51604 15934
rect 51660 15876 51716 15886
rect 51660 15782 51716 15820
rect 52556 15876 52612 15886
rect 51548 15698 51604 15708
rect 51100 15474 51156 15484
rect 50428 15202 50484 15372
rect 52556 15426 52612 15820
rect 52556 15374 52558 15426
rect 52610 15374 52612 15426
rect 52556 15362 52612 15374
rect 52780 15876 52836 15886
rect 50428 15150 50430 15202
rect 50482 15150 50484 15202
rect 50428 15138 50484 15150
rect 52780 15204 52836 15820
rect 53004 15316 53060 16830
rect 53116 15876 53172 20636
rect 53900 19908 53956 25228
rect 54460 22260 54516 22270
rect 54572 22260 54628 26852
rect 54796 25620 54852 25630
rect 54684 24948 54740 24958
rect 54684 24854 54740 24892
rect 54796 24836 54852 25564
rect 54908 25620 54964 27020
rect 55244 27010 55300 27020
rect 55356 26908 55412 28028
rect 55692 27860 55748 27870
rect 55692 27188 55748 27804
rect 55692 27122 55748 27132
rect 56028 27186 56084 28364
rect 56140 27412 56196 28700
rect 56364 28754 56420 31164
rect 56700 31220 56756 31230
rect 56700 31126 56756 31164
rect 58156 30324 58212 30334
rect 58156 30230 58212 30268
rect 57148 29652 57204 29662
rect 57148 29558 57204 29596
rect 57596 29652 57652 29662
rect 57484 29426 57540 29438
rect 57484 29374 57486 29426
rect 57538 29374 57540 29426
rect 56924 29316 56980 29326
rect 57484 29316 57540 29374
rect 56924 29314 57540 29316
rect 56924 29262 56926 29314
rect 56978 29262 57540 29314
rect 56924 29260 57540 29262
rect 56924 29250 56980 29260
rect 57484 28980 57540 29260
rect 57484 28914 57540 28924
rect 56364 28702 56366 28754
rect 56418 28702 56420 28754
rect 56364 28644 56420 28702
rect 57596 28754 57652 29596
rect 58156 29652 58212 29662
rect 58156 29558 58212 29596
rect 57820 29538 57876 29550
rect 57820 29486 57822 29538
rect 57874 29486 57876 29538
rect 57820 29204 57876 29486
rect 57820 29138 57876 29148
rect 57596 28702 57598 28754
rect 57650 28702 57652 28754
rect 57596 28690 57652 28702
rect 57820 28756 57876 28766
rect 56364 28578 56420 28588
rect 57148 28644 57204 28654
rect 57148 28550 57204 28588
rect 57820 28418 57876 28700
rect 57820 28366 57822 28418
rect 57874 28366 57876 28418
rect 57820 28354 57876 28366
rect 58156 28644 58212 28654
rect 58156 28308 58212 28588
rect 58156 28242 58212 28252
rect 57820 27970 57876 27982
rect 57820 27918 57822 27970
rect 57874 27918 57876 27970
rect 56140 27346 56196 27356
rect 57148 27746 57204 27758
rect 57148 27694 57150 27746
rect 57202 27694 57204 27746
rect 56028 27134 56030 27186
rect 56082 27134 56084 27186
rect 56028 27122 56084 27134
rect 55132 26852 55412 26908
rect 57148 26908 57204 27694
rect 57596 27746 57652 27758
rect 57596 27694 57598 27746
rect 57650 27694 57652 27746
rect 57596 27636 57652 27694
rect 57596 27570 57652 27580
rect 57820 27300 57876 27918
rect 58156 27858 58212 27870
rect 58156 27806 58158 27858
rect 58210 27806 58212 27858
rect 58156 27636 58212 27806
rect 58156 27570 58212 27580
rect 57820 27234 57876 27244
rect 58156 27188 58212 27198
rect 58156 27094 58212 27132
rect 57148 26852 57540 26908
rect 55132 26290 55188 26852
rect 55244 26516 55300 26526
rect 55244 26422 55300 26460
rect 57148 26402 57204 26414
rect 57148 26350 57150 26402
rect 57202 26350 57204 26402
rect 55132 26238 55134 26290
rect 55186 26238 55188 26290
rect 55132 26226 55188 26238
rect 55468 26290 55524 26302
rect 55468 26238 55470 26290
rect 55522 26238 55524 26290
rect 55356 26180 55412 26190
rect 55356 26086 55412 26124
rect 55468 25620 55524 26238
rect 54908 25618 55300 25620
rect 54908 25566 54910 25618
rect 54962 25566 55300 25618
rect 54908 25564 55300 25566
rect 54908 25554 54964 25564
rect 54908 24836 54964 24846
rect 54796 24834 54964 24836
rect 54796 24782 54910 24834
rect 54962 24782 54964 24834
rect 54796 24780 54964 24782
rect 54908 24770 54964 24780
rect 54796 24052 54852 24062
rect 55020 24052 55076 25564
rect 55244 25506 55300 25564
rect 55468 25554 55524 25564
rect 55580 26290 55636 26302
rect 55580 26238 55582 26290
rect 55634 26238 55636 26290
rect 55244 25454 55246 25506
rect 55298 25454 55300 25506
rect 55244 25442 55300 25454
rect 55356 25172 55412 25182
rect 55356 24946 55412 25116
rect 55356 24894 55358 24946
rect 55410 24894 55412 24946
rect 54796 24050 55076 24052
rect 54796 23998 54798 24050
rect 54850 23998 55076 24050
rect 54796 23996 55076 23998
rect 54796 23986 54852 23996
rect 55020 23938 55076 23996
rect 55020 23886 55022 23938
rect 55074 23886 55076 23938
rect 55020 23874 55076 23886
rect 55132 24722 55188 24734
rect 55132 24670 55134 24722
rect 55186 24670 55188 24722
rect 54796 23268 54852 23278
rect 54460 22258 54628 22260
rect 54460 22206 54462 22258
rect 54514 22206 54628 22258
rect 54460 22204 54628 22206
rect 54684 23212 54796 23268
rect 54460 22194 54516 22204
rect 54124 22146 54180 22158
rect 54124 22094 54126 22146
rect 54178 22094 54180 22146
rect 54124 22036 54180 22094
rect 54124 21970 54180 21980
rect 54684 21698 54740 23212
rect 54796 23202 54852 23212
rect 55132 22932 55188 24670
rect 55244 24612 55300 24622
rect 55244 24518 55300 24556
rect 55356 24388 55412 24894
rect 55244 24332 55412 24388
rect 55580 24722 55636 26238
rect 56700 26180 56756 26190
rect 56700 26086 56756 26124
rect 56588 26068 56644 26078
rect 56028 26066 56644 26068
rect 56028 26014 56590 26066
rect 56642 26014 56644 26066
rect 56028 26012 56644 26014
rect 56028 25618 56084 26012
rect 56588 26002 56644 26012
rect 57148 26068 57204 26350
rect 57484 26292 57540 26852
rect 57820 26852 57876 26862
rect 57820 26514 57876 26796
rect 57820 26462 57822 26514
rect 57874 26462 57876 26514
rect 57820 26450 57876 26462
rect 58044 26852 58100 26862
rect 57484 26198 57540 26236
rect 58044 26290 58100 26796
rect 58044 26238 58046 26290
rect 58098 26238 58100 26290
rect 57148 26002 57204 26012
rect 56028 25566 56030 25618
rect 56082 25566 56084 25618
rect 56028 25554 56084 25566
rect 56924 25956 56980 25966
rect 56924 24946 56980 25900
rect 58044 25956 58100 26238
rect 58044 25890 58100 25900
rect 57036 25844 57092 25854
rect 57036 25060 57092 25788
rect 58156 25620 58212 25630
rect 58156 25526 58212 25564
rect 57036 24994 57092 25004
rect 57596 25172 57652 25182
rect 56924 24894 56926 24946
rect 56978 24894 56980 24946
rect 56924 24882 56980 24894
rect 57484 24948 57540 24958
rect 57484 24854 57540 24892
rect 55580 24670 55582 24722
rect 55634 24670 55636 24722
rect 55244 24052 55300 24332
rect 55244 23154 55300 23996
rect 55580 23492 55636 24670
rect 57148 24834 57204 24846
rect 57148 24782 57150 24834
rect 57202 24782 57204 24834
rect 56028 24612 56084 24622
rect 56028 24518 56084 24556
rect 55916 24500 55972 24510
rect 55804 24498 55972 24500
rect 55804 24446 55918 24498
rect 55970 24446 55972 24498
rect 55804 24444 55972 24446
rect 55804 24050 55860 24444
rect 55916 24434 55972 24444
rect 57148 24500 57204 24782
rect 57148 24434 57204 24444
rect 55804 23998 55806 24050
rect 55858 23998 55860 24050
rect 55804 23986 55860 23998
rect 57484 23492 57540 23502
rect 55580 23436 55748 23492
rect 55580 23268 55636 23278
rect 55580 23174 55636 23212
rect 55244 23102 55246 23154
rect 55298 23102 55300 23154
rect 55244 23090 55300 23102
rect 55356 23154 55412 23166
rect 55356 23102 55358 23154
rect 55410 23102 55412 23154
rect 55356 22932 55412 23102
rect 55692 23154 55748 23436
rect 55692 23102 55694 23154
rect 55746 23102 55748 23154
rect 55468 23044 55524 23054
rect 55468 22950 55524 22988
rect 54684 21646 54686 21698
rect 54738 21646 54740 21698
rect 54684 21634 54740 21646
rect 54796 22876 55412 22932
rect 53788 19906 53956 19908
rect 53788 19854 53902 19906
rect 53954 19854 53956 19906
rect 53788 19852 53956 19854
rect 53676 19236 53732 19246
rect 53676 19142 53732 19180
rect 53452 19124 53508 19134
rect 53452 19030 53508 19068
rect 53340 19010 53396 19022
rect 53340 18958 53342 19010
rect 53394 18958 53396 19010
rect 53340 17444 53396 18958
rect 53564 19010 53620 19022
rect 53564 18958 53566 19010
rect 53618 18958 53620 19010
rect 53564 18564 53620 18958
rect 53788 19012 53844 19852
rect 53900 19842 53956 19852
rect 54012 21588 54068 21598
rect 54012 20916 54068 21532
rect 54796 21588 54852 22876
rect 55692 22820 55748 23102
rect 57148 23266 57204 23278
rect 57484 23268 57540 23436
rect 57148 23214 57150 23266
rect 57202 23214 57204 23266
rect 56700 23044 56756 23054
rect 56700 22950 56756 22988
rect 56588 22932 56644 22942
rect 55356 22764 55748 22820
rect 56028 22930 56644 22932
rect 56028 22878 56590 22930
rect 56642 22878 56644 22930
rect 56028 22876 56644 22878
rect 54908 22372 54964 22382
rect 55244 22372 55300 22382
rect 54908 22370 55300 22372
rect 54908 22318 54910 22370
rect 54962 22318 55246 22370
rect 55298 22318 55300 22370
rect 54908 22316 55300 22318
rect 54908 21812 54964 22316
rect 55244 22306 55300 22316
rect 54908 21746 54964 21756
rect 55244 22148 55300 22158
rect 55356 22148 55412 22764
rect 56028 22482 56084 22876
rect 56588 22866 56644 22876
rect 57148 22820 57204 23214
rect 57148 22754 57204 22764
rect 57260 23266 57540 23268
rect 57260 23214 57486 23266
rect 57538 23214 57540 23266
rect 57260 23212 57540 23214
rect 56028 22430 56030 22482
rect 56082 22430 56084 22482
rect 56028 22418 56084 22430
rect 57036 22484 57092 22494
rect 55300 22092 55412 22148
rect 55244 21810 55300 22092
rect 55244 21758 55246 21810
rect 55298 21758 55300 21810
rect 55244 21746 55300 21758
rect 55356 21812 55412 21822
rect 54908 21588 54964 21598
rect 54796 21586 54964 21588
rect 54796 21534 54910 21586
rect 54962 21534 54964 21586
rect 54796 21532 54964 21534
rect 54796 21476 54852 21532
rect 54908 21522 54964 21532
rect 55132 21588 55188 21598
rect 55132 21494 55188 21532
rect 53900 19236 53956 19246
rect 54012 19236 54068 20860
rect 53900 19234 54068 19236
rect 53900 19182 53902 19234
rect 53954 19182 54068 19234
rect 53900 19180 54068 19182
rect 54572 21420 54852 21476
rect 55020 21476 55076 21486
rect 54572 19236 54628 21420
rect 55020 21382 55076 21420
rect 53900 19170 53956 19180
rect 54572 19122 54628 19180
rect 54572 19070 54574 19122
rect 54626 19070 54628 19122
rect 54572 19058 54628 19070
rect 54236 19012 54292 19022
rect 53788 19010 54292 19012
rect 53788 18958 54238 19010
rect 54290 18958 54292 19010
rect 53788 18956 54292 18958
rect 53452 18508 53620 18564
rect 53452 17778 53508 18508
rect 53564 18340 53620 18350
rect 53564 17890 53620 18284
rect 53564 17838 53566 17890
rect 53618 17838 53620 17890
rect 53564 17826 53620 17838
rect 53452 17726 53454 17778
rect 53506 17726 53508 17778
rect 53452 17714 53508 17726
rect 53340 15988 53396 17388
rect 53452 15988 53508 15998
rect 53340 15986 53508 15988
rect 53340 15934 53454 15986
rect 53506 15934 53508 15986
rect 53340 15932 53508 15934
rect 53452 15922 53508 15932
rect 53116 15782 53172 15820
rect 53228 15316 53284 15326
rect 53004 15314 53284 15316
rect 53004 15262 53230 15314
rect 53282 15262 53284 15314
rect 53004 15260 53284 15262
rect 53228 15250 53284 15260
rect 52780 15138 52836 15148
rect 51660 14644 51716 14654
rect 51660 14530 51716 14588
rect 51660 14478 51662 14530
rect 51714 14478 51716 14530
rect 51660 14466 51716 14478
rect 50988 14418 51044 14430
rect 50988 14366 50990 14418
rect 51042 14366 51044 14418
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 49812 13916 49924 13972
rect 50764 13972 50820 13982
rect 49756 13878 49812 13916
rect 49644 13794 49700 13804
rect 50092 13860 50148 13870
rect 50092 13766 50148 13804
rect 50764 13858 50820 13916
rect 50876 13972 50932 13982
rect 50988 13972 51044 14366
rect 50876 13970 51044 13972
rect 50876 13918 50878 13970
rect 50930 13918 51044 13970
rect 50876 13916 51044 13918
rect 50876 13906 50932 13916
rect 50764 13806 50766 13858
rect 50818 13806 50820 13858
rect 50764 13794 50820 13806
rect 54236 13860 54292 18956
rect 55244 18452 55300 18462
rect 55356 18452 55412 21756
rect 56812 21812 56868 21822
rect 55692 21476 55748 21486
rect 55692 21382 55748 21420
rect 55804 21364 55860 21374
rect 55804 21362 56196 21364
rect 55804 21310 55806 21362
rect 55858 21310 56196 21362
rect 55804 21308 56196 21310
rect 55804 21298 55860 21308
rect 56140 20914 56196 21308
rect 56140 20862 56142 20914
rect 56194 20862 56196 20914
rect 56140 20850 56196 20862
rect 56812 20802 56868 21756
rect 57036 21812 57092 22428
rect 57036 21746 57092 21756
rect 57148 21812 57204 21822
rect 57260 21812 57316 23212
rect 57484 23202 57540 23212
rect 57148 21810 57316 21812
rect 57148 21758 57150 21810
rect 57202 21758 57316 21810
rect 57148 21756 57316 21758
rect 57596 21810 57652 25116
rect 58156 25172 58212 25182
rect 57820 25060 57876 25070
rect 57820 24946 57876 25004
rect 57820 24894 57822 24946
rect 57874 24894 57876 24946
rect 57820 24882 57876 24894
rect 58156 24946 58212 25116
rect 58156 24894 58158 24946
rect 58210 24894 58212 24946
rect 58156 24882 58212 24894
rect 58156 24276 58212 24286
rect 57932 24052 57988 24062
rect 57932 23958 57988 23996
rect 57820 23380 57876 23390
rect 57820 23286 57876 23324
rect 57932 23268 57988 23278
rect 58156 23268 58212 24220
rect 57988 23212 58100 23268
rect 57932 23202 57988 23212
rect 58044 22484 58100 23212
rect 58156 23266 58324 23268
rect 58156 23214 58158 23266
rect 58210 23214 58324 23266
rect 58156 23212 58324 23214
rect 58156 23202 58212 23212
rect 58156 22484 58212 22494
rect 58044 22482 58212 22484
rect 58044 22430 58158 22482
rect 58210 22430 58212 22482
rect 58044 22428 58212 22430
rect 58156 22418 58212 22428
rect 58156 22260 58212 22270
rect 57596 21758 57598 21810
rect 57650 21758 57652 21810
rect 57148 21746 57204 21756
rect 57596 21746 57652 21758
rect 57820 21812 57876 21822
rect 58156 21812 58212 22204
rect 57820 21718 57876 21756
rect 57932 21810 58212 21812
rect 57932 21758 58158 21810
rect 58210 21758 58212 21810
rect 57932 21756 58212 21758
rect 57820 20916 57876 20926
rect 57932 20916 57988 21756
rect 58156 21746 58212 21756
rect 57820 20914 57988 20916
rect 57820 20862 57822 20914
rect 57874 20862 57988 20914
rect 57820 20860 57988 20862
rect 58268 20914 58324 23212
rect 58268 20862 58270 20914
rect 58322 20862 58324 20914
rect 57820 20850 57876 20860
rect 58268 20850 58324 20862
rect 56812 20750 56814 20802
rect 56866 20750 56868 20802
rect 56812 20738 56868 20750
rect 55300 18396 55412 18452
rect 55244 18358 55300 18396
rect 54460 18340 54516 18350
rect 54460 18246 54516 18284
rect 54236 13794 54292 13804
rect 50316 13746 50372 13758
rect 50316 13694 50318 13746
rect 50370 13694 50372 13746
rect 50316 13636 50372 13694
rect 50316 13570 50372 13580
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 49532 3714 49588 3724
rect 40460 3390 40462 3442
rect 40514 3390 40516 3442
rect 40460 3378 40516 3390
rect 40684 3554 40740 3566
rect 40684 3502 40686 3554
rect 40738 3502 40740 3554
rect 40684 3444 40740 3502
rect 40684 3378 40740 3388
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 39004 2492 39620 2548
rect 39676 2716 39956 2772
rect 39004 800 39060 2492
rect 39676 800 39732 2716
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 24192 0 24304 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 31584 0 31696 800
rect 32256 0 32368 800
rect 32928 0 33040 800
rect 33600 0 33712 800
rect 34272 0 34384 800
rect 34944 0 35056 800
rect 35616 0 35728 800
rect 36288 0 36400 800
rect 36960 0 37072 800
rect 37632 0 37744 800
rect 38304 0 38416 800
rect 38976 0 39088 800
rect 39648 0 39760 800
<< via2 >>
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 20188 56082 20244 56084
rect 20188 56030 20190 56082
rect 20190 56030 20242 56082
rect 20242 56030 20244 56082
rect 20188 56028 20244 56030
rect 20860 56028 20916 56084
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 8764 55132 8820 55188
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 2044 49922 2100 49924
rect 2044 49870 2046 49922
rect 2046 49870 2098 49922
rect 2098 49870 2100 49922
rect 2044 49868 2100 49870
rect 1932 49756 1988 49812
rect 1708 49644 1764 49700
rect 2492 49698 2548 49700
rect 2492 49646 2494 49698
rect 2494 49646 2546 49698
rect 2546 49646 2548 49698
rect 2492 49644 2548 49646
rect 1708 49084 1764 49140
rect 1708 48412 1764 48468
rect 2044 48354 2100 48356
rect 2044 48302 2046 48354
rect 2046 48302 2098 48354
rect 2098 48302 2100 48354
rect 2044 48300 2100 48302
rect 1708 47740 1764 47796
rect 2044 47234 2100 47236
rect 2044 47182 2046 47234
rect 2046 47182 2098 47234
rect 2098 47182 2100 47234
rect 2044 47180 2100 47182
rect 1708 47068 1764 47124
rect 2492 48412 2548 48468
rect 2492 47740 2548 47796
rect 2492 47068 2548 47124
rect 3612 47180 3668 47236
rect 1708 46396 1764 46452
rect 2380 45778 2436 45780
rect 2380 45726 2382 45778
rect 2382 45726 2434 45778
rect 2434 45726 2436 45778
rect 2380 45724 2436 45726
rect 2044 45218 2100 45220
rect 2044 45166 2046 45218
rect 2046 45166 2098 45218
rect 2098 45166 2100 45218
rect 2044 45164 2100 45166
rect 1820 45052 1876 45108
rect 1708 44940 1764 44996
rect 2492 44994 2548 44996
rect 2492 44942 2494 44994
rect 2494 44942 2546 44994
rect 2546 44942 2548 44994
rect 2492 44940 2548 44942
rect 2156 44492 2212 44548
rect 1708 44380 1764 44436
rect 1932 43708 1988 43764
rect 2044 43650 2100 43652
rect 2044 43598 2046 43650
rect 2046 43598 2098 43650
rect 2098 43598 2100 43650
rect 2044 43596 2100 43598
rect 1708 43036 1764 43092
rect 2492 43036 2548 43092
rect 2156 42700 2212 42756
rect 2044 42642 2100 42644
rect 2044 42590 2046 42642
rect 2046 42590 2098 42642
rect 2098 42590 2100 42642
rect 2044 42588 2100 42590
rect 1708 42364 1764 42420
rect 2492 42364 2548 42420
rect 2940 46396 2996 46452
rect 2716 43820 2772 43876
rect 3164 45778 3220 45780
rect 3164 45726 3166 45778
rect 3166 45726 3218 45778
rect 3218 45726 3220 45778
rect 3164 45724 3220 45726
rect 2604 41916 2660 41972
rect 3948 49868 4004 49924
rect 3724 43820 3780 43876
rect 3836 43372 3892 43428
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 5964 48300 6020 48356
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 5292 44492 5348 44548
rect 4284 43484 4340 43540
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 5740 43426 5796 43428
rect 5740 43374 5742 43426
rect 5742 43374 5794 43426
rect 5794 43374 5796 43426
rect 5740 43372 5796 43374
rect 4844 42588 4900 42644
rect 4284 41970 4340 41972
rect 4284 41918 4286 41970
rect 4286 41918 4338 41970
rect 4338 41918 4340 41970
rect 4284 41916 4340 41918
rect 4956 41916 5012 41972
rect 1708 41692 1764 41748
rect 2044 41356 2100 41412
rect 1820 41186 1876 41188
rect 1820 41134 1822 41186
rect 1822 41134 1874 41186
rect 1874 41134 1876 41186
rect 1820 41132 1876 41134
rect 2492 41132 2548 41188
rect 2716 41804 2772 41860
rect 2380 41074 2436 41076
rect 2380 41022 2382 41074
rect 2382 41022 2434 41074
rect 2434 41022 2436 41074
rect 2380 41020 2436 41022
rect 2940 41692 2996 41748
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 3164 41074 3220 41076
rect 3164 41022 3166 41074
rect 3166 41022 3218 41074
rect 3218 41022 3220 41074
rect 3164 41020 3220 41022
rect 1820 40348 1876 40404
rect 5852 42754 5908 42756
rect 5852 42702 5854 42754
rect 5854 42702 5906 42754
rect 5906 42702 5908 42754
rect 5852 42700 5908 42702
rect 5852 42194 5908 42196
rect 5852 42142 5854 42194
rect 5854 42142 5906 42194
rect 5906 42142 5908 42194
rect 5852 42140 5908 42142
rect 8428 46956 8484 47012
rect 6748 45164 6804 45220
rect 6300 41970 6356 41972
rect 6300 41918 6302 41970
rect 6302 41918 6354 41970
rect 6354 41918 6356 41970
rect 6300 41916 6356 41918
rect 1708 40236 1764 40292
rect 4620 40402 4676 40404
rect 4620 40350 4622 40402
rect 4622 40350 4674 40402
rect 4674 40350 4676 40402
rect 4620 40348 4676 40350
rect 2492 40236 2548 40292
rect 2044 40124 2100 40180
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 1932 39730 1988 39732
rect 1932 39678 1934 39730
rect 1934 39678 1986 39730
rect 1986 39678 1988 39730
rect 1932 39676 1988 39678
rect 4284 39618 4340 39620
rect 4284 39566 4286 39618
rect 4286 39566 4338 39618
rect 4338 39566 4340 39618
rect 4284 39564 4340 39566
rect 1708 39004 1764 39060
rect 2044 38946 2100 38948
rect 2044 38894 2046 38946
rect 2046 38894 2098 38946
rect 2098 38894 2100 38946
rect 2044 38892 2100 38894
rect 4620 38946 4676 38948
rect 4620 38894 4622 38946
rect 4622 38894 4674 38946
rect 4674 38894 4676 38946
rect 4620 38892 4676 38894
rect 4732 38834 4788 38836
rect 4732 38782 4734 38834
rect 4734 38782 4786 38834
rect 4786 38782 4788 38834
rect 4732 38780 4788 38782
rect 5292 39116 5348 39172
rect 1708 38332 1764 38388
rect 5180 38610 5236 38612
rect 5180 38558 5182 38610
rect 5182 38558 5234 38610
rect 5234 38558 5236 38610
rect 5180 38556 5236 38558
rect 2492 38332 2548 38388
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 5068 38444 5124 38500
rect 2044 37938 2100 37940
rect 2044 37886 2046 37938
rect 2046 37886 2098 37938
rect 2098 37886 2100 37938
rect 2044 37884 2100 37886
rect 1708 37660 1764 37716
rect 2492 37660 2548 37716
rect 2044 37490 2100 37492
rect 2044 37438 2046 37490
rect 2046 37438 2098 37490
rect 2098 37438 2100 37490
rect 2044 37436 2100 37438
rect 5068 37436 5124 37492
rect 1708 36988 1764 37044
rect 1708 36428 1764 36484
rect 2940 36988 2996 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 2492 36428 2548 36484
rect 2716 36540 2772 36596
rect 2380 36370 2436 36372
rect 2380 36318 2382 36370
rect 2382 36318 2434 36370
rect 2434 36318 2436 36370
rect 2380 36316 2436 36318
rect 3164 36370 3220 36372
rect 3164 36318 3166 36370
rect 3166 36318 3218 36370
rect 3218 36318 3220 36370
rect 3164 36316 3220 36318
rect 2044 36258 2100 36260
rect 2044 36206 2046 36258
rect 2046 36206 2098 36258
rect 2098 36206 2100 36258
rect 2044 36204 2100 36206
rect 5740 38780 5796 38836
rect 5964 38834 6020 38836
rect 5964 38782 5966 38834
rect 5966 38782 6018 38834
rect 6018 38782 6020 38834
rect 5964 38780 6020 38782
rect 5404 37884 5460 37940
rect 5292 36204 5348 36260
rect 5628 38444 5684 38500
rect 5852 38274 5908 38276
rect 5852 38222 5854 38274
rect 5854 38222 5906 38274
rect 5906 38222 5908 38274
rect 5852 38220 5908 38222
rect 6188 39116 6244 39172
rect 6188 38556 6244 38612
rect 6076 38220 6132 38276
rect 6188 38332 6244 38388
rect 6076 37884 6132 37940
rect 6412 37884 6468 37940
rect 6412 37548 6468 37604
rect 6524 37324 6580 37380
rect 14588 54460 14644 54516
rect 17052 54460 17108 54516
rect 15596 53788 15652 53844
rect 14588 53618 14644 53620
rect 14588 53566 14590 53618
rect 14590 53566 14642 53618
rect 14642 53566 14644 53618
rect 14588 53564 14644 53566
rect 15484 53564 15540 53620
rect 16828 53452 16884 53508
rect 17388 53842 17444 53844
rect 17388 53790 17390 53842
rect 17390 53790 17442 53842
rect 17442 53790 17444 53842
rect 17388 53788 17444 53790
rect 17612 54514 17668 54516
rect 17612 54462 17614 54514
rect 17614 54462 17666 54514
rect 17666 54462 17668 54514
rect 17612 54460 17668 54462
rect 17612 53730 17668 53732
rect 17612 53678 17614 53730
rect 17614 53678 17666 53730
rect 17666 53678 17668 53730
rect 17612 53676 17668 53678
rect 16940 52780 16996 52836
rect 12908 50428 12964 50484
rect 10108 49868 10164 49924
rect 12236 49868 12292 49924
rect 14588 51266 14644 51268
rect 14588 51214 14590 51266
rect 14590 51214 14642 51266
rect 14642 51214 14644 51266
rect 14588 51212 14644 51214
rect 14700 50764 14756 50820
rect 13692 50706 13748 50708
rect 13692 50654 13694 50706
rect 13694 50654 13746 50706
rect 13746 50654 13748 50706
rect 13692 50652 13748 50654
rect 13580 50482 13636 50484
rect 13580 50430 13582 50482
rect 13582 50430 13634 50482
rect 13634 50430 13636 50482
rect 13580 50428 13636 50430
rect 13468 49868 13524 49924
rect 14028 49868 14084 49924
rect 13356 49756 13412 49812
rect 12236 48860 12292 48916
rect 9660 46956 9716 47012
rect 11004 46786 11060 46788
rect 11004 46734 11006 46786
rect 11006 46734 11058 46786
rect 11058 46734 11060 46786
rect 11004 46732 11060 46734
rect 12012 48242 12068 48244
rect 12012 48190 12014 48242
rect 12014 48190 12066 48242
rect 12066 48190 12068 48242
rect 12012 48188 12068 48190
rect 13356 48860 13412 48916
rect 12908 48188 12964 48244
rect 12908 47740 12964 47796
rect 11788 46786 11844 46788
rect 11788 46734 11790 46786
rect 11790 46734 11842 46786
rect 11842 46734 11844 46786
rect 11788 46732 11844 46734
rect 9884 46562 9940 46564
rect 9884 46510 9886 46562
rect 9886 46510 9938 46562
rect 9938 46510 9940 46562
rect 9884 46508 9940 46510
rect 11228 46002 11284 46004
rect 11228 45950 11230 46002
rect 11230 45950 11282 46002
rect 11282 45950 11284 46002
rect 11228 45948 11284 45950
rect 11676 46674 11732 46676
rect 11676 46622 11678 46674
rect 11678 46622 11730 46674
rect 11730 46622 11732 46674
rect 11676 46620 11732 46622
rect 9772 44994 9828 44996
rect 9772 44942 9774 44994
rect 9774 44942 9826 44994
rect 9826 44942 9828 44994
rect 9772 44940 9828 44942
rect 10108 44604 10164 44660
rect 6860 43596 6916 43652
rect 8092 43484 8148 43540
rect 7868 42924 7924 42980
rect 7532 42642 7588 42644
rect 7532 42590 7534 42642
rect 7534 42590 7586 42642
rect 7586 42590 7588 42642
rect 7532 42588 7588 42590
rect 8652 43538 8708 43540
rect 8652 43486 8654 43538
rect 8654 43486 8706 43538
rect 8706 43486 8708 43538
rect 8652 43484 8708 43486
rect 8204 43372 8260 43428
rect 8764 42642 8820 42644
rect 8764 42590 8766 42642
rect 8766 42590 8818 42642
rect 8818 42590 8820 42642
rect 8764 42588 8820 42590
rect 7084 42140 7140 42196
rect 8092 41356 8148 41412
rect 8316 40460 8372 40516
rect 7644 40236 7700 40292
rect 7084 39564 7140 39620
rect 6860 38834 6916 38836
rect 6860 38782 6862 38834
rect 6862 38782 6914 38834
rect 6914 38782 6916 38834
rect 6860 38780 6916 38782
rect 6748 38722 6804 38724
rect 6748 38670 6750 38722
rect 6750 38670 6802 38722
rect 6802 38670 6804 38722
rect 6748 38668 6804 38670
rect 7644 37938 7700 37940
rect 7644 37886 7646 37938
rect 7646 37886 7698 37938
rect 7698 37886 7700 37938
rect 7644 37884 7700 37886
rect 7308 37548 7364 37604
rect 7532 37548 7588 37604
rect 6972 37378 7028 37380
rect 6972 37326 6974 37378
rect 6974 37326 7026 37378
rect 7026 37326 7028 37378
rect 6972 37324 7028 37326
rect 6636 36540 6692 36596
rect 7308 36540 7364 36596
rect 1708 35644 1764 35700
rect 4284 35698 4340 35700
rect 4284 35646 4286 35698
rect 4286 35646 4338 35698
rect 4338 35646 4340 35698
rect 4284 35644 4340 35646
rect 7532 35644 7588 35700
rect 7980 35756 8036 35812
rect 5180 35532 5236 35588
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 1932 34972 1988 35028
rect 1932 34076 1988 34132
rect 8764 40124 8820 40180
rect 9100 40908 9156 40964
rect 8540 40012 8596 40068
rect 8988 40012 9044 40068
rect 9548 40236 9604 40292
rect 9548 39564 9604 39620
rect 8764 37938 8820 37940
rect 8764 37886 8766 37938
rect 8766 37886 8818 37938
rect 8818 37886 8820 37938
rect 8764 37884 8820 37886
rect 8428 36594 8484 36596
rect 8428 36542 8430 36594
rect 8430 36542 8482 36594
rect 8482 36542 8484 36594
rect 8428 36540 8484 36542
rect 8316 35756 8372 35812
rect 8428 35586 8484 35588
rect 8428 35534 8430 35586
rect 8430 35534 8482 35586
rect 8482 35534 8484 35586
rect 8428 35532 8484 35534
rect 5068 34076 5124 34132
rect 4284 33852 4340 33908
rect 1708 32284 1764 32340
rect 3052 31836 3108 31892
rect 3388 31836 3444 31892
rect 2940 31666 2996 31668
rect 2940 31614 2942 31666
rect 2942 31614 2994 31666
rect 2994 31614 2996 31666
rect 2940 31612 2996 31614
rect 2044 31554 2100 31556
rect 2044 31502 2046 31554
rect 2046 31502 2098 31554
rect 2098 31502 2100 31554
rect 2044 31500 2100 31502
rect 1820 31164 1876 31220
rect 2044 31106 2100 31108
rect 2044 31054 2046 31106
rect 2046 31054 2098 31106
rect 2098 31054 2100 31106
rect 2044 31052 2100 31054
rect 2380 30994 2436 30996
rect 2380 30942 2382 30994
rect 2382 30942 2434 30994
rect 2434 30942 2436 30994
rect 2380 30940 2436 30942
rect 2716 30716 2772 30772
rect 1708 29426 1764 29428
rect 1708 29374 1710 29426
rect 1710 29374 1762 29426
rect 1762 29374 1764 29426
rect 1708 29372 1764 29374
rect 3164 31554 3220 31556
rect 3164 31502 3166 31554
rect 3166 31502 3218 31554
rect 3218 31502 3220 31554
rect 3164 31500 3220 31502
rect 4060 31836 4116 31892
rect 3724 31724 3780 31780
rect 3836 31666 3892 31668
rect 3836 31614 3838 31666
rect 3838 31614 3890 31666
rect 3890 31614 3892 31666
rect 3836 31612 3892 31614
rect 3052 30828 3108 30884
rect 3052 30268 3108 30324
rect 3164 30940 3220 30996
rect 2828 30156 2884 30212
rect 2492 30098 2548 30100
rect 2492 30046 2494 30098
rect 2494 30046 2546 30098
rect 2546 30046 2548 30098
rect 2492 30044 2548 30046
rect 2044 29650 2100 29652
rect 2044 29598 2046 29650
rect 2046 29598 2098 29650
rect 2098 29598 2100 29650
rect 2044 29596 2100 29598
rect 3388 30380 3444 30436
rect 3612 30044 3668 30100
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4732 33458 4788 33460
rect 4732 33406 4734 33458
rect 4734 33406 4786 33458
rect 4786 33406 4788 33458
rect 4732 33404 4788 33406
rect 4620 32620 4676 32676
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4620 31778 4676 31780
rect 4620 31726 4622 31778
rect 4622 31726 4674 31778
rect 4674 31726 4676 31778
rect 4620 31724 4676 31726
rect 5628 34076 5684 34132
rect 5180 31948 5236 32004
rect 5292 33404 5348 33460
rect 5404 32674 5460 32676
rect 5404 32622 5406 32674
rect 5406 32622 5458 32674
rect 5458 32622 5460 32674
rect 5404 32620 5460 32622
rect 5404 31948 5460 32004
rect 4508 31666 4564 31668
rect 4508 31614 4510 31666
rect 4510 31614 4562 31666
rect 4562 31614 4564 31666
rect 4508 31612 4564 31614
rect 4732 31500 4788 31556
rect 5068 31500 5124 31556
rect 5516 31612 5572 31668
rect 2716 29538 2772 29540
rect 2716 29486 2718 29538
rect 2718 29486 2770 29538
rect 2770 29486 2772 29538
rect 2716 29484 2772 29486
rect 2380 29260 2436 29316
rect 2380 28924 2436 28980
rect 3164 29372 3220 29428
rect 1708 28364 1764 28420
rect 1708 27356 1764 27412
rect 1708 26908 1764 26964
rect 2492 28530 2548 28532
rect 2492 28478 2494 28530
rect 2494 28478 2546 28530
rect 2546 28478 2548 28530
rect 2492 28476 2548 28478
rect 2716 28082 2772 28084
rect 2716 28030 2718 28082
rect 2718 28030 2770 28082
rect 2770 28030 2772 28082
rect 2716 28028 2772 28030
rect 3500 28252 3556 28308
rect 3612 28476 3668 28532
rect 3276 27916 3332 27972
rect 2044 27692 2100 27748
rect 2604 27580 2660 27636
rect 2044 27244 2100 27300
rect 2492 26908 2548 26964
rect 1596 25788 1652 25844
rect 1708 25564 1764 25620
rect 1820 25228 1876 25284
rect 1708 24892 1764 24948
rect 1708 23996 1764 24052
rect 2044 26460 2100 26516
rect 2492 26348 2548 26404
rect 2492 26178 2548 26180
rect 2492 26126 2494 26178
rect 2494 26126 2546 26178
rect 2546 26126 2548 26178
rect 2492 26124 2548 26126
rect 2268 25676 2324 25732
rect 2716 27132 2772 27188
rect 3724 27916 3780 27972
rect 3388 27356 3444 27412
rect 2604 25564 2660 25620
rect 3724 27132 3780 27188
rect 3500 26572 3556 26628
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4508 30044 4564 30100
rect 5852 33852 5908 33908
rect 7196 33852 7252 33908
rect 5740 33404 5796 33460
rect 7084 33404 7140 33460
rect 5852 33122 5908 33124
rect 5852 33070 5854 33122
rect 5854 33070 5906 33122
rect 5906 33070 5908 33122
rect 5852 33068 5908 33070
rect 5740 30210 5796 30212
rect 5740 30158 5742 30210
rect 5742 30158 5794 30210
rect 5794 30158 5796 30210
rect 5740 30156 5796 30158
rect 4508 29148 4564 29204
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 3948 28476 4004 28532
rect 4620 28252 4676 28308
rect 4172 27858 4228 27860
rect 4172 27806 4174 27858
rect 4174 27806 4226 27858
rect 4226 27806 4228 27858
rect 4172 27804 4228 27806
rect 5068 29314 5124 29316
rect 5068 29262 5070 29314
rect 5070 29262 5122 29314
rect 5122 29262 5124 29314
rect 5068 29260 5124 29262
rect 4844 28476 4900 28532
rect 5068 28418 5124 28420
rect 5068 28366 5070 28418
rect 5070 28366 5122 28418
rect 5122 28366 5124 28418
rect 5068 28364 5124 28366
rect 5068 27970 5124 27972
rect 5068 27918 5070 27970
rect 5070 27918 5122 27970
rect 5122 27918 5124 27970
rect 5068 27916 5124 27918
rect 4844 27692 4900 27748
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4508 27132 4564 27188
rect 4060 26850 4116 26852
rect 4060 26798 4062 26850
rect 4062 26798 4114 26850
rect 4114 26798 4116 26850
rect 4060 26796 4116 26798
rect 2716 25394 2772 25396
rect 2716 25342 2718 25394
rect 2718 25342 2770 25394
rect 2770 25342 2772 25394
rect 2716 25340 2772 25342
rect 3164 25340 3220 25396
rect 3948 26572 4004 26628
rect 3500 25116 3556 25172
rect 2716 24946 2772 24948
rect 2716 24894 2718 24946
rect 2718 24894 2770 24946
rect 2770 24894 2772 24946
rect 2716 24892 2772 24894
rect 2380 24722 2436 24724
rect 2380 24670 2382 24722
rect 2382 24670 2434 24722
rect 2434 24670 2436 24722
rect 2380 24668 2436 24670
rect 2380 24220 2436 24276
rect 1708 22876 1764 22932
rect 1708 22428 1764 22484
rect 2940 23154 2996 23156
rect 2940 23102 2942 23154
rect 2942 23102 2994 23154
rect 2994 23102 2996 23154
rect 2940 23100 2996 23102
rect 1708 22204 1764 22260
rect 1708 21810 1764 21812
rect 1708 21758 1710 21810
rect 1710 21758 1762 21810
rect 1762 21758 1764 21810
rect 1708 21756 1764 21758
rect 1708 20860 1764 20916
rect 1708 20188 1764 20244
rect 2268 21474 2324 21476
rect 2268 21422 2270 21474
rect 2270 21422 2322 21474
rect 2322 21422 2324 21474
rect 2268 21420 2324 21422
rect 2492 21756 2548 21812
rect 2940 21980 2996 22036
rect 2604 21586 2660 21588
rect 2604 21534 2606 21586
rect 2606 21534 2658 21586
rect 2658 21534 2660 21586
rect 2604 21532 2660 21534
rect 3836 26124 3892 26180
rect 3724 26012 3780 26068
rect 4060 26236 4116 26292
rect 4060 25676 4116 25732
rect 4508 26348 4564 26404
rect 5068 27074 5124 27076
rect 5068 27022 5070 27074
rect 5070 27022 5122 27074
rect 5122 27022 5124 27074
rect 5068 27020 5124 27022
rect 4732 26796 4788 26852
rect 4620 26178 4676 26180
rect 4620 26126 4622 26178
rect 4622 26126 4674 26178
rect 4674 26126 4676 26178
rect 4620 26124 4676 26126
rect 4844 26348 4900 26404
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 5740 29148 5796 29204
rect 5628 28476 5684 28532
rect 5292 27858 5348 27860
rect 5292 27806 5294 27858
rect 5294 27806 5346 27858
rect 5346 27806 5348 27858
rect 5292 27804 5348 27806
rect 5404 27692 5460 27748
rect 5740 26962 5796 26964
rect 5740 26910 5742 26962
rect 5742 26910 5794 26962
rect 5794 26910 5796 26962
rect 5740 26908 5796 26910
rect 6300 33122 6356 33124
rect 6300 33070 6302 33122
rect 6302 33070 6354 33122
rect 6354 33070 6356 33122
rect 6300 33068 6356 33070
rect 6972 32620 7028 32676
rect 8652 33852 8708 33908
rect 8540 33404 8596 33460
rect 7532 32620 7588 32676
rect 6300 32396 6356 32452
rect 7644 32450 7700 32452
rect 7644 32398 7646 32450
rect 7646 32398 7698 32450
rect 7698 32398 7700 32450
rect 7644 32396 7700 32398
rect 8540 32562 8596 32564
rect 8540 32510 8542 32562
rect 8542 32510 8594 32562
rect 8594 32510 8596 32562
rect 8540 32508 8596 32510
rect 8316 32396 8372 32452
rect 6188 31948 6244 32004
rect 7644 31948 7700 32004
rect 6524 31778 6580 31780
rect 6524 31726 6526 31778
rect 6526 31726 6578 31778
rect 6578 31726 6580 31778
rect 6524 31724 6580 31726
rect 5964 31666 6020 31668
rect 5964 31614 5966 31666
rect 5966 31614 6018 31666
rect 6018 31614 6020 31666
rect 5964 31612 6020 31614
rect 7532 31388 7588 31444
rect 8540 31276 8596 31332
rect 5964 31218 6020 31220
rect 5964 31166 5966 31218
rect 5966 31166 6018 31218
rect 6018 31166 6020 31218
rect 5964 31164 6020 31166
rect 8428 31052 8484 31108
rect 6412 30882 6468 30884
rect 6412 30830 6414 30882
rect 6414 30830 6466 30882
rect 6466 30830 6468 30882
rect 6412 30828 6468 30830
rect 7980 30380 8036 30436
rect 5964 30098 6020 30100
rect 5964 30046 5966 30098
rect 5966 30046 6018 30098
rect 6018 30046 6020 30098
rect 5964 30044 6020 30046
rect 8204 30156 8260 30212
rect 8652 30044 8708 30100
rect 7980 29932 8036 29988
rect 6972 29596 7028 29652
rect 7868 29372 7924 29428
rect 7756 28700 7812 28756
rect 6972 28588 7028 28644
rect 5964 27916 6020 27972
rect 6188 27020 6244 27076
rect 7420 28588 7476 28644
rect 7420 27580 7476 27636
rect 8540 29596 8596 29652
rect 8988 31612 9044 31668
rect 9100 31388 9156 31444
rect 9100 31052 9156 31108
rect 8876 30434 8932 30436
rect 8876 30382 8878 30434
rect 8878 30382 8930 30434
rect 8930 30382 8932 30434
rect 8876 30380 8932 30382
rect 8876 29650 8932 29652
rect 8876 29598 8878 29650
rect 8878 29598 8930 29650
rect 8930 29598 8932 29650
rect 8876 29596 8932 29598
rect 8092 29426 8148 29428
rect 8092 29374 8094 29426
rect 8094 29374 8146 29426
rect 8146 29374 8148 29426
rect 8092 29372 8148 29374
rect 8988 29426 9044 29428
rect 8988 29374 8990 29426
rect 8990 29374 9042 29426
rect 9042 29374 9044 29426
rect 8988 29372 9044 29374
rect 8092 28754 8148 28756
rect 8092 28702 8094 28754
rect 8094 28702 8146 28754
rect 8146 28702 8148 28754
rect 8092 28700 8148 28702
rect 8204 28642 8260 28644
rect 8204 28590 8206 28642
rect 8206 28590 8258 28642
rect 8258 28590 8260 28642
rect 8204 28588 8260 28590
rect 8652 28364 8708 28420
rect 7980 27634 8036 27636
rect 7980 27582 7982 27634
rect 7982 27582 8034 27634
rect 8034 27582 8036 27634
rect 7980 27580 8036 27582
rect 8876 27804 8932 27860
rect 8540 27580 8596 27636
rect 4060 25340 4116 25396
rect 3612 24892 3668 24948
rect 3948 25116 4004 25172
rect 4172 24892 4228 24948
rect 5404 26178 5460 26180
rect 5404 26126 5406 26178
rect 5406 26126 5458 26178
rect 5458 26126 5460 26178
rect 5404 26124 5460 26126
rect 5964 26348 6020 26404
rect 5852 25676 5908 25732
rect 4844 25282 4900 25284
rect 4844 25230 4846 25282
rect 4846 25230 4898 25282
rect 4898 25230 4900 25282
rect 4844 25228 4900 25230
rect 5516 25116 5572 25172
rect 4732 24834 4788 24836
rect 4732 24782 4734 24834
rect 4734 24782 4786 24834
rect 4786 24782 4788 24834
rect 4732 24780 4788 24782
rect 3724 23772 3780 23828
rect 3612 22988 3668 23044
rect 3948 23660 4004 23716
rect 3276 21308 3332 21364
rect 2380 20972 2436 21028
rect 2268 20914 2324 20916
rect 2268 20862 2270 20914
rect 2270 20862 2322 20914
rect 2322 20862 2324 20914
rect 2268 20860 2324 20862
rect 2492 20524 2548 20580
rect 2940 20748 2996 20804
rect 3836 21810 3892 21812
rect 3836 21758 3838 21810
rect 3838 21758 3890 21810
rect 3890 21758 3892 21810
rect 3836 21756 3892 21758
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 3724 21196 3780 21252
rect 2716 20300 2772 20356
rect 2604 20188 2660 20244
rect 1708 19516 1764 19572
rect 1708 18172 1764 18228
rect 1708 17724 1764 17780
rect 2044 19010 2100 19012
rect 2044 18958 2046 19010
rect 2046 18958 2098 19010
rect 2098 18958 2100 19010
rect 2044 18956 2100 18958
rect 2380 18844 2436 18900
rect 3500 20578 3556 20580
rect 3500 20526 3502 20578
rect 3502 20526 3554 20578
rect 3554 20526 3556 20578
rect 3500 20524 3556 20526
rect 4844 23660 4900 23716
rect 4620 22988 4676 23044
rect 4844 23324 4900 23380
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 5068 24050 5124 24052
rect 5068 23998 5070 24050
rect 5070 23998 5122 24050
rect 5122 23998 5124 24050
rect 5068 23996 5124 23998
rect 5404 24610 5460 24612
rect 5404 24558 5406 24610
rect 5406 24558 5458 24610
rect 5458 24558 5460 24610
rect 5404 24556 5460 24558
rect 6188 26012 6244 26068
rect 6188 25730 6244 25732
rect 6188 25678 6190 25730
rect 6190 25678 6242 25730
rect 6242 25678 6244 25730
rect 6188 25676 6244 25678
rect 5964 25228 6020 25284
rect 5852 25116 5908 25172
rect 5740 24444 5796 24500
rect 5292 23772 5348 23828
rect 7980 26962 8036 26964
rect 7980 26910 7982 26962
rect 7982 26910 8034 26962
rect 8034 26910 8036 26962
rect 7980 26908 8036 26910
rect 7308 26178 7364 26180
rect 7308 26126 7310 26178
rect 7310 26126 7362 26178
rect 7362 26126 7364 26178
rect 7308 26124 7364 26126
rect 7980 25618 8036 25620
rect 7980 25566 7982 25618
rect 7982 25566 8034 25618
rect 8034 25566 8036 25618
rect 7980 25564 8036 25566
rect 6412 25116 6468 25172
rect 6188 24834 6244 24836
rect 6188 24782 6190 24834
rect 6190 24782 6242 24834
rect 6242 24782 6244 24834
rect 6188 24780 6244 24782
rect 6300 24498 6356 24500
rect 6300 24446 6302 24498
rect 6302 24446 6354 24498
rect 6354 24446 6356 24498
rect 6300 24444 6356 24446
rect 5740 23772 5796 23828
rect 5740 23548 5796 23604
rect 5292 22988 5348 23044
rect 5964 23714 6020 23716
rect 5964 23662 5966 23714
rect 5966 23662 6018 23714
rect 6018 23662 6020 23714
rect 5964 23660 6020 23662
rect 6636 23996 6692 24052
rect 6300 23548 6356 23604
rect 6636 23772 6692 23828
rect 6300 23154 6356 23156
rect 6300 23102 6302 23154
rect 6302 23102 6354 23154
rect 6354 23102 6356 23154
rect 6300 23100 6356 23102
rect 4172 21196 4228 21252
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 5740 21698 5796 21700
rect 5740 21646 5742 21698
rect 5742 21646 5794 21698
rect 5794 21646 5796 21698
rect 5740 21644 5796 21646
rect 5292 21586 5348 21588
rect 5292 21534 5294 21586
rect 5294 21534 5346 21586
rect 5346 21534 5348 21586
rect 5292 21532 5348 21534
rect 4172 20802 4228 20804
rect 4172 20750 4174 20802
rect 4174 20750 4226 20802
rect 4226 20750 4228 20802
rect 4172 20748 4228 20750
rect 4844 20802 4900 20804
rect 4844 20750 4846 20802
rect 4846 20750 4898 20802
rect 4898 20750 4900 20802
rect 4844 20748 4900 20750
rect 2716 19122 2772 19124
rect 2716 19070 2718 19122
rect 2718 19070 2770 19122
rect 2770 19070 2772 19122
rect 2716 19068 2772 19070
rect 2044 17836 2100 17892
rect 3388 19404 3444 19460
rect 6188 22482 6244 22484
rect 6188 22430 6190 22482
rect 6190 22430 6242 22482
rect 6242 22430 6244 22482
rect 6188 22428 6244 22430
rect 6300 21362 6356 21364
rect 6300 21310 6302 21362
rect 6302 21310 6354 21362
rect 6354 21310 6356 21362
rect 6300 21308 6356 21310
rect 5964 20748 6020 20804
rect 4172 19740 4228 19796
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4844 19628 4900 19684
rect 3164 18844 3220 18900
rect 3836 19234 3892 19236
rect 3836 19182 3838 19234
rect 3838 19182 3890 19234
rect 3890 19182 3892 19234
rect 3836 19180 3892 19182
rect 2940 17612 2996 17668
rect 1596 17276 1652 17332
rect 1708 17500 1764 17556
rect 1708 16156 1764 16212
rect 1708 15596 1764 15652
rect 1708 15036 1764 15092
rect 2380 16882 2436 16884
rect 2380 16830 2382 16882
rect 2382 16830 2434 16882
rect 2434 16830 2436 16882
rect 2380 16828 2436 16830
rect 3164 17106 3220 17108
rect 3164 17054 3166 17106
rect 3166 17054 3218 17106
rect 3218 17054 3220 17106
rect 3164 17052 3220 17054
rect 2492 16716 2548 16772
rect 2044 16604 2100 16660
rect 3276 16716 3332 16772
rect 2716 16268 2772 16324
rect 2380 15484 2436 15540
rect 2044 15426 2100 15428
rect 2044 15374 2046 15426
rect 2046 15374 2098 15426
rect 2098 15374 2100 15426
rect 2044 15372 2100 15374
rect 2716 15538 2772 15540
rect 2716 15486 2718 15538
rect 2718 15486 2770 15538
rect 2770 15486 2772 15538
rect 2716 15484 2772 15486
rect 3052 15314 3108 15316
rect 3052 15262 3054 15314
rect 3054 15262 3106 15314
rect 3106 15262 3108 15314
rect 3052 15260 3108 15262
rect 2044 14700 2100 14756
rect 2716 14588 2772 14644
rect 2492 14530 2548 14532
rect 2492 14478 2494 14530
rect 2494 14478 2546 14530
rect 2546 14478 2548 14530
rect 2492 14476 2548 14478
rect 1708 13356 1764 13412
rect 1708 12572 1764 12628
rect 1708 12178 1764 12180
rect 1708 12126 1710 12178
rect 1710 12126 1762 12178
rect 1762 12126 1764 12178
rect 1708 12124 1764 12126
rect 1708 11452 1764 11508
rect 1708 10722 1764 10724
rect 1708 10670 1710 10722
rect 1710 10670 1762 10722
rect 1762 10670 1764 10722
rect 1708 10668 1764 10670
rect 2716 13692 2772 13748
rect 2492 13020 2548 13076
rect 2380 12962 2436 12964
rect 2380 12910 2382 12962
rect 2382 12910 2434 12962
rect 2434 12910 2436 12962
rect 2380 12908 2436 12910
rect 3276 13468 3332 13524
rect 3612 18396 3668 18452
rect 3724 15708 3780 15764
rect 3612 15372 3668 15428
rect 3948 18396 4004 18452
rect 4060 17052 4116 17108
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 4620 18508 4676 18564
rect 5628 19906 5684 19908
rect 5628 19854 5630 19906
rect 5630 19854 5682 19906
rect 5682 19854 5684 19906
rect 5628 19852 5684 19854
rect 4844 18508 4900 18564
rect 4508 18396 4564 18452
rect 4396 18284 4452 18340
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 6300 20300 6356 20356
rect 6636 23042 6692 23044
rect 6636 22990 6638 23042
rect 6638 22990 6690 23042
rect 6690 22990 6692 23042
rect 6636 22988 6692 22990
rect 6636 22204 6692 22260
rect 7756 25452 7812 25508
rect 7308 24722 7364 24724
rect 7308 24670 7310 24722
rect 7310 24670 7362 24722
rect 7362 24670 7364 24722
rect 7308 24668 7364 24670
rect 7084 24556 7140 24612
rect 6972 23660 7028 23716
rect 8988 27634 9044 27636
rect 8988 27582 8990 27634
rect 8990 27582 9042 27634
rect 9042 27582 9044 27634
rect 8988 27580 9044 27582
rect 8988 26908 9044 26964
rect 8428 26290 8484 26292
rect 8428 26238 8430 26290
rect 8430 26238 8482 26290
rect 8482 26238 8484 26290
rect 8428 26236 8484 26238
rect 9548 35532 9604 35588
rect 9548 31948 9604 32004
rect 9436 31724 9492 31780
rect 9996 42812 10052 42868
rect 9996 39618 10052 39620
rect 9996 39566 9998 39618
rect 9998 39566 10050 39618
rect 10050 39566 10052 39618
rect 9996 39564 10052 39566
rect 9996 39004 10052 39060
rect 10780 45500 10836 45556
rect 11788 46508 11844 46564
rect 13468 48748 13524 48804
rect 13132 47740 13188 47796
rect 12460 46620 12516 46676
rect 13132 46060 13188 46116
rect 13244 46956 13300 47012
rect 11788 45778 11844 45780
rect 11788 45726 11790 45778
rect 11790 45726 11842 45778
rect 11842 45726 11844 45778
rect 11788 45724 11844 45726
rect 11676 45500 11732 45556
rect 12236 45612 12292 45668
rect 11228 45218 11284 45220
rect 11228 45166 11230 45218
rect 11230 45166 11282 45218
rect 11282 45166 11284 45218
rect 11228 45164 11284 45166
rect 10892 44994 10948 44996
rect 10892 44942 10894 44994
rect 10894 44942 10946 44994
rect 10946 44942 10948 44994
rect 10892 44940 10948 44942
rect 11452 44098 11508 44100
rect 11452 44046 11454 44098
rect 11454 44046 11506 44098
rect 11506 44046 11508 44098
rect 11452 44044 11508 44046
rect 12572 45724 12628 45780
rect 12236 45388 12292 45444
rect 12124 45276 12180 45332
rect 12012 44044 12068 44100
rect 12012 43596 12068 43652
rect 10556 43538 10612 43540
rect 10556 43486 10558 43538
rect 10558 43486 10610 43538
rect 10610 43486 10612 43538
rect 10556 43484 10612 43486
rect 11340 43426 11396 43428
rect 11340 43374 11342 43426
rect 11342 43374 11394 43426
rect 11394 43374 11396 43426
rect 11340 43372 11396 43374
rect 11228 42978 11284 42980
rect 11228 42926 11230 42978
rect 11230 42926 11282 42978
rect 11282 42926 11284 42978
rect 11228 42924 11284 42926
rect 12236 43484 12292 43540
rect 13244 45388 13300 45444
rect 13020 44322 13076 44324
rect 13020 44270 13022 44322
rect 13022 44270 13074 44322
rect 13074 44270 13076 44322
rect 13020 44268 13076 44270
rect 12460 43148 12516 43204
rect 10444 42866 10500 42868
rect 10444 42814 10446 42866
rect 10446 42814 10498 42866
rect 10498 42814 10500 42866
rect 10444 42812 10500 42814
rect 11004 42812 11060 42868
rect 10892 41186 10948 41188
rect 10892 41134 10894 41186
rect 10894 41134 10946 41186
rect 10946 41134 10948 41186
rect 10892 41132 10948 41134
rect 10668 40460 10724 40516
rect 10892 39730 10948 39732
rect 10892 39678 10894 39730
rect 10894 39678 10946 39730
rect 10946 39678 10948 39730
rect 10892 39676 10948 39678
rect 10220 39058 10276 39060
rect 10220 39006 10222 39058
rect 10222 39006 10274 39058
rect 10274 39006 10276 39058
rect 10220 39004 10276 39006
rect 10892 37996 10948 38052
rect 11340 42700 11396 42756
rect 12796 42924 12852 42980
rect 13132 44044 13188 44100
rect 12012 42700 12068 42756
rect 11564 42642 11620 42644
rect 11564 42590 11566 42642
rect 11566 42590 11618 42642
rect 11618 42590 11620 42642
rect 11564 42588 11620 42590
rect 11116 41804 11172 41860
rect 12572 42588 12628 42644
rect 11452 40460 11508 40516
rect 11116 39676 11172 39732
rect 11564 39730 11620 39732
rect 11564 39678 11566 39730
rect 11566 39678 11618 39730
rect 11618 39678 11620 39730
rect 11564 39676 11620 39678
rect 12572 42082 12628 42084
rect 12572 42030 12574 42082
rect 12574 42030 12626 42082
rect 12626 42030 12628 42082
rect 12572 42028 12628 42030
rect 12348 41970 12404 41972
rect 12348 41918 12350 41970
rect 12350 41918 12402 41970
rect 12402 41918 12404 41970
rect 12348 41916 12404 41918
rect 12796 41804 12852 41860
rect 12908 40572 12964 40628
rect 11900 39618 11956 39620
rect 11900 39566 11902 39618
rect 11902 39566 11954 39618
rect 11954 39566 11956 39618
rect 11900 39564 11956 39566
rect 12908 39618 12964 39620
rect 12908 39566 12910 39618
rect 12910 39566 12962 39618
rect 12962 39566 12964 39618
rect 12908 39564 12964 39566
rect 11116 39058 11172 39060
rect 11116 39006 11118 39058
rect 11118 39006 11170 39058
rect 11170 39006 11172 39058
rect 11116 39004 11172 39006
rect 12460 39004 12516 39060
rect 11564 37996 11620 38052
rect 11340 37938 11396 37940
rect 11340 37886 11342 37938
rect 11342 37886 11394 37938
rect 11394 37886 11396 37938
rect 11340 37884 11396 37886
rect 12012 38050 12068 38052
rect 12012 37998 12014 38050
rect 12014 37998 12066 38050
rect 12066 37998 12068 38050
rect 12012 37996 12068 37998
rect 12236 37884 12292 37940
rect 11452 37436 11508 37492
rect 12572 38332 12628 38388
rect 11788 36482 11844 36484
rect 11788 36430 11790 36482
rect 11790 36430 11842 36482
rect 11842 36430 11844 36482
rect 11788 36428 11844 36430
rect 11004 35532 11060 35588
rect 11004 35308 11060 35364
rect 11004 34300 11060 34356
rect 10220 33964 10276 34020
rect 10556 33852 10612 33908
rect 11004 34018 11060 34020
rect 11004 33966 11006 34018
rect 11006 33966 11058 34018
rect 11058 33966 11060 34018
rect 11004 33964 11060 33966
rect 10444 33458 10500 33460
rect 10444 33406 10446 33458
rect 10446 33406 10498 33458
rect 10498 33406 10500 33458
rect 10444 33404 10500 33406
rect 9772 32674 9828 32676
rect 9772 32622 9774 32674
rect 9774 32622 9826 32674
rect 9826 32622 9828 32674
rect 9772 32620 9828 32622
rect 9996 32562 10052 32564
rect 9996 32510 9998 32562
rect 9998 32510 10050 32562
rect 10050 32510 10052 32562
rect 9996 32508 10052 32510
rect 10220 31836 10276 31892
rect 9660 31724 9716 31780
rect 9548 31388 9604 31444
rect 10108 31666 10164 31668
rect 10108 31614 10110 31666
rect 10110 31614 10162 31666
rect 10162 31614 10164 31666
rect 10108 31612 10164 31614
rect 10332 31666 10388 31668
rect 10332 31614 10334 31666
rect 10334 31614 10386 31666
rect 10386 31614 10388 31666
rect 10332 31612 10388 31614
rect 10220 31554 10276 31556
rect 10220 31502 10222 31554
rect 10222 31502 10274 31554
rect 10274 31502 10276 31554
rect 10220 31500 10276 31502
rect 12012 35756 12068 35812
rect 11564 33852 11620 33908
rect 11452 33404 11508 33460
rect 10668 31612 10724 31668
rect 9324 30716 9380 30772
rect 9548 30268 9604 30324
rect 9660 30044 9716 30100
rect 9772 29986 9828 29988
rect 9772 29934 9774 29986
rect 9774 29934 9826 29986
rect 9826 29934 9828 29986
rect 9772 29932 9828 29934
rect 9996 30716 10052 30772
rect 10220 30322 10276 30324
rect 10220 30270 10222 30322
rect 10222 30270 10274 30322
rect 10274 30270 10276 30322
rect 10220 30268 10276 30270
rect 10108 29650 10164 29652
rect 10108 29598 10110 29650
rect 10110 29598 10162 29650
rect 10162 29598 10164 29650
rect 10108 29596 10164 29598
rect 9772 27858 9828 27860
rect 9772 27806 9774 27858
rect 9774 27806 9826 27858
rect 9826 27806 9828 27858
rect 9772 27804 9828 27806
rect 9548 27580 9604 27636
rect 9212 25452 9268 25508
rect 9212 23548 9268 23604
rect 9548 26178 9604 26180
rect 9548 26126 9550 26178
rect 9550 26126 9602 26178
rect 9602 26126 9604 26178
rect 9548 26124 9604 26126
rect 9996 28364 10052 28420
rect 10220 27356 10276 27412
rect 10556 30210 10612 30212
rect 10556 30158 10558 30210
rect 10558 30158 10610 30210
rect 10610 30158 10612 30210
rect 10556 30156 10612 30158
rect 10444 30098 10500 30100
rect 10444 30046 10446 30098
rect 10446 30046 10498 30098
rect 10498 30046 10500 30098
rect 10444 30044 10500 30046
rect 10780 30940 10836 30996
rect 10780 29596 10836 29652
rect 10444 27804 10500 27860
rect 11340 31666 11396 31668
rect 11340 31614 11342 31666
rect 11342 31614 11394 31666
rect 11394 31614 11396 31666
rect 11340 31612 11396 31614
rect 11116 31554 11172 31556
rect 11116 31502 11118 31554
rect 11118 31502 11170 31554
rect 11170 31502 11172 31554
rect 11116 31500 11172 31502
rect 11676 33122 11732 33124
rect 11676 33070 11678 33122
rect 11678 33070 11730 33122
rect 11730 33070 11732 33122
rect 11676 33068 11732 33070
rect 11564 31836 11620 31892
rect 13020 37996 13076 38052
rect 12684 37324 12740 37380
rect 12572 37154 12628 37156
rect 12572 37102 12574 37154
rect 12574 37102 12626 37154
rect 12626 37102 12628 37154
rect 12572 37100 12628 37102
rect 13580 46114 13636 46116
rect 13580 46062 13582 46114
rect 13582 46062 13634 46114
rect 13634 46062 13636 46114
rect 13580 46060 13636 46062
rect 13692 45500 13748 45556
rect 13580 44210 13636 44212
rect 13580 44158 13582 44210
rect 13582 44158 13634 44210
rect 13634 44158 13636 44210
rect 13580 44156 13636 44158
rect 13468 43148 13524 43204
rect 13580 43372 13636 43428
rect 13468 42978 13524 42980
rect 13468 42926 13470 42978
rect 13470 42926 13522 42978
rect 13522 42926 13524 42978
rect 13468 42924 13524 42926
rect 13692 42700 13748 42756
rect 13692 42530 13748 42532
rect 13692 42478 13694 42530
rect 13694 42478 13746 42530
rect 13746 42478 13748 42530
rect 13692 42476 13748 42478
rect 13244 41020 13300 41076
rect 15820 50706 15876 50708
rect 15820 50654 15822 50706
rect 15822 50654 15874 50706
rect 15874 50654 15876 50706
rect 15820 50652 15876 50654
rect 16268 51996 16324 52052
rect 16492 51996 16548 52052
rect 16156 51266 16212 51268
rect 16156 51214 16158 51266
rect 16158 51214 16210 51266
rect 16210 51214 16212 51266
rect 16156 51212 16212 51214
rect 15708 50594 15764 50596
rect 15708 50542 15710 50594
rect 15710 50542 15762 50594
rect 15762 50542 15764 50594
rect 15708 50540 15764 50542
rect 15036 49532 15092 49588
rect 14700 48130 14756 48132
rect 14700 48078 14702 48130
rect 14702 48078 14754 48130
rect 14754 48078 14756 48130
rect 14700 48076 14756 48078
rect 14028 46956 14084 47012
rect 13916 45724 13972 45780
rect 14252 45500 14308 45556
rect 14140 45276 14196 45332
rect 13916 44716 13972 44772
rect 13916 44322 13972 44324
rect 13916 44270 13918 44322
rect 13918 44270 13970 44322
rect 13970 44270 13972 44322
rect 13916 44268 13972 44270
rect 14700 46002 14756 46004
rect 14700 45950 14702 46002
rect 14702 45950 14754 46002
rect 14754 45950 14756 46002
rect 14700 45948 14756 45950
rect 14476 45612 14532 45668
rect 14700 45106 14756 45108
rect 14700 45054 14702 45106
rect 14702 45054 14754 45106
rect 14754 45054 14756 45106
rect 14700 45052 14756 45054
rect 15148 49026 15204 49028
rect 15148 48974 15150 49026
rect 15150 48974 15202 49026
rect 15202 48974 15204 49026
rect 15148 48972 15204 48974
rect 15036 48860 15092 48916
rect 14140 44156 14196 44212
rect 13916 43538 13972 43540
rect 13916 43486 13918 43538
rect 13918 43486 13970 43538
rect 13970 43486 13972 43538
rect 13916 43484 13972 43486
rect 14028 42924 14084 42980
rect 13580 42028 13636 42084
rect 13468 41970 13524 41972
rect 13468 41918 13470 41970
rect 13470 41918 13522 41970
rect 13522 41918 13524 41970
rect 13468 41916 13524 41918
rect 13692 41020 13748 41076
rect 13804 41916 13860 41972
rect 14924 44604 14980 44660
rect 15708 49756 15764 49812
rect 17388 53564 17444 53620
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 17948 54460 18004 54516
rect 17836 53564 17892 53620
rect 18956 54514 19012 54516
rect 18956 54462 18958 54514
rect 18958 54462 19010 54514
rect 19010 54462 19012 54514
rect 18956 54460 19012 54462
rect 18396 54402 18452 54404
rect 18396 54350 18398 54402
rect 18398 54350 18450 54402
rect 18450 54350 18452 54402
rect 18396 54348 18452 54350
rect 18956 53788 19012 53844
rect 18396 53676 18452 53732
rect 18172 53564 18228 53620
rect 17388 52108 17444 52164
rect 17500 53506 17556 53508
rect 17500 53454 17502 53506
rect 17502 53454 17554 53506
rect 17554 53454 17556 53506
rect 17500 53452 17556 53454
rect 17724 53058 17780 53060
rect 17724 53006 17726 53058
rect 17726 53006 17778 53058
rect 17778 53006 17780 53058
rect 17724 53004 17780 53006
rect 18172 53058 18228 53060
rect 18172 53006 18174 53058
rect 18174 53006 18226 53058
rect 18226 53006 18228 53058
rect 18172 53004 18228 53006
rect 18172 52780 18228 52836
rect 17724 52332 17780 52388
rect 18060 52332 18116 52388
rect 17836 52162 17892 52164
rect 17836 52110 17838 52162
rect 17838 52110 17890 52162
rect 17890 52110 17892 52162
rect 17836 52108 17892 52110
rect 17052 51660 17108 51716
rect 17948 51660 18004 51716
rect 17052 50764 17108 50820
rect 16380 50540 16436 50596
rect 15932 49756 15988 49812
rect 16492 49980 16548 50036
rect 15820 49532 15876 49588
rect 15820 49026 15876 49028
rect 15820 48974 15822 49026
rect 15822 48974 15874 49026
rect 15874 48974 15876 49026
rect 15820 48972 15876 48974
rect 16156 48860 16212 48916
rect 17612 51548 17668 51604
rect 15148 48748 15204 48804
rect 15260 46844 15316 46900
rect 15148 46002 15204 46004
rect 15148 45950 15150 46002
rect 15150 45950 15202 46002
rect 15202 45950 15204 46002
rect 15148 45948 15204 45950
rect 16044 46844 16100 46900
rect 15708 45890 15764 45892
rect 15708 45838 15710 45890
rect 15710 45838 15762 45890
rect 15762 45838 15764 45890
rect 15708 45836 15764 45838
rect 15372 45164 15428 45220
rect 15260 45106 15316 45108
rect 15260 45054 15262 45106
rect 15262 45054 15314 45106
rect 15314 45054 15316 45106
rect 15260 45052 15316 45054
rect 15148 44492 15204 44548
rect 14476 43596 14532 43652
rect 14364 42978 14420 42980
rect 14364 42926 14366 42978
rect 14366 42926 14418 42978
rect 14418 42926 14420 42978
rect 14364 42924 14420 42926
rect 14028 41244 14084 41300
rect 14252 41132 14308 41188
rect 13804 40908 13860 40964
rect 14028 40460 14084 40516
rect 13468 40290 13524 40292
rect 13468 40238 13470 40290
rect 13470 40238 13522 40290
rect 13522 40238 13524 40290
rect 13468 40236 13524 40238
rect 13580 39618 13636 39620
rect 13580 39566 13582 39618
rect 13582 39566 13634 39618
rect 13634 39566 13636 39618
rect 13580 39564 13636 39566
rect 13580 39058 13636 39060
rect 13580 39006 13582 39058
rect 13582 39006 13634 39058
rect 13634 39006 13636 39058
rect 13580 39004 13636 39006
rect 14252 40236 14308 40292
rect 14140 38108 14196 38164
rect 13804 38050 13860 38052
rect 13804 37998 13806 38050
rect 13806 37998 13858 38050
rect 13858 37998 13860 38050
rect 13804 37996 13860 37998
rect 12460 35756 12516 35812
rect 12572 35420 12628 35476
rect 13356 37100 13412 37156
rect 13356 36428 13412 36484
rect 13804 36482 13860 36484
rect 13804 36430 13806 36482
rect 13806 36430 13858 36482
rect 13858 36430 13860 36482
rect 13804 36428 13860 36430
rect 12908 35586 12964 35588
rect 12908 35534 12910 35586
rect 12910 35534 12962 35586
rect 12962 35534 12964 35586
rect 12908 35532 12964 35534
rect 12236 34354 12292 34356
rect 12236 34302 12238 34354
rect 12238 34302 12290 34354
rect 12290 34302 12292 34354
rect 12236 34300 12292 34302
rect 12684 34300 12740 34356
rect 12348 32396 12404 32452
rect 11004 30716 11060 30772
rect 11564 30380 11620 30436
rect 11004 28252 11060 28308
rect 11564 28252 11620 28308
rect 12124 31612 12180 31668
rect 12908 33346 12964 33348
rect 12908 33294 12910 33346
rect 12910 33294 12962 33346
rect 12962 33294 12964 33346
rect 12908 33292 12964 33294
rect 12012 29986 12068 29988
rect 12012 29934 12014 29986
rect 12014 29934 12066 29986
rect 12066 29934 12068 29986
rect 12012 29932 12068 29934
rect 11788 27858 11844 27860
rect 11788 27806 11790 27858
rect 11790 27806 11842 27858
rect 11842 27806 11844 27858
rect 11788 27804 11844 27806
rect 11788 27356 11844 27412
rect 9996 26460 10052 26516
rect 10444 26012 10500 26068
rect 9660 25116 9716 25172
rect 9548 24050 9604 24052
rect 9548 23998 9550 24050
rect 9550 23998 9602 24050
rect 9602 23998 9604 24050
rect 9548 23996 9604 23998
rect 9436 23436 9492 23492
rect 8764 23378 8820 23380
rect 8764 23326 8766 23378
rect 8766 23326 8818 23378
rect 8818 23326 8820 23378
rect 8764 23324 8820 23326
rect 7420 23266 7476 23268
rect 7420 23214 7422 23266
rect 7422 23214 7474 23266
rect 7474 23214 7476 23266
rect 7420 23212 7476 23214
rect 9660 23266 9716 23268
rect 9660 23214 9662 23266
rect 9662 23214 9714 23266
rect 9714 23214 9716 23266
rect 9660 23212 9716 23214
rect 7532 22316 7588 22372
rect 7308 21868 7364 21924
rect 7308 20860 7364 20916
rect 7420 20802 7476 20804
rect 7420 20750 7422 20802
rect 7422 20750 7474 20802
rect 7474 20750 7476 20802
rect 7420 20748 7476 20750
rect 7308 20524 7364 20580
rect 7532 20300 7588 20356
rect 6748 20188 6804 20244
rect 6412 19404 6468 19460
rect 6972 19740 7028 19796
rect 6188 19292 6244 19348
rect 6076 19068 6132 19124
rect 5740 18396 5796 18452
rect 5068 18338 5124 18340
rect 5068 18286 5070 18338
rect 5070 18286 5122 18338
rect 5122 18286 5124 18338
rect 5068 18284 5124 18286
rect 8876 23154 8932 23156
rect 8876 23102 8878 23154
rect 8878 23102 8930 23154
rect 8930 23102 8932 23154
rect 8876 23100 8932 23102
rect 7868 22258 7924 22260
rect 7868 22206 7870 22258
rect 7870 22206 7922 22258
rect 7922 22206 7924 22258
rect 7868 22204 7924 22206
rect 8316 21868 8372 21924
rect 8092 21420 8148 21476
rect 7980 20972 8036 21028
rect 8204 20972 8260 21028
rect 8540 21532 8596 21588
rect 9436 21980 9492 22036
rect 9436 21586 9492 21588
rect 9436 21534 9438 21586
rect 9438 21534 9490 21586
rect 9490 21534 9492 21586
rect 9436 21532 9492 21534
rect 9436 21308 9492 21364
rect 8876 20972 8932 21028
rect 7420 19852 7476 19908
rect 7532 18956 7588 19012
rect 5068 17778 5124 17780
rect 5068 17726 5070 17778
rect 5070 17726 5122 17778
rect 5122 17726 5124 17778
rect 5068 17724 5124 17726
rect 6972 18172 7028 18228
rect 7308 18508 7364 18564
rect 7868 18396 7924 18452
rect 8092 19068 8148 19124
rect 6188 17666 6244 17668
rect 6188 17614 6190 17666
rect 6190 17614 6242 17666
rect 6242 17614 6244 17666
rect 6188 17612 6244 17614
rect 4284 17106 4340 17108
rect 4284 17054 4286 17106
rect 4286 17054 4338 17106
rect 4338 17054 4340 17106
rect 4284 17052 4340 17054
rect 4060 16156 4116 16212
rect 4284 16716 4340 16772
rect 4060 15314 4116 15316
rect 4060 15262 4062 15314
rect 4062 15262 4114 15314
rect 4114 15262 4116 15314
rect 4060 15260 4116 15262
rect 5068 16716 5124 16772
rect 5180 16828 5236 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4620 16210 4676 16212
rect 4620 16158 4622 16210
rect 4622 16158 4674 16210
rect 4674 16158 4676 16210
rect 4620 16156 4676 16158
rect 4732 15708 4788 15764
rect 4844 15596 4900 15652
rect 4508 15314 4564 15316
rect 4508 15262 4510 15314
rect 4510 15262 4562 15314
rect 4562 15262 4564 15314
rect 4508 15260 4564 15262
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5516 16716 5572 16772
rect 3388 13074 3444 13076
rect 3388 13022 3390 13074
rect 3390 13022 3442 13074
rect 3442 13022 3444 13074
rect 3388 13020 3444 13022
rect 2044 12738 2100 12740
rect 2044 12686 2046 12738
rect 2046 12686 2098 12738
rect 2098 12686 2100 12738
rect 2044 12684 2100 12686
rect 2044 12460 2100 12516
rect 5068 14530 5124 14532
rect 5068 14478 5070 14530
rect 5070 14478 5122 14530
rect 5122 14478 5124 14530
rect 5068 14476 5124 14478
rect 4284 13356 4340 13412
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 3612 12348 3668 12404
rect 2492 11676 2548 11732
rect 2604 12012 2660 12068
rect 2044 11564 2100 11620
rect 4172 12572 4228 12628
rect 3276 12066 3332 12068
rect 3276 12014 3278 12066
rect 3278 12014 3330 12066
rect 3330 12014 3332 12066
rect 3276 12012 3332 12014
rect 3164 11452 3220 11508
rect 3388 11900 3444 11956
rect 2716 11340 2772 11396
rect 2380 10780 2436 10836
rect 3948 11676 4004 11732
rect 4508 12402 4564 12404
rect 4508 12350 4510 12402
rect 4510 12350 4562 12402
rect 4562 12350 4564 12402
rect 4508 12348 4564 12350
rect 5068 13634 5124 13636
rect 5068 13582 5070 13634
rect 5070 13582 5122 13634
rect 5122 13582 5124 13634
rect 5068 13580 5124 13582
rect 4956 13020 5012 13076
rect 6636 16770 6692 16772
rect 6636 16718 6638 16770
rect 6638 16718 6690 16770
rect 6690 16718 6692 16770
rect 6636 16716 6692 16718
rect 7308 17724 7364 17780
rect 6860 17276 6916 17332
rect 6972 16492 7028 16548
rect 6972 16268 7028 16324
rect 5964 15484 6020 15540
rect 7084 15820 7140 15876
rect 6076 15260 6132 15316
rect 6188 15484 6244 15540
rect 6748 15260 6804 15316
rect 5964 15036 6020 15092
rect 7084 15148 7140 15204
rect 6972 15036 7028 15092
rect 5292 13468 5348 13524
rect 5740 12962 5796 12964
rect 5740 12910 5742 12962
rect 5742 12910 5794 12962
rect 5794 12910 5796 12962
rect 5740 12908 5796 12910
rect 4844 12290 4900 12292
rect 4844 12238 4846 12290
rect 4846 12238 4898 12290
rect 4898 12238 4900 12290
rect 4844 12236 4900 12238
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4956 11228 5012 11284
rect 5852 12402 5908 12404
rect 5852 12350 5854 12402
rect 5854 12350 5906 12402
rect 5906 12350 5908 12402
rect 5852 12348 5908 12350
rect 6076 12236 6132 12292
rect 7532 17554 7588 17556
rect 7532 17502 7534 17554
rect 7534 17502 7586 17554
rect 7586 17502 7588 17554
rect 7532 17500 7588 17502
rect 7756 17554 7812 17556
rect 7756 17502 7758 17554
rect 7758 17502 7810 17554
rect 7810 17502 7812 17554
rect 7756 17500 7812 17502
rect 8540 20524 8596 20580
rect 8652 20748 8708 20804
rect 8876 20636 8932 20692
rect 8876 20130 8932 20132
rect 8876 20078 8878 20130
rect 8878 20078 8930 20130
rect 8930 20078 8932 20130
rect 8876 20076 8932 20078
rect 9212 19852 9268 19908
rect 8428 19346 8484 19348
rect 8428 19294 8430 19346
rect 8430 19294 8482 19346
rect 8482 19294 8484 19346
rect 8428 19292 8484 19294
rect 8316 19180 8372 19236
rect 8316 17724 8372 17780
rect 8092 17554 8148 17556
rect 8092 17502 8094 17554
rect 8094 17502 8146 17554
rect 8146 17502 8148 17554
rect 8092 17500 8148 17502
rect 7868 17276 7924 17332
rect 8204 16492 8260 16548
rect 8092 16268 8148 16324
rect 8540 18396 8596 18452
rect 8652 18956 8708 19012
rect 8988 18732 9044 18788
rect 8876 18674 8932 18676
rect 8876 18622 8878 18674
rect 8878 18622 8930 18674
rect 8930 18622 8932 18674
rect 8876 18620 8932 18622
rect 8764 18284 8820 18340
rect 10108 25116 10164 25172
rect 10556 24668 10612 24724
rect 9884 23660 9940 23716
rect 9884 23324 9940 23380
rect 9996 23154 10052 23156
rect 9996 23102 9998 23154
rect 9998 23102 10050 23154
rect 10050 23102 10052 23154
rect 9996 23100 10052 23102
rect 10556 22876 10612 22932
rect 9996 22428 10052 22484
rect 10556 22428 10612 22484
rect 9660 20300 9716 20356
rect 9548 20018 9604 20020
rect 9548 19966 9550 20018
rect 9550 19966 9602 20018
rect 9602 19966 9604 20018
rect 9548 19964 9604 19966
rect 9884 19964 9940 20020
rect 9212 18620 9268 18676
rect 9324 18732 9380 18788
rect 8876 17948 8932 18004
rect 8876 17666 8932 17668
rect 8876 17614 8878 17666
rect 8878 17614 8930 17666
rect 8930 17614 8932 17666
rect 8876 17612 8932 17614
rect 9324 17948 9380 18004
rect 8764 16322 8820 16324
rect 8764 16270 8766 16322
rect 8766 16270 8818 16322
rect 8818 16270 8820 16322
rect 8764 16268 8820 16270
rect 8316 15596 8372 15652
rect 8092 15260 8148 15316
rect 7420 15036 7476 15092
rect 7756 14530 7812 14532
rect 7756 14478 7758 14530
rect 7758 14478 7810 14530
rect 7810 14478 7812 14530
rect 7756 14476 7812 14478
rect 7308 14364 7364 14420
rect 7756 14140 7812 14196
rect 7196 14028 7252 14084
rect 6972 13356 7028 13412
rect 6412 12460 6468 12516
rect 5292 12178 5348 12180
rect 5292 12126 5294 12178
rect 5294 12126 5346 12178
rect 5346 12126 5348 12178
rect 5292 12124 5348 12126
rect 6860 12290 6916 12292
rect 6860 12238 6862 12290
rect 6862 12238 6914 12290
rect 6914 12238 6916 12290
rect 6860 12236 6916 12238
rect 3948 10834 4004 10836
rect 3948 10782 3950 10834
rect 3950 10782 4002 10834
rect 4002 10782 4004 10834
rect 3948 10780 4004 10782
rect 2044 9826 2100 9828
rect 2044 9774 2046 9826
rect 2046 9774 2098 9826
rect 2098 9774 2100 9826
rect 2044 9772 2100 9774
rect 2492 10668 2548 10724
rect 4396 10722 4452 10724
rect 4396 10670 4398 10722
rect 4398 10670 4450 10722
rect 4450 10670 4452 10722
rect 4396 10668 4452 10670
rect 4956 10668 5012 10724
rect 3052 10108 3108 10164
rect 3836 10108 3892 10164
rect 2716 9714 2772 9716
rect 2716 9662 2718 9714
rect 2718 9662 2770 9714
rect 2770 9662 2772 9714
rect 2716 9660 2772 9662
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4284 9884 4340 9940
rect 5740 11506 5796 11508
rect 5740 11454 5742 11506
rect 5742 11454 5794 11506
rect 5794 11454 5796 11506
rect 5740 11452 5796 11454
rect 5628 11282 5684 11284
rect 5628 11230 5630 11282
rect 5630 11230 5682 11282
rect 5682 11230 5684 11282
rect 5628 11228 5684 11230
rect 5516 10834 5572 10836
rect 5516 10782 5518 10834
rect 5518 10782 5570 10834
rect 5570 10782 5572 10834
rect 5516 10780 5572 10782
rect 5628 10444 5684 10500
rect 5180 10332 5236 10388
rect 5068 9772 5124 9828
rect 5516 9884 5572 9940
rect 5964 10668 6020 10724
rect 7644 13858 7700 13860
rect 7644 13806 7646 13858
rect 7646 13806 7698 13858
rect 7698 13806 7700 13858
rect 7644 13804 7700 13806
rect 6860 11900 6916 11956
rect 7980 14252 8036 14308
rect 7980 14028 8036 14084
rect 8204 14476 8260 14532
rect 8652 15260 8708 15316
rect 8428 15148 8484 15204
rect 8316 14364 8372 14420
rect 8092 13356 8148 13412
rect 8988 15874 9044 15876
rect 8988 15822 8990 15874
rect 8990 15822 9042 15874
rect 9042 15822 9044 15874
rect 8988 15820 9044 15822
rect 9436 15596 9492 15652
rect 9884 19234 9940 19236
rect 9884 19182 9886 19234
rect 9886 19182 9938 19234
rect 9938 19182 9940 19234
rect 9884 19180 9940 19182
rect 9660 18956 9716 19012
rect 10108 20636 10164 20692
rect 11004 26460 11060 26516
rect 11676 26066 11732 26068
rect 11676 26014 11678 26066
rect 11678 26014 11730 26066
rect 11730 26014 11732 26066
rect 11676 26012 11732 26014
rect 11116 25116 11172 25172
rect 11564 23436 11620 23492
rect 12572 31500 12628 31556
rect 12460 30994 12516 30996
rect 12460 30942 12462 30994
rect 12462 30942 12514 30994
rect 12514 30942 12516 30994
rect 12460 30940 12516 30942
rect 12796 30828 12852 30884
rect 12572 29986 12628 29988
rect 12572 29934 12574 29986
rect 12574 29934 12626 29986
rect 12626 29934 12628 29986
rect 12572 29932 12628 29934
rect 12796 28530 12852 28532
rect 12796 28478 12798 28530
rect 12798 28478 12850 28530
rect 12850 28478 12852 28530
rect 12796 28476 12852 28478
rect 12572 28364 12628 28420
rect 12684 28252 12740 28308
rect 12460 27356 12516 27412
rect 12124 26908 12180 26964
rect 12796 27970 12852 27972
rect 12796 27918 12798 27970
rect 12798 27918 12850 27970
rect 12850 27918 12852 27970
rect 12796 27916 12852 27918
rect 13356 34636 13412 34692
rect 13580 33292 13636 33348
rect 13692 35420 13748 35476
rect 13468 33122 13524 33124
rect 13468 33070 13470 33122
rect 13470 33070 13522 33122
rect 13522 33070 13524 33122
rect 13468 33068 13524 33070
rect 13356 32060 13412 32116
rect 14252 37826 14308 37828
rect 14252 37774 14254 37826
rect 14254 37774 14306 37826
rect 14306 37774 14308 37826
rect 14252 37772 14308 37774
rect 14364 37266 14420 37268
rect 14364 37214 14366 37266
rect 14366 37214 14418 37266
rect 14418 37214 14420 37266
rect 14364 37212 14420 37214
rect 14700 42476 14756 42532
rect 14812 42700 14868 42756
rect 14588 41074 14644 41076
rect 14588 41022 14590 41074
rect 14590 41022 14642 41074
rect 14642 41022 14644 41074
rect 14588 41020 14644 41022
rect 14700 40908 14756 40964
rect 15148 42530 15204 42532
rect 15148 42478 15150 42530
rect 15150 42478 15202 42530
rect 15202 42478 15204 42530
rect 15148 42476 15204 42478
rect 15036 41916 15092 41972
rect 14924 41244 14980 41300
rect 15036 41186 15092 41188
rect 15036 41134 15038 41186
rect 15038 41134 15090 41186
rect 15090 41134 15092 41186
rect 15036 41132 15092 41134
rect 17500 49810 17556 49812
rect 17500 49758 17502 49810
rect 17502 49758 17554 49810
rect 17554 49758 17556 49810
rect 17500 49756 17556 49758
rect 17052 49644 17108 49700
rect 16716 48748 16772 48804
rect 16492 48300 16548 48356
rect 16380 48076 16436 48132
rect 16380 46674 16436 46676
rect 16380 46622 16382 46674
rect 16382 46622 16434 46674
rect 16434 46622 16436 46674
rect 16380 46620 16436 46622
rect 15484 44716 15540 44772
rect 15820 44604 15876 44660
rect 15484 44492 15540 44548
rect 15596 44268 15652 44324
rect 16380 44268 16436 44324
rect 15484 43708 15540 43764
rect 14924 40572 14980 40628
rect 14812 38162 14868 38164
rect 14812 38110 14814 38162
rect 14814 38110 14866 38162
rect 14866 38110 14868 38162
rect 14812 38108 14868 38110
rect 14812 37378 14868 37380
rect 14812 37326 14814 37378
rect 14814 37326 14866 37378
rect 14866 37326 14868 37378
rect 14812 37324 14868 37326
rect 14700 37212 14756 37268
rect 14476 36428 14532 36484
rect 15484 40236 15540 40292
rect 16044 42476 16100 42532
rect 15820 41186 15876 41188
rect 15820 41134 15822 41186
rect 15822 41134 15874 41186
rect 15874 41134 15876 41186
rect 15820 41132 15876 41134
rect 16380 41020 16436 41076
rect 15932 40962 15988 40964
rect 15932 40910 15934 40962
rect 15934 40910 15986 40962
rect 15986 40910 15988 40962
rect 15932 40908 15988 40910
rect 16380 40348 16436 40404
rect 16716 46786 16772 46788
rect 16716 46734 16718 46786
rect 16718 46734 16770 46786
rect 16770 46734 16772 46786
rect 16716 46732 16772 46734
rect 17388 49644 17444 49700
rect 17276 49532 17332 49588
rect 17164 48802 17220 48804
rect 17164 48750 17166 48802
rect 17166 48750 17218 48802
rect 17218 48750 17220 48802
rect 17164 48748 17220 48750
rect 17164 47458 17220 47460
rect 17164 47406 17166 47458
rect 17166 47406 17218 47458
rect 17218 47406 17220 47458
rect 17164 47404 17220 47406
rect 18844 53730 18900 53732
rect 18844 53678 18846 53730
rect 18846 53678 18898 53730
rect 18898 53678 18900 53730
rect 18844 53676 18900 53678
rect 18956 53618 19012 53620
rect 18956 53566 18958 53618
rect 18958 53566 19010 53618
rect 19010 53566 19012 53618
rect 18956 53564 19012 53566
rect 18396 53340 18452 53396
rect 19180 53618 19236 53620
rect 19180 53566 19182 53618
rect 19182 53566 19234 53618
rect 19234 53566 19236 53618
rect 19180 53564 19236 53566
rect 18956 53116 19012 53172
rect 19292 53340 19348 53396
rect 19852 54348 19908 54404
rect 19740 53730 19796 53732
rect 19740 53678 19742 53730
rect 19742 53678 19794 53730
rect 19794 53678 19796 53730
rect 19740 53676 19796 53678
rect 19964 53676 20020 53732
rect 22988 55244 23044 55300
rect 23324 54684 23380 54740
rect 20300 53676 20356 53732
rect 20188 53618 20244 53620
rect 20188 53566 20190 53618
rect 20190 53566 20242 53618
rect 20242 53566 20244 53618
rect 20188 53564 20244 53566
rect 19964 53506 20020 53508
rect 19964 53454 19966 53506
rect 19966 53454 20018 53506
rect 20018 53454 20020 53506
rect 19964 53452 20020 53454
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 18620 52834 18676 52836
rect 18620 52782 18622 52834
rect 18622 52782 18674 52834
rect 18674 52782 18676 52834
rect 18620 52780 18676 52782
rect 20412 52556 20468 52612
rect 18172 52108 18228 52164
rect 17836 49980 17892 50036
rect 17724 49586 17780 49588
rect 17724 49534 17726 49586
rect 17726 49534 17778 49586
rect 17778 49534 17780 49586
rect 17724 49532 17780 49534
rect 17836 48354 17892 48356
rect 17836 48302 17838 48354
rect 17838 48302 17890 48354
rect 17890 48302 17892 48354
rect 17836 48300 17892 48302
rect 17612 47404 17668 47460
rect 17948 46844 18004 46900
rect 18060 48300 18116 48356
rect 17948 46674 18004 46676
rect 17948 46622 17950 46674
rect 17950 46622 18002 46674
rect 18002 46622 18004 46674
rect 17948 46620 18004 46622
rect 16828 45612 16884 45668
rect 17276 44716 17332 44772
rect 16828 43260 16884 43316
rect 17612 45836 17668 45892
rect 17948 46060 18004 46116
rect 17500 45106 17556 45108
rect 17500 45054 17502 45106
rect 17502 45054 17554 45106
rect 17554 45054 17556 45106
rect 17500 45052 17556 45054
rect 19180 52162 19236 52164
rect 19180 52110 19182 52162
rect 19182 52110 19234 52162
rect 19234 52110 19236 52162
rect 19180 52108 19236 52110
rect 19740 52108 19796 52164
rect 18732 51772 18788 51828
rect 19516 51660 19572 51716
rect 19404 51212 19460 51268
rect 19068 50594 19124 50596
rect 19068 50542 19070 50594
rect 19070 50542 19122 50594
rect 19122 50542 19124 50594
rect 19068 50540 19124 50542
rect 18396 50034 18452 50036
rect 18396 49982 18398 50034
rect 18398 49982 18450 50034
rect 18450 49982 18452 50034
rect 18396 49980 18452 49982
rect 18508 49756 18564 49812
rect 20412 52162 20468 52164
rect 20412 52110 20414 52162
rect 20414 52110 20466 52162
rect 20466 52110 20468 52162
rect 20412 52108 20468 52110
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 20748 53788 20804 53844
rect 21980 53676 22036 53732
rect 21644 53340 21700 53396
rect 20636 52274 20692 52276
rect 20636 52222 20638 52274
rect 20638 52222 20690 52274
rect 20690 52222 20692 52274
rect 20636 52220 20692 52222
rect 20748 52162 20804 52164
rect 20748 52110 20750 52162
rect 20750 52110 20802 52162
rect 20802 52110 20804 52162
rect 20748 52108 20804 52110
rect 20188 50540 20244 50596
rect 19740 50316 19796 50372
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19516 49810 19572 49812
rect 19516 49758 19518 49810
rect 19518 49758 19570 49810
rect 19570 49758 19572 49810
rect 19516 49756 19572 49758
rect 19628 49698 19684 49700
rect 19628 49646 19630 49698
rect 19630 49646 19682 49698
rect 19682 49646 19684 49698
rect 19628 49644 19684 49646
rect 18284 46060 18340 46116
rect 18620 46844 18676 46900
rect 18396 44210 18452 44212
rect 18396 44158 18398 44210
rect 18398 44158 18450 44210
rect 18450 44158 18452 44210
rect 18396 44156 18452 44158
rect 17500 43650 17556 43652
rect 17500 43598 17502 43650
rect 17502 43598 17554 43650
rect 17554 43598 17556 43650
rect 17500 43596 17556 43598
rect 16604 40962 16660 40964
rect 16604 40910 16606 40962
rect 16606 40910 16658 40962
rect 16658 40910 16660 40962
rect 16604 40908 16660 40910
rect 16940 40460 16996 40516
rect 16828 40290 16884 40292
rect 16828 40238 16830 40290
rect 16830 40238 16882 40290
rect 16882 40238 16884 40290
rect 16828 40236 16884 40238
rect 16828 39564 16884 39620
rect 15484 37938 15540 37940
rect 15484 37886 15486 37938
rect 15486 37886 15538 37938
rect 15538 37886 15540 37938
rect 15484 37884 15540 37886
rect 16044 38892 16100 38948
rect 15820 38050 15876 38052
rect 15820 37998 15822 38050
rect 15822 37998 15874 38050
rect 15874 37998 15876 38050
rect 15820 37996 15876 37998
rect 15708 37042 15764 37044
rect 15708 36990 15710 37042
rect 15710 36990 15762 37042
rect 15762 36990 15764 37042
rect 15708 36988 15764 36990
rect 16156 37212 16212 37268
rect 14588 35868 14644 35924
rect 14364 35756 14420 35812
rect 14140 35698 14196 35700
rect 14140 35646 14142 35698
rect 14142 35646 14194 35698
rect 14194 35646 14196 35698
rect 14140 35644 14196 35646
rect 16044 36258 16100 36260
rect 16044 36206 16046 36258
rect 16046 36206 16098 36258
rect 16098 36206 16100 36258
rect 16044 36204 16100 36206
rect 16604 37938 16660 37940
rect 16604 37886 16606 37938
rect 16606 37886 16658 37938
rect 16658 37886 16660 37938
rect 16604 37884 16660 37886
rect 17836 43260 17892 43316
rect 17724 43148 17780 43204
rect 18956 43596 19012 43652
rect 20076 48860 20132 48916
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19516 48242 19572 48244
rect 19516 48190 19518 48242
rect 19518 48190 19570 48242
rect 19570 48190 19572 48242
rect 19516 48188 19572 48190
rect 21644 52780 21700 52836
rect 22092 53506 22148 53508
rect 22092 53454 22094 53506
rect 22094 53454 22146 53506
rect 22146 53454 22148 53506
rect 22092 53452 22148 53454
rect 22092 53004 22148 53060
rect 22652 53676 22708 53732
rect 22988 53564 23044 53620
rect 22316 53340 22372 53396
rect 22204 53116 22260 53172
rect 21420 52220 21476 52276
rect 21868 52444 21924 52500
rect 21980 52162 22036 52164
rect 21980 52110 21982 52162
rect 21982 52110 22034 52162
rect 22034 52110 22036 52162
rect 21980 52108 22036 52110
rect 23212 53452 23268 53508
rect 22988 53004 23044 53060
rect 22428 52162 22484 52164
rect 22428 52110 22430 52162
rect 22430 52110 22482 52162
rect 22482 52110 22484 52162
rect 22428 52108 22484 52110
rect 23548 52108 23604 52164
rect 23324 51548 23380 51604
rect 23660 51490 23716 51492
rect 23660 51438 23662 51490
rect 23662 51438 23714 51490
rect 23714 51438 23716 51490
rect 23660 51436 23716 51438
rect 20636 50316 20692 50372
rect 20636 50034 20692 50036
rect 20636 49982 20638 50034
rect 20638 49982 20690 50034
rect 20690 49982 20692 50034
rect 20636 49980 20692 49982
rect 20412 49698 20468 49700
rect 20412 49646 20414 49698
rect 20414 49646 20466 49698
rect 20466 49646 20468 49698
rect 20412 49644 20468 49646
rect 19516 47404 19572 47460
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19628 46060 19684 46116
rect 20188 46620 20244 46676
rect 19852 45948 19908 46004
rect 20524 46674 20580 46676
rect 20524 46622 20526 46674
rect 20526 46622 20578 46674
rect 20578 46622 20580 46674
rect 20524 46620 20580 46622
rect 20636 46508 20692 46564
rect 19964 45612 20020 45668
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19404 44210 19460 44212
rect 19404 44158 19406 44210
rect 19406 44158 19458 44210
rect 19458 44158 19460 44210
rect 19404 44156 19460 44158
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19964 43708 20020 43764
rect 19068 43148 19124 43204
rect 19852 43650 19908 43652
rect 19852 43598 19854 43650
rect 19854 43598 19906 43650
rect 19906 43598 19908 43650
rect 19852 43596 19908 43598
rect 20524 45948 20580 46004
rect 20412 45890 20468 45892
rect 20412 45838 20414 45890
rect 20414 45838 20466 45890
rect 20466 45838 20468 45890
rect 20412 45836 20468 45838
rect 20748 46002 20804 46004
rect 20748 45950 20750 46002
rect 20750 45950 20802 46002
rect 20802 45950 20804 46002
rect 20748 45948 20804 45950
rect 20300 45612 20356 45668
rect 20748 45052 20804 45108
rect 21756 50204 21812 50260
rect 21308 49756 21364 49812
rect 21756 50034 21812 50036
rect 21756 49982 21758 50034
rect 21758 49982 21810 50034
rect 21810 49982 21812 50034
rect 21756 49980 21812 49982
rect 22092 50482 22148 50484
rect 22092 50430 22094 50482
rect 22094 50430 22146 50482
rect 22146 50430 22148 50482
rect 22092 50428 22148 50430
rect 22988 51266 23044 51268
rect 22988 51214 22990 51266
rect 22990 51214 23042 51266
rect 23042 51214 23044 51266
rect 22988 51212 23044 51214
rect 23436 51212 23492 51268
rect 24108 53564 24164 53620
rect 24444 53058 24500 53060
rect 24444 53006 24446 53058
rect 24446 53006 24498 53058
rect 24498 53006 24500 53058
rect 24444 53004 24500 53006
rect 24220 52556 24276 52612
rect 24220 52332 24276 52388
rect 24668 52668 24724 52724
rect 24668 52274 24724 52276
rect 24668 52222 24670 52274
rect 24670 52222 24722 52274
rect 24722 52222 24724 52274
rect 24668 52220 24724 52222
rect 23772 50540 23828 50596
rect 24556 50594 24612 50596
rect 24556 50542 24558 50594
rect 24558 50542 24610 50594
rect 24610 50542 24612 50594
rect 24556 50540 24612 50542
rect 21868 48188 21924 48244
rect 21084 46844 21140 46900
rect 21420 45500 21476 45556
rect 22204 48860 22260 48916
rect 22092 46620 22148 46676
rect 21868 45890 21924 45892
rect 21868 45838 21870 45890
rect 21870 45838 21922 45890
rect 21922 45838 21924 45890
rect 21868 45836 21924 45838
rect 21644 45388 21700 45444
rect 21868 45612 21924 45668
rect 20188 43484 20244 43540
rect 20524 43596 20580 43652
rect 18172 42978 18228 42980
rect 18172 42926 18174 42978
rect 18174 42926 18226 42978
rect 18226 42926 18228 42978
rect 18172 42924 18228 42926
rect 18284 42866 18340 42868
rect 18284 42814 18286 42866
rect 18286 42814 18338 42866
rect 18338 42814 18340 42866
rect 18284 42812 18340 42814
rect 17836 42642 17892 42644
rect 17836 42590 17838 42642
rect 17838 42590 17890 42642
rect 17890 42590 17892 42642
rect 17836 42588 17892 42590
rect 17724 38892 17780 38948
rect 16492 36988 16548 37044
rect 16940 37100 16996 37156
rect 16716 36482 16772 36484
rect 16716 36430 16718 36482
rect 16718 36430 16770 36482
rect 16770 36430 16772 36482
rect 16716 36428 16772 36430
rect 15596 35922 15652 35924
rect 15596 35870 15598 35922
rect 15598 35870 15650 35922
rect 15650 35870 15652 35922
rect 15596 35868 15652 35870
rect 15036 35756 15092 35812
rect 14252 35308 14308 35364
rect 14140 34690 14196 34692
rect 14140 34638 14142 34690
rect 14142 34638 14194 34690
rect 14194 34638 14196 34690
rect 14140 34636 14196 34638
rect 14252 33404 14308 33460
rect 14028 33292 14084 33348
rect 14252 32956 14308 33012
rect 14364 33068 14420 33124
rect 14476 32844 14532 32900
rect 15148 35586 15204 35588
rect 15148 35534 15150 35586
rect 15150 35534 15202 35586
rect 15202 35534 15204 35586
rect 15148 35532 15204 35534
rect 15148 34300 15204 34356
rect 14924 33068 14980 33124
rect 14588 32732 14644 32788
rect 13916 32284 13972 32340
rect 14140 32338 14196 32340
rect 14140 32286 14142 32338
rect 14142 32286 14194 32338
rect 14194 32286 14196 32338
rect 14140 32284 14196 32286
rect 15148 33122 15204 33124
rect 15148 33070 15150 33122
rect 15150 33070 15202 33122
rect 15202 33070 15204 33122
rect 15148 33068 15204 33070
rect 15148 32844 15204 32900
rect 14364 32284 14420 32340
rect 13804 32060 13860 32116
rect 14140 32060 14196 32116
rect 13916 31388 13972 31444
rect 13244 30882 13300 30884
rect 13244 30830 13246 30882
rect 13246 30830 13298 30882
rect 13298 30830 13300 30882
rect 13244 30828 13300 30830
rect 13020 30268 13076 30324
rect 13804 30098 13860 30100
rect 13804 30046 13806 30098
rect 13806 30046 13858 30098
rect 13858 30046 13860 30098
rect 13804 30044 13860 30046
rect 13580 28476 13636 28532
rect 14028 28418 14084 28420
rect 14028 28366 14030 28418
rect 14030 28366 14082 28418
rect 14082 28366 14084 28418
rect 14028 28364 14084 28366
rect 12908 27020 12964 27076
rect 11900 25116 11956 25172
rect 12236 24610 12292 24612
rect 12236 24558 12238 24610
rect 12238 24558 12290 24610
rect 12290 24558 12292 24610
rect 12236 24556 12292 24558
rect 12460 24332 12516 24388
rect 12908 24050 12964 24052
rect 12908 23998 12910 24050
rect 12910 23998 12962 24050
rect 12962 23998 12964 24050
rect 12908 23996 12964 23998
rect 12572 23548 12628 23604
rect 11788 23324 11844 23380
rect 12012 23324 12068 23380
rect 11900 22988 11956 23044
rect 11564 22764 11620 22820
rect 11564 22540 11620 22596
rect 11340 22428 11396 22484
rect 10780 21420 10836 21476
rect 10220 19740 10276 19796
rect 10556 20076 10612 20132
rect 10332 18732 10388 18788
rect 10220 18620 10276 18676
rect 11116 19010 11172 19012
rect 11116 18958 11118 19010
rect 11118 18958 11170 19010
rect 11170 18958 11172 19010
rect 11116 18956 11172 18958
rect 11004 18620 11060 18676
rect 10332 18172 10388 18228
rect 11452 19740 11508 19796
rect 11340 18450 11396 18452
rect 11340 18398 11342 18450
rect 11342 18398 11394 18450
rect 11394 18398 11396 18450
rect 11340 18396 11396 18398
rect 10220 17052 10276 17108
rect 9884 16492 9940 16548
rect 9660 15596 9716 15652
rect 9884 15596 9940 15652
rect 10444 15538 10500 15540
rect 10444 15486 10446 15538
rect 10446 15486 10498 15538
rect 10498 15486 10500 15538
rect 10444 15484 10500 15486
rect 9884 15314 9940 15316
rect 9884 15262 9886 15314
rect 9886 15262 9938 15314
rect 9938 15262 9940 15314
rect 9884 15260 9940 15262
rect 7756 12460 7812 12516
rect 7644 11564 7700 11620
rect 7308 10834 7364 10836
rect 7308 10782 7310 10834
rect 7310 10782 7362 10834
rect 7362 10782 7364 10834
rect 7308 10780 7364 10782
rect 7868 10780 7924 10836
rect 6524 10610 6580 10612
rect 6524 10558 6526 10610
rect 6526 10558 6578 10610
rect 6578 10558 6580 10610
rect 6524 10556 6580 10558
rect 7084 10556 7140 10612
rect 6188 10444 6244 10500
rect 6076 9714 6132 9716
rect 6076 9662 6078 9714
rect 6078 9662 6130 9714
rect 6130 9662 6132 9714
rect 6076 9660 6132 9662
rect 5964 9212 6020 9268
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 5068 8428 5124 8484
rect 10892 17388 10948 17444
rect 11340 17276 11396 17332
rect 11340 17106 11396 17108
rect 11340 17054 11342 17106
rect 11342 17054 11394 17106
rect 11394 17054 11396 17106
rect 11340 17052 11396 17054
rect 11004 15596 11060 15652
rect 10108 15148 10164 15204
rect 10444 14476 10500 14532
rect 9996 13746 10052 13748
rect 9996 13694 9998 13746
rect 9998 13694 10050 13746
rect 10050 13694 10052 13746
rect 9996 13692 10052 13694
rect 11676 18620 11732 18676
rect 13132 27804 13188 27860
rect 13916 27970 13972 27972
rect 13916 27918 13918 27970
rect 13918 27918 13970 27970
rect 13970 27918 13972 27970
rect 13916 27916 13972 27918
rect 13692 27132 13748 27188
rect 13244 27020 13300 27076
rect 14028 27132 14084 27188
rect 14700 31666 14756 31668
rect 14700 31614 14702 31666
rect 14702 31614 14754 31666
rect 14754 31614 14756 31666
rect 14700 31612 14756 31614
rect 16156 34242 16212 34244
rect 16156 34190 16158 34242
rect 16158 34190 16210 34242
rect 16210 34190 16212 34242
rect 16156 34188 16212 34190
rect 15484 33458 15540 33460
rect 15484 33406 15486 33458
rect 15486 33406 15538 33458
rect 15538 33406 15540 33458
rect 15484 33404 15540 33406
rect 15484 33234 15540 33236
rect 15484 33182 15486 33234
rect 15486 33182 15538 33234
rect 15538 33182 15540 33234
rect 15484 33180 15540 33182
rect 15372 32562 15428 32564
rect 15372 32510 15374 32562
rect 15374 32510 15426 32562
rect 15426 32510 15428 32562
rect 15372 32508 15428 32510
rect 15932 32508 15988 32564
rect 14924 31836 14980 31892
rect 14924 31612 14980 31668
rect 14364 30828 14420 30884
rect 14700 29708 14756 29764
rect 14588 27356 14644 27412
rect 14700 27020 14756 27076
rect 14028 26684 14084 26740
rect 13468 25228 13524 25284
rect 13132 24332 13188 24388
rect 12796 23100 12852 23156
rect 12684 22988 12740 23044
rect 12012 22482 12068 22484
rect 12012 22430 12014 22482
rect 12014 22430 12066 22482
rect 12066 22430 12068 22482
rect 12012 22428 12068 22430
rect 11676 18450 11732 18452
rect 11676 18398 11678 18450
rect 11678 18398 11730 18450
rect 11730 18398 11732 18450
rect 11676 18396 11732 18398
rect 11676 16268 11732 16324
rect 11788 16098 11844 16100
rect 11788 16046 11790 16098
rect 11790 16046 11842 16098
rect 11842 16046 11844 16098
rect 11788 16044 11844 16046
rect 11676 14700 11732 14756
rect 13132 23042 13188 23044
rect 13132 22990 13134 23042
rect 13134 22990 13186 23042
rect 13186 22990 13188 23042
rect 13132 22988 13188 22990
rect 12348 21868 12404 21924
rect 12012 20524 12068 20580
rect 12012 20130 12068 20132
rect 12012 20078 12014 20130
rect 12014 20078 12066 20130
rect 12066 20078 12068 20130
rect 12012 20076 12068 20078
rect 12012 19180 12068 19236
rect 12124 16156 12180 16212
rect 11900 14588 11956 14644
rect 11116 13916 11172 13972
rect 11452 13692 11508 13748
rect 10444 12684 10500 12740
rect 10668 12738 10724 12740
rect 10668 12686 10670 12738
rect 10670 12686 10722 12738
rect 10722 12686 10724 12738
rect 10668 12684 10724 12686
rect 8652 11900 8708 11956
rect 9100 11900 9156 11956
rect 8988 11788 9044 11844
rect 8540 10780 8596 10836
rect 7868 10556 7924 10612
rect 7532 9324 7588 9380
rect 8428 10444 8484 10500
rect 8764 9772 8820 9828
rect 9996 12012 10052 12068
rect 10108 11788 10164 11844
rect 11340 11506 11396 11508
rect 11340 11454 11342 11506
rect 11342 11454 11394 11506
rect 11394 11454 11396 11506
rect 11340 11452 11396 11454
rect 11452 11340 11508 11396
rect 10668 11116 10724 11172
rect 13020 21868 13076 21924
rect 12684 21756 12740 21812
rect 13468 22540 13524 22596
rect 13468 22316 13524 22372
rect 13468 21868 13524 21924
rect 13356 21810 13412 21812
rect 13356 21758 13358 21810
rect 13358 21758 13410 21810
rect 13410 21758 13412 21810
rect 13356 21756 13412 21758
rect 13916 25730 13972 25732
rect 13916 25678 13918 25730
rect 13918 25678 13970 25730
rect 13970 25678 13972 25730
rect 13916 25676 13972 25678
rect 14476 26460 14532 26516
rect 14588 26684 14644 26740
rect 14252 26236 14308 26292
rect 15260 31666 15316 31668
rect 15260 31614 15262 31666
rect 15262 31614 15314 31666
rect 15314 31614 15316 31666
rect 15260 31612 15316 31614
rect 15148 30828 15204 30884
rect 15372 30268 15428 30324
rect 15036 26572 15092 26628
rect 14476 26012 14532 26068
rect 13692 24668 13748 24724
rect 13916 24332 13972 24388
rect 13804 23324 13860 23380
rect 13692 21810 13748 21812
rect 13692 21758 13694 21810
rect 13694 21758 13746 21810
rect 13746 21758 13748 21810
rect 13692 21756 13748 21758
rect 13692 21420 13748 21476
rect 13244 19740 13300 19796
rect 12908 19346 12964 19348
rect 12908 19294 12910 19346
rect 12910 19294 12962 19346
rect 12962 19294 12964 19346
rect 12908 19292 12964 19294
rect 12460 18732 12516 18788
rect 12460 18508 12516 18564
rect 12348 16098 12404 16100
rect 12348 16046 12350 16098
rect 12350 16046 12402 16098
rect 12402 16046 12404 16098
rect 12348 16044 12404 16046
rect 13020 18060 13076 18116
rect 13356 17724 13412 17780
rect 13132 16994 13188 16996
rect 13132 16942 13134 16994
rect 13134 16942 13186 16994
rect 13186 16942 13188 16994
rect 13132 16940 13188 16942
rect 12796 15932 12852 15988
rect 13132 15596 13188 15652
rect 13020 15314 13076 15316
rect 13020 15262 13022 15314
rect 13022 15262 13074 15314
rect 13074 15262 13076 15314
rect 13020 15260 13076 15262
rect 13580 19292 13636 19348
rect 14028 20076 14084 20132
rect 14364 24668 14420 24724
rect 14700 25282 14756 25284
rect 14700 25230 14702 25282
rect 14702 25230 14754 25282
rect 14754 25230 14756 25282
rect 14700 25228 14756 25230
rect 15036 25564 15092 25620
rect 14924 25116 14980 25172
rect 15148 25228 15204 25284
rect 14812 24610 14868 24612
rect 14812 24558 14814 24610
rect 14814 24558 14866 24610
rect 14866 24558 14868 24610
rect 14812 24556 14868 24558
rect 14700 24332 14756 24388
rect 14812 23324 14868 23380
rect 14252 21868 14308 21924
rect 14700 22146 14756 22148
rect 14700 22094 14702 22146
rect 14702 22094 14754 22146
rect 14754 22094 14756 22146
rect 14700 22092 14756 22094
rect 14252 21586 14308 21588
rect 14252 21534 14254 21586
rect 14254 21534 14306 21586
rect 14306 21534 14308 21586
rect 14252 21532 14308 21534
rect 14588 21420 14644 21476
rect 15260 22258 15316 22260
rect 15260 22206 15262 22258
rect 15262 22206 15314 22258
rect 15314 22206 15316 22258
rect 15260 22204 15316 22206
rect 15148 22146 15204 22148
rect 15148 22094 15150 22146
rect 15150 22094 15202 22146
rect 15202 22094 15204 22146
rect 15148 22092 15204 22094
rect 14924 21532 14980 21588
rect 15148 21474 15204 21476
rect 15148 21422 15150 21474
rect 15150 21422 15202 21474
rect 15202 21422 15204 21474
rect 15148 21420 15204 21422
rect 15596 31612 15652 31668
rect 15820 31890 15876 31892
rect 15820 31838 15822 31890
rect 15822 31838 15874 31890
rect 15874 31838 15876 31890
rect 15820 31836 15876 31838
rect 15708 31276 15764 31332
rect 15596 30882 15652 30884
rect 15596 30830 15598 30882
rect 15598 30830 15650 30882
rect 15650 30830 15652 30882
rect 15596 30828 15652 30830
rect 16380 34130 16436 34132
rect 16380 34078 16382 34130
rect 16382 34078 16434 34130
rect 16434 34078 16436 34130
rect 16380 34076 16436 34078
rect 16156 33068 16212 33124
rect 16492 33180 16548 33236
rect 16828 33068 16884 33124
rect 16828 32396 16884 32452
rect 16380 31554 16436 31556
rect 16380 31502 16382 31554
rect 16382 31502 16434 31554
rect 16434 31502 16436 31554
rect 16380 31500 16436 31502
rect 16380 30940 16436 30996
rect 17500 36988 17556 37044
rect 17164 36652 17220 36708
rect 17388 36370 17444 36372
rect 17388 36318 17390 36370
rect 17390 36318 17442 36370
rect 17442 36318 17444 36370
rect 17388 36316 17444 36318
rect 17164 36204 17220 36260
rect 17052 34300 17108 34356
rect 17836 36428 17892 36484
rect 19404 42642 19460 42644
rect 19404 42590 19406 42642
rect 19406 42590 19458 42642
rect 19458 42590 19460 42642
rect 19404 42588 19460 42590
rect 19068 41916 19124 41972
rect 20076 43036 20132 43092
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 21420 43708 21476 43764
rect 20972 43596 21028 43652
rect 20748 43538 20804 43540
rect 20748 43486 20750 43538
rect 20750 43486 20802 43538
rect 20802 43486 20804 43538
rect 20748 43484 20804 43486
rect 20748 41970 20804 41972
rect 20748 41918 20750 41970
rect 20750 41918 20802 41970
rect 20802 41918 20804 41970
rect 20748 41916 20804 41918
rect 21308 42476 21364 42532
rect 19628 41468 19684 41524
rect 20188 41468 20244 41524
rect 19852 41074 19908 41076
rect 19852 41022 19854 41074
rect 19854 41022 19906 41074
rect 19906 41022 19908 41074
rect 19852 41020 19908 41022
rect 18732 40460 18788 40516
rect 19836 40794 19892 40796
rect 18844 40402 18900 40404
rect 18844 40350 18846 40402
rect 18846 40350 18898 40402
rect 18898 40350 18900 40402
rect 18844 40348 18900 40350
rect 19404 40684 19460 40740
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 18396 39618 18452 39620
rect 18396 39566 18398 39618
rect 18398 39566 18450 39618
rect 18450 39566 18452 39618
rect 18396 39564 18452 39566
rect 21420 42028 21476 42084
rect 21420 41244 21476 41300
rect 21196 40402 21252 40404
rect 21196 40350 21198 40402
rect 21198 40350 21250 40402
rect 21250 40350 21252 40402
rect 21196 40348 21252 40350
rect 21308 40572 21364 40628
rect 19068 39506 19124 39508
rect 19068 39454 19070 39506
rect 19070 39454 19122 39506
rect 19122 39454 19124 39506
rect 19068 39452 19124 39454
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 18732 38444 18788 38500
rect 18060 37548 18116 37604
rect 17948 36316 18004 36372
rect 18508 36428 18564 36484
rect 19964 38050 20020 38052
rect 19964 37998 19966 38050
rect 19966 37998 20018 38050
rect 20018 37998 20020 38050
rect 19964 37996 20020 37998
rect 19516 36540 19572 36596
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20860 37938 20916 37940
rect 20860 37886 20862 37938
rect 20862 37886 20914 37938
rect 20914 37886 20916 37938
rect 20860 37884 20916 37886
rect 20188 37324 20244 37380
rect 20524 37212 20580 37268
rect 21196 37996 21252 38052
rect 21420 38556 21476 38612
rect 21308 37826 21364 37828
rect 21308 37774 21310 37826
rect 21310 37774 21362 37826
rect 21362 37774 21364 37826
rect 21308 37772 21364 37774
rect 21756 44828 21812 44884
rect 22092 45276 22148 45332
rect 22540 48914 22596 48916
rect 22540 48862 22542 48914
rect 22542 48862 22594 48914
rect 22594 48862 22596 48914
rect 22540 48860 22596 48862
rect 23548 48748 23604 48804
rect 24668 49922 24724 49924
rect 24668 49870 24670 49922
rect 24670 49870 24722 49922
rect 24722 49870 24724 49922
rect 24668 49868 24724 49870
rect 24108 48188 24164 48244
rect 24332 48748 24388 48804
rect 24668 47740 24724 47796
rect 22764 45778 22820 45780
rect 22764 45726 22766 45778
rect 22766 45726 22818 45778
rect 22818 45726 22820 45778
rect 22764 45724 22820 45726
rect 22764 45388 22820 45444
rect 22652 44210 22708 44212
rect 22652 44158 22654 44210
rect 22654 44158 22706 44210
rect 22706 44158 22708 44210
rect 22652 44156 22708 44158
rect 23212 45052 23268 45108
rect 23884 46002 23940 46004
rect 23884 45950 23886 46002
rect 23886 45950 23938 46002
rect 23938 45950 23940 46002
rect 23884 45948 23940 45950
rect 24332 45724 24388 45780
rect 23660 45276 23716 45332
rect 23772 45500 23828 45556
rect 23548 44940 23604 44996
rect 23884 44940 23940 44996
rect 22316 43820 22372 43876
rect 22540 43314 22596 43316
rect 22540 43262 22542 43314
rect 22542 43262 22594 43314
rect 22594 43262 22596 43314
rect 22540 43260 22596 43262
rect 22316 42530 22372 42532
rect 22316 42478 22318 42530
rect 22318 42478 22370 42530
rect 22370 42478 22372 42530
rect 22316 42476 22372 42478
rect 24892 47964 24948 48020
rect 24892 47458 24948 47460
rect 24892 47406 24894 47458
rect 24894 47406 24946 47458
rect 24946 47406 24948 47458
rect 24892 47404 24948 47406
rect 24220 44380 24276 44436
rect 22764 42754 22820 42756
rect 22764 42702 22766 42754
rect 22766 42702 22818 42754
rect 22818 42702 22820 42754
rect 22764 42700 22820 42702
rect 22092 41298 22148 41300
rect 22092 41246 22094 41298
rect 22094 41246 22146 41298
rect 22146 41246 22148 41298
rect 22092 41244 22148 41246
rect 22428 41186 22484 41188
rect 22428 41134 22430 41186
rect 22430 41134 22482 41186
rect 22482 41134 22484 41186
rect 22428 41132 22484 41134
rect 21868 40796 21924 40852
rect 22204 40572 22260 40628
rect 21644 40348 21700 40404
rect 22540 40514 22596 40516
rect 22540 40462 22542 40514
rect 22542 40462 22594 40514
rect 22594 40462 22596 40514
rect 22540 40460 22596 40462
rect 22764 40962 22820 40964
rect 22764 40910 22766 40962
rect 22766 40910 22818 40962
rect 22818 40910 22820 40962
rect 22764 40908 22820 40910
rect 22764 40684 22820 40740
rect 21980 39228 22036 39284
rect 21756 38556 21812 38612
rect 21756 37884 21812 37940
rect 21420 37266 21476 37268
rect 21420 37214 21422 37266
rect 21422 37214 21474 37266
rect 21474 37214 21476 37266
rect 21420 37212 21476 37214
rect 21308 37100 21364 37156
rect 20636 36594 20692 36596
rect 20636 36542 20638 36594
rect 20638 36542 20690 36594
rect 20690 36542 20692 36594
rect 20636 36540 20692 36542
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 17612 34300 17668 34356
rect 18396 34354 18452 34356
rect 18396 34302 18398 34354
rect 18398 34302 18450 34354
rect 18450 34302 18452 34354
rect 18396 34300 18452 34302
rect 17948 34076 18004 34132
rect 17724 34018 17780 34020
rect 17724 33966 17726 34018
rect 17726 33966 17778 34018
rect 17778 33966 17780 34018
rect 17724 33964 17780 33966
rect 18508 34018 18564 34020
rect 18508 33966 18510 34018
rect 18510 33966 18562 34018
rect 18562 33966 18564 34018
rect 18508 33964 18564 33966
rect 18284 33628 18340 33684
rect 18508 33740 18564 33796
rect 17612 33068 17668 33124
rect 17276 32956 17332 33012
rect 16940 31388 16996 31444
rect 17164 31612 17220 31668
rect 17164 31164 17220 31220
rect 17388 31666 17444 31668
rect 17388 31614 17390 31666
rect 17390 31614 17442 31666
rect 17442 31614 17444 31666
rect 17388 31612 17444 31614
rect 16492 30492 16548 30548
rect 15932 27356 15988 27412
rect 15484 25618 15540 25620
rect 15484 25566 15486 25618
rect 15486 25566 15538 25618
rect 15538 25566 15540 25618
rect 15484 25564 15540 25566
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 21644 37324 21700 37380
rect 21644 34802 21700 34804
rect 21644 34750 21646 34802
rect 21646 34750 21698 34802
rect 21698 34750 21700 34802
rect 21644 34748 21700 34750
rect 18844 33516 18900 33572
rect 19068 33628 19124 33684
rect 18620 32732 18676 32788
rect 17724 31276 17780 31332
rect 17724 30994 17780 30996
rect 17724 30942 17726 30994
rect 17726 30942 17778 30994
rect 17778 30942 17780 30994
rect 17724 30940 17780 30942
rect 17164 30492 17220 30548
rect 16940 30210 16996 30212
rect 16940 30158 16942 30210
rect 16942 30158 16994 30210
rect 16994 30158 16996 30210
rect 16940 30156 16996 30158
rect 17388 30380 17444 30436
rect 18060 30492 18116 30548
rect 17836 30210 17892 30212
rect 17836 30158 17838 30210
rect 17838 30158 17890 30210
rect 17890 30158 17892 30210
rect 17836 30156 17892 30158
rect 18732 31666 18788 31668
rect 18732 31614 18734 31666
rect 18734 31614 18786 31666
rect 18786 31614 18788 31666
rect 18732 31612 18788 31614
rect 20300 33458 20356 33460
rect 20300 33406 20302 33458
rect 20302 33406 20354 33458
rect 20354 33406 20356 33458
rect 20300 33404 20356 33406
rect 19516 33292 19572 33348
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19740 32732 19796 32788
rect 18844 31218 18900 31220
rect 18844 31166 18846 31218
rect 18846 31166 18898 31218
rect 18898 31166 18900 31218
rect 18844 31164 18900 31166
rect 18620 30940 18676 30996
rect 19068 30940 19124 30996
rect 17724 30044 17780 30100
rect 17612 29986 17668 29988
rect 17612 29934 17614 29986
rect 17614 29934 17666 29986
rect 17666 29934 17668 29986
rect 17612 29932 17668 29934
rect 17836 29202 17892 29204
rect 17836 29150 17838 29202
rect 17838 29150 17890 29202
rect 17890 29150 17892 29202
rect 17836 29148 17892 29150
rect 18732 30492 18788 30548
rect 18956 30156 19012 30212
rect 19180 30716 19236 30772
rect 20524 31666 20580 31668
rect 20524 31614 20526 31666
rect 20526 31614 20578 31666
rect 20578 31614 20580 31666
rect 20524 31612 20580 31614
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20300 31218 20356 31220
rect 20300 31166 20302 31218
rect 20302 31166 20354 31218
rect 20354 31166 20356 31218
rect 20300 31164 20356 31166
rect 19628 30940 19684 30996
rect 19852 30994 19908 30996
rect 19852 30942 19854 30994
rect 19854 30942 19906 30994
rect 19906 30942 19908 30994
rect 19852 30940 19908 30942
rect 16716 26290 16772 26292
rect 16716 26238 16718 26290
rect 16718 26238 16770 26290
rect 16770 26238 16772 26290
rect 16716 26236 16772 26238
rect 15596 25116 15652 25172
rect 16492 23996 16548 24052
rect 16604 24834 16660 24836
rect 16604 24782 16606 24834
rect 16606 24782 16658 24834
rect 16658 24782 16660 24834
rect 16604 24780 16660 24782
rect 16492 23266 16548 23268
rect 16492 23214 16494 23266
rect 16494 23214 16546 23266
rect 16546 23214 16548 23266
rect 16492 23212 16548 23214
rect 15932 21362 15988 21364
rect 15932 21310 15934 21362
rect 15934 21310 15986 21362
rect 15986 21310 15988 21362
rect 15932 21308 15988 21310
rect 16156 21868 16212 21924
rect 16828 23378 16884 23380
rect 16828 23326 16830 23378
rect 16830 23326 16882 23378
rect 16882 23326 16884 23378
rect 16828 23324 16884 23326
rect 16604 21756 16660 21812
rect 16716 21698 16772 21700
rect 16716 21646 16718 21698
rect 16718 21646 16770 21698
rect 16770 21646 16772 21698
rect 16716 21644 16772 21646
rect 16604 21196 16660 21252
rect 14812 19964 14868 20020
rect 15036 20076 15092 20132
rect 14364 19794 14420 19796
rect 14364 19742 14366 19794
rect 14366 19742 14418 19794
rect 14418 19742 14420 19794
rect 14364 19740 14420 19742
rect 13692 19122 13748 19124
rect 13692 19070 13694 19122
rect 13694 19070 13746 19122
rect 13746 19070 13748 19122
rect 13692 19068 13748 19070
rect 13804 18508 13860 18564
rect 13916 18172 13972 18228
rect 12572 14588 12628 14644
rect 13020 13970 13076 13972
rect 13020 13918 13022 13970
rect 13022 13918 13074 13970
rect 13074 13918 13076 13970
rect 13020 13916 13076 13918
rect 12572 13132 12628 13188
rect 11788 12124 11844 12180
rect 9548 10780 9604 10836
rect 10220 10780 10276 10836
rect 9660 10722 9716 10724
rect 9660 10670 9662 10722
rect 9662 10670 9714 10722
rect 9714 10670 9716 10722
rect 9660 10668 9716 10670
rect 9548 10610 9604 10612
rect 9548 10558 9550 10610
rect 9550 10558 9602 10610
rect 9602 10558 9604 10610
rect 9548 10556 9604 10558
rect 8428 9324 8484 9380
rect 10444 10332 10500 10388
rect 9772 9266 9828 9268
rect 9772 9214 9774 9266
rect 9774 9214 9826 9266
rect 9826 9214 9828 9266
rect 9772 9212 9828 9214
rect 8092 8876 8148 8932
rect 7308 8316 7364 8372
rect 7980 8316 8036 8372
rect 9660 8930 9716 8932
rect 9660 8878 9662 8930
rect 9662 8878 9714 8930
rect 9714 8878 9716 8930
rect 9660 8876 9716 8878
rect 9772 8428 9828 8484
rect 8764 8316 8820 8372
rect 8988 7698 9044 7700
rect 8988 7646 8990 7698
rect 8990 7646 9042 7698
rect 9042 7646 9044 7698
rect 8988 7644 9044 7646
rect 11900 11170 11956 11172
rect 11900 11118 11902 11170
rect 11902 11118 11954 11170
rect 11954 11118 11956 11170
rect 11900 11116 11956 11118
rect 11564 10780 11620 10836
rect 12348 11788 12404 11844
rect 12236 11394 12292 11396
rect 12236 11342 12238 11394
rect 12238 11342 12290 11394
rect 12290 11342 12292 11394
rect 12236 11340 12292 11342
rect 12124 10892 12180 10948
rect 9884 8204 9940 8260
rect 10780 8316 10836 8372
rect 11788 9826 11844 9828
rect 11788 9774 11790 9826
rect 11790 9774 11842 9826
rect 11842 9774 11844 9826
rect 11788 9772 11844 9774
rect 12460 11004 12516 11060
rect 12460 10332 12516 10388
rect 12572 10892 12628 10948
rect 13692 17778 13748 17780
rect 13692 17726 13694 17778
rect 13694 17726 13746 17778
rect 13746 17726 13748 17778
rect 13692 17724 13748 17726
rect 13916 17500 13972 17556
rect 13692 15986 13748 15988
rect 13692 15934 13694 15986
rect 13694 15934 13746 15986
rect 13746 15934 13748 15986
rect 13692 15932 13748 15934
rect 14028 16604 14084 16660
rect 13580 13244 13636 13300
rect 13468 13186 13524 13188
rect 13468 13134 13470 13186
rect 13470 13134 13522 13186
rect 13522 13134 13524 13186
rect 13468 13132 13524 13134
rect 14476 19122 14532 19124
rect 14476 19070 14478 19122
rect 14478 19070 14530 19122
rect 14530 19070 14532 19122
rect 14476 19068 14532 19070
rect 15372 19964 15428 20020
rect 15036 18674 15092 18676
rect 15036 18622 15038 18674
rect 15038 18622 15090 18674
rect 15090 18622 15092 18674
rect 15036 18620 15092 18622
rect 15484 18844 15540 18900
rect 16156 20300 16212 20356
rect 16044 19234 16100 19236
rect 16044 19182 16046 19234
rect 16046 19182 16098 19234
rect 16098 19182 16100 19234
rect 16044 19180 16100 19182
rect 15708 19122 15764 19124
rect 15708 19070 15710 19122
rect 15710 19070 15762 19122
rect 15762 19070 15764 19122
rect 15708 19068 15764 19070
rect 15596 18732 15652 18788
rect 16156 18844 16212 18900
rect 15484 18508 15540 18564
rect 15820 18508 15876 18564
rect 15260 18396 15316 18452
rect 15036 18226 15092 18228
rect 15036 18174 15038 18226
rect 15038 18174 15090 18226
rect 15090 18174 15092 18226
rect 15036 18172 15092 18174
rect 15932 18396 15988 18452
rect 16156 17948 16212 18004
rect 14476 17500 14532 17556
rect 16492 19068 16548 19124
rect 16604 18620 16660 18676
rect 19292 30044 19348 30100
rect 18620 29148 18676 29204
rect 18508 28700 18564 28756
rect 19516 29986 19572 29988
rect 19516 29934 19518 29986
rect 19518 29934 19570 29986
rect 19570 29934 19572 29986
rect 19516 29932 19572 29934
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19292 28754 19348 28756
rect 19292 28702 19294 28754
rect 19294 28702 19346 28754
rect 19346 28702 19348 28754
rect 19292 28700 19348 28702
rect 19068 28028 19124 28084
rect 17836 27804 17892 27860
rect 18284 27858 18340 27860
rect 18284 27806 18286 27858
rect 18286 27806 18338 27858
rect 18338 27806 18340 27858
rect 18284 27804 18340 27806
rect 17500 26460 17556 26516
rect 17612 27692 17668 27748
rect 17500 26290 17556 26292
rect 17500 26238 17502 26290
rect 17502 26238 17554 26290
rect 17554 26238 17556 26290
rect 17500 26236 17556 26238
rect 18172 27746 18228 27748
rect 18172 27694 18174 27746
rect 18174 27694 18226 27746
rect 18226 27694 18228 27746
rect 18172 27692 18228 27694
rect 18284 27468 18340 27524
rect 18060 26460 18116 26516
rect 18732 27132 18788 27188
rect 18508 26684 18564 26740
rect 18956 27132 19012 27188
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19628 28028 19684 28084
rect 20076 27746 20132 27748
rect 20076 27694 20078 27746
rect 20078 27694 20130 27746
rect 20130 27694 20132 27746
rect 20076 27692 20132 27694
rect 19852 27244 19908 27300
rect 19628 27020 19684 27076
rect 18956 26684 19012 26740
rect 18396 25618 18452 25620
rect 18396 25566 18398 25618
rect 18398 25566 18450 25618
rect 18450 25566 18452 25618
rect 18396 25564 18452 25566
rect 17612 25452 17668 25508
rect 17388 23378 17444 23380
rect 17388 23326 17390 23378
rect 17390 23326 17442 23378
rect 17442 23326 17444 23378
rect 17388 23324 17444 23326
rect 20412 27074 20468 27076
rect 20412 27022 20414 27074
rect 20414 27022 20466 27074
rect 20466 27022 20468 27074
rect 20412 27020 20468 27022
rect 20188 26908 20244 26964
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20972 34188 21028 34244
rect 20860 32786 20916 32788
rect 20860 32734 20862 32786
rect 20862 32734 20914 32786
rect 20914 32734 20916 32786
rect 20860 32732 20916 32734
rect 21868 37266 21924 37268
rect 21868 37214 21870 37266
rect 21870 37214 21922 37266
rect 21922 37214 21924 37266
rect 21868 37212 21924 37214
rect 21756 33740 21812 33796
rect 21084 33404 21140 33460
rect 21868 33404 21924 33460
rect 21532 31388 21588 31444
rect 21868 30994 21924 30996
rect 21868 30942 21870 30994
rect 21870 30942 21922 30994
rect 21922 30942 21924 30994
rect 21868 30940 21924 30942
rect 22428 38892 22484 38948
rect 22764 38892 22820 38948
rect 22316 37884 22372 37940
rect 23100 42700 23156 42756
rect 22988 42530 23044 42532
rect 22988 42478 22990 42530
rect 22990 42478 23042 42530
rect 23042 42478 23044 42530
rect 22988 42476 23044 42478
rect 22988 41804 23044 41860
rect 23996 43538 24052 43540
rect 23996 43486 23998 43538
rect 23998 43486 24050 43538
rect 24050 43486 24052 43538
rect 23996 43484 24052 43486
rect 23436 42700 23492 42756
rect 23996 43036 24052 43092
rect 23884 42754 23940 42756
rect 23884 42702 23886 42754
rect 23886 42702 23938 42754
rect 23938 42702 23940 42754
rect 23884 42700 23940 42702
rect 23772 42642 23828 42644
rect 23772 42590 23774 42642
rect 23774 42590 23826 42642
rect 23826 42590 23828 42642
rect 23772 42588 23828 42590
rect 24332 42812 24388 42868
rect 24220 42476 24276 42532
rect 23660 41916 23716 41972
rect 23100 41132 23156 41188
rect 24108 41916 24164 41972
rect 23996 41244 24052 41300
rect 23212 41020 23268 41076
rect 23436 40460 23492 40516
rect 23212 40236 23268 40292
rect 25676 54738 25732 54740
rect 25676 54686 25678 54738
rect 25678 54686 25730 54738
rect 25730 54686 25732 54738
rect 25676 54684 25732 54686
rect 25340 53564 25396 53620
rect 25116 52556 25172 52612
rect 25228 53228 25284 53284
rect 25676 53058 25732 53060
rect 25676 53006 25678 53058
rect 25678 53006 25730 53058
rect 25730 53006 25732 53058
rect 25676 53004 25732 53006
rect 25228 52332 25284 52388
rect 25452 52668 25508 52724
rect 25900 53452 25956 53508
rect 26796 55356 26852 55412
rect 27020 53676 27076 53732
rect 26684 53452 26740 53508
rect 26572 52668 26628 52724
rect 26908 53116 26964 53172
rect 26348 52556 26404 52612
rect 25788 52332 25844 52388
rect 26796 52386 26852 52388
rect 26796 52334 26798 52386
rect 26798 52334 26850 52386
rect 26850 52334 26852 52386
rect 26796 52332 26852 52334
rect 25340 52220 25396 52276
rect 25452 52108 25508 52164
rect 25452 50204 25508 50260
rect 25452 49756 25508 49812
rect 25228 49698 25284 49700
rect 25228 49646 25230 49698
rect 25230 49646 25282 49698
rect 25282 49646 25284 49698
rect 25228 49644 25284 49646
rect 25452 48466 25508 48468
rect 25452 48414 25454 48466
rect 25454 48414 25506 48466
rect 25506 48414 25508 48466
rect 25452 48412 25508 48414
rect 26236 52162 26292 52164
rect 26236 52110 26238 52162
rect 26238 52110 26290 52162
rect 26290 52110 26292 52162
rect 26236 52108 26292 52110
rect 25676 51996 25732 52052
rect 26908 51996 26964 52052
rect 27020 52108 27076 52164
rect 26796 51212 26852 51268
rect 26572 49922 26628 49924
rect 26572 49870 26574 49922
rect 26574 49870 26626 49922
rect 26626 49870 26628 49922
rect 26572 49868 26628 49870
rect 26124 49810 26180 49812
rect 26124 49758 26126 49810
rect 26126 49758 26178 49810
rect 26178 49758 26180 49810
rect 26124 49756 26180 49758
rect 26796 50092 26852 50148
rect 25788 49084 25844 49140
rect 25004 44604 25060 44660
rect 25116 48188 25172 48244
rect 25004 44434 25060 44436
rect 25004 44382 25006 44434
rect 25006 44382 25058 44434
rect 25058 44382 25060 44434
rect 25004 44380 25060 44382
rect 25564 48076 25620 48132
rect 25340 47852 25396 47908
rect 25564 47740 25620 47796
rect 25676 47404 25732 47460
rect 25340 46844 25396 46900
rect 25340 45500 25396 45556
rect 25340 45330 25396 45332
rect 25340 45278 25342 45330
rect 25342 45278 25394 45330
rect 25394 45278 25396 45330
rect 25340 45276 25396 45278
rect 24556 43596 24612 43652
rect 26572 47852 26628 47908
rect 26460 47404 26516 47460
rect 26236 47180 26292 47236
rect 26348 46956 26404 47012
rect 26796 48412 26852 48468
rect 27020 49138 27076 49140
rect 27020 49086 27022 49138
rect 27022 49086 27074 49138
rect 27074 49086 27076 49138
rect 27020 49084 27076 49086
rect 26908 48188 26964 48244
rect 29484 56082 29540 56084
rect 29484 56030 29486 56082
rect 29486 56030 29538 56082
rect 29538 56030 29540 56082
rect 29484 56028 29540 56030
rect 27580 55244 27636 55300
rect 28476 55186 28532 55188
rect 28476 55134 28478 55186
rect 28478 55134 28530 55186
rect 28530 55134 28532 55186
rect 28476 55132 28532 55134
rect 29260 55132 29316 55188
rect 27804 53618 27860 53620
rect 27804 53566 27806 53618
rect 27806 53566 27858 53618
rect 27858 53566 27860 53618
rect 27804 53564 27860 53566
rect 27916 53506 27972 53508
rect 27916 53454 27918 53506
rect 27918 53454 27970 53506
rect 27970 53454 27972 53506
rect 27916 53452 27972 53454
rect 28364 53730 28420 53732
rect 28364 53678 28366 53730
rect 28366 53678 28418 53730
rect 28418 53678 28420 53730
rect 28364 53676 28420 53678
rect 29372 53730 29428 53732
rect 29372 53678 29374 53730
rect 29374 53678 29426 53730
rect 29426 53678 29428 53730
rect 29372 53676 29428 53678
rect 29148 53564 29204 53620
rect 29596 55356 29652 55412
rect 29820 54236 29876 54292
rect 29484 53564 29540 53620
rect 28140 53228 28196 53284
rect 29596 53228 29652 53284
rect 28028 53116 28084 53172
rect 29596 52780 29652 52836
rect 29708 53452 29764 53508
rect 30156 53170 30212 53172
rect 30156 53118 30158 53170
rect 30158 53118 30210 53170
rect 30210 53118 30212 53170
rect 30156 53116 30212 53118
rect 29260 52668 29316 52724
rect 28812 52444 28868 52500
rect 28364 51436 28420 51492
rect 27580 50706 27636 50708
rect 27580 50654 27582 50706
rect 27582 50654 27634 50706
rect 27634 50654 27636 50706
rect 27580 50652 27636 50654
rect 28588 51266 28644 51268
rect 28588 51214 28590 51266
rect 28590 51214 28642 51266
rect 28642 51214 28644 51266
rect 28588 51212 28644 51214
rect 28364 50540 28420 50596
rect 28476 50482 28532 50484
rect 28476 50430 28478 50482
rect 28478 50430 28530 50482
rect 28530 50430 28532 50482
rect 28476 50428 28532 50430
rect 27244 50204 27300 50260
rect 27356 50092 27412 50148
rect 27580 49922 27636 49924
rect 27580 49870 27582 49922
rect 27582 49870 27634 49922
rect 27634 49870 27636 49922
rect 27580 49868 27636 49870
rect 27468 49698 27524 49700
rect 27468 49646 27470 49698
rect 27470 49646 27522 49698
rect 27522 49646 27524 49698
rect 27468 49644 27524 49646
rect 29148 51602 29204 51604
rect 29148 51550 29150 51602
rect 29150 51550 29202 51602
rect 29202 51550 29204 51602
rect 29148 51548 29204 51550
rect 29484 52556 29540 52612
rect 29372 52444 29428 52500
rect 29260 49980 29316 50036
rect 28812 49810 28868 49812
rect 28812 49758 28814 49810
rect 28814 49758 28866 49810
rect 28866 49758 28868 49810
rect 28812 49756 28868 49758
rect 29708 52220 29764 52276
rect 30604 56028 30660 56084
rect 30492 53676 30548 53732
rect 31612 56252 31668 56308
rect 30492 53004 30548 53060
rect 30716 53228 30772 53284
rect 30268 52332 30324 52388
rect 30492 52220 30548 52276
rect 30044 52050 30100 52052
rect 30044 51998 30046 52050
rect 30046 51998 30098 52050
rect 30098 51998 30100 52050
rect 30044 51996 30100 51998
rect 29708 51548 29764 51604
rect 30716 50540 30772 50596
rect 29932 50482 29988 50484
rect 29932 50430 29934 50482
rect 29934 50430 29986 50482
rect 29986 50430 29988 50482
rect 29932 50428 29988 50430
rect 29484 49922 29540 49924
rect 29484 49870 29486 49922
rect 29486 49870 29538 49922
rect 29538 49870 29540 49922
rect 29484 49868 29540 49870
rect 28588 49084 28644 49140
rect 27580 48076 27636 48132
rect 27804 48076 27860 48132
rect 26908 47964 26964 48020
rect 25228 45164 25284 45220
rect 24556 43372 24612 43428
rect 24556 42754 24612 42756
rect 24556 42702 24558 42754
rect 24558 42702 24610 42754
rect 24610 42702 24612 42754
rect 24556 42700 24612 42702
rect 24780 42530 24836 42532
rect 24780 42478 24782 42530
rect 24782 42478 24834 42530
rect 24834 42478 24836 42530
rect 24780 42476 24836 42478
rect 24668 41858 24724 41860
rect 24668 41806 24670 41858
rect 24670 41806 24722 41858
rect 24722 41806 24724 41858
rect 24668 41804 24724 41806
rect 24108 41020 24164 41076
rect 23996 40348 24052 40404
rect 23772 39900 23828 39956
rect 24108 40124 24164 40180
rect 23772 38162 23828 38164
rect 23772 38110 23774 38162
rect 23774 38110 23826 38162
rect 23826 38110 23828 38162
rect 23772 38108 23828 38110
rect 22316 37266 22372 37268
rect 22316 37214 22318 37266
rect 22318 37214 22370 37266
rect 22370 37214 22372 37266
rect 22316 37212 22372 37214
rect 23100 37100 23156 37156
rect 23548 37212 23604 37268
rect 22988 36204 23044 36260
rect 22652 35308 22708 35364
rect 23324 36092 23380 36148
rect 23436 35532 23492 35588
rect 25116 42754 25172 42756
rect 25116 42702 25118 42754
rect 25118 42702 25170 42754
rect 25170 42702 25172 42754
rect 25116 42700 25172 42702
rect 24892 41356 24948 41412
rect 24332 41186 24388 41188
rect 24332 41134 24334 41186
rect 24334 41134 24386 41186
rect 24386 41134 24388 41186
rect 24332 41132 24388 41134
rect 24444 41020 24500 41076
rect 25004 41074 25060 41076
rect 25004 41022 25006 41074
rect 25006 41022 25058 41074
rect 25058 41022 25060 41074
rect 25004 41020 25060 41022
rect 24556 40908 24612 40964
rect 24332 40012 24388 40068
rect 24444 40572 24500 40628
rect 24332 39340 24388 39396
rect 26460 46002 26516 46004
rect 26460 45950 26462 46002
rect 26462 45950 26514 46002
rect 26514 45950 26516 46002
rect 26460 45948 26516 45950
rect 25564 44492 25620 44548
rect 26236 45052 26292 45108
rect 27020 47404 27076 47460
rect 27692 47234 27748 47236
rect 27692 47182 27694 47234
rect 27694 47182 27746 47234
rect 27746 47182 27748 47234
rect 27692 47180 27748 47182
rect 27916 47234 27972 47236
rect 27916 47182 27918 47234
rect 27918 47182 27970 47234
rect 27970 47182 27972 47234
rect 27916 47180 27972 47182
rect 27804 47068 27860 47124
rect 27580 46674 27636 46676
rect 27580 46622 27582 46674
rect 27582 46622 27634 46674
rect 27634 46622 27636 46674
rect 27580 46620 27636 46622
rect 26460 44828 26516 44884
rect 25900 44546 25956 44548
rect 25900 44494 25902 44546
rect 25902 44494 25954 44546
rect 25954 44494 25956 44546
rect 25900 44492 25956 44494
rect 25900 44268 25956 44324
rect 25676 43596 25732 43652
rect 25788 42924 25844 42980
rect 25676 42812 25732 42868
rect 26124 44492 26180 44548
rect 27132 45164 27188 45220
rect 27020 45052 27076 45108
rect 26796 44492 26852 44548
rect 27132 44322 27188 44324
rect 27132 44270 27134 44322
rect 27134 44270 27186 44322
rect 27186 44270 27188 44322
rect 27132 44268 27188 44270
rect 27468 43762 27524 43764
rect 27468 43710 27470 43762
rect 27470 43710 27522 43762
rect 27522 43710 27524 43762
rect 27468 43708 27524 43710
rect 26572 43596 26628 43652
rect 27020 43650 27076 43652
rect 27020 43598 27022 43650
rect 27022 43598 27074 43650
rect 27074 43598 27076 43650
rect 27020 43596 27076 43598
rect 26460 43426 26516 43428
rect 26460 43374 26462 43426
rect 26462 43374 26514 43426
rect 26514 43374 26516 43426
rect 26460 43372 26516 43374
rect 27132 43426 27188 43428
rect 27132 43374 27134 43426
rect 27134 43374 27186 43426
rect 27186 43374 27188 43426
rect 27132 43372 27188 43374
rect 26572 43314 26628 43316
rect 26572 43262 26574 43314
rect 26574 43262 26626 43314
rect 26626 43262 26628 43314
rect 26572 43260 26628 43262
rect 25340 42642 25396 42644
rect 25340 42590 25342 42642
rect 25342 42590 25394 42642
rect 25394 42590 25396 42642
rect 25340 42588 25396 42590
rect 25228 40572 25284 40628
rect 24780 40460 24836 40516
rect 25228 40348 25284 40404
rect 24332 36092 24388 36148
rect 24108 35922 24164 35924
rect 24108 35870 24110 35922
rect 24110 35870 24162 35922
rect 24162 35870 24164 35922
rect 24108 35868 24164 35870
rect 23660 35698 23716 35700
rect 23660 35646 23662 35698
rect 23662 35646 23714 35698
rect 23714 35646 23716 35698
rect 23660 35644 23716 35646
rect 23548 35196 23604 35252
rect 23212 34914 23268 34916
rect 23212 34862 23214 34914
rect 23214 34862 23266 34914
rect 23266 34862 23268 34914
rect 23212 34860 23268 34862
rect 22428 34690 22484 34692
rect 22428 34638 22430 34690
rect 22430 34638 22482 34690
rect 22482 34638 22484 34690
rect 22428 34636 22484 34638
rect 22876 34748 22932 34804
rect 23212 34636 23268 34692
rect 22764 33740 22820 33796
rect 22988 33346 23044 33348
rect 22988 33294 22990 33346
rect 22990 33294 23042 33346
rect 23042 33294 23044 33346
rect 22988 33292 23044 33294
rect 22540 33234 22596 33236
rect 22540 33182 22542 33234
rect 22542 33182 22594 33234
rect 22594 33182 22596 33234
rect 22540 33180 22596 33182
rect 22540 32732 22596 32788
rect 23212 32060 23268 32116
rect 22876 31612 22932 31668
rect 22316 31164 22372 31220
rect 22540 31276 22596 31332
rect 21532 30380 21588 30436
rect 21756 30492 21812 30548
rect 21644 29596 21700 29652
rect 20636 25900 20692 25956
rect 21644 27858 21700 27860
rect 21644 27806 21646 27858
rect 21646 27806 21698 27858
rect 21698 27806 21700 27858
rect 21644 27804 21700 27806
rect 21084 26908 21140 26964
rect 19404 25452 19460 25508
rect 17948 25282 18004 25284
rect 17948 25230 17950 25282
rect 17950 25230 18002 25282
rect 18002 25230 18004 25282
rect 17948 25228 18004 25230
rect 19292 25228 19348 25284
rect 18732 25004 18788 25060
rect 19068 24780 19124 24836
rect 17724 24050 17780 24052
rect 17724 23998 17726 24050
rect 17726 23998 17778 24050
rect 17778 23998 17780 24050
rect 17724 23996 17780 23998
rect 17500 21868 17556 21924
rect 17612 21810 17668 21812
rect 17612 21758 17614 21810
rect 17614 21758 17666 21810
rect 17666 21758 17668 21810
rect 17612 21756 17668 21758
rect 17500 21698 17556 21700
rect 17500 21646 17502 21698
rect 17502 21646 17554 21698
rect 17554 21646 17556 21698
rect 17500 21644 17556 21646
rect 17388 21586 17444 21588
rect 17388 21534 17390 21586
rect 17390 21534 17442 21586
rect 17442 21534 17444 21586
rect 17388 21532 17444 21534
rect 18956 24108 19012 24164
rect 18060 23324 18116 23380
rect 17948 22482 18004 22484
rect 17948 22430 17950 22482
rect 17950 22430 18002 22482
rect 18002 22430 18004 22482
rect 17948 22428 18004 22430
rect 20300 25506 20356 25508
rect 20300 25454 20302 25506
rect 20302 25454 20354 25506
rect 20354 25454 20356 25506
rect 20300 25452 20356 25454
rect 19404 25004 19460 25060
rect 19516 25340 19572 25396
rect 19068 23772 19124 23828
rect 18284 21980 18340 22036
rect 17724 20748 17780 20804
rect 18172 21308 18228 21364
rect 17276 19122 17332 19124
rect 17276 19070 17278 19122
rect 17278 19070 17330 19122
rect 17330 19070 17332 19122
rect 17276 19068 17332 19070
rect 16940 18508 16996 18564
rect 18732 22258 18788 22260
rect 18732 22206 18734 22258
rect 18734 22206 18786 22258
rect 18786 22206 18788 22258
rect 18732 22204 18788 22206
rect 18844 21532 18900 21588
rect 18956 22988 19012 23044
rect 19852 25282 19908 25284
rect 19852 25230 19854 25282
rect 19854 25230 19906 25282
rect 19906 25230 19908 25282
rect 19852 25228 19908 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20300 24332 20356 24388
rect 19964 24050 20020 24052
rect 19964 23998 19966 24050
rect 19966 23998 20018 24050
rect 20018 23998 20020 24050
rect 19964 23996 20020 23998
rect 19180 22428 19236 22484
rect 19180 21756 19236 21812
rect 18508 21196 18564 21252
rect 18508 20802 18564 20804
rect 18508 20750 18510 20802
rect 18510 20750 18562 20802
rect 18562 20750 18564 20802
rect 18508 20748 18564 20750
rect 15596 17442 15652 17444
rect 15596 17390 15598 17442
rect 15598 17390 15650 17442
rect 15650 17390 15652 17442
rect 15596 17388 15652 17390
rect 14028 15596 14084 15652
rect 14364 16156 14420 16212
rect 13804 15314 13860 15316
rect 13804 15262 13806 15314
rect 13806 15262 13858 15314
rect 13858 15262 13860 15314
rect 13804 15260 13860 15262
rect 13916 14530 13972 14532
rect 13916 14478 13918 14530
rect 13918 14478 13970 14530
rect 13970 14478 13972 14530
rect 13916 14476 13972 14478
rect 13804 13746 13860 13748
rect 13804 13694 13806 13746
rect 13806 13694 13858 13746
rect 13858 13694 13860 13746
rect 13804 13692 13860 13694
rect 13916 13244 13972 13300
rect 13692 12738 13748 12740
rect 13692 12686 13694 12738
rect 13694 12686 13746 12738
rect 13746 12686 13748 12738
rect 13692 12684 13748 12686
rect 13580 12460 13636 12516
rect 13132 12402 13188 12404
rect 13132 12350 13134 12402
rect 13134 12350 13186 12402
rect 13186 12350 13188 12402
rect 13132 12348 13188 12350
rect 13020 12236 13076 12292
rect 13692 12236 13748 12292
rect 13244 12178 13300 12180
rect 13244 12126 13246 12178
rect 13246 12126 13298 12178
rect 13298 12126 13300 12178
rect 13244 12124 13300 12126
rect 12908 11564 12964 11620
rect 13020 11900 13076 11956
rect 12796 11452 12852 11508
rect 12796 10668 12852 10724
rect 13580 11788 13636 11844
rect 13244 10834 13300 10836
rect 13244 10782 13246 10834
rect 13246 10782 13298 10834
rect 13298 10782 13300 10834
rect 13244 10780 13300 10782
rect 13020 9436 13076 9492
rect 11228 8428 11284 8484
rect 10220 8092 10276 8148
rect 10668 8146 10724 8148
rect 10668 8094 10670 8146
rect 10670 8094 10722 8146
rect 10722 8094 10724 8146
rect 10668 8092 10724 8094
rect 9772 7644 9828 7700
rect 10556 7980 10612 8036
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 12236 8258 12292 8260
rect 12236 8206 12238 8258
rect 12238 8206 12290 8258
rect 12290 8206 12292 8258
rect 12236 8204 12292 8206
rect 12684 8428 12740 8484
rect 12124 8034 12180 8036
rect 12124 7982 12126 8034
rect 12126 7982 12178 8034
rect 12178 7982 12180 8034
rect 12124 7980 12180 7982
rect 12572 7980 12628 8036
rect 13916 11676 13972 11732
rect 14364 15314 14420 15316
rect 14364 15262 14366 15314
rect 14366 15262 14418 15314
rect 14418 15262 14420 15314
rect 14364 15260 14420 15262
rect 14700 16940 14756 16996
rect 15036 16994 15092 16996
rect 15036 16942 15038 16994
rect 15038 16942 15090 16994
rect 15090 16942 15092 16994
rect 15036 16940 15092 16942
rect 14812 16604 14868 16660
rect 15708 16604 15764 16660
rect 14700 15372 14756 15428
rect 15260 15596 15316 15652
rect 14140 12348 14196 12404
rect 15596 15036 15652 15092
rect 14812 14530 14868 14532
rect 14812 14478 14814 14530
rect 14814 14478 14866 14530
rect 14866 14478 14868 14530
rect 14812 14476 14868 14478
rect 15036 13692 15092 13748
rect 14700 12684 14756 12740
rect 14700 12402 14756 12404
rect 14700 12350 14702 12402
rect 14702 12350 14754 12402
rect 14754 12350 14756 12402
rect 14700 12348 14756 12350
rect 15484 12348 15540 12404
rect 15372 11676 15428 11732
rect 14028 11394 14084 11396
rect 14028 11342 14030 11394
rect 14030 11342 14082 11394
rect 14082 11342 14084 11394
rect 14028 11340 14084 11342
rect 13804 10892 13860 10948
rect 14700 11116 14756 11172
rect 13916 10668 13972 10724
rect 13692 9660 13748 9716
rect 13804 10108 13860 10164
rect 13692 8258 13748 8260
rect 13692 8206 13694 8258
rect 13694 8206 13746 8258
rect 13746 8206 13748 8258
rect 13692 8204 13748 8206
rect 13580 8034 13636 8036
rect 13580 7982 13582 8034
rect 13582 7982 13634 8034
rect 13634 7982 13636 8034
rect 13580 7980 13636 7982
rect 16156 16492 16212 16548
rect 16156 15314 16212 15316
rect 16156 15262 16158 15314
rect 16158 15262 16210 15314
rect 16210 15262 16212 15314
rect 16156 15260 16212 15262
rect 16156 14924 16212 14980
rect 15708 10780 15764 10836
rect 16716 17442 16772 17444
rect 16716 17390 16718 17442
rect 16718 17390 16770 17442
rect 16770 17390 16772 17442
rect 16716 17388 16772 17390
rect 16716 16492 16772 16548
rect 17052 16268 17108 16324
rect 17164 17948 17220 18004
rect 17948 18396 18004 18452
rect 18844 20748 18900 20804
rect 19404 20802 19460 20804
rect 19404 20750 19406 20802
rect 19406 20750 19458 20802
rect 19458 20750 19460 20802
rect 19404 20748 19460 20750
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19852 23042 19908 23044
rect 19852 22990 19854 23042
rect 19854 22990 19906 23042
rect 19906 22990 19908 23042
rect 19852 22988 19908 22990
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19964 20802 20020 20804
rect 19964 20750 19966 20802
rect 19966 20750 20018 20802
rect 20018 20750 20020 20802
rect 19964 20748 20020 20750
rect 19628 20412 19684 20468
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 18620 19234 18676 19236
rect 18620 19182 18622 19234
rect 18622 19182 18674 19234
rect 18674 19182 18676 19234
rect 18620 19180 18676 19182
rect 19628 19180 19684 19236
rect 17388 17778 17444 17780
rect 17388 17726 17390 17778
rect 17390 17726 17442 17778
rect 17442 17726 17444 17778
rect 17388 17724 17444 17726
rect 18844 18508 18900 18564
rect 18284 17724 18340 17780
rect 19404 18732 19460 18788
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19292 18396 19348 18452
rect 19740 18172 19796 18228
rect 18956 17052 19012 17108
rect 19404 17052 19460 17108
rect 17276 16604 17332 16660
rect 18396 16268 18452 16324
rect 16604 15314 16660 15316
rect 16604 15262 16606 15314
rect 16606 15262 16658 15314
rect 16658 15262 16660 15314
rect 16604 15260 16660 15262
rect 16716 15202 16772 15204
rect 16716 15150 16718 15202
rect 16718 15150 16770 15202
rect 16770 15150 16772 15202
rect 16716 15148 16772 15150
rect 16380 15036 16436 15092
rect 16380 13580 16436 13636
rect 16492 13468 16548 13524
rect 17612 15202 17668 15204
rect 17612 15150 17614 15202
rect 17614 15150 17666 15202
rect 17666 15150 17668 15202
rect 17612 15148 17668 15150
rect 17052 14418 17108 14420
rect 17052 14366 17054 14418
rect 17054 14366 17106 14418
rect 17106 14366 17108 14418
rect 17052 14364 17108 14366
rect 16828 13916 16884 13972
rect 17948 15260 18004 15316
rect 18396 15148 18452 15204
rect 17276 13580 17332 13636
rect 16604 11788 16660 11844
rect 16604 11340 16660 11396
rect 16268 10332 16324 10388
rect 14812 10108 14868 10164
rect 16044 10108 16100 10164
rect 14476 9436 14532 9492
rect 15148 9660 15204 9716
rect 14588 8316 14644 8372
rect 17052 11564 17108 11620
rect 16940 11394 16996 11396
rect 16940 11342 16942 11394
rect 16942 11342 16994 11394
rect 16994 11342 16996 11394
rect 16940 11340 16996 11342
rect 16604 10610 16660 10612
rect 16604 10558 16606 10610
rect 16606 10558 16658 10610
rect 16658 10558 16660 10610
rect 16604 10556 16660 10558
rect 16380 9884 16436 9940
rect 17164 11170 17220 11172
rect 17164 11118 17166 11170
rect 17166 11118 17218 11170
rect 17218 11118 17220 11170
rect 17164 11116 17220 11118
rect 17052 10108 17108 10164
rect 16828 9938 16884 9940
rect 16828 9886 16830 9938
rect 16830 9886 16882 9938
rect 16882 9886 16884 9938
rect 16828 9884 16884 9886
rect 16716 9772 16772 9828
rect 16380 9324 16436 9380
rect 16268 9266 16324 9268
rect 16268 9214 16270 9266
rect 16270 9214 16322 9266
rect 16322 9214 16324 9266
rect 16268 9212 16324 9214
rect 17052 9212 17108 9268
rect 15932 8428 15988 8484
rect 16380 7474 16436 7476
rect 16380 7422 16382 7474
rect 16382 7422 16434 7474
rect 16434 7422 16436 7474
rect 16380 7420 16436 7422
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 17388 11788 17444 11844
rect 17836 13916 17892 13972
rect 18060 14364 18116 14420
rect 18508 14476 18564 14532
rect 18956 15148 19012 15204
rect 18396 14418 18452 14420
rect 18396 14366 18398 14418
rect 18398 14366 18450 14418
rect 18450 14366 18452 14418
rect 18396 14364 18452 14366
rect 18060 13580 18116 13636
rect 17612 13522 17668 13524
rect 17612 13470 17614 13522
rect 17614 13470 17666 13522
rect 17666 13470 17668 13522
rect 17612 13468 17668 13470
rect 17388 10556 17444 10612
rect 17724 11676 17780 11732
rect 18396 13634 18452 13636
rect 18396 13582 18398 13634
rect 18398 13582 18450 13634
rect 18450 13582 18452 13634
rect 18396 13580 18452 13582
rect 18844 14588 18900 14644
rect 18732 14530 18788 14532
rect 18732 14478 18734 14530
rect 18734 14478 18786 14530
rect 18786 14478 18788 14530
rect 18732 14476 18788 14478
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20076 17106 20132 17108
rect 20076 17054 20078 17106
rect 20078 17054 20130 17106
rect 20130 17054 20132 17106
rect 20076 17052 20132 17054
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19628 14588 19684 14644
rect 19740 15148 19796 15204
rect 19516 14476 19572 14532
rect 19404 14418 19460 14420
rect 19404 14366 19406 14418
rect 19406 14366 19458 14418
rect 19458 14366 19460 14418
rect 19404 14364 19460 14366
rect 18620 12236 18676 12292
rect 17724 9826 17780 9828
rect 17724 9774 17726 9826
rect 17726 9774 17778 9826
rect 17778 9774 17780 9826
rect 17724 9772 17780 9774
rect 17500 9714 17556 9716
rect 17500 9662 17502 9714
rect 17502 9662 17554 9714
rect 17554 9662 17556 9714
rect 17500 9660 17556 9662
rect 18172 9660 18228 9716
rect 18060 9100 18116 9156
rect 18396 10780 18452 10836
rect 18396 10556 18452 10612
rect 21420 27692 21476 27748
rect 21308 27074 21364 27076
rect 21308 27022 21310 27074
rect 21310 27022 21362 27074
rect 21362 27022 21364 27074
rect 21308 27020 21364 27022
rect 21532 26962 21588 26964
rect 21532 26910 21534 26962
rect 21534 26910 21586 26962
rect 21586 26910 21588 26962
rect 21532 26908 21588 26910
rect 21196 26460 21252 26516
rect 21308 25394 21364 25396
rect 21308 25342 21310 25394
rect 21310 25342 21362 25394
rect 21362 25342 21364 25394
rect 21308 25340 21364 25342
rect 20860 24332 20916 24388
rect 21532 23938 21588 23940
rect 21532 23886 21534 23938
rect 21534 23886 21586 23938
rect 21586 23886 21588 23938
rect 21532 23884 21588 23886
rect 21308 23772 21364 23828
rect 20636 22988 20692 23044
rect 20972 21980 21028 22036
rect 21196 21810 21252 21812
rect 21196 21758 21198 21810
rect 21198 21758 21250 21810
rect 21250 21758 21252 21810
rect 21196 21756 21252 21758
rect 21420 21698 21476 21700
rect 21420 21646 21422 21698
rect 21422 21646 21474 21698
rect 21474 21646 21476 21698
rect 21420 21644 21476 21646
rect 20860 20748 20916 20804
rect 20524 20300 20580 20356
rect 20748 20636 20804 20692
rect 22988 31164 23044 31220
rect 22316 30380 22372 30436
rect 22428 30268 22484 30324
rect 22876 30434 22932 30436
rect 22876 30382 22878 30434
rect 22878 30382 22930 30434
rect 22930 30382 22932 30434
rect 22876 30380 22932 30382
rect 23100 30940 23156 30996
rect 22428 29650 22484 29652
rect 22428 29598 22430 29650
rect 22430 29598 22482 29650
rect 22482 29598 22484 29650
rect 22428 29596 22484 29598
rect 22316 29484 22372 29540
rect 21980 29148 22036 29204
rect 22204 28754 22260 28756
rect 22204 28702 22206 28754
rect 22206 28702 22258 28754
rect 22258 28702 22260 28754
rect 22204 28700 22260 28702
rect 21980 28364 22036 28420
rect 25116 39228 25172 39284
rect 25340 40236 25396 40292
rect 25900 42476 25956 42532
rect 26236 42476 26292 42532
rect 27244 42700 27300 42756
rect 26572 42642 26628 42644
rect 26572 42590 26574 42642
rect 26574 42590 26626 42642
rect 26626 42590 26628 42642
rect 26572 42588 26628 42590
rect 26572 42364 26628 42420
rect 26684 42140 26740 42196
rect 25676 41356 25732 41412
rect 25788 40684 25844 40740
rect 27356 41858 27412 41860
rect 27356 41806 27358 41858
rect 27358 41806 27410 41858
rect 27410 41806 27412 41858
rect 27356 41804 27412 41806
rect 26684 40626 26740 40628
rect 26684 40574 26686 40626
rect 26686 40574 26738 40626
rect 26738 40574 26740 40626
rect 26684 40572 26740 40574
rect 27020 41020 27076 41076
rect 25116 38444 25172 38500
rect 25788 38834 25844 38836
rect 25788 38782 25790 38834
rect 25790 38782 25842 38834
rect 25842 38782 25844 38834
rect 25788 38780 25844 38782
rect 25676 38108 25732 38164
rect 24780 36764 24836 36820
rect 24780 36316 24836 36372
rect 24668 35922 24724 35924
rect 24668 35870 24670 35922
rect 24670 35870 24722 35922
rect 24722 35870 24724 35922
rect 24668 35868 24724 35870
rect 24108 34914 24164 34916
rect 24108 34862 24110 34914
rect 24110 34862 24162 34914
rect 24162 34862 24164 34914
rect 24108 34860 24164 34862
rect 23884 34802 23940 34804
rect 23884 34750 23886 34802
rect 23886 34750 23938 34802
rect 23938 34750 23940 34802
rect 23884 34748 23940 34750
rect 23772 34636 23828 34692
rect 23548 33964 23604 34020
rect 24444 34690 24500 34692
rect 24444 34638 24446 34690
rect 24446 34638 24498 34690
rect 24498 34638 24500 34690
rect 24444 34636 24500 34638
rect 25116 36092 25172 36148
rect 25676 37266 25732 37268
rect 25676 37214 25678 37266
rect 25678 37214 25730 37266
rect 25730 37214 25732 37266
rect 25676 37212 25732 37214
rect 25564 36258 25620 36260
rect 25564 36206 25566 36258
rect 25566 36206 25618 36258
rect 25618 36206 25620 36258
rect 25564 36204 25620 36206
rect 25452 35532 25508 35588
rect 24220 33292 24276 33348
rect 24892 33346 24948 33348
rect 24892 33294 24894 33346
rect 24894 33294 24946 33346
rect 24946 33294 24948 33346
rect 24892 33292 24948 33294
rect 25340 33292 25396 33348
rect 23548 33068 23604 33124
rect 24556 33234 24612 33236
rect 24556 33182 24558 33234
rect 24558 33182 24610 33234
rect 24610 33182 24612 33234
rect 24556 33180 24612 33182
rect 24444 32732 24500 32788
rect 25228 32674 25284 32676
rect 25228 32622 25230 32674
rect 25230 32622 25282 32674
rect 25282 32622 25284 32674
rect 25228 32620 25284 32622
rect 23660 32060 23716 32116
rect 23996 31890 24052 31892
rect 23996 31838 23998 31890
rect 23998 31838 24050 31890
rect 24050 31838 24052 31890
rect 23996 31836 24052 31838
rect 24668 31836 24724 31892
rect 25676 33234 25732 33236
rect 25676 33182 25678 33234
rect 25678 33182 25730 33234
rect 25730 33182 25732 33234
rect 25676 33180 25732 33182
rect 25676 32844 25732 32900
rect 25564 32786 25620 32788
rect 25564 32734 25566 32786
rect 25566 32734 25618 32786
rect 25618 32734 25620 32786
rect 25564 32732 25620 32734
rect 25452 32562 25508 32564
rect 25452 32510 25454 32562
rect 25454 32510 25506 32562
rect 25506 32510 25508 32562
rect 25452 32508 25508 32510
rect 23884 31666 23940 31668
rect 23884 31614 23886 31666
rect 23886 31614 23938 31666
rect 23938 31614 23940 31666
rect 23884 31612 23940 31614
rect 24556 31612 24612 31668
rect 23772 30994 23828 30996
rect 23772 30942 23774 30994
rect 23774 30942 23826 30994
rect 23826 30942 23828 30994
rect 23772 30940 23828 30942
rect 23660 30828 23716 30884
rect 23548 30322 23604 30324
rect 23548 30270 23550 30322
rect 23550 30270 23602 30322
rect 23602 30270 23604 30322
rect 23548 30268 23604 30270
rect 24444 31276 24500 31332
rect 24780 31500 24836 31556
rect 24668 31164 24724 31220
rect 25452 31218 25508 31220
rect 25452 31166 25454 31218
rect 25454 31166 25506 31218
rect 25506 31166 25508 31218
rect 25452 31164 25508 31166
rect 24444 30994 24500 30996
rect 24444 30942 24446 30994
rect 24446 30942 24498 30994
rect 24498 30942 24500 30994
rect 24444 30940 24500 30942
rect 25340 30882 25396 30884
rect 25340 30830 25342 30882
rect 25342 30830 25394 30882
rect 25394 30830 25396 30882
rect 25340 30828 25396 30830
rect 24332 30716 24388 30772
rect 26236 40290 26292 40292
rect 26236 40238 26238 40290
rect 26238 40238 26290 40290
rect 26290 40238 26292 40290
rect 26236 40236 26292 40238
rect 26236 39900 26292 39956
rect 26124 39676 26180 39732
rect 26124 38108 26180 38164
rect 26012 37772 26068 37828
rect 26460 39564 26516 39620
rect 28028 45666 28084 45668
rect 28028 45614 28030 45666
rect 28030 45614 28082 45666
rect 28082 45614 28084 45666
rect 28028 45612 28084 45614
rect 28364 43820 28420 43876
rect 27916 43596 27972 43652
rect 28140 43260 28196 43316
rect 28252 42642 28308 42644
rect 28252 42590 28254 42642
rect 28254 42590 28306 42642
rect 28306 42590 28308 42642
rect 28252 42588 28308 42590
rect 27916 41132 27972 41188
rect 28924 48860 28980 48916
rect 28812 45612 28868 45668
rect 28700 42588 28756 42644
rect 27916 40684 27972 40740
rect 27580 39676 27636 39732
rect 28476 40684 28532 40740
rect 27692 39618 27748 39620
rect 27692 39566 27694 39618
rect 27694 39566 27746 39618
rect 27746 39566 27748 39618
rect 27692 39564 27748 39566
rect 27132 39004 27188 39060
rect 26908 38780 26964 38836
rect 28252 39676 28308 39732
rect 28028 39394 28084 39396
rect 28028 39342 28030 39394
rect 28030 39342 28082 39394
rect 28082 39342 28084 39394
rect 28028 39340 28084 39342
rect 28140 39004 28196 39060
rect 27692 38668 27748 38724
rect 26348 36652 26404 36708
rect 26796 36482 26852 36484
rect 26796 36430 26798 36482
rect 26798 36430 26850 36482
rect 26850 36430 26852 36482
rect 26796 36428 26852 36430
rect 26572 36204 26628 36260
rect 26908 36204 26964 36260
rect 27020 36876 27076 36932
rect 27804 37826 27860 37828
rect 27804 37774 27806 37826
rect 27806 37774 27858 37826
rect 27858 37774 27860 37826
rect 27804 37772 27860 37774
rect 27580 36764 27636 36820
rect 28588 37826 28644 37828
rect 28588 37774 28590 37826
rect 28590 37774 28642 37826
rect 28642 37774 28644 37826
rect 28588 37772 28644 37774
rect 28812 41132 28868 41188
rect 29260 48188 29316 48244
rect 29372 48130 29428 48132
rect 29372 48078 29374 48130
rect 29374 48078 29426 48130
rect 29426 48078 29428 48130
rect 29372 48076 29428 48078
rect 31388 54738 31444 54740
rect 31388 54686 31390 54738
rect 31390 54686 31442 54738
rect 31442 54686 31444 54738
rect 31388 54684 31444 54686
rect 31612 54460 31668 54516
rect 31276 53228 31332 53284
rect 30940 53116 30996 53172
rect 31836 53058 31892 53060
rect 31836 53006 31838 53058
rect 31838 53006 31890 53058
rect 31890 53006 31892 53058
rect 31836 53004 31892 53006
rect 31500 52946 31556 52948
rect 31500 52894 31502 52946
rect 31502 52894 31554 52946
rect 31554 52894 31556 52946
rect 31500 52892 31556 52894
rect 33180 56306 33236 56308
rect 33180 56254 33182 56306
rect 33182 56254 33234 56306
rect 33234 56254 33236 56306
rect 33180 56252 33236 56254
rect 32284 53452 32340 53508
rect 31388 52386 31444 52388
rect 31388 52334 31390 52386
rect 31390 52334 31442 52386
rect 31442 52334 31444 52386
rect 31388 52332 31444 52334
rect 31724 51996 31780 52052
rect 29932 48860 29988 48916
rect 30044 49980 30100 50036
rect 30156 49756 30212 49812
rect 30044 48748 30100 48804
rect 29148 47068 29204 47124
rect 30156 47068 30212 47124
rect 30156 46732 30212 46788
rect 29148 46620 29204 46676
rect 30492 50092 30548 50148
rect 30940 50092 30996 50148
rect 31500 49756 31556 49812
rect 31388 48802 31444 48804
rect 31388 48750 31390 48802
rect 31390 48750 31442 48802
rect 31442 48750 31444 48802
rect 31388 48748 31444 48750
rect 30380 48242 30436 48244
rect 30380 48190 30382 48242
rect 30382 48190 30434 48242
rect 30434 48190 30436 48242
rect 30380 48188 30436 48190
rect 30940 48300 30996 48356
rect 30828 46732 30884 46788
rect 30940 46674 30996 46676
rect 30940 46622 30942 46674
rect 30942 46622 30994 46674
rect 30994 46622 30996 46674
rect 30940 46620 30996 46622
rect 29260 45666 29316 45668
rect 29260 45614 29262 45666
rect 29262 45614 29314 45666
rect 29314 45614 29316 45666
rect 29260 45612 29316 45614
rect 29484 45106 29540 45108
rect 29484 45054 29486 45106
rect 29486 45054 29538 45106
rect 29538 45054 29540 45106
rect 29484 45052 29540 45054
rect 30380 45106 30436 45108
rect 30380 45054 30382 45106
rect 30382 45054 30434 45106
rect 30434 45054 30436 45106
rect 30380 45052 30436 45054
rect 29932 44716 29988 44772
rect 29148 44322 29204 44324
rect 29148 44270 29150 44322
rect 29150 44270 29202 44322
rect 29202 44270 29204 44322
rect 29148 44268 29204 44270
rect 30380 43708 30436 43764
rect 29036 43650 29092 43652
rect 29036 43598 29038 43650
rect 29038 43598 29090 43650
rect 29090 43598 29092 43650
rect 29036 43596 29092 43598
rect 29036 41692 29092 41748
rect 29596 43538 29652 43540
rect 29596 43486 29598 43538
rect 29598 43486 29650 43538
rect 29650 43486 29652 43538
rect 29596 43484 29652 43486
rect 29820 42812 29876 42868
rect 29260 42642 29316 42644
rect 29260 42590 29262 42642
rect 29262 42590 29314 42642
rect 29314 42590 29316 42642
rect 29260 42588 29316 42590
rect 29372 42364 29428 42420
rect 29148 40684 29204 40740
rect 29484 40684 29540 40740
rect 29260 40236 29316 40292
rect 29260 39730 29316 39732
rect 29260 39678 29262 39730
rect 29262 39678 29314 39730
rect 29314 39678 29316 39730
rect 29260 39676 29316 39678
rect 29596 38668 29652 38724
rect 28924 38444 28980 38500
rect 28028 37266 28084 37268
rect 28028 37214 28030 37266
rect 28030 37214 28082 37266
rect 28082 37214 28084 37266
rect 28028 37212 28084 37214
rect 27916 36876 27972 36932
rect 28140 36764 28196 36820
rect 28476 36988 28532 37044
rect 27580 36428 27636 36484
rect 27804 36370 27860 36372
rect 27804 36318 27806 36370
rect 27806 36318 27858 36370
rect 27858 36318 27860 36370
rect 27804 36316 27860 36318
rect 28028 36370 28084 36372
rect 28028 36318 28030 36370
rect 28030 36318 28082 36370
rect 28082 36318 28084 36370
rect 28028 36316 28084 36318
rect 27804 35756 27860 35812
rect 27580 34860 27636 34916
rect 26460 34636 26516 34692
rect 27244 34690 27300 34692
rect 27244 34638 27246 34690
rect 27246 34638 27298 34690
rect 27298 34638 27300 34690
rect 27244 34636 27300 34638
rect 25900 33516 25956 33572
rect 25900 32620 25956 32676
rect 24220 30156 24276 30212
rect 26012 31612 26068 31668
rect 23996 29986 24052 29988
rect 23996 29934 23998 29986
rect 23998 29934 24050 29986
rect 24050 29934 24052 29986
rect 23996 29932 24052 29934
rect 23436 29596 23492 29652
rect 23324 29538 23380 29540
rect 23324 29486 23326 29538
rect 23326 29486 23378 29538
rect 23378 29486 23380 29538
rect 23324 29484 23380 29486
rect 24892 29986 24948 29988
rect 24892 29934 24894 29986
rect 24894 29934 24946 29986
rect 24946 29934 24948 29986
rect 24892 29932 24948 29934
rect 24892 29260 24948 29316
rect 25676 28924 25732 28980
rect 25228 28812 25284 28868
rect 22428 27858 22484 27860
rect 22428 27806 22430 27858
rect 22430 27806 22482 27858
rect 22482 27806 22484 27858
rect 22428 27804 22484 27806
rect 24668 28700 24724 28756
rect 24220 28476 24276 28532
rect 23996 28418 24052 28420
rect 23996 28366 23998 28418
rect 23998 28366 24050 28418
rect 24050 28366 24052 28418
rect 23996 28364 24052 28366
rect 22764 27356 22820 27412
rect 23100 27020 23156 27076
rect 21756 26290 21812 26292
rect 21756 26238 21758 26290
rect 21758 26238 21810 26290
rect 21810 26238 21812 26290
rect 21756 26236 21812 26238
rect 21980 25900 22036 25956
rect 21756 25676 21812 25732
rect 21980 23212 22036 23268
rect 21756 21756 21812 21812
rect 21756 20636 21812 20692
rect 21868 22988 21924 23044
rect 21868 22428 21924 22484
rect 22764 26514 22820 26516
rect 22764 26462 22766 26514
rect 22766 26462 22818 26514
rect 22818 26462 22820 26514
rect 22764 26460 22820 26462
rect 22428 26348 22484 26404
rect 23436 27074 23492 27076
rect 23436 27022 23438 27074
rect 23438 27022 23490 27074
rect 23490 27022 23492 27074
rect 23436 27020 23492 27022
rect 23884 27074 23940 27076
rect 23884 27022 23886 27074
rect 23886 27022 23938 27074
rect 23938 27022 23940 27074
rect 23884 27020 23940 27022
rect 22988 26012 23044 26068
rect 23324 26124 23380 26180
rect 22876 25452 22932 25508
rect 22428 25228 22484 25284
rect 22428 25004 22484 25060
rect 22204 23884 22260 23940
rect 24108 26178 24164 26180
rect 24108 26126 24110 26178
rect 24110 26126 24162 26178
rect 24162 26126 24164 26178
rect 24108 26124 24164 26126
rect 23548 26012 23604 26068
rect 23996 24834 24052 24836
rect 23996 24782 23998 24834
rect 23998 24782 24050 24834
rect 24050 24782 24052 24834
rect 23996 24780 24052 24782
rect 22428 23042 22484 23044
rect 22428 22990 22430 23042
rect 22430 22990 22482 23042
rect 22482 22990 22484 23042
rect 22428 22988 22484 22990
rect 21980 21980 22036 22036
rect 21868 20860 21924 20916
rect 21196 20018 21252 20020
rect 21196 19966 21198 20018
rect 21198 19966 21250 20018
rect 21250 19966 21252 20018
rect 21196 19964 21252 19966
rect 21084 19180 21140 19236
rect 20412 19010 20468 19012
rect 20412 18958 20414 19010
rect 20414 18958 20466 19010
rect 20466 18958 20468 19010
rect 20412 18956 20468 18958
rect 20860 18956 20916 19012
rect 20300 18060 20356 18116
rect 21196 19068 21252 19124
rect 21084 18956 21140 19012
rect 20524 17612 20580 17668
rect 20412 17106 20468 17108
rect 20412 17054 20414 17106
rect 20414 17054 20466 17106
rect 20466 17054 20468 17106
rect 20412 17052 20468 17054
rect 20748 17106 20804 17108
rect 20748 17054 20750 17106
rect 20750 17054 20802 17106
rect 20802 17054 20804 17106
rect 20748 17052 20804 17054
rect 22092 21644 22148 21700
rect 21980 20802 22036 20804
rect 21980 20750 21982 20802
rect 21982 20750 22034 20802
rect 22034 20750 22036 20802
rect 21980 20748 22036 20750
rect 22428 20748 22484 20804
rect 22316 20690 22372 20692
rect 22316 20638 22318 20690
rect 22318 20638 22370 20690
rect 22370 20638 22372 20690
rect 22316 20636 22372 20638
rect 21644 19234 21700 19236
rect 21644 19182 21646 19234
rect 21646 19182 21698 19234
rect 21698 19182 21700 19234
rect 21644 19180 21700 19182
rect 22204 19852 22260 19908
rect 21420 17666 21476 17668
rect 21420 17614 21422 17666
rect 21422 17614 21474 17666
rect 21474 17614 21476 17666
rect 21420 17612 21476 17614
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20188 14140 20244 14196
rect 20300 14476 20356 14532
rect 20044 14084 20100 14086
rect 20188 13580 20244 13636
rect 19068 12572 19124 12628
rect 19180 12290 19236 12292
rect 19180 12238 19182 12290
rect 19182 12238 19234 12290
rect 19234 12238 19236 12290
rect 19180 12236 19236 12238
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19740 12402 19796 12404
rect 19740 12350 19742 12402
rect 19742 12350 19794 12402
rect 19794 12350 19796 12402
rect 19740 12348 19796 12350
rect 20636 12290 20692 12292
rect 20636 12238 20638 12290
rect 20638 12238 20690 12290
rect 20690 12238 20692 12290
rect 20636 12236 20692 12238
rect 20860 11676 20916 11732
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19068 9826 19124 9828
rect 19068 9774 19070 9826
rect 19070 9774 19122 9826
rect 19122 9774 19124 9826
rect 19068 9772 19124 9774
rect 18956 8258 19012 8260
rect 18956 8206 18958 8258
rect 18958 8206 19010 8258
rect 19010 8206 19012 8258
rect 18956 8204 19012 8206
rect 19852 9826 19908 9828
rect 19852 9774 19854 9826
rect 19854 9774 19906 9826
rect 19906 9774 19908 9826
rect 19852 9772 19908 9774
rect 19404 9714 19460 9716
rect 19404 9662 19406 9714
rect 19406 9662 19458 9714
rect 19458 9662 19460 9714
rect 19404 9660 19460 9662
rect 20748 10444 20804 10500
rect 20076 9660 20132 9716
rect 20748 9548 20804 9604
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19516 9154 19572 9156
rect 19516 9102 19518 9154
rect 19518 9102 19570 9154
rect 19570 9102 19572 9154
rect 19516 9100 19572 9102
rect 21532 16044 21588 16100
rect 21756 17052 21812 17108
rect 22316 19740 22372 19796
rect 22316 19068 22372 19124
rect 22540 19180 22596 19236
rect 22092 17836 22148 17892
rect 22428 17052 22484 17108
rect 22876 18284 22932 18340
rect 22876 17612 22932 17668
rect 21980 16828 22036 16884
rect 22204 16098 22260 16100
rect 22204 16046 22206 16098
rect 22206 16046 22258 16098
rect 22258 16046 22260 16098
rect 22204 16044 22260 16046
rect 22428 15260 22484 15316
rect 23436 20914 23492 20916
rect 23436 20862 23438 20914
rect 23438 20862 23490 20914
rect 23490 20862 23492 20914
rect 23436 20860 23492 20862
rect 23660 19906 23716 19908
rect 23660 19854 23662 19906
rect 23662 19854 23714 19906
rect 23714 19854 23716 19906
rect 23660 19852 23716 19854
rect 23548 19794 23604 19796
rect 23548 19742 23550 19794
rect 23550 19742 23602 19794
rect 23602 19742 23604 19794
rect 23548 19740 23604 19742
rect 23884 23042 23940 23044
rect 23884 22990 23886 23042
rect 23886 22990 23938 23042
rect 23938 22990 23940 23042
rect 23884 22988 23940 22990
rect 23884 20860 23940 20916
rect 23884 19740 23940 19796
rect 24556 26460 24612 26516
rect 24668 26348 24724 26404
rect 24556 25788 24612 25844
rect 25900 28588 25956 28644
rect 26012 28476 26068 28532
rect 25228 27020 25284 27076
rect 25900 27858 25956 27860
rect 25900 27806 25902 27858
rect 25902 27806 25954 27858
rect 25954 27806 25956 27858
rect 25900 27804 25956 27806
rect 27916 34300 27972 34356
rect 28140 34914 28196 34916
rect 28140 34862 28142 34914
rect 28142 34862 28194 34914
rect 28194 34862 28196 34914
rect 28140 34860 28196 34862
rect 28028 34188 28084 34244
rect 30044 42028 30100 42084
rect 30044 41468 30100 41524
rect 30268 42812 30324 42868
rect 31836 48748 31892 48804
rect 31388 45276 31444 45332
rect 32172 50316 32228 50372
rect 32172 49810 32228 49812
rect 32172 49758 32174 49810
rect 32174 49758 32226 49810
rect 32226 49758 32228 49810
rect 32172 49756 32228 49758
rect 31948 47740 32004 47796
rect 31836 46956 31892 47012
rect 32172 46956 32228 47012
rect 32284 46786 32340 46788
rect 32284 46734 32286 46786
rect 32286 46734 32338 46786
rect 32338 46734 32340 46786
rect 32284 46732 32340 46734
rect 31724 46060 31780 46116
rect 31724 45106 31780 45108
rect 31724 45054 31726 45106
rect 31726 45054 31778 45106
rect 31778 45054 31780 45106
rect 31724 45052 31780 45054
rect 31500 44994 31556 44996
rect 31500 44942 31502 44994
rect 31502 44942 31554 44994
rect 31554 44942 31556 44994
rect 31500 44940 31556 44942
rect 30716 42082 30772 42084
rect 30716 42030 30718 42082
rect 30718 42030 30770 42082
rect 30770 42030 30772 42082
rect 30716 42028 30772 42030
rect 31276 42028 31332 42084
rect 30492 41970 30548 41972
rect 30492 41918 30494 41970
rect 30494 41918 30546 41970
rect 30546 41918 30548 41970
rect 30492 41916 30548 41918
rect 30940 41970 30996 41972
rect 30940 41918 30942 41970
rect 30942 41918 30994 41970
rect 30994 41918 30996 41970
rect 30940 41916 30996 41918
rect 30268 41692 30324 41748
rect 30716 41692 30772 41748
rect 30044 40796 30100 40852
rect 29932 40236 29988 40292
rect 30156 39900 30212 39956
rect 31388 41858 31444 41860
rect 31388 41806 31390 41858
rect 31390 41806 31442 41858
rect 31442 41806 31444 41858
rect 31388 41804 31444 41806
rect 30716 41186 30772 41188
rect 30716 41134 30718 41186
rect 30718 41134 30770 41186
rect 30770 41134 30772 41186
rect 30716 41132 30772 41134
rect 30940 40796 30996 40852
rect 30268 39676 30324 39732
rect 31612 40796 31668 40852
rect 31052 40178 31108 40180
rect 31052 40126 31054 40178
rect 31054 40126 31106 40178
rect 31106 40126 31108 40178
rect 31052 40124 31108 40126
rect 30828 39788 30884 39844
rect 31164 39676 31220 39732
rect 30268 39004 30324 39060
rect 30156 38108 30212 38164
rect 30828 38162 30884 38164
rect 30828 38110 30830 38162
rect 30830 38110 30882 38162
rect 30882 38110 30884 38162
rect 30828 38108 30884 38110
rect 30716 37996 30772 38052
rect 30492 37884 30548 37940
rect 29036 37772 29092 37828
rect 29148 37324 29204 37380
rect 28812 37266 28868 37268
rect 28812 37214 28814 37266
rect 28814 37214 28866 37266
rect 28866 37214 28868 37266
rect 28812 37212 28868 37214
rect 29260 36988 29316 37044
rect 30044 36876 30100 36932
rect 28700 36204 28756 36260
rect 29708 36258 29764 36260
rect 29708 36206 29710 36258
rect 29710 36206 29762 36258
rect 29762 36206 29764 36258
rect 29708 36204 29764 36206
rect 29036 35532 29092 35588
rect 28812 34636 28868 34692
rect 28924 35308 28980 35364
rect 27804 32844 27860 32900
rect 28588 33234 28644 33236
rect 28588 33182 28590 33234
rect 28590 33182 28642 33234
rect 28642 33182 28644 33234
rect 28588 33180 28644 33182
rect 28476 32732 28532 32788
rect 26684 31948 26740 32004
rect 26684 28812 26740 28868
rect 26348 28700 26404 28756
rect 26572 28700 26628 28756
rect 26460 28642 26516 28644
rect 26460 28590 26462 28642
rect 26462 28590 26514 28642
rect 26514 28590 26516 28642
rect 26460 28588 26516 28590
rect 26684 27804 26740 27860
rect 26796 28924 26852 28980
rect 27244 32284 27300 32340
rect 28588 31890 28644 31892
rect 28588 31838 28590 31890
rect 28590 31838 28642 31890
rect 28642 31838 28644 31890
rect 28588 31836 28644 31838
rect 27804 30604 27860 30660
rect 27244 29484 27300 29540
rect 27916 29596 27972 29652
rect 25452 26684 25508 26740
rect 25340 26514 25396 26516
rect 25340 26462 25342 26514
rect 25342 26462 25394 26514
rect 25394 26462 25396 26514
rect 25340 26460 25396 26462
rect 24780 26124 24836 26180
rect 24892 25788 24948 25844
rect 25452 25788 25508 25844
rect 24780 24556 24836 24612
rect 24780 22988 24836 23044
rect 24668 21474 24724 21476
rect 24668 21422 24670 21474
rect 24670 21422 24722 21474
rect 24722 21422 24724 21474
rect 24668 21420 24724 21422
rect 24668 20860 24724 20916
rect 24556 20690 24612 20692
rect 24556 20638 24558 20690
rect 24558 20638 24610 20690
rect 24610 20638 24612 20690
rect 24556 20636 24612 20638
rect 24108 19964 24164 20020
rect 24444 19346 24500 19348
rect 24444 19294 24446 19346
rect 24446 19294 24498 19346
rect 24498 19294 24500 19346
rect 24444 19292 24500 19294
rect 23884 18338 23940 18340
rect 23884 18286 23886 18338
rect 23886 18286 23938 18338
rect 23938 18286 23940 18338
rect 23884 18284 23940 18286
rect 22764 16716 22820 16772
rect 24220 17948 24276 18004
rect 21532 13634 21588 13636
rect 21532 13582 21534 13634
rect 21534 13582 21586 13634
rect 21586 13582 21588 13634
rect 21532 13580 21588 13582
rect 23996 16604 24052 16660
rect 22988 16098 23044 16100
rect 22988 16046 22990 16098
rect 22990 16046 23042 16098
rect 23042 16046 23044 16098
rect 22988 16044 23044 16046
rect 23660 16098 23716 16100
rect 23660 16046 23662 16098
rect 23662 16046 23714 16098
rect 23714 16046 23716 16098
rect 23660 16044 23716 16046
rect 23772 15932 23828 15988
rect 22988 15148 23044 15204
rect 23100 15820 23156 15876
rect 23324 15202 23380 15204
rect 23324 15150 23326 15202
rect 23326 15150 23378 15202
rect 23378 15150 23380 15202
rect 23324 15148 23380 15150
rect 23100 14028 23156 14084
rect 22876 13916 22932 13972
rect 22540 12684 22596 12740
rect 24444 18284 24500 18340
rect 24780 17500 24836 17556
rect 24668 16716 24724 16772
rect 24556 15986 24612 15988
rect 24556 15934 24558 15986
rect 24558 15934 24610 15986
rect 24610 15934 24612 15986
rect 24556 15932 24612 15934
rect 24668 13970 24724 13972
rect 24668 13918 24670 13970
rect 24670 13918 24722 13970
rect 24722 13918 24724 13970
rect 24668 13916 24724 13918
rect 24108 12850 24164 12852
rect 24108 12798 24110 12850
rect 24110 12798 24162 12850
rect 24162 12798 24164 12850
rect 24108 12796 24164 12798
rect 24668 12850 24724 12852
rect 24668 12798 24670 12850
rect 24670 12798 24722 12850
rect 24722 12798 24724 12850
rect 24668 12796 24724 12798
rect 24220 12738 24276 12740
rect 24220 12686 24222 12738
rect 24222 12686 24274 12738
rect 24274 12686 24276 12738
rect 24220 12684 24276 12686
rect 24668 11452 24724 11508
rect 25900 26290 25956 26292
rect 25900 26238 25902 26290
rect 25902 26238 25954 26290
rect 25954 26238 25956 26290
rect 25900 26236 25956 26238
rect 25900 25788 25956 25844
rect 25452 24556 25508 24612
rect 25900 24220 25956 24276
rect 26236 25788 26292 25844
rect 26236 25506 26292 25508
rect 26236 25454 26238 25506
rect 26238 25454 26290 25506
rect 26290 25454 26292 25506
rect 26236 25452 26292 25454
rect 26124 25228 26180 25284
rect 26236 24332 26292 24388
rect 25676 23884 25732 23940
rect 25340 21868 25396 21924
rect 26012 21756 26068 21812
rect 26012 21420 26068 21476
rect 25340 20860 25396 20916
rect 25564 21308 25620 21364
rect 25228 19180 25284 19236
rect 25228 18450 25284 18452
rect 25228 18398 25230 18450
rect 25230 18398 25282 18450
rect 25282 18398 25284 18450
rect 25228 18396 25284 18398
rect 25228 17948 25284 18004
rect 25676 19292 25732 19348
rect 26236 21420 26292 21476
rect 26796 25506 26852 25508
rect 26796 25454 26798 25506
rect 26798 25454 26850 25506
rect 26850 25454 26852 25506
rect 26796 25452 26852 25454
rect 26908 25394 26964 25396
rect 26908 25342 26910 25394
rect 26910 25342 26962 25394
rect 26962 25342 26964 25394
rect 26908 25340 26964 25342
rect 28364 28588 28420 28644
rect 28364 28082 28420 28084
rect 28364 28030 28366 28082
rect 28366 28030 28418 28082
rect 28418 28030 28420 28082
rect 28364 28028 28420 28030
rect 28588 27970 28644 27972
rect 28588 27918 28590 27970
rect 28590 27918 28642 27970
rect 28642 27918 28644 27970
rect 28588 27916 28644 27918
rect 27580 27804 27636 27860
rect 30044 36092 30100 36148
rect 30716 36876 30772 36932
rect 31388 38332 31444 38388
rect 33180 55356 33236 55412
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35756 55522 35812 55524
rect 35756 55470 35758 55522
rect 35758 55470 35810 55522
rect 35810 55470 35812 55522
rect 35756 55468 35812 55470
rect 33740 55410 33796 55412
rect 33740 55358 33742 55410
rect 33742 55358 33794 55410
rect 33794 55358 33796 55410
rect 33740 55356 33796 55358
rect 35980 55356 36036 55412
rect 36764 55468 36820 55524
rect 33628 54796 33684 54852
rect 33292 54572 33348 54628
rect 33516 54402 33572 54404
rect 33516 54350 33518 54402
rect 33518 54350 33570 54402
rect 33570 54350 33572 54402
rect 33516 54348 33572 54350
rect 33964 54402 34020 54404
rect 33964 54350 33966 54402
rect 33966 54350 34018 54402
rect 34018 54350 34020 54402
rect 33964 54348 34020 54350
rect 33292 54236 33348 54292
rect 33180 53788 33236 53844
rect 32732 53228 32788 53284
rect 34636 55074 34692 55076
rect 34636 55022 34638 55074
rect 34638 55022 34690 55074
rect 34690 55022 34692 55074
rect 34636 55020 34692 55022
rect 34412 54796 34468 54852
rect 34188 54738 34244 54740
rect 34188 54686 34190 54738
rect 34190 54686 34242 54738
rect 34242 54686 34244 54738
rect 34188 54684 34244 54686
rect 34188 54402 34244 54404
rect 34188 54350 34190 54402
rect 34190 54350 34242 54402
rect 34242 54350 34244 54402
rect 34188 54348 34244 54350
rect 33628 53676 33684 53732
rect 34188 53788 34244 53844
rect 33516 53228 33572 53284
rect 32508 53170 32564 53172
rect 32508 53118 32510 53170
rect 32510 53118 32562 53170
rect 32562 53118 32564 53170
rect 32508 53116 32564 53118
rect 33292 53116 33348 53172
rect 33068 51996 33124 52052
rect 32732 50316 32788 50372
rect 32060 46060 32116 46116
rect 32508 49922 32564 49924
rect 32508 49870 32510 49922
rect 32510 49870 32562 49922
rect 32562 49870 32564 49922
rect 32508 49868 32564 49870
rect 31948 45164 32004 45220
rect 31836 44380 31892 44436
rect 33068 48860 33124 48916
rect 33180 48636 33236 48692
rect 32844 47740 32900 47796
rect 32844 46396 32900 46452
rect 32284 45276 32340 45332
rect 32508 45164 32564 45220
rect 33404 48860 33460 48916
rect 32508 44322 32564 44324
rect 32508 44270 32510 44322
rect 32510 44270 32562 44322
rect 32562 44270 32564 44322
rect 32508 44268 32564 44270
rect 33180 45052 33236 45108
rect 33404 45890 33460 45892
rect 33404 45838 33406 45890
rect 33406 45838 33458 45890
rect 33458 45838 33460 45890
rect 33404 45836 33460 45838
rect 33404 45500 33460 45556
rect 33404 45276 33460 45332
rect 33292 44716 33348 44772
rect 33628 50428 33684 50484
rect 34076 53452 34132 53508
rect 33964 51548 34020 51604
rect 34636 53116 34692 53172
rect 34412 52892 34468 52948
rect 34412 51996 34468 52052
rect 34076 50428 34132 50484
rect 34300 50204 34356 50260
rect 34300 49980 34356 50036
rect 34860 52892 34916 52948
rect 34636 51602 34692 51604
rect 34636 51550 34638 51602
rect 34638 51550 34690 51602
rect 34690 51550 34692 51602
rect 34636 51548 34692 51550
rect 34524 51378 34580 51380
rect 34524 51326 34526 51378
rect 34526 51326 34578 51378
rect 34578 51326 34580 51378
rect 34524 51324 34580 51326
rect 34748 51212 34804 51268
rect 35644 55186 35700 55188
rect 35644 55134 35646 55186
rect 35646 55134 35698 55186
rect 35698 55134 35700 55186
rect 35644 55132 35700 55134
rect 35084 55074 35140 55076
rect 35084 55022 35086 55074
rect 35086 55022 35138 55074
rect 35138 55022 35140 55074
rect 35084 55020 35140 55022
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 38332 55916 38388 55972
rect 37100 55410 37156 55412
rect 37100 55358 37102 55410
rect 37102 55358 37154 55410
rect 37154 55358 37156 55410
rect 37100 55356 37156 55358
rect 37660 55356 37716 55412
rect 36988 55244 37044 55300
rect 36428 55020 36484 55076
rect 37884 54684 37940 54740
rect 38332 55132 38388 55188
rect 38780 54908 38836 54964
rect 38220 54626 38276 54628
rect 38220 54574 38222 54626
rect 38222 54574 38274 54626
rect 38274 54574 38276 54626
rect 38220 54572 38276 54574
rect 37772 54236 37828 54292
rect 37884 54348 37940 54404
rect 37660 54012 37716 54068
rect 36316 53788 36372 53844
rect 37660 53842 37716 53844
rect 37660 53790 37662 53842
rect 37662 53790 37714 53842
rect 37714 53790 37716 53842
rect 37660 53788 37716 53790
rect 36988 53676 37044 53732
rect 35420 53618 35476 53620
rect 35420 53566 35422 53618
rect 35422 53566 35474 53618
rect 35474 53566 35476 53618
rect 35420 53564 35476 53566
rect 35868 53228 35924 53284
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 34972 51490 35028 51492
rect 34972 51438 34974 51490
rect 34974 51438 35026 51490
rect 35026 51438 35028 51490
rect 34972 51436 35028 51438
rect 34748 50092 34804 50148
rect 33964 49084 34020 49140
rect 33740 48636 33796 48692
rect 34860 47964 34916 48020
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35308 50482 35364 50484
rect 35308 50430 35310 50482
rect 35310 50430 35362 50482
rect 35362 50430 35364 50482
rect 35308 50428 35364 50430
rect 35980 52946 36036 52948
rect 35980 52894 35982 52946
rect 35982 52894 36034 52946
rect 36034 52894 36036 52946
rect 35980 52892 36036 52894
rect 37996 54124 38052 54180
rect 38444 54124 38500 54180
rect 39116 54908 39172 54964
rect 40124 54626 40180 54628
rect 40124 54574 40126 54626
rect 40126 54574 40178 54626
rect 40178 54574 40180 54626
rect 40124 54572 40180 54574
rect 38780 54460 38836 54516
rect 38556 54012 38612 54068
rect 38556 53788 38612 53844
rect 38668 54236 38724 54292
rect 38220 53618 38276 53620
rect 38220 53566 38222 53618
rect 38222 53566 38274 53618
rect 38274 53566 38276 53618
rect 38220 53564 38276 53566
rect 37324 53004 37380 53060
rect 38668 53116 38724 53172
rect 37996 52780 38052 52836
rect 39564 54348 39620 54404
rect 39900 54514 39956 54516
rect 39900 54462 39902 54514
rect 39902 54462 39954 54514
rect 39954 54462 39956 54514
rect 39900 54460 39956 54462
rect 39900 53788 39956 53844
rect 39116 53730 39172 53732
rect 39116 53678 39118 53730
rect 39118 53678 39170 53730
rect 39170 53678 39172 53730
rect 39116 53676 39172 53678
rect 40012 53564 40068 53620
rect 37212 51772 37268 51828
rect 36988 51436 37044 51492
rect 35980 51324 36036 51380
rect 35980 50540 36036 50596
rect 36540 50540 36596 50596
rect 35980 50034 36036 50036
rect 35980 49982 35982 50034
rect 35982 49982 36034 50034
rect 36034 49982 36036 50034
rect 35980 49980 36036 49982
rect 36316 50034 36372 50036
rect 36316 49982 36318 50034
rect 36318 49982 36370 50034
rect 36370 49982 36372 50034
rect 36316 49980 36372 49982
rect 36092 49810 36148 49812
rect 36092 49758 36094 49810
rect 36094 49758 36146 49810
rect 36146 49758 36148 49810
rect 36092 49756 36148 49758
rect 39228 51996 39284 52052
rect 39452 51996 39508 52052
rect 38780 51378 38836 51380
rect 38780 51326 38782 51378
rect 38782 51326 38834 51378
rect 38834 51326 38836 51378
rect 38780 51324 38836 51326
rect 37212 51212 37268 51268
rect 37100 50652 37156 50708
rect 37212 49980 37268 50036
rect 36204 49698 36260 49700
rect 36204 49646 36206 49698
rect 36206 49646 36258 49698
rect 36258 49646 36260 49698
rect 36204 49644 36260 49646
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35084 48636 35140 48692
rect 36316 48802 36372 48804
rect 36316 48750 36318 48802
rect 36318 48750 36370 48802
rect 36370 48750 36372 48802
rect 36316 48748 36372 48750
rect 35644 48188 35700 48244
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35532 47628 35588 47684
rect 34300 47234 34356 47236
rect 34300 47182 34302 47234
rect 34302 47182 34354 47234
rect 34354 47182 34356 47234
rect 34300 47180 34356 47182
rect 34076 46786 34132 46788
rect 34076 46734 34078 46786
rect 34078 46734 34130 46786
rect 34130 46734 34132 46786
rect 34076 46732 34132 46734
rect 33964 46396 34020 46452
rect 33964 46002 34020 46004
rect 33964 45950 33966 46002
rect 33966 45950 34018 46002
rect 34018 45950 34020 46002
rect 33964 45948 34020 45950
rect 33852 45276 33908 45332
rect 33628 44940 33684 44996
rect 33068 43708 33124 43764
rect 33628 44044 33684 44100
rect 33404 43708 33460 43764
rect 33516 43650 33572 43652
rect 33516 43598 33518 43650
rect 33518 43598 33570 43650
rect 33570 43598 33572 43650
rect 33516 43596 33572 43598
rect 33852 44940 33908 44996
rect 34524 47234 34580 47236
rect 34524 47182 34526 47234
rect 34526 47182 34578 47234
rect 34578 47182 34580 47234
rect 34524 47180 34580 47182
rect 34412 45218 34468 45220
rect 34412 45166 34414 45218
rect 34414 45166 34466 45218
rect 34466 45166 34468 45218
rect 34412 45164 34468 45166
rect 34524 45052 34580 45108
rect 33964 44268 34020 44324
rect 34076 44604 34132 44660
rect 33852 44210 33908 44212
rect 33852 44158 33854 44210
rect 33854 44158 33906 44210
rect 33906 44158 33908 44210
rect 33852 44156 33908 44158
rect 32396 41916 32452 41972
rect 32284 40124 32340 40180
rect 32508 41020 32564 41076
rect 32508 40402 32564 40404
rect 32508 40350 32510 40402
rect 32510 40350 32562 40402
rect 32562 40350 32564 40402
rect 32508 40348 32564 40350
rect 32508 39564 32564 39620
rect 32396 39394 32452 39396
rect 32396 39342 32398 39394
rect 32398 39342 32450 39394
rect 32450 39342 32452 39394
rect 32396 39340 32452 39342
rect 32508 39228 32564 39284
rect 32732 42642 32788 42644
rect 32732 42590 32734 42642
rect 32734 42590 32786 42642
rect 32786 42590 32788 42642
rect 32732 42588 32788 42590
rect 32844 42028 32900 42084
rect 34188 43596 34244 43652
rect 33740 42812 33796 42868
rect 34188 42476 34244 42532
rect 33740 42194 33796 42196
rect 33740 42142 33742 42194
rect 33742 42142 33794 42194
rect 33794 42142 33796 42194
rect 33740 42140 33796 42142
rect 33740 41692 33796 41748
rect 32844 39676 32900 39732
rect 31836 38332 31892 38388
rect 31388 37884 31444 37940
rect 31612 36428 31668 36484
rect 30268 36092 30324 36148
rect 30492 35980 30548 36036
rect 31052 36258 31108 36260
rect 31052 36206 31054 36258
rect 31054 36206 31106 36258
rect 31106 36206 31108 36258
rect 31052 36204 31108 36206
rect 30716 36092 30772 36148
rect 29708 35308 29764 35364
rect 30604 35532 30660 35588
rect 30492 35420 30548 35476
rect 29484 34636 29540 34692
rect 29932 34242 29988 34244
rect 29932 34190 29934 34242
rect 29934 34190 29986 34242
rect 29986 34190 29988 34242
rect 29932 34188 29988 34190
rect 29484 32844 29540 32900
rect 29820 32786 29876 32788
rect 29820 32734 29822 32786
rect 29822 32734 29874 32786
rect 29874 32734 29876 32786
rect 29820 32732 29876 32734
rect 29148 32284 29204 32340
rect 29260 32396 29316 32452
rect 29148 31836 29204 31892
rect 28476 26684 28532 26740
rect 27580 26460 27636 26516
rect 28140 26460 28196 26516
rect 27692 26236 27748 26292
rect 27244 25394 27300 25396
rect 27244 25342 27246 25394
rect 27246 25342 27298 25394
rect 27298 25342 27300 25394
rect 27244 25340 27300 25342
rect 27468 25394 27524 25396
rect 27468 25342 27470 25394
rect 27470 25342 27522 25394
rect 27522 25342 27524 25394
rect 27468 25340 27524 25342
rect 27356 25282 27412 25284
rect 27356 25230 27358 25282
rect 27358 25230 27410 25282
rect 27410 25230 27412 25282
rect 27356 25228 27412 25230
rect 27020 25004 27076 25060
rect 26460 23938 26516 23940
rect 26460 23886 26462 23938
rect 26462 23886 26514 23938
rect 26514 23886 26516 23938
rect 26460 23884 26516 23886
rect 26908 23212 26964 23268
rect 26572 21756 26628 21812
rect 26908 21698 26964 21700
rect 26908 21646 26910 21698
rect 26910 21646 26962 21698
rect 26962 21646 26964 21698
rect 26908 21644 26964 21646
rect 26684 21474 26740 21476
rect 26684 21422 26686 21474
rect 26686 21422 26738 21474
rect 26738 21422 26740 21474
rect 26684 21420 26740 21422
rect 27580 24892 27636 24948
rect 27804 25340 27860 25396
rect 29708 32284 29764 32340
rect 31164 35810 31220 35812
rect 31164 35758 31166 35810
rect 31166 35758 31218 35810
rect 31218 35758 31220 35810
rect 31164 35756 31220 35758
rect 30828 35308 30884 35364
rect 30268 34690 30324 34692
rect 30268 34638 30270 34690
rect 30270 34638 30322 34690
rect 30322 34638 30324 34690
rect 30268 34636 30324 34638
rect 30492 34188 30548 34244
rect 30044 32674 30100 32676
rect 30044 32622 30046 32674
rect 30046 32622 30098 32674
rect 30098 32622 30100 32674
rect 30044 32620 30100 32622
rect 29484 31778 29540 31780
rect 29484 31726 29486 31778
rect 29486 31726 29538 31778
rect 29538 31726 29540 31778
rect 29484 31724 29540 31726
rect 29820 31554 29876 31556
rect 29820 31502 29822 31554
rect 29822 31502 29874 31554
rect 29874 31502 29876 31554
rect 29820 31500 29876 31502
rect 29932 31164 29988 31220
rect 29484 30994 29540 30996
rect 29484 30942 29486 30994
rect 29486 30942 29538 30994
rect 29538 30942 29540 30994
rect 29484 30940 29540 30942
rect 29820 30994 29876 30996
rect 29820 30942 29822 30994
rect 29822 30942 29874 30994
rect 29874 30942 29876 30994
rect 29820 30940 29876 30942
rect 29708 30268 29764 30324
rect 30380 31836 30436 31892
rect 30156 31778 30212 31780
rect 30156 31726 30158 31778
rect 30158 31726 30210 31778
rect 30210 31726 30212 31778
rect 30156 31724 30212 31726
rect 30268 31500 30324 31556
rect 30268 31052 30324 31108
rect 30156 30322 30212 30324
rect 30156 30270 30158 30322
rect 30158 30270 30210 30322
rect 30210 30270 30212 30322
rect 30156 30268 30212 30270
rect 29484 29372 29540 29428
rect 29260 28082 29316 28084
rect 29260 28030 29262 28082
rect 29262 28030 29314 28082
rect 29314 28030 29316 28082
rect 29260 28028 29316 28030
rect 29372 27916 29428 27972
rect 29932 29372 29988 29428
rect 30492 30604 30548 30660
rect 29596 28588 29652 28644
rect 30716 31164 30772 31220
rect 31612 35810 31668 35812
rect 31612 35758 31614 35810
rect 31614 35758 31666 35810
rect 31666 35758 31668 35810
rect 31612 35756 31668 35758
rect 31276 35644 31332 35700
rect 31052 33516 31108 33572
rect 29708 28028 29764 28084
rect 30268 28082 30324 28084
rect 30268 28030 30270 28082
rect 30270 28030 30322 28082
rect 30322 28030 30324 28082
rect 30268 28028 30324 28030
rect 28924 26684 28980 26740
rect 28476 25618 28532 25620
rect 28476 25566 28478 25618
rect 28478 25566 28530 25618
rect 28530 25566 28532 25618
rect 28476 25564 28532 25566
rect 28140 25452 28196 25508
rect 27804 25004 27860 25060
rect 28028 24892 28084 24948
rect 27356 23938 27412 23940
rect 27356 23886 27358 23938
rect 27358 23886 27410 23938
rect 27410 23886 27412 23938
rect 27356 23884 27412 23886
rect 29148 26290 29204 26292
rect 29148 26238 29150 26290
rect 29150 26238 29202 26290
rect 29202 26238 29204 26290
rect 29148 26236 29204 26238
rect 28700 24556 28756 24612
rect 27580 23884 27636 23940
rect 27020 21084 27076 21140
rect 26684 20524 26740 20580
rect 27132 20076 27188 20132
rect 26124 19122 26180 19124
rect 26124 19070 26126 19122
rect 26126 19070 26178 19122
rect 26178 19070 26180 19122
rect 26124 19068 26180 19070
rect 27132 19068 27188 19124
rect 26796 18956 26852 19012
rect 26572 18732 26628 18788
rect 26348 18172 26404 18228
rect 25004 17836 25060 17892
rect 25228 16828 25284 16884
rect 25340 17500 25396 17556
rect 25228 15260 25284 15316
rect 25004 13916 25060 13972
rect 25004 13244 25060 13300
rect 25116 12850 25172 12852
rect 25116 12798 25118 12850
rect 25118 12798 25170 12850
rect 25170 12798 25172 12850
rect 25116 12796 25172 12798
rect 27132 18732 27188 18788
rect 26684 18450 26740 18452
rect 26684 18398 26686 18450
rect 26686 18398 26738 18450
rect 26738 18398 26740 18450
rect 26684 18396 26740 18398
rect 27020 18284 27076 18340
rect 25452 16380 25508 16436
rect 26012 17388 26068 17444
rect 25788 17106 25844 17108
rect 25788 17054 25790 17106
rect 25790 17054 25842 17106
rect 25842 17054 25844 17106
rect 25788 17052 25844 17054
rect 25564 16716 25620 16772
rect 25676 16828 25732 16884
rect 26908 17500 26964 17556
rect 26796 16716 26852 16772
rect 25564 16044 25620 16100
rect 25900 15260 25956 15316
rect 25340 14812 25396 14868
rect 26012 14418 26068 14420
rect 26012 14366 26014 14418
rect 26014 14366 26066 14418
rect 26066 14366 26068 14418
rect 26012 14364 26068 14366
rect 26012 14140 26068 14196
rect 25564 13970 25620 13972
rect 25564 13918 25566 13970
rect 25566 13918 25618 13970
rect 25618 13918 25620 13970
rect 25564 13916 25620 13918
rect 25340 13692 25396 13748
rect 22092 10498 22148 10500
rect 22092 10446 22094 10498
rect 22094 10446 22146 10498
rect 22146 10446 22148 10498
rect 22092 10444 22148 10446
rect 23660 10108 23716 10164
rect 22652 9772 22708 9828
rect 21868 9602 21924 9604
rect 21868 9550 21870 9602
rect 21870 9550 21922 9602
rect 21922 9550 21924 9602
rect 21868 9548 21924 9550
rect 21084 9324 21140 9380
rect 22988 9266 23044 9268
rect 22988 9214 22990 9266
rect 22990 9214 23042 9266
rect 23042 9214 23044 9266
rect 22988 9212 23044 9214
rect 23436 9212 23492 9268
rect 19292 8204 19348 8260
rect 23884 9772 23940 9828
rect 24668 9548 24724 9604
rect 24108 9154 24164 9156
rect 24108 9102 24110 9154
rect 24110 9102 24162 9154
rect 24162 9102 24164 9154
rect 24108 9100 24164 9102
rect 20076 8204 20132 8260
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 18508 7420 18564 7476
rect 18284 6524 18340 6580
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 17836 3948 17892 4004
rect 18396 3948 18452 4004
rect 18060 3724 18116 3780
rect 18172 3388 18228 3444
rect 25340 11452 25396 11508
rect 27580 23266 27636 23268
rect 27580 23214 27582 23266
rect 27582 23214 27634 23266
rect 27634 23214 27636 23266
rect 27580 23212 27636 23214
rect 27692 23100 27748 23156
rect 29484 25004 29540 25060
rect 30492 27580 30548 27636
rect 30492 27356 30548 27412
rect 29708 25676 29764 25732
rect 29820 25228 29876 25284
rect 30940 33404 30996 33460
rect 30828 30044 30884 30100
rect 31500 35196 31556 35252
rect 31388 34802 31444 34804
rect 31388 34750 31390 34802
rect 31390 34750 31442 34802
rect 31442 34750 31444 34802
rect 31388 34748 31444 34750
rect 32508 36988 32564 37044
rect 32732 36652 32788 36708
rect 32172 36428 32228 36484
rect 31836 36258 31892 36260
rect 31836 36206 31838 36258
rect 31838 36206 31890 36258
rect 31890 36206 31892 36258
rect 31836 36204 31892 36206
rect 33180 40236 33236 40292
rect 33852 40402 33908 40404
rect 33852 40350 33854 40402
rect 33854 40350 33906 40402
rect 33906 40350 33908 40402
rect 33852 40348 33908 40350
rect 34412 44604 34468 44660
rect 34972 47404 35028 47460
rect 35196 47068 35252 47124
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 36092 48524 36148 48580
rect 36988 49698 37044 49700
rect 36988 49646 36990 49698
rect 36990 49646 37042 49698
rect 37042 49646 37044 49698
rect 36988 49644 37044 49646
rect 36764 48636 36820 48692
rect 36428 48076 36484 48132
rect 35756 47516 35812 47572
rect 36092 47458 36148 47460
rect 36092 47406 36094 47458
rect 36094 47406 36146 47458
rect 36146 47406 36148 47458
rect 36092 47404 36148 47406
rect 36876 48300 36932 48356
rect 37548 50652 37604 50708
rect 39564 51266 39620 51268
rect 39564 51214 39566 51266
rect 39566 51214 39618 51266
rect 39618 51214 39620 51266
rect 39564 51212 39620 51214
rect 39004 51100 39060 51156
rect 38332 50652 38388 50708
rect 38892 50764 38948 50820
rect 38220 50428 38276 50484
rect 37548 49756 37604 49812
rect 38332 49532 38388 49588
rect 38108 49026 38164 49028
rect 38108 48974 38110 49026
rect 38110 48974 38162 49026
rect 38162 48974 38164 49026
rect 38108 48972 38164 48974
rect 37436 48748 37492 48804
rect 37996 48636 38052 48692
rect 37660 48300 37716 48356
rect 36988 48130 37044 48132
rect 36988 48078 36990 48130
rect 36990 48078 37042 48130
rect 37042 48078 37044 48130
rect 36988 48076 37044 48078
rect 36876 47628 36932 47684
rect 38444 48748 38500 48804
rect 37436 47628 37492 47684
rect 36428 47404 36484 47460
rect 36316 47346 36372 47348
rect 36316 47294 36318 47346
rect 36318 47294 36370 47346
rect 36370 47294 36372 47346
rect 36316 47292 36372 47294
rect 35756 47068 35812 47124
rect 36092 47180 36148 47236
rect 35868 45836 35924 45892
rect 35532 45724 35588 45780
rect 34860 45612 34916 45668
rect 34748 45276 34804 45332
rect 35084 45106 35140 45108
rect 35084 45054 35086 45106
rect 35086 45054 35138 45106
rect 35138 45054 35140 45106
rect 35084 45052 35140 45054
rect 34748 44940 34804 44996
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35756 44716 35812 44772
rect 35404 44660 35460 44662
rect 34524 44268 34580 44324
rect 34412 43708 34468 43764
rect 34412 43484 34468 43540
rect 34860 44156 34916 44212
rect 34748 44044 34804 44100
rect 35308 43708 35364 43764
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35532 42812 35588 42868
rect 34748 42700 34804 42756
rect 35420 42754 35476 42756
rect 35420 42702 35422 42754
rect 35422 42702 35474 42754
rect 35474 42702 35476 42754
rect 35420 42700 35476 42702
rect 34748 42530 34804 42532
rect 34748 42478 34750 42530
rect 34750 42478 34802 42530
rect 34802 42478 34804 42530
rect 34748 42476 34804 42478
rect 34524 42140 34580 42196
rect 33516 39900 33572 39956
rect 33964 39506 34020 39508
rect 33964 39454 33966 39506
rect 33966 39454 34018 39506
rect 34018 39454 34020 39506
rect 33964 39452 34020 39454
rect 34188 39116 34244 39172
rect 33964 39058 34020 39060
rect 33964 39006 33966 39058
rect 33966 39006 34018 39058
rect 34018 39006 34020 39058
rect 33964 39004 34020 39006
rect 34300 39058 34356 39060
rect 34300 39006 34302 39058
rect 34302 39006 34354 39058
rect 34354 39006 34356 39058
rect 34300 39004 34356 39006
rect 33516 37996 33572 38052
rect 33964 37826 34020 37828
rect 33964 37774 33966 37826
rect 33966 37774 34018 37826
rect 34018 37774 34020 37826
rect 33964 37772 34020 37774
rect 33068 37548 33124 37604
rect 33180 37436 33236 37492
rect 33404 37548 33460 37604
rect 33852 37548 33908 37604
rect 33292 36988 33348 37044
rect 33404 36540 33460 36596
rect 32732 35644 32788 35700
rect 32508 35196 32564 35252
rect 32956 35532 33012 35588
rect 31724 35084 31780 35140
rect 33740 35196 33796 35252
rect 31612 34018 31668 34020
rect 31612 33966 31614 34018
rect 31614 33966 31666 34018
rect 31666 33966 31668 34018
rect 31612 33964 31668 33966
rect 33740 34636 33796 34692
rect 32284 33964 32340 34020
rect 31276 33404 31332 33460
rect 33628 33852 33684 33908
rect 31276 33234 31332 33236
rect 31276 33182 31278 33234
rect 31278 33182 31330 33234
rect 31330 33182 31332 33234
rect 31276 33180 31332 33182
rect 31724 33180 31780 33236
rect 32508 33234 32564 33236
rect 32508 33182 32510 33234
rect 32510 33182 32562 33234
rect 32562 33182 32564 33234
rect 32508 33180 32564 33182
rect 32060 33068 32116 33124
rect 31388 32620 31444 32676
rect 31052 32284 31108 32340
rect 31164 30882 31220 30884
rect 31164 30830 31166 30882
rect 31166 30830 31218 30882
rect 31218 30830 31220 30882
rect 31164 30828 31220 30830
rect 31500 30604 31556 30660
rect 30940 29426 30996 29428
rect 30940 29374 30942 29426
rect 30942 29374 30994 29426
rect 30994 29374 30996 29426
rect 30940 29372 30996 29374
rect 31052 29314 31108 29316
rect 31052 29262 31054 29314
rect 31054 29262 31106 29314
rect 31106 29262 31108 29314
rect 31052 29260 31108 29262
rect 30828 28754 30884 28756
rect 30828 28702 30830 28754
rect 30830 28702 30882 28754
rect 30882 28702 30884 28754
rect 30828 28700 30884 28702
rect 31836 32284 31892 32340
rect 32172 31666 32228 31668
rect 32172 31614 32174 31666
rect 32174 31614 32226 31666
rect 32226 31614 32228 31666
rect 32172 31612 32228 31614
rect 31948 31164 32004 31220
rect 31724 31106 31780 31108
rect 31724 31054 31726 31106
rect 31726 31054 31778 31106
rect 31778 31054 31780 31106
rect 31724 31052 31780 31054
rect 31836 30994 31892 30996
rect 31836 30942 31838 30994
rect 31838 30942 31890 30994
rect 31890 30942 31892 30994
rect 31836 30940 31892 30942
rect 31948 30716 32004 30772
rect 31612 30380 31668 30436
rect 31612 30210 31668 30212
rect 31612 30158 31614 30210
rect 31614 30158 31666 30210
rect 31666 30158 31668 30210
rect 31612 30156 31668 30158
rect 31836 30044 31892 30100
rect 32956 33122 33012 33124
rect 32956 33070 32958 33122
rect 32958 33070 33010 33122
rect 33010 33070 33012 33122
rect 32956 33068 33012 33070
rect 32956 32508 33012 32564
rect 33180 31164 33236 31220
rect 33068 30044 33124 30100
rect 33516 30770 33572 30772
rect 33516 30718 33518 30770
rect 33518 30718 33570 30770
rect 33570 30718 33572 30770
rect 33516 30716 33572 30718
rect 34076 36540 34132 36596
rect 35084 42140 35140 42196
rect 35084 41970 35140 41972
rect 35084 41918 35086 41970
rect 35086 41918 35138 41970
rect 35138 41918 35140 41970
rect 35084 41916 35140 41918
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35868 42252 35924 42308
rect 35644 40962 35700 40964
rect 35644 40910 35646 40962
rect 35646 40910 35698 40962
rect 35698 40910 35700 40962
rect 35644 40908 35700 40910
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34860 39394 34916 39396
rect 34860 39342 34862 39394
rect 34862 39342 34914 39394
rect 34914 39342 34916 39394
rect 34860 39340 34916 39342
rect 34300 37938 34356 37940
rect 34300 37886 34302 37938
rect 34302 37886 34354 37938
rect 34354 37886 34356 37938
rect 34300 37884 34356 37886
rect 34636 37826 34692 37828
rect 34636 37774 34638 37826
rect 34638 37774 34690 37826
rect 34690 37774 34692 37826
rect 34636 37772 34692 37774
rect 34412 37490 34468 37492
rect 34412 37438 34414 37490
rect 34414 37438 34466 37490
rect 34466 37438 34468 37490
rect 34412 37436 34468 37438
rect 34412 36988 34468 37044
rect 34300 36370 34356 36372
rect 34300 36318 34302 36370
rect 34302 36318 34354 36370
rect 34354 36318 34356 36370
rect 34300 36316 34356 36318
rect 34524 36652 34580 36708
rect 34636 36482 34692 36484
rect 34636 36430 34638 36482
rect 34638 36430 34690 36482
rect 34690 36430 34692 36482
rect 34636 36428 34692 36430
rect 35308 39340 35364 39396
rect 35868 40908 35924 40964
rect 35868 39618 35924 39620
rect 35868 39566 35870 39618
rect 35870 39566 35922 39618
rect 35922 39566 35924 39618
rect 35868 39564 35924 39566
rect 37436 47404 37492 47460
rect 36764 47180 36820 47236
rect 36652 46674 36708 46676
rect 36652 46622 36654 46674
rect 36654 46622 36706 46674
rect 36706 46622 36708 46674
rect 36652 46620 36708 46622
rect 36204 46562 36260 46564
rect 36204 46510 36206 46562
rect 36206 46510 36258 46562
rect 36258 46510 36260 46562
rect 36204 46508 36260 46510
rect 37100 46508 37156 46564
rect 36204 45948 36260 46004
rect 37324 46396 37380 46452
rect 36316 43484 36372 43540
rect 37772 47346 37828 47348
rect 37772 47294 37774 47346
rect 37774 47294 37826 47346
rect 37826 47294 37828 47346
rect 37772 47292 37828 47294
rect 37884 47180 37940 47236
rect 37996 46956 38052 47012
rect 37884 46674 37940 46676
rect 37884 46622 37886 46674
rect 37886 46622 37938 46674
rect 37938 46622 37940 46674
rect 37884 46620 37940 46622
rect 38332 46508 38388 46564
rect 37996 46060 38052 46116
rect 37772 43708 37828 43764
rect 37660 43538 37716 43540
rect 37660 43486 37662 43538
rect 37662 43486 37714 43538
rect 37714 43486 37716 43538
rect 37660 43484 37716 43486
rect 36428 41916 36484 41972
rect 37436 41356 37492 41412
rect 36092 40572 36148 40628
rect 36204 40908 36260 40964
rect 36988 40962 37044 40964
rect 36988 40910 36990 40962
rect 36990 40910 37042 40962
rect 37042 40910 37044 40962
rect 36988 40908 37044 40910
rect 38108 44546 38164 44548
rect 38108 44494 38110 44546
rect 38110 44494 38162 44546
rect 38162 44494 38164 44546
rect 38108 44492 38164 44494
rect 38780 47628 38836 47684
rect 38668 46060 38724 46116
rect 38668 44492 38724 44548
rect 37660 40908 37716 40964
rect 38556 44322 38612 44324
rect 38556 44270 38558 44322
rect 38558 44270 38610 44322
rect 38610 44270 38612 44322
rect 38556 44268 38612 44270
rect 36652 40796 36708 40852
rect 37100 40796 37156 40852
rect 37100 40348 37156 40404
rect 36652 40012 36708 40068
rect 35420 38946 35476 38948
rect 35420 38894 35422 38946
rect 35422 38894 35474 38946
rect 35474 38894 35476 38946
rect 35420 38892 35476 38894
rect 35420 38668 35476 38724
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34972 38108 35028 38164
rect 35644 38332 35700 38388
rect 35084 37884 35140 37940
rect 35196 37436 35252 37492
rect 35308 37324 35364 37380
rect 35308 36988 35364 37044
rect 35644 36988 35700 37044
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35980 38946 36036 38948
rect 35980 38894 35982 38946
rect 35982 38894 36034 38946
rect 36034 38894 36036 38946
rect 35980 38892 36036 38894
rect 35980 38108 36036 38164
rect 35980 37324 36036 37380
rect 36540 39340 36596 39396
rect 36652 38946 36708 38948
rect 36652 38894 36654 38946
rect 36654 38894 36706 38946
rect 36706 38894 36708 38946
rect 36652 38892 36708 38894
rect 36988 38946 37044 38948
rect 36988 38894 36990 38946
rect 36990 38894 37042 38946
rect 37042 38894 37044 38946
rect 36988 38892 37044 38894
rect 36204 38332 36260 38388
rect 37212 39618 37268 39620
rect 37212 39566 37214 39618
rect 37214 39566 37266 39618
rect 37266 39566 37268 39618
rect 37212 39564 37268 39566
rect 37548 39676 37604 39732
rect 38668 43708 38724 43764
rect 39116 50594 39172 50596
rect 39116 50542 39118 50594
rect 39118 50542 39170 50594
rect 39170 50542 39172 50594
rect 39116 50540 39172 50542
rect 39004 48524 39060 48580
rect 38892 47404 38948 47460
rect 40124 53788 40180 53844
rect 40236 53058 40292 53060
rect 40236 53006 40238 53058
rect 40238 53006 40290 53058
rect 40290 53006 40292 53058
rect 40236 53004 40292 53006
rect 40236 52220 40292 52276
rect 41132 54572 41188 54628
rect 40908 54348 40964 54404
rect 42140 55244 42196 55300
rect 43260 56028 43316 56084
rect 42476 54684 42532 54740
rect 41020 53170 41076 53172
rect 41020 53118 41022 53170
rect 41022 53118 41074 53170
rect 41074 53118 41076 53170
rect 41020 53116 41076 53118
rect 41356 54514 41412 54516
rect 41356 54462 41358 54514
rect 41358 54462 41410 54514
rect 41410 54462 41412 54514
rect 41356 54460 41412 54462
rect 41468 53676 41524 53732
rect 42252 54124 42308 54180
rect 41916 53842 41972 53844
rect 41916 53790 41918 53842
rect 41918 53790 41970 53842
rect 41970 53790 41972 53842
rect 41916 53788 41972 53790
rect 42028 53004 42084 53060
rect 40796 51100 40852 51156
rect 41356 51324 41412 51380
rect 40908 50764 40964 50820
rect 41132 51212 41188 51268
rect 40796 50540 40852 50596
rect 41244 50482 41300 50484
rect 41244 50430 41246 50482
rect 41246 50430 41298 50482
rect 41298 50430 41300 50482
rect 41244 50428 41300 50430
rect 40348 49698 40404 49700
rect 40348 49646 40350 49698
rect 40350 49646 40402 49698
rect 40402 49646 40404 49698
rect 40348 49644 40404 49646
rect 39900 49084 39956 49140
rect 41020 49644 41076 49700
rect 39900 47628 39956 47684
rect 40460 48076 40516 48132
rect 40124 47964 40180 48020
rect 40124 47458 40180 47460
rect 40124 47406 40126 47458
rect 40126 47406 40178 47458
rect 40178 47406 40180 47458
rect 40124 47404 40180 47406
rect 40012 47180 40068 47236
rect 39004 46508 39060 46564
rect 38892 44604 38948 44660
rect 40012 46562 40068 46564
rect 40012 46510 40014 46562
rect 40014 46510 40066 46562
rect 40066 46510 40068 46562
rect 40012 46508 40068 46510
rect 40236 46002 40292 46004
rect 40236 45950 40238 46002
rect 40238 45950 40290 46002
rect 40290 45950 40292 46002
rect 40236 45948 40292 45950
rect 40124 45890 40180 45892
rect 40124 45838 40126 45890
rect 40126 45838 40178 45890
rect 40178 45838 40180 45890
rect 40124 45836 40180 45838
rect 39900 45666 39956 45668
rect 39900 45614 39902 45666
rect 39902 45614 39954 45666
rect 39954 45614 39956 45666
rect 39900 45612 39956 45614
rect 40460 47516 40516 47572
rect 40460 47234 40516 47236
rect 40460 47182 40462 47234
rect 40462 47182 40514 47234
rect 40514 47182 40516 47234
rect 40460 47180 40516 47182
rect 40908 46732 40964 46788
rect 40460 46620 40516 46676
rect 40460 46060 40516 46116
rect 42588 54514 42644 54516
rect 42588 54462 42590 54514
rect 42590 54462 42642 54514
rect 42642 54462 42644 54514
rect 42588 54460 42644 54462
rect 42588 53788 42644 53844
rect 42924 54348 42980 54404
rect 42924 54012 42980 54068
rect 42588 53506 42644 53508
rect 42588 53454 42590 53506
rect 42590 53454 42642 53506
rect 42642 53454 42644 53506
rect 42588 53452 42644 53454
rect 43148 53452 43204 53508
rect 42588 51324 42644 51380
rect 41916 50594 41972 50596
rect 41916 50542 41918 50594
rect 41918 50542 41970 50594
rect 41970 50542 41972 50594
rect 41916 50540 41972 50542
rect 41468 50316 41524 50372
rect 41692 49810 41748 49812
rect 41692 49758 41694 49810
rect 41694 49758 41746 49810
rect 41746 49758 41748 49810
rect 41692 49756 41748 49758
rect 42028 48860 42084 48916
rect 41804 48748 41860 48804
rect 42140 48412 42196 48468
rect 41356 48076 41412 48132
rect 41244 47404 41300 47460
rect 41468 47180 41524 47236
rect 43820 55468 43876 55524
rect 49532 56082 49588 56084
rect 49532 56030 49534 56082
rect 49534 56030 49586 56082
rect 49586 56030 49588 56082
rect 49532 56028 49588 56030
rect 50428 56082 50484 56084
rect 50428 56030 50430 56082
rect 50430 56030 50482 56082
rect 50482 56030 50484 56082
rect 50428 56028 50484 56030
rect 47628 55970 47684 55972
rect 47628 55918 47630 55970
rect 47630 55918 47682 55970
rect 47682 55918 47684 55970
rect 47628 55916 47684 55918
rect 43932 55186 43988 55188
rect 43932 55134 43934 55186
rect 43934 55134 43986 55186
rect 43986 55134 43988 55186
rect 43932 55132 43988 55134
rect 45052 54460 45108 54516
rect 43820 54012 43876 54068
rect 43596 53730 43652 53732
rect 43596 53678 43598 53730
rect 43598 53678 43650 53730
rect 43650 53678 43652 53730
rect 43596 53676 43652 53678
rect 45052 53676 45108 53732
rect 44156 53618 44212 53620
rect 44156 53566 44158 53618
rect 44158 53566 44210 53618
rect 44210 53566 44212 53618
rect 44156 53564 44212 53566
rect 43708 53004 43764 53060
rect 44044 53004 44100 53060
rect 43260 49532 43316 49588
rect 44156 51772 44212 51828
rect 43820 51378 43876 51380
rect 43820 51326 43822 51378
rect 43822 51326 43874 51378
rect 43874 51326 43876 51378
rect 43820 51324 43876 51326
rect 43372 50428 43428 50484
rect 44940 50482 44996 50484
rect 44940 50430 44942 50482
rect 44942 50430 44994 50482
rect 44994 50430 44996 50482
rect 44940 50428 44996 50430
rect 45052 50370 45108 50372
rect 45052 50318 45054 50370
rect 45054 50318 45106 50370
rect 45106 50318 45108 50370
rect 45052 50316 45108 50318
rect 44716 50092 44772 50148
rect 44604 49980 44660 50036
rect 42924 48860 42980 48916
rect 42476 48802 42532 48804
rect 42476 48750 42478 48802
rect 42478 48750 42530 48802
rect 42530 48750 42532 48802
rect 42476 48748 42532 48750
rect 42812 48466 42868 48468
rect 42812 48414 42814 48466
rect 42814 48414 42866 48466
rect 42866 48414 42868 48466
rect 42812 48412 42868 48414
rect 43596 48914 43652 48916
rect 43596 48862 43598 48914
rect 43598 48862 43650 48914
rect 43650 48862 43652 48914
rect 43596 48860 43652 48862
rect 44492 48860 44548 48916
rect 43036 48748 43092 48804
rect 41132 46674 41188 46676
rect 41132 46622 41134 46674
rect 41134 46622 41186 46674
rect 41186 46622 41188 46674
rect 41132 46620 41188 46622
rect 41916 46450 41972 46452
rect 41916 46398 41918 46450
rect 41918 46398 41970 46450
rect 41970 46398 41972 46450
rect 41916 46396 41972 46398
rect 41020 46284 41076 46340
rect 40796 46002 40852 46004
rect 40796 45950 40798 46002
rect 40798 45950 40850 46002
rect 40850 45950 40852 46002
rect 40796 45948 40852 45950
rect 42140 46284 42196 46340
rect 42140 46060 42196 46116
rect 41580 45836 41636 45892
rect 39340 44210 39396 44212
rect 39340 44158 39342 44210
rect 39342 44158 39394 44210
rect 39394 44158 39396 44210
rect 39340 44156 39396 44158
rect 38444 42530 38500 42532
rect 38444 42478 38446 42530
rect 38446 42478 38498 42530
rect 38498 42478 38500 42530
rect 38444 42476 38500 42478
rect 38892 42530 38948 42532
rect 38892 42478 38894 42530
rect 38894 42478 38946 42530
rect 38946 42478 38948 42530
rect 38892 42476 38948 42478
rect 42364 45836 42420 45892
rect 40236 44156 40292 44212
rect 40124 43650 40180 43652
rect 40124 43598 40126 43650
rect 40126 43598 40178 43650
rect 40178 43598 40180 43650
rect 40124 43596 40180 43598
rect 41020 43596 41076 43652
rect 40124 42140 40180 42196
rect 38220 41804 38276 41860
rect 38780 41804 38836 41860
rect 38444 41580 38500 41636
rect 38108 40684 38164 40740
rect 39676 41580 39732 41636
rect 38668 40684 38724 40740
rect 37772 39564 37828 39620
rect 37324 38892 37380 38948
rect 36204 37660 36260 37716
rect 35084 36258 35140 36260
rect 35084 36206 35086 36258
rect 35086 36206 35138 36258
rect 35138 36206 35140 36258
rect 35084 36204 35140 36206
rect 34188 35698 34244 35700
rect 34188 35646 34190 35698
rect 34190 35646 34242 35698
rect 34242 35646 34244 35698
rect 34188 35644 34244 35646
rect 34076 35532 34132 35588
rect 34300 34690 34356 34692
rect 34300 34638 34302 34690
rect 34302 34638 34354 34690
rect 34354 34638 34356 34690
rect 34300 34636 34356 34638
rect 33964 34524 34020 34580
rect 35532 36370 35588 36372
rect 35532 36318 35534 36370
rect 35534 36318 35586 36370
rect 35586 36318 35588 36370
rect 35532 36316 35588 36318
rect 35756 36316 35812 36372
rect 35644 36258 35700 36260
rect 35644 36206 35646 36258
rect 35646 36206 35698 36258
rect 35698 36206 35700 36258
rect 35644 36204 35700 36206
rect 35196 35532 35252 35588
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34412 34300 34468 34356
rect 34524 34972 34580 35028
rect 34412 34076 34468 34132
rect 34188 34018 34244 34020
rect 34188 33966 34190 34018
rect 34190 33966 34242 34018
rect 34242 33966 34244 34018
rect 34188 33964 34244 33966
rect 34748 34524 34804 34580
rect 35532 34636 35588 34692
rect 34972 34412 35028 34468
rect 34748 34018 34804 34020
rect 34748 33966 34750 34018
rect 34750 33966 34802 34018
rect 34802 33966 34804 34018
rect 34748 33964 34804 33966
rect 34972 33906 35028 33908
rect 34972 33854 34974 33906
rect 34974 33854 35026 33906
rect 35026 33854 35028 33906
rect 34972 33852 35028 33854
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 33852 33122 33908 33124
rect 33852 33070 33854 33122
rect 33854 33070 33906 33122
rect 33906 33070 33908 33122
rect 33852 33068 33908 33070
rect 33740 32508 33796 32564
rect 34300 33122 34356 33124
rect 34300 33070 34302 33122
rect 34302 33070 34354 33122
rect 34354 33070 34356 33122
rect 34300 33068 34356 33070
rect 33852 32396 33908 32452
rect 33964 31388 34020 31444
rect 34300 31388 34356 31444
rect 34188 30994 34244 30996
rect 34188 30942 34190 30994
rect 34190 30942 34242 30994
rect 34242 30942 34244 30994
rect 34188 30940 34244 30942
rect 33740 30156 33796 30212
rect 33852 30882 33908 30884
rect 33852 30830 33854 30882
rect 33854 30830 33906 30882
rect 33906 30830 33908 30882
rect 33852 30828 33908 30830
rect 32172 29708 32228 29764
rect 31836 29260 31892 29316
rect 31836 28700 31892 28756
rect 31164 27074 31220 27076
rect 31164 27022 31166 27074
rect 31166 27022 31218 27074
rect 31218 27022 31220 27074
rect 31164 27020 31220 27022
rect 30940 26962 30996 26964
rect 30940 26910 30942 26962
rect 30942 26910 30994 26962
rect 30994 26910 30996 26962
rect 30940 26908 30996 26910
rect 30604 26684 30660 26740
rect 33292 29538 33348 29540
rect 33292 29486 33294 29538
rect 33294 29486 33346 29538
rect 33346 29486 33348 29538
rect 33292 29484 33348 29486
rect 32956 29036 33012 29092
rect 32396 28754 32452 28756
rect 32396 28702 32398 28754
rect 32398 28702 32450 28754
rect 32450 28702 32452 28754
rect 32396 28700 32452 28702
rect 32060 28642 32116 28644
rect 32060 28590 32062 28642
rect 32062 28590 32114 28642
rect 32114 28590 32116 28642
rect 32060 28588 32116 28590
rect 31948 27858 32004 27860
rect 31948 27806 31950 27858
rect 31950 27806 32002 27858
rect 32002 27806 32004 27858
rect 31948 27804 32004 27806
rect 33292 29260 33348 29316
rect 33404 29148 33460 29204
rect 33404 28754 33460 28756
rect 33404 28702 33406 28754
rect 33406 28702 33458 28754
rect 33458 28702 33460 28754
rect 33404 28700 33460 28702
rect 33292 28588 33348 28644
rect 33628 28476 33684 28532
rect 32060 27468 32116 27524
rect 33180 27244 33236 27300
rect 32620 27132 32676 27188
rect 31612 27020 31668 27076
rect 32060 27074 32116 27076
rect 32060 27022 32062 27074
rect 32062 27022 32114 27074
rect 32114 27022 32116 27074
rect 32060 27020 32116 27022
rect 32284 27020 32340 27076
rect 31836 26962 31892 26964
rect 31836 26910 31838 26962
rect 31838 26910 31890 26962
rect 31890 26910 31892 26962
rect 31836 26908 31892 26910
rect 32956 26962 33012 26964
rect 32956 26910 32958 26962
rect 32958 26910 33010 26962
rect 33010 26910 33012 26962
rect 32956 26908 33012 26910
rect 33628 27186 33684 27188
rect 33628 27134 33630 27186
rect 33630 27134 33682 27186
rect 33682 27134 33684 27186
rect 33628 27132 33684 27134
rect 33852 29596 33908 29652
rect 35308 33068 35364 33124
rect 35420 32620 35476 32676
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35644 33628 35700 33684
rect 35868 34972 35924 35028
rect 36092 36652 36148 36708
rect 36316 36988 36372 37044
rect 36204 34130 36260 34132
rect 36204 34078 36206 34130
rect 36206 34078 36258 34130
rect 36258 34078 36260 34130
rect 36204 34076 36260 34078
rect 35980 33068 36036 33124
rect 35980 32396 36036 32452
rect 35868 31612 35924 31668
rect 37100 37996 37156 38052
rect 36988 37660 37044 37716
rect 36540 37324 36596 37380
rect 36428 34524 36484 34580
rect 36988 36652 37044 36708
rect 37772 38108 37828 38164
rect 38444 39618 38500 39620
rect 38444 39566 38446 39618
rect 38446 39566 38498 39618
rect 38498 39566 38500 39618
rect 38444 39564 38500 39566
rect 38444 39340 38500 39396
rect 37436 37378 37492 37380
rect 37436 37326 37438 37378
rect 37438 37326 37490 37378
rect 37490 37326 37492 37378
rect 37436 37324 37492 37326
rect 37100 36594 37156 36596
rect 37100 36542 37102 36594
rect 37102 36542 37154 36594
rect 37154 36542 37156 36594
rect 37100 36540 37156 36542
rect 36988 35868 37044 35924
rect 37772 37266 37828 37268
rect 37772 37214 37774 37266
rect 37774 37214 37826 37266
rect 37826 37214 37828 37266
rect 37772 37212 37828 37214
rect 38780 40348 38836 40404
rect 38892 39394 38948 39396
rect 38892 39342 38894 39394
rect 38894 39342 38946 39394
rect 38946 39342 38948 39394
rect 38892 39340 38948 39342
rect 38556 37212 38612 37268
rect 38220 37100 38276 37156
rect 39228 38444 39284 38500
rect 39004 36092 39060 36148
rect 37548 35532 37604 35588
rect 36540 34412 36596 34468
rect 37660 35084 37716 35140
rect 38108 35586 38164 35588
rect 38108 35534 38110 35586
rect 38110 35534 38162 35586
rect 38162 35534 38164 35586
rect 38108 35532 38164 35534
rect 37100 35026 37156 35028
rect 37100 34974 37102 35026
rect 37102 34974 37154 35026
rect 37154 34974 37156 35026
rect 37100 34972 37156 34974
rect 37100 34354 37156 34356
rect 37100 34302 37102 34354
rect 37102 34302 37154 34354
rect 37154 34302 37156 34354
rect 37100 34300 37156 34302
rect 36652 33964 36708 34020
rect 36540 33628 36596 33684
rect 36316 32620 36372 32676
rect 35868 30882 35924 30884
rect 35868 30830 35870 30882
rect 35870 30830 35922 30882
rect 35922 30830 35924 30882
rect 35868 30828 35924 30830
rect 35644 30770 35700 30772
rect 35644 30718 35646 30770
rect 35646 30718 35698 30770
rect 35698 30718 35700 30770
rect 35644 30716 35700 30718
rect 34636 30492 34692 30548
rect 36316 30604 36372 30660
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34412 30322 34468 30324
rect 34412 30270 34414 30322
rect 34414 30270 34466 30322
rect 34466 30270 34468 30322
rect 34412 30268 34468 30270
rect 35084 30268 35140 30324
rect 34524 30156 34580 30212
rect 34188 30044 34244 30100
rect 34300 29650 34356 29652
rect 34300 29598 34302 29650
rect 34302 29598 34354 29650
rect 34354 29598 34356 29650
rect 34300 29596 34356 29598
rect 34524 29484 34580 29540
rect 34412 29426 34468 29428
rect 34412 29374 34414 29426
rect 34414 29374 34466 29426
rect 34466 29374 34468 29426
rect 34412 29372 34468 29374
rect 33852 29148 33908 29204
rect 34412 28700 34468 28756
rect 34076 28588 34132 28644
rect 33964 27244 34020 27300
rect 30380 26124 30436 26180
rect 31500 26290 31556 26292
rect 31500 26238 31502 26290
rect 31502 26238 31554 26290
rect 31554 26238 31556 26290
rect 31500 26236 31556 26238
rect 29372 24332 29428 24388
rect 28812 22988 28868 23044
rect 29036 23266 29092 23268
rect 29036 23214 29038 23266
rect 29038 23214 29090 23266
rect 29090 23214 29092 23266
rect 29036 23212 29092 23214
rect 29148 22988 29204 23044
rect 29036 22876 29092 22932
rect 28364 22652 28420 22708
rect 29820 24610 29876 24612
rect 29820 24558 29822 24610
rect 29822 24558 29874 24610
rect 29874 24558 29876 24610
rect 29820 24556 29876 24558
rect 30268 24722 30324 24724
rect 30268 24670 30270 24722
rect 30270 24670 30322 24722
rect 30322 24670 30324 24722
rect 30268 24668 30324 24670
rect 30604 24050 30660 24052
rect 30604 23998 30606 24050
rect 30606 23998 30658 24050
rect 30658 23998 30660 24050
rect 30604 23996 30660 23998
rect 29372 22652 29428 22708
rect 28140 22540 28196 22596
rect 28588 22204 28644 22260
rect 28028 22092 28084 22148
rect 28252 21868 28308 21924
rect 29148 22092 29204 22148
rect 29148 21810 29204 21812
rect 29148 21758 29150 21810
rect 29150 21758 29202 21810
rect 29202 21758 29204 21810
rect 29148 21756 29204 21758
rect 28476 21698 28532 21700
rect 28476 21646 28478 21698
rect 28478 21646 28530 21698
rect 28530 21646 28532 21698
rect 28476 21644 28532 21646
rect 28028 21586 28084 21588
rect 28028 21534 28030 21586
rect 28030 21534 28082 21586
rect 28082 21534 28084 21586
rect 28028 21532 28084 21534
rect 28028 21196 28084 21252
rect 28364 21586 28420 21588
rect 28364 21534 28366 21586
rect 28366 21534 28418 21586
rect 28418 21534 28420 21586
rect 28364 21532 28420 21534
rect 28140 20748 28196 20804
rect 28476 21420 28532 21476
rect 28476 20860 28532 20916
rect 28364 20524 28420 20580
rect 28588 20578 28644 20580
rect 28588 20526 28590 20578
rect 28590 20526 28642 20578
rect 28642 20526 28644 20578
rect 28588 20524 28644 20526
rect 27916 20076 27972 20132
rect 29596 22988 29652 23044
rect 29708 22540 29764 22596
rect 29820 22876 29876 22932
rect 29596 22092 29652 22148
rect 30044 23154 30100 23156
rect 30044 23102 30046 23154
rect 30046 23102 30098 23154
rect 30098 23102 30100 23154
rect 30044 23100 30100 23102
rect 30044 22540 30100 22596
rect 29484 21586 29540 21588
rect 29484 21534 29486 21586
rect 29486 21534 29538 21586
rect 29538 21534 29540 21586
rect 29484 21532 29540 21534
rect 30044 20802 30100 20804
rect 30044 20750 30046 20802
rect 30046 20750 30098 20802
rect 30098 20750 30100 20802
rect 30044 20748 30100 20750
rect 29932 20690 29988 20692
rect 29932 20638 29934 20690
rect 29934 20638 29986 20690
rect 29986 20638 29988 20690
rect 29932 20636 29988 20638
rect 29484 20578 29540 20580
rect 29484 20526 29486 20578
rect 29486 20526 29538 20578
rect 29538 20526 29540 20578
rect 29484 20524 29540 20526
rect 28028 19234 28084 19236
rect 28028 19182 28030 19234
rect 28030 19182 28082 19234
rect 28082 19182 28084 19234
rect 28028 19180 28084 19182
rect 28588 19234 28644 19236
rect 28588 19182 28590 19234
rect 28590 19182 28642 19234
rect 28642 19182 28644 19234
rect 28588 19180 28644 19182
rect 27580 17666 27636 17668
rect 27580 17614 27582 17666
rect 27582 17614 27634 17666
rect 27634 17614 27636 17666
rect 27580 17612 27636 17614
rect 27468 17442 27524 17444
rect 27468 17390 27470 17442
rect 27470 17390 27522 17442
rect 27522 17390 27524 17442
rect 27468 17388 27524 17390
rect 28028 18226 28084 18228
rect 28028 18174 28030 18226
rect 28030 18174 28082 18226
rect 28082 18174 28084 18226
rect 28028 18172 28084 18174
rect 27692 16940 27748 16996
rect 27804 17612 27860 17668
rect 27356 16716 27412 16772
rect 27356 16492 27412 16548
rect 26348 14812 26404 14868
rect 26572 16098 26628 16100
rect 26572 16046 26574 16098
rect 26574 16046 26626 16098
rect 26626 16046 26628 16098
rect 26572 16044 26628 16046
rect 27020 16044 27076 16100
rect 26908 15314 26964 15316
rect 26908 15262 26910 15314
rect 26910 15262 26962 15314
rect 26962 15262 26964 15314
rect 26908 15260 26964 15262
rect 26908 14812 26964 14868
rect 26684 14530 26740 14532
rect 26684 14478 26686 14530
rect 26686 14478 26738 14530
rect 26738 14478 26740 14530
rect 26684 14476 26740 14478
rect 26796 14418 26852 14420
rect 26796 14366 26798 14418
rect 26798 14366 26850 14418
rect 26850 14366 26852 14418
rect 26796 14364 26852 14366
rect 27020 13916 27076 13972
rect 26012 13746 26068 13748
rect 26012 13694 26014 13746
rect 26014 13694 26066 13746
rect 26066 13694 26068 13746
rect 26012 13692 26068 13694
rect 26236 13356 26292 13412
rect 26572 13356 26628 13412
rect 26460 13020 26516 13076
rect 26012 12738 26068 12740
rect 26012 12686 26014 12738
rect 26014 12686 26066 12738
rect 26066 12686 26068 12738
rect 26012 12684 26068 12686
rect 26796 13020 26852 13076
rect 26908 12962 26964 12964
rect 26908 12910 26910 12962
rect 26910 12910 26962 12962
rect 26962 12910 26964 12962
rect 26908 12908 26964 12910
rect 27692 15986 27748 15988
rect 27692 15934 27694 15986
rect 27694 15934 27746 15986
rect 27746 15934 27748 15986
rect 27692 15932 27748 15934
rect 29036 18732 29092 18788
rect 29820 20578 29876 20580
rect 29820 20526 29822 20578
rect 29822 20526 29874 20578
rect 29874 20526 29876 20578
rect 29820 20524 29876 20526
rect 30492 23266 30548 23268
rect 30492 23214 30494 23266
rect 30494 23214 30546 23266
rect 30546 23214 30548 23266
rect 30492 23212 30548 23214
rect 30940 23212 30996 23268
rect 30492 22204 30548 22260
rect 31276 23996 31332 24052
rect 31388 23212 31444 23268
rect 31052 23100 31108 23156
rect 31500 23154 31556 23156
rect 31500 23102 31502 23154
rect 31502 23102 31554 23154
rect 31554 23102 31556 23154
rect 31500 23100 31556 23102
rect 31724 26684 31780 26740
rect 33964 26908 34020 26964
rect 33068 24722 33124 24724
rect 33068 24670 33070 24722
rect 33070 24670 33122 24722
rect 33122 24670 33124 24722
rect 33068 24668 33124 24670
rect 32284 24220 32340 24276
rect 33516 24722 33572 24724
rect 33516 24670 33518 24722
rect 33518 24670 33570 24722
rect 33570 24670 33572 24722
rect 33516 24668 33572 24670
rect 32060 23436 32116 23492
rect 32844 23660 32900 23716
rect 32508 23212 32564 23268
rect 31724 22988 31780 23044
rect 32060 22876 32116 22932
rect 30940 22316 30996 22372
rect 31500 22316 31556 22372
rect 30716 22092 30772 22148
rect 30492 21308 30548 21364
rect 31052 21868 31108 21924
rect 30828 21644 30884 21700
rect 31500 21810 31556 21812
rect 31500 21758 31502 21810
rect 31502 21758 31554 21810
rect 31554 21758 31556 21810
rect 31500 21756 31556 21758
rect 31836 22316 31892 22372
rect 33180 23436 33236 23492
rect 33068 23154 33124 23156
rect 33068 23102 33070 23154
rect 33070 23102 33122 23154
rect 33122 23102 33124 23154
rect 33068 23100 33124 23102
rect 32956 22876 33012 22932
rect 32284 22204 32340 22260
rect 32396 22316 32452 22372
rect 31836 22146 31892 22148
rect 31836 22094 31838 22146
rect 31838 22094 31890 22146
rect 31890 22094 31892 22146
rect 31836 22092 31892 22094
rect 31724 21756 31780 21812
rect 30716 21196 30772 21252
rect 30380 20300 30436 20356
rect 29708 19234 29764 19236
rect 29708 19182 29710 19234
rect 29710 19182 29762 19234
rect 29762 19182 29764 19234
rect 29708 19180 29764 19182
rect 28252 17948 28308 18004
rect 29372 17948 29428 18004
rect 28364 17666 28420 17668
rect 28364 17614 28366 17666
rect 28366 17614 28418 17666
rect 28418 17614 28420 17666
rect 28364 17612 28420 17614
rect 28588 17554 28644 17556
rect 28588 17502 28590 17554
rect 28590 17502 28642 17554
rect 28642 17502 28644 17554
rect 28588 17500 28644 17502
rect 28476 17442 28532 17444
rect 28476 17390 28478 17442
rect 28478 17390 28530 17442
rect 28530 17390 28532 17442
rect 28476 17388 28532 17390
rect 29148 17554 29204 17556
rect 29148 17502 29150 17554
rect 29150 17502 29202 17554
rect 29202 17502 29204 17554
rect 29148 17500 29204 17502
rect 28588 17276 28644 17332
rect 28476 16940 28532 16996
rect 28364 16716 28420 16772
rect 28028 15372 28084 15428
rect 27132 13858 27188 13860
rect 27132 13806 27134 13858
rect 27134 13806 27186 13858
rect 27186 13806 27188 13858
rect 27132 13804 27188 13806
rect 27244 15036 27300 15092
rect 26908 12684 26964 12740
rect 27580 14476 27636 14532
rect 27468 14364 27524 14420
rect 27916 14812 27972 14868
rect 29484 17164 29540 17220
rect 29484 16994 29540 16996
rect 29484 16942 29486 16994
rect 29486 16942 29538 16994
rect 29538 16942 29540 16994
rect 29484 16940 29540 16942
rect 28588 16658 28644 16660
rect 28588 16606 28590 16658
rect 28590 16606 28642 16658
rect 28642 16606 28644 16658
rect 28588 16604 28644 16606
rect 28812 15426 28868 15428
rect 28812 15374 28814 15426
rect 28814 15374 28866 15426
rect 28866 15374 28868 15426
rect 28812 15372 28868 15374
rect 27804 13522 27860 13524
rect 27804 13470 27806 13522
rect 27806 13470 27858 13522
rect 27858 13470 27860 13522
rect 27804 13468 27860 13470
rect 28924 13468 28980 13524
rect 28252 13356 28308 13412
rect 30156 18508 30212 18564
rect 30156 17948 30212 18004
rect 30268 17666 30324 17668
rect 30268 17614 30270 17666
rect 30270 17614 30322 17666
rect 30322 17614 30324 17666
rect 30268 17612 30324 17614
rect 30044 17276 30100 17332
rect 30492 17442 30548 17444
rect 30492 17390 30494 17442
rect 30494 17390 30546 17442
rect 30546 17390 30548 17442
rect 30492 17388 30548 17390
rect 29708 14364 29764 14420
rect 29372 13858 29428 13860
rect 29372 13806 29374 13858
rect 29374 13806 29426 13858
rect 29426 13806 29428 13858
rect 29372 13804 29428 13806
rect 29932 13580 29988 13636
rect 27356 12684 27412 12740
rect 28364 12962 28420 12964
rect 28364 12910 28366 12962
rect 28366 12910 28418 12962
rect 28418 12910 28420 12962
rect 28364 12908 28420 12910
rect 28140 12348 28196 12404
rect 28252 12236 28308 12292
rect 29148 12962 29204 12964
rect 29148 12910 29150 12962
rect 29150 12910 29202 12962
rect 29202 12910 29204 12962
rect 29148 12908 29204 12910
rect 28924 12348 28980 12404
rect 25900 11676 25956 11732
rect 27356 12178 27412 12180
rect 27356 12126 27358 12178
rect 27358 12126 27410 12178
rect 27410 12126 27412 12178
rect 27356 12124 27412 12126
rect 26012 11394 26068 11396
rect 26012 11342 26014 11394
rect 26014 11342 26066 11394
rect 26066 11342 26068 11394
rect 26012 11340 26068 11342
rect 26796 11676 26852 11732
rect 27580 11676 27636 11732
rect 27132 11506 27188 11508
rect 27132 11454 27134 11506
rect 27134 11454 27186 11506
rect 27186 11454 27188 11506
rect 27132 11452 27188 11454
rect 28364 11676 28420 11732
rect 26124 10668 26180 10724
rect 27244 10722 27300 10724
rect 27244 10670 27246 10722
rect 27246 10670 27298 10722
rect 27298 10670 27300 10722
rect 27244 10668 27300 10670
rect 25116 10108 25172 10164
rect 26796 10444 26852 10500
rect 25228 9548 25284 9604
rect 25228 9042 25284 9044
rect 25228 8990 25230 9042
rect 25230 8990 25282 9042
rect 25282 8990 25284 9042
rect 25228 8988 25284 8990
rect 26684 9212 26740 9268
rect 27244 9996 27300 10052
rect 27020 9826 27076 9828
rect 27020 9774 27022 9826
rect 27022 9774 27074 9826
rect 27074 9774 27076 9826
rect 27020 9772 27076 9774
rect 26796 9100 26852 9156
rect 27020 8988 27076 9044
rect 27804 9996 27860 10052
rect 29820 12402 29876 12404
rect 29820 12350 29822 12402
rect 29822 12350 29874 12402
rect 29874 12350 29876 12402
rect 29820 12348 29876 12350
rect 29148 12236 29204 12292
rect 29596 12290 29652 12292
rect 29596 12238 29598 12290
rect 29598 12238 29650 12290
rect 29650 12238 29652 12290
rect 29596 12236 29652 12238
rect 29484 12178 29540 12180
rect 29484 12126 29486 12178
rect 29486 12126 29538 12178
rect 29538 12126 29540 12178
rect 29484 12124 29540 12126
rect 29148 11228 29204 11284
rect 29932 11282 29988 11284
rect 29932 11230 29934 11282
rect 29934 11230 29986 11282
rect 29986 11230 29988 11282
rect 29932 11228 29988 11230
rect 28812 9996 28868 10052
rect 28028 9826 28084 9828
rect 28028 9774 28030 9826
rect 28030 9774 28082 9826
rect 28082 9774 28084 9826
rect 28028 9772 28084 9774
rect 27916 9602 27972 9604
rect 27916 9550 27918 9602
rect 27918 9550 27970 9602
rect 27970 9550 27972 9602
rect 27916 9548 27972 9550
rect 28252 9436 28308 9492
rect 28588 9548 28644 9604
rect 27692 9212 27748 9268
rect 30044 9996 30100 10052
rect 29484 9042 29540 9044
rect 29484 8990 29486 9042
rect 29486 8990 29538 9042
rect 29538 8990 29540 9042
rect 29484 8988 29540 8990
rect 18620 3388 18676 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 29596 3330 29652 3332
rect 29596 3278 29598 3330
rect 29598 3278 29650 3330
rect 29650 3278 29652 3330
rect 29596 3276 29652 3278
rect 30268 16994 30324 16996
rect 30268 16942 30270 16994
rect 30270 16942 30322 16994
rect 30322 16942 30324 16994
rect 30268 16940 30324 16942
rect 31052 20914 31108 20916
rect 31052 20862 31054 20914
rect 31054 20862 31106 20914
rect 31106 20862 31108 20914
rect 31052 20860 31108 20862
rect 31388 20860 31444 20916
rect 31500 21420 31556 21476
rect 31164 20524 31220 20580
rect 30940 18450 30996 18452
rect 30940 18398 30942 18450
rect 30942 18398 30994 18450
rect 30994 18398 30996 18450
rect 30940 18396 30996 18398
rect 30940 18060 30996 18116
rect 31052 17948 31108 18004
rect 30940 17724 30996 17780
rect 31052 17164 31108 17220
rect 31500 20412 31556 20468
rect 31276 19346 31332 19348
rect 31276 19294 31278 19346
rect 31278 19294 31330 19346
rect 31330 19294 31332 19346
rect 31276 19292 31332 19294
rect 33740 25900 33796 25956
rect 33964 26178 34020 26180
rect 33964 26126 33966 26178
rect 33966 26126 34018 26178
rect 34018 26126 34020 26178
rect 33964 26124 34020 26126
rect 34188 27244 34244 27300
rect 34412 25900 34468 25956
rect 34076 25228 34132 25284
rect 34188 25788 34244 25844
rect 33964 24668 34020 24724
rect 33628 23324 33684 23380
rect 33404 22594 33460 22596
rect 33404 22542 33406 22594
rect 33406 22542 33458 22594
rect 33458 22542 33460 22594
rect 33404 22540 33460 22542
rect 33628 22370 33684 22372
rect 33628 22318 33630 22370
rect 33630 22318 33682 22370
rect 33682 22318 33684 22370
rect 33628 22316 33684 22318
rect 32620 22092 32676 22148
rect 32956 22258 33012 22260
rect 32956 22206 32958 22258
rect 32958 22206 33010 22258
rect 33010 22206 33012 22258
rect 32956 22204 33012 22206
rect 32396 21980 32452 22036
rect 32172 21756 32228 21812
rect 32284 21362 32340 21364
rect 32284 21310 32286 21362
rect 32286 21310 32338 21362
rect 32338 21310 32340 21362
rect 32284 21308 32340 21310
rect 31612 19292 31668 19348
rect 33180 21868 33236 21924
rect 33180 20914 33236 20916
rect 33180 20862 33182 20914
rect 33182 20862 33234 20914
rect 33234 20862 33236 20914
rect 33180 20860 33236 20862
rect 32956 20300 33012 20356
rect 33292 19740 33348 19796
rect 32844 19234 32900 19236
rect 32844 19182 32846 19234
rect 32846 19182 32898 19234
rect 32898 19182 32900 19234
rect 32844 19180 32900 19182
rect 32060 18396 32116 18452
rect 31948 18338 32004 18340
rect 31948 18286 31950 18338
rect 31950 18286 32002 18338
rect 32002 18286 32004 18338
rect 31948 18284 32004 18286
rect 31388 17724 31444 17780
rect 31612 18172 31668 18228
rect 31276 16268 31332 16324
rect 31052 15372 31108 15428
rect 31276 15372 31332 15428
rect 30604 15090 30660 15092
rect 30604 15038 30606 15090
rect 30606 15038 30658 15090
rect 30658 15038 30660 15090
rect 30604 15036 30660 15038
rect 31164 13916 31220 13972
rect 31052 13804 31108 13860
rect 30940 13356 30996 13412
rect 30716 12908 30772 12964
rect 30940 12348 30996 12404
rect 30492 12236 30548 12292
rect 30268 11394 30324 11396
rect 30268 11342 30270 11394
rect 30270 11342 30322 11394
rect 30322 11342 30324 11394
rect 30268 11340 30324 11342
rect 30268 9042 30324 9044
rect 30268 8990 30270 9042
rect 30270 8990 30322 9042
rect 30322 8990 30324 9042
rect 30268 8988 30324 8990
rect 32060 17724 32116 17780
rect 31724 17554 31780 17556
rect 31724 17502 31726 17554
rect 31726 17502 31778 17554
rect 31778 17502 31780 17554
rect 31724 17500 31780 17502
rect 31836 15484 31892 15540
rect 31948 15372 32004 15428
rect 31612 15148 31668 15204
rect 32060 15036 32116 15092
rect 31612 13916 31668 13972
rect 31612 12962 31668 12964
rect 31612 12910 31614 12962
rect 31614 12910 31666 12962
rect 31666 12910 31668 12962
rect 31612 12908 31668 12910
rect 31388 12850 31444 12852
rect 31388 12798 31390 12850
rect 31390 12798 31442 12850
rect 31442 12798 31444 12850
rect 31388 12796 31444 12798
rect 31500 12572 31556 12628
rect 31612 12348 31668 12404
rect 31276 11394 31332 11396
rect 31276 11342 31278 11394
rect 31278 11342 31330 11394
rect 31330 11342 31332 11394
rect 31276 11340 31332 11342
rect 31500 11282 31556 11284
rect 31500 11230 31502 11282
rect 31502 11230 31554 11282
rect 31554 11230 31556 11282
rect 31500 11228 31556 11230
rect 31836 13356 31892 13412
rect 31948 12572 32004 12628
rect 32956 19010 33012 19012
rect 32956 18958 32958 19010
rect 32958 18958 33010 19010
rect 33010 18958 33012 19010
rect 32956 18956 33012 18958
rect 33068 18450 33124 18452
rect 33068 18398 33070 18450
rect 33070 18398 33122 18450
rect 33122 18398 33124 18450
rect 33068 18396 33124 18398
rect 32620 18284 32676 18340
rect 33180 18338 33236 18340
rect 33180 18286 33182 18338
rect 33182 18286 33234 18338
rect 33234 18286 33236 18338
rect 33180 18284 33236 18286
rect 32396 17666 32452 17668
rect 32396 17614 32398 17666
rect 32398 17614 32450 17666
rect 32450 17614 32452 17666
rect 32396 17612 32452 17614
rect 33292 17666 33348 17668
rect 33292 17614 33294 17666
rect 33294 17614 33346 17666
rect 33346 17614 33348 17666
rect 33292 17612 33348 17614
rect 33180 17388 33236 17444
rect 32508 16828 32564 16884
rect 32732 15986 32788 15988
rect 32732 15934 32734 15986
rect 32734 15934 32786 15986
rect 32786 15934 32788 15986
rect 32732 15932 32788 15934
rect 33180 16828 33236 16884
rect 33068 16322 33124 16324
rect 33068 16270 33070 16322
rect 33070 16270 33122 16322
rect 33122 16270 33124 16322
rect 33068 16268 33124 16270
rect 33628 22092 33684 22148
rect 33852 23212 33908 23268
rect 34076 23100 34132 23156
rect 33964 23042 34020 23044
rect 33964 22990 33966 23042
rect 33966 22990 34018 23042
rect 34018 22990 34020 23042
rect 33964 22988 34020 22990
rect 34076 22652 34132 22708
rect 33852 22540 33908 22596
rect 34076 22146 34132 22148
rect 34076 22094 34078 22146
rect 34078 22094 34130 22146
rect 34130 22094 34132 22146
rect 34076 22092 34132 22094
rect 33740 21644 33796 21700
rect 33964 21868 34020 21924
rect 33516 19234 33572 19236
rect 33516 19182 33518 19234
rect 33518 19182 33570 19234
rect 33570 19182 33572 19234
rect 33516 19180 33572 19182
rect 33516 18396 33572 18452
rect 33628 20076 33684 20132
rect 33628 16716 33684 16772
rect 33292 16492 33348 16548
rect 33068 15986 33124 15988
rect 33068 15934 33070 15986
rect 33070 15934 33122 15986
rect 33122 15934 33124 15986
rect 33068 15932 33124 15934
rect 33292 15820 33348 15876
rect 32620 15484 32676 15540
rect 32284 15426 32340 15428
rect 32284 15374 32286 15426
rect 32286 15374 32338 15426
rect 32338 15374 32340 15426
rect 32284 15372 32340 15374
rect 32396 15202 32452 15204
rect 32396 15150 32398 15202
rect 32398 15150 32450 15202
rect 32450 15150 32452 15202
rect 32396 15148 32452 15150
rect 31836 12348 31892 12404
rect 32060 12348 32116 12404
rect 32060 12066 32116 12068
rect 32060 12014 32062 12066
rect 32062 12014 32114 12066
rect 32114 12014 32116 12066
rect 32060 12012 32116 12014
rect 32508 12684 32564 12740
rect 32508 12290 32564 12292
rect 32508 12238 32510 12290
rect 32510 12238 32562 12290
rect 32562 12238 32564 12290
rect 32508 12236 32564 12238
rect 32172 11394 32228 11396
rect 32172 11342 32174 11394
rect 32174 11342 32226 11394
rect 32226 11342 32228 11394
rect 32172 11340 32228 11342
rect 31388 9660 31444 9716
rect 30268 3388 30324 3444
rect 31836 9714 31892 9716
rect 31836 9662 31838 9714
rect 31838 9662 31890 9714
rect 31890 9662 31892 9714
rect 31836 9660 31892 9662
rect 31500 8258 31556 8260
rect 31500 8206 31502 8258
rect 31502 8206 31554 8258
rect 31554 8206 31556 8258
rect 31500 8204 31556 8206
rect 32396 10556 32452 10612
rect 33068 15426 33124 15428
rect 33068 15374 33070 15426
rect 33070 15374 33122 15426
rect 33122 15374 33124 15426
rect 33068 15372 33124 15374
rect 33292 15036 33348 15092
rect 33292 14530 33348 14532
rect 33292 14478 33294 14530
rect 33294 14478 33346 14530
rect 33346 14478 33348 14530
rect 33292 14476 33348 14478
rect 33964 20802 34020 20804
rect 33964 20750 33966 20802
rect 33966 20750 34018 20802
rect 34018 20750 34020 20802
rect 33964 20748 34020 20750
rect 33964 17442 34020 17444
rect 33964 17390 33966 17442
rect 33966 17390 34018 17442
rect 34018 17390 34020 17442
rect 33964 17388 34020 17390
rect 34860 30210 34916 30212
rect 34860 30158 34862 30210
rect 34862 30158 34914 30210
rect 34914 30158 34916 30210
rect 34860 30156 34916 30158
rect 34860 29986 34916 29988
rect 34860 29934 34862 29986
rect 34862 29934 34914 29986
rect 34914 29934 34916 29986
rect 34860 29932 34916 29934
rect 35532 30156 35588 30212
rect 36764 33906 36820 33908
rect 36764 33854 36766 33906
rect 36766 33854 36818 33906
rect 36818 33854 36820 33906
rect 36764 33852 36820 33854
rect 37436 33628 37492 33684
rect 39564 38444 39620 38500
rect 41580 42924 41636 42980
rect 42140 45052 42196 45108
rect 42140 44268 42196 44324
rect 42140 43708 42196 43764
rect 42028 43314 42084 43316
rect 42028 43262 42030 43314
rect 42030 43262 42082 43314
rect 42082 43262 42084 43314
rect 42028 43260 42084 43262
rect 41580 42194 41636 42196
rect 41580 42142 41582 42194
rect 41582 42142 41634 42194
rect 41634 42142 41636 42194
rect 41580 42140 41636 42142
rect 41020 41356 41076 41412
rect 41580 41804 41636 41860
rect 41468 41356 41524 41412
rect 41468 40796 41524 40852
rect 40348 39900 40404 39956
rect 40348 38108 40404 38164
rect 41356 40514 41412 40516
rect 41356 40462 41358 40514
rect 41358 40462 41410 40514
rect 41410 40462 41412 40514
rect 41356 40460 41412 40462
rect 41692 41468 41748 41524
rect 41692 40626 41748 40628
rect 41692 40574 41694 40626
rect 41694 40574 41746 40626
rect 41746 40574 41748 40626
rect 41692 40572 41748 40574
rect 41580 40348 41636 40404
rect 41020 39788 41076 39844
rect 41244 39452 41300 39508
rect 40908 38108 40964 38164
rect 40572 37938 40628 37940
rect 40572 37886 40574 37938
rect 40574 37886 40626 37938
rect 40626 37886 40628 37938
rect 40572 37884 40628 37886
rect 40012 37548 40068 37604
rect 39340 37154 39396 37156
rect 39340 37102 39342 37154
rect 39342 37102 39394 37154
rect 39394 37102 39396 37154
rect 39340 37100 39396 37102
rect 39788 37266 39844 37268
rect 39788 37214 39790 37266
rect 39790 37214 39842 37266
rect 39842 37214 39844 37266
rect 39788 37212 39844 37214
rect 40348 37324 40404 37380
rect 41132 37378 41188 37380
rect 41132 37326 41134 37378
rect 41134 37326 41186 37378
rect 41186 37326 41188 37378
rect 41132 37324 41188 37326
rect 40908 37266 40964 37268
rect 40908 37214 40910 37266
rect 40910 37214 40962 37266
rect 40962 37214 40964 37266
rect 40908 37212 40964 37214
rect 39564 36482 39620 36484
rect 39564 36430 39566 36482
rect 39566 36430 39618 36482
rect 39618 36430 39620 36482
rect 39564 36428 39620 36430
rect 39676 35980 39732 36036
rect 40236 36482 40292 36484
rect 40236 36430 40238 36482
rect 40238 36430 40290 36482
rect 40290 36430 40292 36482
rect 40236 36428 40292 36430
rect 41020 37154 41076 37156
rect 41020 37102 41022 37154
rect 41022 37102 41074 37154
rect 41074 37102 41076 37154
rect 41020 37100 41076 37102
rect 40908 36876 40964 36932
rect 40236 35980 40292 36036
rect 37772 33852 37828 33908
rect 37100 33122 37156 33124
rect 37100 33070 37102 33122
rect 37102 33070 37154 33122
rect 37154 33070 37156 33122
rect 37100 33068 37156 33070
rect 39452 34914 39508 34916
rect 39452 34862 39454 34914
rect 39454 34862 39506 34914
rect 39506 34862 39508 34914
rect 39452 34860 39508 34862
rect 39228 34748 39284 34804
rect 38780 34690 38836 34692
rect 38780 34638 38782 34690
rect 38782 34638 38834 34690
rect 38834 34638 38836 34690
rect 38780 34636 38836 34638
rect 39004 33628 39060 33684
rect 37212 32450 37268 32452
rect 37212 32398 37214 32450
rect 37214 32398 37266 32450
rect 37266 32398 37268 32450
rect 37212 32396 37268 32398
rect 36764 32060 36820 32116
rect 36652 31164 36708 31220
rect 36764 30940 36820 30996
rect 36876 31724 36932 31780
rect 36540 30770 36596 30772
rect 36540 30718 36542 30770
rect 36542 30718 36594 30770
rect 36594 30718 36596 30770
rect 36540 30716 36596 30718
rect 35420 29820 35476 29876
rect 36092 29820 36148 29876
rect 36316 30156 36372 30212
rect 36428 29820 36484 29876
rect 35644 29708 35700 29764
rect 35196 29426 35252 29428
rect 35196 29374 35198 29426
rect 35198 29374 35250 29426
rect 35250 29374 35252 29426
rect 35196 29372 35252 29374
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34860 28700 34916 28756
rect 36652 29708 36708 29764
rect 35756 29036 35812 29092
rect 36316 29426 36372 29428
rect 36316 29374 36318 29426
rect 36318 29374 36370 29426
rect 36370 29374 36372 29426
rect 36316 29372 36372 29374
rect 36428 29314 36484 29316
rect 36428 29262 36430 29314
rect 36430 29262 36482 29314
rect 36482 29262 36484 29314
rect 36428 29260 36484 29262
rect 36988 31388 37044 31444
rect 36988 30492 37044 30548
rect 37100 31164 37156 31220
rect 37212 30882 37268 30884
rect 37212 30830 37214 30882
rect 37214 30830 37266 30882
rect 37266 30830 37268 30882
rect 37212 30828 37268 30830
rect 37212 30322 37268 30324
rect 37212 30270 37214 30322
rect 37214 30270 37266 30322
rect 37266 30270 37268 30322
rect 37212 30268 37268 30270
rect 36876 29260 36932 29316
rect 38332 32396 38388 32452
rect 38108 31164 38164 31220
rect 38108 30994 38164 30996
rect 38108 30942 38110 30994
rect 38110 30942 38162 30994
rect 38162 30942 38164 30994
rect 38108 30940 38164 30942
rect 37884 30716 37940 30772
rect 37436 30044 37492 30100
rect 37548 30492 37604 30548
rect 37548 29708 37604 29764
rect 36652 29036 36708 29092
rect 37548 29426 37604 29428
rect 37548 29374 37550 29426
rect 37550 29374 37602 29426
rect 37602 29374 37604 29426
rect 37548 29372 37604 29374
rect 35980 28924 36036 28980
rect 36428 28924 36484 28980
rect 36428 28700 36484 28756
rect 36764 28700 36820 28756
rect 35532 28642 35588 28644
rect 35532 28590 35534 28642
rect 35534 28590 35586 28642
rect 35586 28590 35588 28642
rect 35532 28588 35588 28590
rect 35084 28530 35140 28532
rect 35084 28478 35086 28530
rect 35086 28478 35138 28530
rect 35138 28478 35140 28530
rect 35084 28476 35140 28478
rect 36316 28588 36372 28644
rect 35756 28476 35812 28532
rect 36204 28530 36260 28532
rect 36204 28478 36206 28530
rect 36206 28478 36258 28530
rect 36258 28478 36260 28530
rect 36204 28476 36260 28478
rect 36540 28642 36596 28644
rect 36540 28590 36542 28642
rect 36542 28590 36594 28642
rect 36594 28590 36596 28642
rect 36540 28588 36596 28590
rect 35868 28364 35924 28420
rect 36652 28364 36708 28420
rect 34748 27468 34804 27524
rect 35980 27692 36036 27748
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35308 27244 35364 27300
rect 34748 27132 34804 27188
rect 35756 27020 35812 27076
rect 34748 26962 34804 26964
rect 34748 26910 34750 26962
rect 34750 26910 34802 26962
rect 34802 26910 34804 26962
rect 34748 26908 34804 26910
rect 34636 26460 34692 26516
rect 35532 26460 35588 26516
rect 35084 26012 35140 26068
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34636 25116 34692 25172
rect 36316 27244 36372 27300
rect 36428 27074 36484 27076
rect 36428 27022 36430 27074
rect 36430 27022 36482 27074
rect 36482 27022 36484 27074
rect 36428 27020 36484 27022
rect 36428 26796 36484 26852
rect 36428 26514 36484 26516
rect 36428 26462 36430 26514
rect 36430 26462 36482 26514
rect 36482 26462 36484 26514
rect 36428 26460 36484 26462
rect 35980 26012 36036 26068
rect 35756 25676 35812 25732
rect 35084 24946 35140 24948
rect 35084 24894 35086 24946
rect 35086 24894 35138 24946
rect 35138 24894 35140 24946
rect 35084 24892 35140 24894
rect 34748 24834 34804 24836
rect 34748 24782 34750 24834
rect 34750 24782 34802 24834
rect 34802 24782 34804 24834
rect 34748 24780 34804 24782
rect 36092 24946 36148 24948
rect 36092 24894 36094 24946
rect 36094 24894 36146 24946
rect 36146 24894 36148 24946
rect 36092 24892 36148 24894
rect 35420 24834 35476 24836
rect 35420 24782 35422 24834
rect 35422 24782 35474 24834
rect 35474 24782 35476 24834
rect 35420 24780 35476 24782
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 36428 24834 36484 24836
rect 36428 24782 36430 24834
rect 36430 24782 36482 24834
rect 36482 24782 36484 24834
rect 36428 24780 36484 24782
rect 35756 24668 35812 24724
rect 34748 23714 34804 23716
rect 34748 23662 34750 23714
rect 34750 23662 34802 23714
rect 34802 23662 34804 23714
rect 34748 23660 34804 23662
rect 34636 23154 34692 23156
rect 34636 23102 34638 23154
rect 34638 23102 34690 23154
rect 34690 23102 34692 23154
rect 34636 23100 34692 23102
rect 34524 22988 34580 23044
rect 34412 22930 34468 22932
rect 34412 22878 34414 22930
rect 34414 22878 34466 22930
rect 34466 22878 34468 22930
rect 34412 22876 34468 22878
rect 34972 23042 35028 23044
rect 34972 22990 34974 23042
rect 34974 22990 35026 23042
rect 35026 22990 35028 23042
rect 34972 22988 35028 22990
rect 35196 23212 35252 23268
rect 34524 22652 34580 22708
rect 34300 22204 34356 22260
rect 34412 21868 34468 21924
rect 34300 21644 34356 21700
rect 34412 21196 34468 21252
rect 34300 17948 34356 18004
rect 34300 17388 34356 17444
rect 34412 20802 34468 20804
rect 34412 20750 34414 20802
rect 34414 20750 34466 20802
rect 34466 20750 34468 20802
rect 34412 20748 34468 20750
rect 34524 17276 34580 17332
rect 34412 17052 34468 17108
rect 33852 16044 33908 16100
rect 33852 15596 33908 15652
rect 33964 16716 34020 16772
rect 33516 15036 33572 15092
rect 33292 13858 33348 13860
rect 33292 13806 33294 13858
rect 33294 13806 33346 13858
rect 33346 13806 33348 13858
rect 33292 13804 33348 13806
rect 33404 12850 33460 12852
rect 33404 12798 33406 12850
rect 33406 12798 33458 12850
rect 33458 12798 33460 12850
rect 33404 12796 33460 12798
rect 33180 12402 33236 12404
rect 33180 12350 33182 12402
rect 33182 12350 33234 12402
rect 33234 12350 33236 12402
rect 33180 12348 33236 12350
rect 33404 12572 33460 12628
rect 33180 10610 33236 10612
rect 33180 10558 33182 10610
rect 33182 10558 33234 10610
rect 33234 10558 33236 10610
rect 33180 10556 33236 10558
rect 33068 9996 33124 10052
rect 33180 8204 33236 8260
rect 33180 7644 33236 7700
rect 33852 15148 33908 15204
rect 34300 15874 34356 15876
rect 34300 15822 34302 15874
rect 34302 15822 34354 15874
rect 34354 15822 34356 15874
rect 34300 15820 34356 15822
rect 34748 22540 34804 22596
rect 34860 22092 34916 22148
rect 34860 21810 34916 21812
rect 34860 21758 34862 21810
rect 34862 21758 34914 21810
rect 34914 21758 34916 21810
rect 34860 21756 34916 21758
rect 34748 20524 34804 20580
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35756 23042 35812 23044
rect 35756 22990 35758 23042
rect 35758 22990 35810 23042
rect 35810 22990 35812 23042
rect 35756 22988 35812 22990
rect 35868 22540 35924 22596
rect 35756 22204 35812 22260
rect 36204 22316 36260 22372
rect 35532 22146 35588 22148
rect 35532 22094 35534 22146
rect 35534 22094 35586 22146
rect 35586 22094 35588 22146
rect 35532 22092 35588 22094
rect 35868 21980 35924 22036
rect 35308 21308 35364 21364
rect 35868 21474 35924 21476
rect 35868 21422 35870 21474
rect 35870 21422 35922 21474
rect 35922 21422 35924 21474
rect 35868 21420 35924 21422
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 36204 21308 36260 21364
rect 36316 21868 36372 21924
rect 35196 20578 35252 20580
rect 35196 20526 35198 20578
rect 35198 20526 35250 20578
rect 35250 20526 35252 20578
rect 35196 20524 35252 20526
rect 35308 20188 35364 20244
rect 34972 20130 35028 20132
rect 34972 20078 34974 20130
rect 34974 20078 35026 20130
rect 35026 20078 35028 20130
rect 34972 20076 35028 20078
rect 34860 20018 34916 20020
rect 34860 19966 34862 20018
rect 34862 19966 34914 20018
rect 34914 19966 34916 20018
rect 34860 19964 34916 19966
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35868 20524 35924 20580
rect 36092 20802 36148 20804
rect 36092 20750 36094 20802
rect 36094 20750 36146 20802
rect 36146 20750 36148 20802
rect 36092 20748 36148 20750
rect 36092 20188 36148 20244
rect 36540 20412 36596 20468
rect 36316 20018 36372 20020
rect 36316 19966 36318 20018
rect 36318 19966 36370 20018
rect 36370 19966 36372 20018
rect 36316 19964 36372 19966
rect 35868 19292 35924 19348
rect 35756 18956 35812 19012
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 34748 17442 34804 17444
rect 34748 17390 34750 17442
rect 34750 17390 34802 17442
rect 34802 17390 34804 17442
rect 34748 17388 34804 17390
rect 34972 17276 35028 17332
rect 34860 16716 34916 16772
rect 34748 16098 34804 16100
rect 34748 16046 34750 16098
rect 34750 16046 34802 16098
rect 34802 16046 34804 16098
rect 34748 16044 34804 16046
rect 34188 15090 34244 15092
rect 34188 15038 34190 15090
rect 34190 15038 34242 15090
rect 34242 15038 34244 15090
rect 34188 15036 34244 15038
rect 34076 14924 34132 14980
rect 34076 14476 34132 14532
rect 34076 13746 34132 13748
rect 34076 13694 34078 13746
rect 34078 13694 34130 13746
rect 34130 13694 34132 13746
rect 34076 13692 34132 13694
rect 34524 13804 34580 13860
rect 33964 12290 34020 12292
rect 33964 12238 33966 12290
rect 33966 12238 34018 12290
rect 34018 12238 34020 12290
rect 33964 12236 34020 12238
rect 33628 11394 33684 11396
rect 33628 11342 33630 11394
rect 33630 11342 33682 11394
rect 33682 11342 33684 11394
rect 33628 11340 33684 11342
rect 32956 3500 33012 3556
rect 34300 12738 34356 12740
rect 34300 12686 34302 12738
rect 34302 12686 34354 12738
rect 34354 12686 34356 12738
rect 34300 12684 34356 12686
rect 34748 13468 34804 13524
rect 34188 12012 34244 12068
rect 34076 11788 34132 11844
rect 34524 11788 34580 11844
rect 34636 12124 34692 12180
rect 34300 11506 34356 11508
rect 34300 11454 34302 11506
rect 34302 11454 34354 11506
rect 34354 11454 34356 11506
rect 34300 11452 34356 11454
rect 34748 12012 34804 12068
rect 34524 10556 34580 10612
rect 34076 10332 34132 10388
rect 33740 9324 33796 9380
rect 33964 8428 34020 8484
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 36204 18732 36260 18788
rect 35868 18620 35924 18676
rect 36428 18620 36484 18676
rect 36428 18172 36484 18228
rect 36428 17276 36484 17332
rect 35756 16380 35812 16436
rect 35532 16098 35588 16100
rect 35532 16046 35534 16098
rect 35534 16046 35586 16098
rect 35586 16046 35588 16098
rect 35532 16044 35588 16046
rect 35196 15484 35252 15540
rect 35644 15932 35700 15988
rect 34972 14530 35028 14532
rect 34972 14478 34974 14530
rect 34974 14478 35026 14530
rect 35026 14478 35028 14530
rect 34972 14476 35028 14478
rect 35420 15202 35476 15204
rect 35420 15150 35422 15202
rect 35422 15150 35474 15202
rect 35474 15150 35476 15202
rect 35420 15148 35476 15150
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34972 14252 35028 14308
rect 34972 12290 35028 12292
rect 34972 12238 34974 12290
rect 34974 12238 35026 12290
rect 35026 12238 35028 12290
rect 34972 12236 35028 12238
rect 35980 15874 36036 15876
rect 35980 15822 35982 15874
rect 35982 15822 36034 15874
rect 36034 15822 36036 15874
rect 35980 15820 36036 15822
rect 35980 15538 36036 15540
rect 35980 15486 35982 15538
rect 35982 15486 36034 15538
rect 36034 15486 36036 15538
rect 35980 15484 36036 15486
rect 35756 15148 35812 15204
rect 35868 14812 35924 14868
rect 36092 14700 36148 14756
rect 35980 14140 36036 14196
rect 35420 13692 35476 13748
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 12684 35252 12740
rect 34972 12012 35028 12068
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 11506 35252 11508
rect 35196 11454 35198 11506
rect 35198 11454 35250 11506
rect 35250 11454 35252 11506
rect 35196 11452 35252 11454
rect 34860 11340 34916 11396
rect 35420 10668 35476 10724
rect 34524 9660 34580 9716
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 36316 14812 36372 14868
rect 36204 13468 36260 13524
rect 35868 10892 35924 10948
rect 35756 10610 35812 10612
rect 35756 10558 35758 10610
rect 35758 10558 35810 10610
rect 35810 10558 35812 10610
rect 35756 10556 35812 10558
rect 36876 26962 36932 26964
rect 36876 26910 36878 26962
rect 36878 26910 36930 26962
rect 36930 26910 36932 26962
rect 36876 26908 36932 26910
rect 36988 24332 37044 24388
rect 36988 23548 37044 23604
rect 37324 28924 37380 28980
rect 37436 28700 37492 28756
rect 37548 28588 37604 28644
rect 37772 30156 37828 30212
rect 38108 30380 38164 30436
rect 38220 30210 38276 30212
rect 38220 30158 38222 30210
rect 38222 30158 38274 30210
rect 38274 30158 38276 30210
rect 38220 30156 38276 30158
rect 38108 30044 38164 30100
rect 37996 29986 38052 29988
rect 37996 29934 37998 29986
rect 37998 29934 38050 29986
rect 38050 29934 38052 29986
rect 37996 29932 38052 29934
rect 38108 29820 38164 29876
rect 37884 29708 37940 29764
rect 37212 27580 37268 27636
rect 37324 27244 37380 27300
rect 37212 27020 37268 27076
rect 37212 26796 37268 26852
rect 37324 23436 37380 23492
rect 37100 22930 37156 22932
rect 37100 22878 37102 22930
rect 37102 22878 37154 22930
rect 37154 22878 37156 22930
rect 37100 22876 37156 22878
rect 36764 21474 36820 21476
rect 36764 21422 36766 21474
rect 36766 21422 36818 21474
rect 36818 21422 36820 21474
rect 36764 21420 36820 21422
rect 36764 19180 36820 19236
rect 36652 18956 36708 19012
rect 36652 18732 36708 18788
rect 38220 27746 38276 27748
rect 38220 27694 38222 27746
rect 38222 27694 38274 27746
rect 38274 27694 38276 27746
rect 38220 27692 38276 27694
rect 38108 27244 38164 27300
rect 37772 27074 37828 27076
rect 37772 27022 37774 27074
rect 37774 27022 37826 27074
rect 37826 27022 37828 27074
rect 37772 27020 37828 27022
rect 37772 26796 37828 26852
rect 39452 33180 39508 33236
rect 38892 32786 38948 32788
rect 38892 32734 38894 32786
rect 38894 32734 38946 32786
rect 38946 32734 38948 32786
rect 38892 32732 38948 32734
rect 39340 32786 39396 32788
rect 39340 32734 39342 32786
rect 39342 32734 39394 32786
rect 39394 32734 39396 32786
rect 39340 32732 39396 32734
rect 38444 31724 38500 31780
rect 38556 31836 38612 31892
rect 38556 30882 38612 30884
rect 38556 30830 38558 30882
rect 38558 30830 38610 30882
rect 38610 30830 38612 30882
rect 38556 30828 38612 30830
rect 39452 32172 39508 32228
rect 39452 31836 39508 31892
rect 39788 34748 39844 34804
rect 40012 35084 40068 35140
rect 39676 34636 39732 34692
rect 40124 34914 40180 34916
rect 40124 34862 40126 34914
rect 40126 34862 40178 34914
rect 40178 34862 40180 34914
rect 40124 34860 40180 34862
rect 40572 36092 40628 36148
rect 41580 39116 41636 39172
rect 42812 45106 42868 45108
rect 42812 45054 42814 45106
rect 42814 45054 42866 45106
rect 42866 45054 42868 45106
rect 42812 45052 42868 45054
rect 43708 46396 43764 46452
rect 44380 46284 44436 46340
rect 43708 45890 43764 45892
rect 43708 45838 43710 45890
rect 43710 45838 43762 45890
rect 43762 45838 43764 45890
rect 43708 45836 43764 45838
rect 43372 45612 43428 45668
rect 43148 45106 43204 45108
rect 43148 45054 43150 45106
rect 43150 45054 43202 45106
rect 43202 45054 43204 45106
rect 43148 45052 43204 45054
rect 43260 44994 43316 44996
rect 43260 44942 43262 44994
rect 43262 44942 43314 44994
rect 43314 44942 43316 44994
rect 43260 44940 43316 44942
rect 43260 44380 43316 44436
rect 42476 42700 42532 42756
rect 43036 44322 43092 44324
rect 43036 44270 43038 44322
rect 43038 44270 43090 44322
rect 43090 44270 43092 44322
rect 43036 44268 43092 44270
rect 42812 44098 42868 44100
rect 42812 44046 42814 44098
rect 42814 44046 42866 44098
rect 42866 44046 42868 44098
rect 42812 44044 42868 44046
rect 43484 45164 43540 45220
rect 43932 45164 43988 45220
rect 43708 45052 43764 45108
rect 43820 44994 43876 44996
rect 43820 44942 43822 44994
rect 43822 44942 43874 44994
rect 43874 44942 43876 44994
rect 43820 44940 43876 44942
rect 43820 44434 43876 44436
rect 43820 44382 43822 44434
rect 43822 44382 43874 44434
rect 43874 44382 43876 44434
rect 43820 44380 43876 44382
rect 43932 44044 43988 44100
rect 42364 42642 42420 42644
rect 42364 42590 42366 42642
rect 42366 42590 42418 42642
rect 42418 42590 42420 42642
rect 42364 42588 42420 42590
rect 42364 41804 42420 41860
rect 42028 40796 42084 40852
rect 42252 40572 42308 40628
rect 42588 40514 42644 40516
rect 42588 40462 42590 40514
rect 42590 40462 42642 40514
rect 42642 40462 42644 40514
rect 42588 40460 42644 40462
rect 42364 39340 42420 39396
rect 42028 37938 42084 37940
rect 42028 37886 42030 37938
rect 42030 37886 42082 37938
rect 42082 37886 42084 37938
rect 42028 37884 42084 37886
rect 41356 37490 41412 37492
rect 41356 37438 41358 37490
rect 41358 37438 41410 37490
rect 41410 37438 41412 37490
rect 41356 37436 41412 37438
rect 40908 35644 40964 35700
rect 41804 36988 41860 37044
rect 42364 38556 42420 38612
rect 41916 36876 41972 36932
rect 40908 35196 40964 35252
rect 40348 34690 40404 34692
rect 40348 34638 40350 34690
rect 40350 34638 40402 34690
rect 40402 34638 40404 34690
rect 40348 34636 40404 34638
rect 40348 33628 40404 33684
rect 40012 33068 40068 33124
rect 40684 32284 40740 32340
rect 40348 32060 40404 32116
rect 39676 31388 39732 31444
rect 39340 30716 39396 30772
rect 39676 30828 39732 30884
rect 40124 31052 40180 31108
rect 38668 30210 38724 30212
rect 38668 30158 38670 30210
rect 38670 30158 38722 30210
rect 38722 30158 38724 30210
rect 38668 30156 38724 30158
rect 38444 29708 38500 29764
rect 39452 29986 39508 29988
rect 39452 29934 39454 29986
rect 39454 29934 39506 29986
rect 39506 29934 39508 29986
rect 39452 29932 39508 29934
rect 38556 29596 38612 29652
rect 39004 29820 39060 29876
rect 39228 29708 39284 29764
rect 38780 29426 38836 29428
rect 38780 29374 38782 29426
rect 38782 29374 38834 29426
rect 38834 29374 38836 29426
rect 38780 29372 38836 29374
rect 39452 29426 39508 29428
rect 39452 29374 39454 29426
rect 39454 29374 39506 29426
rect 39506 29374 39508 29426
rect 39452 29372 39508 29374
rect 38556 29314 38612 29316
rect 38556 29262 38558 29314
rect 38558 29262 38610 29314
rect 38610 29262 38612 29314
rect 38556 29260 38612 29262
rect 39004 29260 39060 29316
rect 38444 28364 38500 28420
rect 37996 26348 38052 26404
rect 37772 25282 37828 25284
rect 37772 25230 37774 25282
rect 37774 25230 37826 25282
rect 37826 25230 37828 25282
rect 37772 25228 37828 25230
rect 37660 24780 37716 24836
rect 37548 22930 37604 22932
rect 37548 22878 37550 22930
rect 37550 22878 37602 22930
rect 37602 22878 37604 22930
rect 37548 22876 37604 22878
rect 37324 22092 37380 22148
rect 37100 19852 37156 19908
rect 37212 19964 37268 20020
rect 36764 18562 36820 18564
rect 36764 18510 36766 18562
rect 36766 18510 36818 18562
rect 36818 18510 36820 18562
rect 36764 18508 36820 18510
rect 36652 18060 36708 18116
rect 36876 16716 36932 16772
rect 38444 26796 38500 26852
rect 38668 27804 38724 27860
rect 38780 27746 38836 27748
rect 38780 27694 38782 27746
rect 38782 27694 38834 27746
rect 38834 27694 38836 27746
rect 38780 27692 38836 27694
rect 39004 28418 39060 28420
rect 39004 28366 39006 28418
rect 39006 28366 39058 28418
rect 39058 28366 39060 28418
rect 39004 28364 39060 28366
rect 39228 27858 39284 27860
rect 39228 27806 39230 27858
rect 39230 27806 39282 27858
rect 39282 27806 39284 27858
rect 39228 27804 39284 27806
rect 40236 30156 40292 30212
rect 40012 29986 40068 29988
rect 40012 29934 40014 29986
rect 40014 29934 40066 29986
rect 40066 29934 40068 29986
rect 40012 29932 40068 29934
rect 39900 27132 39956 27188
rect 38556 26348 38612 26404
rect 39228 25900 39284 25956
rect 39116 25788 39172 25844
rect 38780 25676 38836 25732
rect 38556 25394 38612 25396
rect 38556 25342 38558 25394
rect 38558 25342 38610 25394
rect 38610 25342 38612 25394
rect 38556 25340 38612 25342
rect 38332 25282 38388 25284
rect 38332 25230 38334 25282
rect 38334 25230 38386 25282
rect 38386 25230 38388 25282
rect 38332 25228 38388 25230
rect 37772 23324 37828 23380
rect 37436 20802 37492 20804
rect 37436 20750 37438 20802
rect 37438 20750 37490 20802
rect 37490 20750 37492 20802
rect 37436 20748 37492 20750
rect 37100 16268 37156 16324
rect 37324 18060 37380 18116
rect 37660 21474 37716 21476
rect 37660 21422 37662 21474
rect 37662 21422 37714 21474
rect 37714 21422 37716 21474
rect 37660 21420 37716 21422
rect 37660 21026 37716 21028
rect 37660 20974 37662 21026
rect 37662 20974 37714 21026
rect 37714 20974 37716 21026
rect 37660 20972 37716 20974
rect 37884 24668 37940 24724
rect 37996 23938 38052 23940
rect 37996 23886 37998 23938
rect 37998 23886 38050 23938
rect 38050 23886 38052 23938
rect 37996 23884 38052 23886
rect 37884 21980 37940 22036
rect 37996 23548 38052 23604
rect 38444 24498 38500 24500
rect 38444 24446 38446 24498
rect 38446 24446 38498 24498
rect 38498 24446 38500 24498
rect 38444 24444 38500 24446
rect 38220 23436 38276 23492
rect 38108 23324 38164 23380
rect 38108 22540 38164 22596
rect 38220 22092 38276 22148
rect 38108 21586 38164 21588
rect 38108 21534 38110 21586
rect 38110 21534 38162 21586
rect 38162 21534 38164 21586
rect 38108 21532 38164 21534
rect 38332 20972 38388 21028
rect 38108 19906 38164 19908
rect 38108 19854 38110 19906
rect 38110 19854 38162 19906
rect 38162 19854 38164 19906
rect 38108 19852 38164 19854
rect 37772 19292 37828 19348
rect 38108 19234 38164 19236
rect 38108 19182 38110 19234
rect 38110 19182 38162 19234
rect 38162 19182 38164 19234
rect 38108 19180 38164 19182
rect 37772 18732 37828 18788
rect 37548 18172 37604 18228
rect 37436 17276 37492 17332
rect 36988 15986 37044 15988
rect 36988 15934 36990 15986
rect 36990 15934 37042 15986
rect 37042 15934 37044 15986
rect 36988 15932 37044 15934
rect 37100 15484 37156 15540
rect 37548 16492 37604 16548
rect 37436 15932 37492 15988
rect 37324 15874 37380 15876
rect 37324 15822 37326 15874
rect 37326 15822 37378 15874
rect 37378 15822 37380 15874
rect 37324 15820 37380 15822
rect 37212 14530 37268 14532
rect 37212 14478 37214 14530
rect 37214 14478 37266 14530
rect 37266 14478 37268 14530
rect 37212 14476 37268 14478
rect 36988 14306 37044 14308
rect 36988 14254 36990 14306
rect 36990 14254 37042 14306
rect 37042 14254 37044 14306
rect 36988 14252 37044 14254
rect 36652 14140 36708 14196
rect 36764 13746 36820 13748
rect 36764 13694 36766 13746
rect 36766 13694 36818 13746
rect 36818 13694 36820 13746
rect 36764 13692 36820 13694
rect 36204 10834 36260 10836
rect 36204 10782 36206 10834
rect 36206 10782 36258 10834
rect 36258 10782 36260 10834
rect 36204 10780 36260 10782
rect 36652 13468 36708 13524
rect 36092 10610 36148 10612
rect 36092 10558 36094 10610
rect 36094 10558 36146 10610
rect 36146 10558 36148 10610
rect 36092 10556 36148 10558
rect 35980 10444 36036 10500
rect 35756 9714 35812 9716
rect 35756 9662 35758 9714
rect 35758 9662 35810 9714
rect 35810 9662 35812 9714
rect 35756 9660 35812 9662
rect 35084 9436 35140 9492
rect 34972 9266 35028 9268
rect 34972 9214 34974 9266
rect 34974 9214 35026 9266
rect 35026 9214 35028 9266
rect 34972 9212 35028 9214
rect 35196 9212 35252 9268
rect 35308 9154 35364 9156
rect 35308 9102 35310 9154
rect 35310 9102 35362 9154
rect 35362 9102 35364 9154
rect 35308 9100 35364 9102
rect 35868 9266 35924 9268
rect 35868 9214 35870 9266
rect 35870 9214 35922 9266
rect 35922 9214 35924 9266
rect 35868 9212 35924 9214
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35420 8428 35476 8484
rect 35532 7644 35588 7700
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35084 4956 35140 5012
rect 33516 3554 33572 3556
rect 33516 3502 33518 3554
rect 33518 3502 33570 3554
rect 33570 3502 33572 3554
rect 33516 3500 33572 3502
rect 34748 3724 34804 3780
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35420 3612 35476 3668
rect 35196 3388 35252 3444
rect 35756 3388 35812 3444
rect 36540 10780 36596 10836
rect 39116 25228 39172 25284
rect 39340 25788 39396 25844
rect 38780 23714 38836 23716
rect 38780 23662 38782 23714
rect 38782 23662 38834 23714
rect 38834 23662 38836 23714
rect 38780 23660 38836 23662
rect 38556 23436 38612 23492
rect 39116 23938 39172 23940
rect 39116 23886 39118 23938
rect 39118 23886 39170 23938
rect 39170 23886 39172 23938
rect 39116 23884 39172 23886
rect 38556 21980 38612 22036
rect 38668 21474 38724 21476
rect 38668 21422 38670 21474
rect 38670 21422 38722 21474
rect 38722 21422 38724 21474
rect 38668 21420 38724 21422
rect 38892 23154 38948 23156
rect 38892 23102 38894 23154
rect 38894 23102 38946 23154
rect 38946 23102 38948 23154
rect 38892 23100 38948 23102
rect 38892 22258 38948 22260
rect 38892 22206 38894 22258
rect 38894 22206 38946 22258
rect 38946 22206 38948 22258
rect 38892 22204 38948 22206
rect 39340 23154 39396 23156
rect 39340 23102 39342 23154
rect 39342 23102 39394 23154
rect 39394 23102 39396 23154
rect 39340 23100 39396 23102
rect 39116 22988 39172 23044
rect 39116 22540 39172 22596
rect 39228 22876 39284 22932
rect 40012 26460 40068 26516
rect 40124 27858 40180 27860
rect 40124 27806 40126 27858
rect 40126 27806 40178 27858
rect 40178 27806 40180 27858
rect 40124 27804 40180 27806
rect 40012 26236 40068 26292
rect 39788 25506 39844 25508
rect 39788 25454 39790 25506
rect 39790 25454 39842 25506
rect 39842 25454 39844 25506
rect 39788 25452 39844 25454
rect 40236 27468 40292 27524
rect 41916 36370 41972 36372
rect 41916 36318 41918 36370
rect 41918 36318 41970 36370
rect 41970 36318 41972 36370
rect 41916 36316 41972 36318
rect 41132 36092 41188 36148
rect 41804 36204 41860 36260
rect 41244 35922 41300 35924
rect 41244 35870 41246 35922
rect 41246 35870 41298 35922
rect 41298 35870 41300 35922
rect 41244 35868 41300 35870
rect 41468 35196 41524 35252
rect 41916 36092 41972 36148
rect 42252 36092 42308 36148
rect 42028 35698 42084 35700
rect 42028 35646 42030 35698
rect 42030 35646 42082 35698
rect 42082 35646 42084 35698
rect 42028 35644 42084 35646
rect 42028 34860 42084 34916
rect 42588 36652 42644 36708
rect 43820 43260 43876 43316
rect 42812 40124 42868 40180
rect 43148 39788 43204 39844
rect 42812 37996 42868 38052
rect 42812 36482 42868 36484
rect 42812 36430 42814 36482
rect 42814 36430 42866 36482
rect 42866 36430 42868 36482
rect 42812 36428 42868 36430
rect 42476 36258 42532 36260
rect 42476 36206 42478 36258
rect 42478 36206 42530 36258
rect 42530 36206 42532 36258
rect 42476 36204 42532 36206
rect 42364 34860 42420 34916
rect 41132 34300 41188 34356
rect 41692 34690 41748 34692
rect 41692 34638 41694 34690
rect 41694 34638 41746 34690
rect 41746 34638 41748 34690
rect 41692 34636 41748 34638
rect 42028 34300 42084 34356
rect 42028 33964 42084 34020
rect 41244 32284 41300 32340
rect 41020 31052 41076 31108
rect 40796 30828 40852 30884
rect 41020 30828 41076 30884
rect 40684 30210 40740 30212
rect 40684 30158 40686 30210
rect 40686 30158 40738 30210
rect 40738 30158 40740 30210
rect 40684 30156 40740 30158
rect 40684 29372 40740 29428
rect 40796 29036 40852 29092
rect 40908 27634 40964 27636
rect 40908 27582 40910 27634
rect 40910 27582 40962 27634
rect 40962 27582 40964 27634
rect 40908 27580 40964 27582
rect 40796 27020 40852 27076
rect 41244 28252 41300 28308
rect 41692 32562 41748 32564
rect 41692 32510 41694 32562
rect 41694 32510 41746 32562
rect 41746 32510 41748 32562
rect 41692 32508 41748 32510
rect 42812 35532 42868 35588
rect 42700 35308 42756 35364
rect 42924 34914 42980 34916
rect 42924 34862 42926 34914
rect 42926 34862 42978 34914
rect 42978 34862 42980 34914
rect 42924 34860 42980 34862
rect 43484 40460 43540 40516
rect 43932 40684 43988 40740
rect 44380 40908 44436 40964
rect 43372 40290 43428 40292
rect 43372 40238 43374 40290
rect 43374 40238 43426 40290
rect 43426 40238 43428 40290
rect 43372 40236 43428 40238
rect 43260 38668 43316 38724
rect 43260 36652 43316 36708
rect 43932 40290 43988 40292
rect 43932 40238 43934 40290
rect 43934 40238 43986 40290
rect 43986 40238 43988 40290
rect 43932 40236 43988 40238
rect 44268 40236 44324 40292
rect 43820 40124 43876 40180
rect 44940 49810 44996 49812
rect 44940 49758 44942 49810
rect 44942 49758 44994 49810
rect 44994 49758 44996 49810
rect 44940 49756 44996 49758
rect 49644 55356 49700 55412
rect 46396 55132 46452 55188
rect 45500 53788 45556 53844
rect 45388 53452 45444 53508
rect 45388 51324 45444 51380
rect 45724 53788 45780 53844
rect 45612 53452 45668 53508
rect 46396 54348 46452 54404
rect 46060 53564 46116 53620
rect 46172 53452 46228 53508
rect 46508 54012 46564 54068
rect 46060 51996 46116 52052
rect 46508 53564 46564 53620
rect 47292 53788 47348 53844
rect 47740 54514 47796 54516
rect 47740 54462 47742 54514
rect 47742 54462 47794 54514
rect 47794 54462 47796 54514
rect 47740 54460 47796 54462
rect 48188 54402 48244 54404
rect 48188 54350 48190 54402
rect 48190 54350 48242 54402
rect 48242 54350 48244 54402
rect 48188 54348 48244 54350
rect 51660 55410 51716 55412
rect 51660 55358 51662 55410
rect 51662 55358 51714 55410
rect 51714 55358 51716 55410
rect 51660 55356 51716 55358
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 49644 54460 49700 54516
rect 48412 53730 48468 53732
rect 48412 53678 48414 53730
rect 48414 53678 48466 53730
rect 48466 53678 48468 53730
rect 48412 53676 48468 53678
rect 47516 53564 47572 53620
rect 49532 53506 49588 53508
rect 49532 53454 49534 53506
rect 49534 53454 49586 53506
rect 49586 53454 49588 53506
rect 49532 53452 49588 53454
rect 47180 52780 47236 52836
rect 46620 52274 46676 52276
rect 46620 52222 46622 52274
rect 46622 52222 46674 52274
rect 46674 52222 46676 52274
rect 46620 52220 46676 52222
rect 48188 52834 48244 52836
rect 48188 52782 48190 52834
rect 48190 52782 48242 52834
rect 48242 52782 48244 52834
rect 48188 52780 48244 52782
rect 48748 52780 48804 52836
rect 47180 52220 47236 52276
rect 46060 51490 46116 51492
rect 46060 51438 46062 51490
rect 46062 51438 46114 51490
rect 46114 51438 46116 51490
rect 46060 51436 46116 51438
rect 46620 51378 46676 51380
rect 46620 51326 46622 51378
rect 46622 51326 46674 51378
rect 46674 51326 46676 51378
rect 46620 51324 46676 51326
rect 45276 49980 45332 50036
rect 45388 49810 45444 49812
rect 45388 49758 45390 49810
rect 45390 49758 45442 49810
rect 45442 49758 45444 49810
rect 45388 49756 45444 49758
rect 45164 48802 45220 48804
rect 45164 48750 45166 48802
rect 45166 48750 45218 48802
rect 45218 48750 45220 48802
rect 45164 48748 45220 48750
rect 46396 48748 46452 48804
rect 44940 47234 44996 47236
rect 44940 47182 44942 47234
rect 44942 47182 44994 47234
rect 44994 47182 44996 47234
rect 44940 47180 44996 47182
rect 46060 47068 46116 47124
rect 45052 46284 45108 46340
rect 45164 45890 45220 45892
rect 45164 45838 45166 45890
rect 45166 45838 45218 45890
rect 45218 45838 45220 45890
rect 45164 45836 45220 45838
rect 45836 46172 45892 46228
rect 45388 45778 45444 45780
rect 45388 45726 45390 45778
rect 45390 45726 45442 45778
rect 45442 45726 45444 45778
rect 45388 45724 45444 45726
rect 45164 45218 45220 45220
rect 45164 45166 45166 45218
rect 45166 45166 45218 45218
rect 45218 45166 45220 45218
rect 45164 45164 45220 45166
rect 45164 44882 45220 44884
rect 45164 44830 45166 44882
rect 45166 44830 45218 44882
rect 45218 44830 45220 44882
rect 45164 44828 45220 44830
rect 45388 44716 45444 44772
rect 45052 41916 45108 41972
rect 46956 51996 47012 52052
rect 49308 51996 49364 52052
rect 47852 51490 47908 51492
rect 47852 51438 47854 51490
rect 47854 51438 47906 51490
rect 47906 51438 47908 51490
rect 47852 51436 47908 51438
rect 47068 49756 47124 49812
rect 46620 46732 46676 46788
rect 46844 46060 46900 46116
rect 48076 49980 48132 50036
rect 48748 51324 48804 51380
rect 49196 51266 49252 51268
rect 49196 51214 49198 51266
rect 49198 51214 49250 51266
rect 49250 51214 49252 51266
rect 49196 51212 49252 51214
rect 49420 51772 49476 51828
rect 49308 50540 49364 50596
rect 48860 50034 48916 50036
rect 48860 49982 48862 50034
rect 48862 49982 48914 50034
rect 48914 49982 48916 50034
rect 48860 49980 48916 49982
rect 49084 49922 49140 49924
rect 49084 49870 49086 49922
rect 49086 49870 49138 49922
rect 49138 49870 49140 49922
rect 49084 49868 49140 49870
rect 47404 48076 47460 48132
rect 47292 47180 47348 47236
rect 48188 48130 48244 48132
rect 48188 48078 48190 48130
rect 48190 48078 48242 48130
rect 48242 48078 48244 48130
rect 48188 48076 48244 48078
rect 47740 47068 47796 47124
rect 47068 46844 47124 46900
rect 46172 45836 46228 45892
rect 45836 45666 45892 45668
rect 45836 45614 45838 45666
rect 45838 45614 45890 45666
rect 45890 45614 45892 45666
rect 45836 45612 45892 45614
rect 46284 44940 46340 44996
rect 49196 48972 49252 49028
rect 48748 48242 48804 48244
rect 48748 48190 48750 48242
rect 48750 48190 48802 48242
rect 48802 48190 48804 48242
rect 48748 48188 48804 48190
rect 49868 53676 49924 53732
rect 49980 53564 50036 53620
rect 51548 54348 51604 54404
rect 50092 53116 50148 53172
rect 50876 53618 50932 53620
rect 50876 53566 50878 53618
rect 50878 53566 50930 53618
rect 50930 53566 50932 53618
rect 50876 53564 50932 53566
rect 50428 53452 50484 53508
rect 50652 53506 50708 53508
rect 50652 53454 50654 53506
rect 50654 53454 50706 53506
rect 50706 53454 50708 53506
rect 50652 53452 50708 53454
rect 50988 53452 51044 53508
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 49756 52892 49812 52948
rect 50540 52892 50596 52948
rect 49756 51996 49812 52052
rect 50316 52162 50372 52164
rect 50316 52110 50318 52162
rect 50318 52110 50370 52162
rect 50370 52110 50372 52162
rect 50316 52108 50372 52110
rect 50988 53116 51044 53172
rect 50876 52946 50932 52948
rect 50876 52894 50878 52946
rect 50878 52894 50930 52946
rect 50930 52894 50932 52946
rect 50876 52892 50932 52894
rect 50652 52108 50708 52164
rect 50764 51996 50820 52052
rect 49980 51772 50036 51828
rect 50092 50652 50148 50708
rect 50204 51772 50260 51828
rect 50204 51212 50260 51268
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 51324 52946 51380 52948
rect 51324 52894 51326 52946
rect 51326 52894 51378 52946
rect 51378 52894 51380 52946
rect 51324 52892 51380 52894
rect 52332 54402 52388 54404
rect 52332 54350 52334 54402
rect 52334 54350 52386 54402
rect 52386 54350 52388 54402
rect 52332 54348 52388 54350
rect 52444 52946 52500 52948
rect 52444 52894 52446 52946
rect 52446 52894 52498 52946
rect 52498 52894 52500 52946
rect 52444 52892 52500 52894
rect 51660 52780 51716 52836
rect 51324 52162 51380 52164
rect 51324 52110 51326 52162
rect 51326 52110 51378 52162
rect 51378 52110 51380 52162
rect 51324 52108 51380 52110
rect 50988 51548 51044 51604
rect 50876 50988 50932 51044
rect 53564 52108 53620 52164
rect 52444 51490 52500 51492
rect 52444 51438 52446 51490
rect 52446 51438 52498 51490
rect 52498 51438 52500 51490
rect 52444 51436 52500 51438
rect 50876 50540 50932 50596
rect 50316 50428 50372 50484
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 49756 49922 49812 49924
rect 49756 49870 49758 49922
rect 49758 49870 49810 49922
rect 49810 49870 49812 49922
rect 49756 49868 49812 49870
rect 50764 49084 50820 49140
rect 50204 48972 50260 49028
rect 50876 48914 50932 48916
rect 50876 48862 50878 48914
rect 50878 48862 50930 48914
rect 50930 48862 50932 48914
rect 50876 48860 50932 48862
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50428 48412 50484 48468
rect 49532 48188 49588 48244
rect 50204 48188 50260 48244
rect 49868 48130 49924 48132
rect 49868 48078 49870 48130
rect 49870 48078 49922 48130
rect 49922 48078 49924 48130
rect 49868 48076 49924 48078
rect 48748 46898 48804 46900
rect 48748 46846 48750 46898
rect 48750 46846 48802 46898
rect 48802 46846 48804 46898
rect 48748 46844 48804 46846
rect 48300 46114 48356 46116
rect 48300 46062 48302 46114
rect 48302 46062 48354 46114
rect 48354 46062 48356 46114
rect 48300 46060 48356 46062
rect 47292 45836 47348 45892
rect 47964 45778 48020 45780
rect 47964 45726 47966 45778
rect 47966 45726 48018 45778
rect 48018 45726 48020 45778
rect 47964 45724 48020 45726
rect 50428 47964 50484 48020
rect 49196 47180 49252 47236
rect 48972 46060 49028 46116
rect 49644 47180 49700 47236
rect 49756 47068 49812 47124
rect 49420 46786 49476 46788
rect 49420 46734 49422 46786
rect 49422 46734 49474 46786
rect 49474 46734 49476 46786
rect 49420 46732 49476 46734
rect 51212 50540 51268 50596
rect 51436 50988 51492 51044
rect 51996 51100 52052 51156
rect 52556 50988 52612 51044
rect 53116 51378 53172 51380
rect 53116 51326 53118 51378
rect 53118 51326 53170 51378
rect 53170 51326 53172 51378
rect 53116 51324 53172 51326
rect 52668 51100 52724 51156
rect 51996 50706 52052 50708
rect 51996 50654 51998 50706
rect 51998 50654 52050 50706
rect 52050 50654 52052 50706
rect 51996 50652 52052 50654
rect 51884 50540 51940 50596
rect 51996 50428 52052 50484
rect 51884 48860 51940 48916
rect 51324 48412 51380 48468
rect 54572 52108 54628 52164
rect 54684 51436 54740 51492
rect 53900 51378 53956 51380
rect 53900 51326 53902 51378
rect 53902 51326 53954 51378
rect 53954 51326 53956 51378
rect 53900 51324 53956 51326
rect 53564 50652 53620 50708
rect 52892 49868 52948 49924
rect 54124 50034 54180 50036
rect 54124 49982 54126 50034
rect 54126 49982 54178 50034
rect 54178 49982 54180 50034
rect 54124 49980 54180 49982
rect 53900 49922 53956 49924
rect 53900 49870 53902 49922
rect 53902 49870 53954 49922
rect 53954 49870 53956 49922
rect 53900 49868 53956 49870
rect 51772 48076 51828 48132
rect 51212 47740 51268 47796
rect 49644 45836 49700 45892
rect 47068 44940 47124 44996
rect 46508 44828 46564 44884
rect 46060 43538 46116 43540
rect 46060 43486 46062 43538
rect 46062 43486 46114 43538
rect 46114 43486 46116 43538
rect 46060 43484 46116 43486
rect 45276 41858 45332 41860
rect 45276 41806 45278 41858
rect 45278 41806 45330 41858
rect 45330 41806 45332 41858
rect 45276 41804 45332 41806
rect 45500 41804 45556 41860
rect 45724 42924 45780 42980
rect 47852 44882 47908 44884
rect 47852 44830 47854 44882
rect 47854 44830 47906 44882
rect 47906 44830 47908 44882
rect 47852 44828 47908 44830
rect 47628 43484 47684 43540
rect 46508 42700 46564 42756
rect 45612 41468 45668 41524
rect 45836 41580 45892 41636
rect 45836 41132 45892 41188
rect 45052 41020 45108 41076
rect 45276 41074 45332 41076
rect 45276 41022 45278 41074
rect 45278 41022 45330 41074
rect 45330 41022 45332 41074
rect 45276 41020 45332 41022
rect 44940 40348 44996 40404
rect 44604 40124 44660 40180
rect 45276 40402 45332 40404
rect 45276 40350 45278 40402
rect 45278 40350 45330 40402
rect 45330 40350 45332 40402
rect 45276 40348 45332 40350
rect 45612 40908 45668 40964
rect 44828 39564 44884 39620
rect 44268 38780 44324 38836
rect 44156 38722 44212 38724
rect 44156 38670 44158 38722
rect 44158 38670 44210 38722
rect 44210 38670 44212 38722
rect 44156 38668 44212 38670
rect 45948 40962 46004 40964
rect 45948 40910 45950 40962
rect 45950 40910 46002 40962
rect 46002 40910 46004 40962
rect 45948 40908 46004 40910
rect 46508 41858 46564 41860
rect 46508 41806 46510 41858
rect 46510 41806 46562 41858
rect 46562 41806 46564 41858
rect 46508 41804 46564 41806
rect 46396 40684 46452 40740
rect 46508 40460 46564 40516
rect 46732 41804 46788 41860
rect 45836 39618 45892 39620
rect 45836 39566 45838 39618
rect 45838 39566 45890 39618
rect 45890 39566 45892 39618
rect 45836 39564 45892 39566
rect 45500 38946 45556 38948
rect 45500 38894 45502 38946
rect 45502 38894 45554 38946
rect 45554 38894 45556 38946
rect 45500 38892 45556 38894
rect 45500 38668 45556 38724
rect 45836 37490 45892 37492
rect 45836 37438 45838 37490
rect 45838 37438 45890 37490
rect 45890 37438 45892 37490
rect 45836 37436 45892 37438
rect 46620 38610 46676 38612
rect 46620 38558 46622 38610
rect 46622 38558 46674 38610
rect 46674 38558 46676 38610
rect 46620 38556 46676 38558
rect 46620 38050 46676 38052
rect 46620 37998 46622 38050
rect 46622 37998 46674 38050
rect 46674 37998 46676 38050
rect 46620 37996 46676 37998
rect 46284 37378 46340 37380
rect 46284 37326 46286 37378
rect 46286 37326 46338 37378
rect 46338 37326 46340 37378
rect 46284 37324 46340 37326
rect 46060 37266 46116 37268
rect 46060 37214 46062 37266
rect 46062 37214 46114 37266
rect 46114 37214 46116 37266
rect 46060 37212 46116 37214
rect 43708 36204 43764 36260
rect 44940 36258 44996 36260
rect 44940 36206 44942 36258
rect 44942 36206 44994 36258
rect 44994 36206 44996 36258
rect 44940 36204 44996 36206
rect 45276 35756 45332 35812
rect 45500 35868 45556 35924
rect 43484 35644 43540 35700
rect 43260 35308 43316 35364
rect 45836 36204 45892 36260
rect 43484 35084 43540 35140
rect 44940 35084 44996 35140
rect 44044 34690 44100 34692
rect 44044 34638 44046 34690
rect 44046 34638 44098 34690
rect 44098 34638 44100 34690
rect 44044 34636 44100 34638
rect 46396 37212 46452 37268
rect 46508 37324 46564 37380
rect 46172 36258 46228 36260
rect 46172 36206 46174 36258
rect 46174 36206 46226 36258
rect 46226 36206 46228 36258
rect 46172 36204 46228 36206
rect 46060 36092 46116 36148
rect 45948 35586 46004 35588
rect 45948 35534 45950 35586
rect 45950 35534 46002 35586
rect 46002 35534 46004 35586
rect 45948 35532 46004 35534
rect 45836 34524 45892 34580
rect 45948 34690 46004 34692
rect 45948 34638 45950 34690
rect 45950 34638 46002 34690
rect 46002 34638 46004 34690
rect 45948 34636 46004 34638
rect 43708 34018 43764 34020
rect 43708 33966 43710 34018
rect 43710 33966 43762 34018
rect 43762 33966 43764 34018
rect 43708 33964 43764 33966
rect 42812 32508 42868 32564
rect 42140 32284 42196 32340
rect 41468 32172 41524 32228
rect 43596 31890 43652 31892
rect 43596 31838 43598 31890
rect 43598 31838 43650 31890
rect 43650 31838 43652 31890
rect 43596 31836 43652 31838
rect 41692 31164 41748 31220
rect 43148 31554 43204 31556
rect 43148 31502 43150 31554
rect 43150 31502 43202 31554
rect 43202 31502 43204 31554
rect 43148 31500 43204 31502
rect 43596 31388 43652 31444
rect 42700 31164 42756 31220
rect 43036 30882 43092 30884
rect 43036 30830 43038 30882
rect 43038 30830 43090 30882
rect 43090 30830 43092 30882
rect 43036 30828 43092 30830
rect 44268 33234 44324 33236
rect 44268 33182 44270 33234
rect 44270 33182 44322 33234
rect 44322 33182 44324 33234
rect 44268 33180 44324 33182
rect 45052 32562 45108 32564
rect 45052 32510 45054 32562
rect 45054 32510 45106 32562
rect 45106 32510 45108 32562
rect 45052 32508 45108 32510
rect 44604 32172 44660 32228
rect 44156 31554 44212 31556
rect 44156 31502 44158 31554
rect 44158 31502 44210 31554
rect 44210 31502 44212 31554
rect 44156 31500 44212 31502
rect 44604 31106 44660 31108
rect 44604 31054 44606 31106
rect 44606 31054 44658 31106
rect 44658 31054 44660 31106
rect 44604 31052 44660 31054
rect 44044 30828 44100 30884
rect 43708 30492 43764 30548
rect 45052 30828 45108 30884
rect 44380 30044 44436 30100
rect 41916 29596 41972 29652
rect 41468 29036 41524 29092
rect 42700 29426 42756 29428
rect 42700 29374 42702 29426
rect 42702 29374 42754 29426
rect 42754 29374 42756 29426
rect 42700 29372 42756 29374
rect 42476 29314 42532 29316
rect 42476 29262 42478 29314
rect 42478 29262 42530 29314
rect 42530 29262 42532 29314
rect 42476 29260 42532 29262
rect 42476 28924 42532 28980
rect 42588 29148 42644 29204
rect 41468 28028 41524 28084
rect 40348 25900 40404 25956
rect 40236 25394 40292 25396
rect 40236 25342 40238 25394
rect 40238 25342 40290 25394
rect 40290 25342 40292 25394
rect 40236 25340 40292 25342
rect 40348 24668 40404 24724
rect 39788 24498 39844 24500
rect 39788 24446 39790 24498
rect 39790 24446 39842 24498
rect 39842 24446 39844 24498
rect 39788 24444 39844 24446
rect 39564 24332 39620 24388
rect 40348 24050 40404 24052
rect 40348 23998 40350 24050
rect 40350 23998 40402 24050
rect 40402 23998 40404 24050
rect 40348 23996 40404 23998
rect 39564 23772 39620 23828
rect 41356 27858 41412 27860
rect 41356 27806 41358 27858
rect 41358 27806 41410 27858
rect 41410 27806 41412 27858
rect 41356 27804 41412 27806
rect 41804 28028 41860 28084
rect 43036 28924 43092 28980
rect 43708 29538 43764 29540
rect 43708 29486 43710 29538
rect 43710 29486 43762 29538
rect 43762 29486 43764 29538
rect 43708 29484 43764 29486
rect 44156 29484 44212 29540
rect 43372 29426 43428 29428
rect 43372 29374 43374 29426
rect 43374 29374 43426 29426
rect 43426 29374 43428 29426
rect 43372 29372 43428 29374
rect 43260 29260 43316 29316
rect 43820 29260 43876 29316
rect 42364 28082 42420 28084
rect 42364 28030 42366 28082
rect 42366 28030 42418 28082
rect 42418 28030 42420 28082
rect 42364 28028 42420 28030
rect 43260 28642 43316 28644
rect 43260 28590 43262 28642
rect 43262 28590 43314 28642
rect 43314 28590 43316 28642
rect 43260 28588 43316 28590
rect 43596 28588 43652 28644
rect 43708 28530 43764 28532
rect 43708 28478 43710 28530
rect 43710 28478 43762 28530
rect 43762 28478 43764 28530
rect 43708 28476 43764 28478
rect 44940 29202 44996 29204
rect 44940 29150 44942 29202
rect 44942 29150 44994 29202
rect 44994 29150 44996 29202
rect 44940 29148 44996 29150
rect 44268 28924 44324 28980
rect 43932 28812 43988 28868
rect 43484 28252 43540 28308
rect 43036 28028 43092 28084
rect 42588 27970 42644 27972
rect 42588 27918 42590 27970
rect 42590 27918 42642 27970
rect 42642 27918 42644 27970
rect 42588 27916 42644 27918
rect 41468 27074 41524 27076
rect 41468 27022 41470 27074
rect 41470 27022 41522 27074
rect 41522 27022 41524 27074
rect 41468 27020 41524 27022
rect 40572 25506 40628 25508
rect 40572 25454 40574 25506
rect 40574 25454 40626 25506
rect 40626 25454 40628 25506
rect 40572 25452 40628 25454
rect 41468 25900 41524 25956
rect 41132 25788 41188 25844
rect 40684 24556 40740 24612
rect 40572 24444 40628 24500
rect 41020 24834 41076 24836
rect 41020 24782 41022 24834
rect 41022 24782 41074 24834
rect 41074 24782 41076 24834
rect 41020 24780 41076 24782
rect 40908 24722 40964 24724
rect 40908 24670 40910 24722
rect 40910 24670 40962 24722
rect 40962 24670 40964 24722
rect 40908 24668 40964 24670
rect 40236 23154 40292 23156
rect 40236 23102 40238 23154
rect 40238 23102 40290 23154
rect 40290 23102 40292 23154
rect 40236 23100 40292 23102
rect 39452 22540 39508 22596
rect 39564 22204 39620 22260
rect 39788 22258 39844 22260
rect 39788 22206 39790 22258
rect 39790 22206 39842 22258
rect 39842 22206 39844 22258
rect 39788 22204 39844 22206
rect 40460 22764 40516 22820
rect 40236 22428 40292 22484
rect 40012 21810 40068 21812
rect 40012 21758 40014 21810
rect 40014 21758 40066 21810
rect 40066 21758 40068 21810
rect 40012 21756 40068 21758
rect 40684 22482 40740 22484
rect 40684 22430 40686 22482
rect 40686 22430 40738 22482
rect 40738 22430 40740 22482
rect 40684 22428 40740 22430
rect 40236 22258 40292 22260
rect 40236 22206 40238 22258
rect 40238 22206 40290 22258
rect 40290 22206 40292 22258
rect 40236 22204 40292 22206
rect 40684 21868 40740 21924
rect 39900 21644 39956 21700
rect 38892 21586 38948 21588
rect 38892 21534 38894 21586
rect 38894 21534 38946 21586
rect 38946 21534 38948 21586
rect 38892 21532 38948 21534
rect 39004 21420 39060 21476
rect 39004 20412 39060 20468
rect 39788 21586 39844 21588
rect 39788 21534 39790 21586
rect 39790 21534 39842 21586
rect 39842 21534 39844 21586
rect 39788 21532 39844 21534
rect 39340 20636 39396 20692
rect 39116 20524 39172 20580
rect 39340 20412 39396 20468
rect 38668 19740 38724 19796
rect 39116 19628 39172 19684
rect 38556 19346 38612 19348
rect 38556 19294 38558 19346
rect 38558 19294 38610 19346
rect 38610 19294 38612 19346
rect 38556 19292 38612 19294
rect 39452 20300 39508 20356
rect 38556 18956 38612 19012
rect 39676 19852 39732 19908
rect 40348 20860 40404 20916
rect 39900 20300 39956 20356
rect 39564 19740 39620 19796
rect 40460 20748 40516 20804
rect 39788 19740 39844 19796
rect 39564 18844 39620 18900
rect 38556 18450 38612 18452
rect 38556 18398 38558 18450
rect 38558 18398 38610 18450
rect 38610 18398 38612 18450
rect 38556 18396 38612 18398
rect 39228 18450 39284 18452
rect 39228 18398 39230 18450
rect 39230 18398 39282 18450
rect 39282 18398 39284 18450
rect 39228 18396 39284 18398
rect 37884 17666 37940 17668
rect 37884 17614 37886 17666
rect 37886 17614 37938 17666
rect 37938 17614 37940 17666
rect 37884 17612 37940 17614
rect 40572 20524 40628 20580
rect 40236 19740 40292 19796
rect 40124 18620 40180 18676
rect 39676 18450 39732 18452
rect 39676 18398 39678 18450
rect 39678 18398 39730 18450
rect 39730 18398 39732 18450
rect 39676 18396 39732 18398
rect 40348 18450 40404 18452
rect 40348 18398 40350 18450
rect 40350 18398 40402 18450
rect 40402 18398 40404 18450
rect 40348 18396 40404 18398
rect 39788 17948 39844 18004
rect 39676 17666 39732 17668
rect 39676 17614 39678 17666
rect 39678 17614 39730 17666
rect 39730 17614 39732 17666
rect 39676 17612 39732 17614
rect 37772 17106 37828 17108
rect 37772 17054 37774 17106
rect 37774 17054 37826 17106
rect 37826 17054 37828 17106
rect 37772 17052 37828 17054
rect 37996 16716 38052 16772
rect 38220 16380 38276 16436
rect 38108 16044 38164 16100
rect 37884 15986 37940 15988
rect 37884 15934 37886 15986
rect 37886 15934 37938 15986
rect 37938 15934 37940 15986
rect 37884 15932 37940 15934
rect 39004 16940 39060 16996
rect 39116 16828 39172 16884
rect 39228 16716 39284 16772
rect 38108 15596 38164 15652
rect 38220 15260 38276 15316
rect 37996 14924 38052 14980
rect 37548 14252 37604 14308
rect 37884 14028 37940 14084
rect 37772 13970 37828 13972
rect 37772 13918 37774 13970
rect 37774 13918 37826 13970
rect 37826 13918 37828 13970
rect 37772 13916 37828 13918
rect 37548 12124 37604 12180
rect 37100 11394 37156 11396
rect 37100 11342 37102 11394
rect 37102 11342 37154 11394
rect 37154 11342 37156 11394
rect 37100 11340 37156 11342
rect 36988 10780 37044 10836
rect 37100 10444 37156 10500
rect 37324 10556 37380 10612
rect 37772 12684 37828 12740
rect 37772 12290 37828 12292
rect 37772 12238 37774 12290
rect 37774 12238 37826 12290
rect 37826 12238 37828 12290
rect 37772 12236 37828 12238
rect 37772 11228 37828 11284
rect 37884 10444 37940 10500
rect 37884 10108 37940 10164
rect 36428 7698 36484 7700
rect 36428 7646 36430 7698
rect 36430 7646 36482 7698
rect 36482 7646 36484 7698
rect 36428 7644 36484 7646
rect 36876 7644 36932 7700
rect 36652 4956 36708 5012
rect 36092 3612 36148 3668
rect 36204 3388 36260 3444
rect 36316 3500 36372 3556
rect 37100 3500 37156 3556
rect 37548 7980 37604 8036
rect 38444 15260 38500 15316
rect 38892 15596 38948 15652
rect 39452 16994 39508 16996
rect 39452 16942 39454 16994
rect 39454 16942 39506 16994
rect 39506 16942 39508 16994
rect 39452 16940 39508 16942
rect 39676 16828 39732 16884
rect 39228 15538 39284 15540
rect 39228 15486 39230 15538
rect 39230 15486 39282 15538
rect 39282 15486 39284 15538
rect 39228 15484 39284 15486
rect 38780 15148 38836 15204
rect 39564 14476 39620 14532
rect 39340 13916 39396 13972
rect 39452 14364 39508 14420
rect 38780 13692 38836 13748
rect 38108 12012 38164 12068
rect 38556 12738 38612 12740
rect 38556 12686 38558 12738
rect 38558 12686 38610 12738
rect 38610 12686 38612 12738
rect 38556 12684 38612 12686
rect 38556 12460 38612 12516
rect 38444 12178 38500 12180
rect 38444 12126 38446 12178
rect 38446 12126 38498 12178
rect 38498 12126 38500 12178
rect 38444 12124 38500 12126
rect 38780 12402 38836 12404
rect 38780 12350 38782 12402
rect 38782 12350 38834 12402
rect 38834 12350 38836 12402
rect 38780 12348 38836 12350
rect 38668 12290 38724 12292
rect 38668 12238 38670 12290
rect 38670 12238 38722 12290
rect 38722 12238 38724 12290
rect 38668 12236 38724 12238
rect 38332 11676 38388 11732
rect 38220 11618 38276 11620
rect 38220 11566 38222 11618
rect 38222 11566 38274 11618
rect 38274 11566 38276 11618
rect 38220 11564 38276 11566
rect 38332 11340 38388 11396
rect 38556 11340 38612 11396
rect 38220 10892 38276 10948
rect 38444 11116 38500 11172
rect 38108 10556 38164 10612
rect 38220 10668 38276 10724
rect 38780 11452 38836 11508
rect 39116 12066 39172 12068
rect 39116 12014 39118 12066
rect 39118 12014 39170 12066
rect 39170 12014 39172 12066
rect 39116 12012 39172 12014
rect 39004 11452 39060 11508
rect 39452 13692 39508 13748
rect 39564 13580 39620 13636
rect 39452 12236 39508 12292
rect 38780 10780 38836 10836
rect 38444 10386 38500 10388
rect 38444 10334 38446 10386
rect 38446 10334 38498 10386
rect 38498 10334 38500 10386
rect 38444 10332 38500 10334
rect 38220 9042 38276 9044
rect 38220 8990 38222 9042
rect 38222 8990 38274 9042
rect 38274 8990 38276 9042
rect 38220 8988 38276 8990
rect 38332 8876 38388 8932
rect 38220 8034 38276 8036
rect 38220 7982 38222 8034
rect 38222 7982 38274 8034
rect 38274 7982 38276 8034
rect 38220 7980 38276 7982
rect 37548 3554 37604 3556
rect 37548 3502 37550 3554
rect 37550 3502 37602 3554
rect 37602 3502 37604 3554
rect 37548 3500 37604 3502
rect 37884 3500 37940 3556
rect 38668 10108 38724 10164
rect 40348 17948 40404 18004
rect 40012 15148 40068 15204
rect 39900 11788 39956 11844
rect 39788 11394 39844 11396
rect 39788 11342 39790 11394
rect 39790 11342 39842 11394
rect 39842 11342 39844 11394
rect 39788 11340 39844 11342
rect 39676 11282 39732 11284
rect 39676 11230 39678 11282
rect 39678 11230 39730 11282
rect 39730 11230 39732 11282
rect 39676 11228 39732 11230
rect 39900 11170 39956 11172
rect 39900 11118 39902 11170
rect 39902 11118 39954 11170
rect 39954 11118 39956 11170
rect 39900 11116 39956 11118
rect 39004 10556 39060 10612
rect 39788 10444 39844 10500
rect 39228 10220 39284 10276
rect 39452 9772 39508 9828
rect 40012 10108 40068 10164
rect 40124 9660 40180 9716
rect 39788 9154 39844 9156
rect 39788 9102 39790 9154
rect 39790 9102 39842 9154
rect 39842 9102 39844 9154
rect 39788 9100 39844 9102
rect 38892 8988 38948 9044
rect 39564 8428 39620 8484
rect 39676 8988 39732 9044
rect 39900 8930 39956 8932
rect 39900 8878 39902 8930
rect 39902 8878 39954 8930
rect 39954 8878 39956 8930
rect 39900 8876 39956 8878
rect 40124 7698 40180 7700
rect 40124 7646 40126 7698
rect 40126 7646 40178 7698
rect 40178 7646 40180 7698
rect 40124 7644 40180 7646
rect 38668 3948 38724 4004
rect 39004 3554 39060 3556
rect 39004 3502 39006 3554
rect 39006 3502 39058 3554
rect 39058 3502 39060 3554
rect 39004 3500 39060 3502
rect 39900 3388 39956 3444
rect 40348 12684 40404 12740
rect 41468 23938 41524 23940
rect 41468 23886 41470 23938
rect 41470 23886 41522 23938
rect 41522 23886 41524 23938
rect 41468 23884 41524 23886
rect 40908 23100 40964 23156
rect 42140 27858 42196 27860
rect 42140 27806 42142 27858
rect 42142 27806 42194 27858
rect 42194 27806 42196 27858
rect 42140 27804 42196 27806
rect 42588 27468 42644 27524
rect 42028 26684 42084 26740
rect 42700 26684 42756 26740
rect 42812 27804 42868 27860
rect 42028 26460 42084 26516
rect 41916 24444 41972 24500
rect 41804 23772 41860 23828
rect 41468 22764 41524 22820
rect 41692 22594 41748 22596
rect 41692 22542 41694 22594
rect 41694 22542 41746 22594
rect 41746 22542 41748 22594
rect 41692 22540 41748 22542
rect 41244 22482 41300 22484
rect 41244 22430 41246 22482
rect 41246 22430 41298 22482
rect 41298 22430 41300 22482
rect 41244 22428 41300 22430
rect 41916 22428 41972 22484
rect 41020 21810 41076 21812
rect 41020 21758 41022 21810
rect 41022 21758 41074 21810
rect 41074 21758 41076 21810
rect 41020 21756 41076 21758
rect 41468 21698 41524 21700
rect 41468 21646 41470 21698
rect 41470 21646 41522 21698
rect 41522 21646 41524 21698
rect 41468 21644 41524 21646
rect 40908 20690 40964 20692
rect 40908 20638 40910 20690
rect 40910 20638 40962 20690
rect 40962 20638 40964 20690
rect 40908 20636 40964 20638
rect 41356 20972 41412 21028
rect 41020 20578 41076 20580
rect 41020 20526 41022 20578
rect 41022 20526 41074 20578
rect 41074 20526 41076 20578
rect 41020 20524 41076 20526
rect 41020 20300 41076 20356
rect 41468 20300 41524 20356
rect 41020 19404 41076 19460
rect 41356 18508 41412 18564
rect 41244 17724 41300 17780
rect 41244 17500 41300 17556
rect 40684 13074 40740 13076
rect 40684 13022 40686 13074
rect 40686 13022 40738 13074
rect 40738 13022 40740 13074
rect 40684 13020 40740 13022
rect 40572 11900 40628 11956
rect 41132 13858 41188 13860
rect 41132 13806 41134 13858
rect 41134 13806 41186 13858
rect 41186 13806 41188 13858
rect 41132 13804 41188 13806
rect 41132 13580 41188 13636
rect 40908 12124 40964 12180
rect 41020 13468 41076 13524
rect 41132 12850 41188 12852
rect 41132 12798 41134 12850
rect 41134 12798 41186 12850
rect 41186 12798 41188 12850
rect 41132 12796 41188 12798
rect 41468 18060 41524 18116
rect 43820 27858 43876 27860
rect 43820 27806 43822 27858
rect 43822 27806 43874 27858
rect 43874 27806 43876 27858
rect 43820 27804 43876 27806
rect 44380 28700 44436 28756
rect 44156 28588 44212 28644
rect 44604 28476 44660 28532
rect 44044 27692 44100 27748
rect 43036 26908 43092 26964
rect 43260 26908 43316 26964
rect 42588 26402 42644 26404
rect 42588 26350 42590 26402
rect 42590 26350 42642 26402
rect 42642 26350 42644 26402
rect 42588 26348 42644 26350
rect 42476 26290 42532 26292
rect 42476 26238 42478 26290
rect 42478 26238 42530 26290
rect 42530 26238 42532 26290
rect 42476 26236 42532 26238
rect 43148 26402 43204 26404
rect 43148 26350 43150 26402
rect 43150 26350 43202 26402
rect 43202 26350 43204 26402
rect 43148 26348 43204 26350
rect 42252 25564 42308 25620
rect 43372 26514 43428 26516
rect 43372 26462 43374 26514
rect 43374 26462 43426 26514
rect 43426 26462 43428 26514
rect 43372 26460 43428 26462
rect 43820 26684 43876 26740
rect 44044 26962 44100 26964
rect 44044 26910 44046 26962
rect 44046 26910 44098 26962
rect 44098 26910 44100 26962
rect 44044 26908 44100 26910
rect 44156 27020 44212 27076
rect 43932 26460 43988 26516
rect 44044 26348 44100 26404
rect 42924 24722 42980 24724
rect 42924 24670 42926 24722
rect 42926 24670 42978 24722
rect 42978 24670 42980 24722
rect 42924 24668 42980 24670
rect 42140 23996 42196 24052
rect 42364 23378 42420 23380
rect 42364 23326 42366 23378
rect 42366 23326 42418 23378
rect 42418 23326 42420 23378
rect 42364 23324 42420 23326
rect 43148 24444 43204 24500
rect 44716 27746 44772 27748
rect 44716 27694 44718 27746
rect 44718 27694 44770 27746
rect 44770 27694 44772 27746
rect 44716 27692 44772 27694
rect 44828 27132 44884 27188
rect 45836 33516 45892 33572
rect 45612 33234 45668 33236
rect 45612 33182 45614 33234
rect 45614 33182 45666 33234
rect 45666 33182 45668 33234
rect 45612 33180 45668 33182
rect 45388 31836 45444 31892
rect 45836 31948 45892 32004
rect 45724 31106 45780 31108
rect 45724 31054 45726 31106
rect 45726 31054 45778 31106
rect 45778 31054 45780 31106
rect 45724 31052 45780 31054
rect 45948 31612 46004 31668
rect 46060 31052 46116 31108
rect 46060 30380 46116 30436
rect 45948 29484 46004 29540
rect 46172 28812 46228 28868
rect 45276 28418 45332 28420
rect 45276 28366 45278 28418
rect 45278 28366 45330 28418
rect 45330 28366 45332 28418
rect 45276 28364 45332 28366
rect 45388 27916 45444 27972
rect 45388 27468 45444 27524
rect 46172 28140 46228 28196
rect 46620 37212 46676 37268
rect 47404 42754 47460 42756
rect 47404 42702 47406 42754
rect 47406 42702 47458 42754
rect 47458 42702 47460 42754
rect 47404 42700 47460 42702
rect 47516 41970 47572 41972
rect 47516 41918 47518 41970
rect 47518 41918 47570 41970
rect 47570 41918 47572 41970
rect 47516 41916 47572 41918
rect 47628 41580 47684 41636
rect 47068 41356 47124 41412
rect 47628 41186 47684 41188
rect 47628 41134 47630 41186
rect 47630 41134 47682 41186
rect 47682 41134 47684 41186
rect 47628 41132 47684 41134
rect 47516 41074 47572 41076
rect 47516 41022 47518 41074
rect 47518 41022 47570 41074
rect 47570 41022 47572 41074
rect 47516 41020 47572 41022
rect 47068 40236 47124 40292
rect 47180 38668 47236 38724
rect 46844 38220 46900 38276
rect 46956 38556 47012 38612
rect 47292 38220 47348 38276
rect 47068 38050 47124 38052
rect 47068 37998 47070 38050
rect 47070 37998 47122 38050
rect 47122 37998 47124 38050
rect 47068 37996 47124 37998
rect 47068 37266 47124 37268
rect 47068 37214 47070 37266
rect 47070 37214 47122 37266
rect 47122 37214 47124 37266
rect 47068 37212 47124 37214
rect 46732 36652 46788 36708
rect 47516 36482 47572 36484
rect 47516 36430 47518 36482
rect 47518 36430 47570 36482
rect 47570 36430 47572 36482
rect 47516 36428 47572 36430
rect 47852 43596 47908 43652
rect 48860 43650 48916 43652
rect 48860 43598 48862 43650
rect 48862 43598 48914 43650
rect 48914 43598 48916 43650
rect 48860 43596 48916 43598
rect 47852 42140 47908 42196
rect 48860 42530 48916 42532
rect 48860 42478 48862 42530
rect 48862 42478 48914 42530
rect 48914 42478 48916 42530
rect 48860 42476 48916 42478
rect 49308 42530 49364 42532
rect 49308 42478 49310 42530
rect 49310 42478 49362 42530
rect 49362 42478 49364 42530
rect 49308 42476 49364 42478
rect 47964 41916 48020 41972
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50540 46562 50596 46564
rect 50540 46510 50542 46562
rect 50542 46510 50594 46562
rect 50594 46510 50596 46562
rect 50540 46508 50596 46510
rect 50428 46002 50484 46004
rect 50428 45950 50430 46002
rect 50430 45950 50482 46002
rect 50482 45950 50484 46002
rect 50428 45948 50484 45950
rect 51772 47516 51828 47572
rect 52332 47516 52388 47572
rect 51996 46732 52052 46788
rect 50988 45948 51044 46004
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50764 45276 50820 45332
rect 51996 45666 52052 45668
rect 51996 45614 51998 45666
rect 51998 45614 52050 45666
rect 52050 45614 52052 45666
rect 51996 45612 52052 45614
rect 51660 45388 51716 45444
rect 51212 44994 51268 44996
rect 51212 44942 51214 44994
rect 51214 44942 51266 44994
rect 51266 44942 51268 44994
rect 51212 44940 51268 44942
rect 51100 44492 51156 44548
rect 51212 44210 51268 44212
rect 51212 44158 51214 44210
rect 51214 44158 51266 44210
rect 51266 44158 51268 44210
rect 51212 44156 51268 44158
rect 50764 44044 50820 44100
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50988 43932 51044 43988
rect 49980 43650 50036 43652
rect 49980 43598 49982 43650
rect 49982 43598 50034 43650
rect 50034 43598 50036 43650
rect 49980 43596 50036 43598
rect 52220 45388 52276 45444
rect 52108 44940 52164 44996
rect 51884 44434 51940 44436
rect 51884 44382 51886 44434
rect 51886 44382 51938 44434
rect 51938 44382 51940 44434
rect 51884 44380 51940 44382
rect 51660 43932 51716 43988
rect 49868 43314 49924 43316
rect 49868 43262 49870 43314
rect 49870 43262 49922 43314
rect 49922 43262 49924 43314
rect 49868 43260 49924 43262
rect 51772 43538 51828 43540
rect 51772 43486 51774 43538
rect 51774 43486 51826 43538
rect 51826 43486 51828 43538
rect 51772 43484 51828 43486
rect 49756 42924 49812 42980
rect 50652 42924 50708 42980
rect 50988 42812 51044 42868
rect 50764 42754 50820 42756
rect 50764 42702 50766 42754
rect 50766 42702 50818 42754
rect 50818 42702 50820 42754
rect 50764 42700 50820 42702
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50988 42252 51044 42308
rect 50876 41858 50932 41860
rect 50876 41806 50878 41858
rect 50878 41806 50930 41858
rect 50930 41806 50932 41858
rect 50876 41804 50932 41806
rect 49644 41692 49700 41748
rect 49308 41580 49364 41636
rect 48412 40348 48468 40404
rect 48748 41132 48804 41188
rect 48076 40124 48132 40180
rect 49084 41074 49140 41076
rect 49084 41022 49086 41074
rect 49086 41022 49138 41074
rect 49138 41022 49140 41074
rect 49084 41020 49140 41022
rect 48748 39900 48804 39956
rect 48860 40402 48916 40404
rect 48860 40350 48862 40402
rect 48862 40350 48914 40402
rect 48914 40350 48916 40402
rect 48860 40348 48916 40350
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 49308 40402 49364 40404
rect 49308 40350 49310 40402
rect 49310 40350 49362 40402
rect 49362 40350 49364 40402
rect 49308 40348 49364 40350
rect 50316 39394 50372 39396
rect 50316 39342 50318 39394
rect 50318 39342 50370 39394
rect 50370 39342 50372 39394
rect 50316 39340 50372 39342
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 51436 43036 51492 43092
rect 51436 42194 51492 42196
rect 51436 42142 51438 42194
rect 51438 42142 51490 42194
rect 51490 42142 51492 42194
rect 51436 42140 51492 42142
rect 51324 41916 51380 41972
rect 51212 40348 51268 40404
rect 51212 39730 51268 39732
rect 51212 39678 51214 39730
rect 51214 39678 51266 39730
rect 51266 39678 51268 39730
rect 51212 39676 51268 39678
rect 52668 48860 52724 48916
rect 54124 48860 54180 48916
rect 53340 48748 53396 48804
rect 53116 48130 53172 48132
rect 53116 48078 53118 48130
rect 53118 48078 53170 48130
rect 53170 48078 53172 48130
rect 53116 48076 53172 48078
rect 52668 46786 52724 46788
rect 52668 46734 52670 46786
rect 52670 46734 52722 46786
rect 52722 46734 52724 46786
rect 52668 46732 52724 46734
rect 52668 45890 52724 45892
rect 52668 45838 52670 45890
rect 52670 45838 52722 45890
rect 52722 45838 52724 45890
rect 52668 45836 52724 45838
rect 52556 44492 52612 44548
rect 51884 42140 51940 42196
rect 51884 41970 51940 41972
rect 51884 41918 51886 41970
rect 51886 41918 51938 41970
rect 51938 41918 51940 41970
rect 51884 41916 51940 41918
rect 51660 40962 51716 40964
rect 51660 40910 51662 40962
rect 51662 40910 51714 40962
rect 51714 40910 51716 40962
rect 51660 40908 51716 40910
rect 51660 40348 51716 40404
rect 51772 39394 51828 39396
rect 51772 39342 51774 39394
rect 51774 39342 51826 39394
rect 51826 39342 51828 39394
rect 51772 39340 51828 39342
rect 50876 38892 50932 38948
rect 47852 37884 47908 37940
rect 49532 38722 49588 38724
rect 49532 38670 49534 38722
rect 49534 38670 49586 38722
rect 49586 38670 49588 38722
rect 49532 38668 49588 38670
rect 53004 45612 53060 45668
rect 55580 51436 55636 51492
rect 54796 50034 54852 50036
rect 54796 49982 54798 50034
rect 54798 49982 54850 50034
rect 54850 49982 54852 50034
rect 54796 49980 54852 49982
rect 55468 48748 55524 48804
rect 55244 46172 55300 46228
rect 54684 45330 54740 45332
rect 54684 45278 54686 45330
rect 54686 45278 54738 45330
rect 54738 45278 54740 45330
rect 54684 45276 54740 45278
rect 53116 43650 53172 43652
rect 53116 43598 53118 43650
rect 53118 43598 53170 43650
rect 53170 43598 53172 43650
rect 53116 43596 53172 43598
rect 52668 42028 52724 42084
rect 53004 43148 53060 43204
rect 54460 43596 54516 43652
rect 53116 42700 53172 42756
rect 52668 41186 52724 41188
rect 52668 41134 52670 41186
rect 52670 41134 52722 41186
rect 52722 41134 52724 41186
rect 52668 41132 52724 41134
rect 52108 40962 52164 40964
rect 52108 40910 52110 40962
rect 52110 40910 52162 40962
rect 52162 40910 52164 40962
rect 52108 40908 52164 40910
rect 53452 41356 53508 41412
rect 53116 40572 53172 40628
rect 53228 41132 53284 41188
rect 52220 40290 52276 40292
rect 52220 40238 52222 40290
rect 52222 40238 52274 40290
rect 52274 40238 52276 40290
rect 52220 40236 52276 40238
rect 52780 39730 52836 39732
rect 52780 39678 52782 39730
rect 52782 39678 52834 39730
rect 52834 39678 52836 39730
rect 52780 39676 52836 39678
rect 52444 38946 52500 38948
rect 52444 38894 52446 38946
rect 52446 38894 52498 38946
rect 52498 38894 52500 38946
rect 52444 38892 52500 38894
rect 48412 37436 48468 37492
rect 48076 37266 48132 37268
rect 48076 37214 48078 37266
rect 48078 37214 48130 37266
rect 48130 37214 48132 37266
rect 48076 37212 48132 37214
rect 48860 37266 48916 37268
rect 48860 37214 48862 37266
rect 48862 37214 48914 37266
rect 48914 37214 48916 37266
rect 48860 37212 48916 37214
rect 50876 38108 50932 38164
rect 49532 37938 49588 37940
rect 49532 37886 49534 37938
rect 49534 37886 49586 37938
rect 49586 37886 49588 37938
rect 49532 37884 49588 37886
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50428 37490 50484 37492
rect 50428 37438 50430 37490
rect 50430 37438 50482 37490
rect 50482 37438 50484 37490
rect 50428 37436 50484 37438
rect 51212 37378 51268 37380
rect 51212 37326 51214 37378
rect 51214 37326 51266 37378
rect 51266 37326 51268 37378
rect 51212 37324 51268 37326
rect 51548 37266 51604 37268
rect 51548 37214 51550 37266
rect 51550 37214 51602 37266
rect 51602 37214 51604 37266
rect 51548 37212 51604 37214
rect 51324 36988 51380 37044
rect 46956 36092 47012 36148
rect 47180 36258 47236 36260
rect 47180 36206 47182 36258
rect 47182 36206 47234 36258
rect 47234 36206 47236 36258
rect 47180 36204 47236 36206
rect 47180 35756 47236 35812
rect 48076 36258 48132 36260
rect 48076 36206 48078 36258
rect 48078 36206 48130 36258
rect 48130 36206 48132 36258
rect 48076 36204 48132 36206
rect 47852 35810 47908 35812
rect 47852 35758 47854 35810
rect 47854 35758 47906 35810
rect 47906 35758 47908 35810
rect 47852 35756 47908 35758
rect 48076 35756 48132 35812
rect 46508 35420 46564 35476
rect 46620 35084 46676 35140
rect 46620 33628 46676 33684
rect 46396 27804 46452 27860
rect 46508 31612 46564 31668
rect 45836 27132 45892 27188
rect 46396 27580 46452 27636
rect 46060 26684 46116 26740
rect 44604 26402 44660 26404
rect 44604 26350 44606 26402
rect 44606 26350 44658 26402
rect 44658 26350 44660 26402
rect 44604 26348 44660 26350
rect 42812 23436 42868 23492
rect 42924 22988 42980 23044
rect 42476 22876 42532 22932
rect 42028 22316 42084 22372
rect 41804 22204 41860 22260
rect 42364 22092 42420 22148
rect 41916 21420 41972 21476
rect 41804 20802 41860 20804
rect 41804 20750 41806 20802
rect 41806 20750 41858 20802
rect 41858 20750 41860 20802
rect 41804 20748 41860 20750
rect 42588 21980 42644 22036
rect 43148 23436 43204 23492
rect 43484 23714 43540 23716
rect 43484 23662 43486 23714
rect 43486 23662 43538 23714
rect 43538 23662 43540 23714
rect 43484 23660 43540 23662
rect 43484 23378 43540 23380
rect 43484 23326 43486 23378
rect 43486 23326 43538 23378
rect 43538 23326 43540 23378
rect 43484 23324 43540 23326
rect 43372 23100 43428 23156
rect 44492 24722 44548 24724
rect 44492 24670 44494 24722
rect 44494 24670 44546 24722
rect 44546 24670 44548 24722
rect 44492 24668 44548 24670
rect 44604 24556 44660 24612
rect 44380 24108 44436 24164
rect 45948 25116 46004 25172
rect 43820 23548 43876 23604
rect 43708 23212 43764 23268
rect 43932 23042 43988 23044
rect 43932 22990 43934 23042
rect 43934 22990 43986 23042
rect 43986 22990 43988 23042
rect 43932 22988 43988 22990
rect 45052 23436 45108 23492
rect 44380 23042 44436 23044
rect 44380 22990 44382 23042
rect 44382 22990 44434 23042
rect 44434 22990 44436 23042
rect 44380 22988 44436 22990
rect 42924 21868 42980 21924
rect 43036 22370 43092 22372
rect 43036 22318 43038 22370
rect 43038 22318 43090 22370
rect 43090 22318 43092 22370
rect 43036 22316 43092 22318
rect 42700 21474 42756 21476
rect 42700 21422 42702 21474
rect 42702 21422 42754 21474
rect 42754 21422 42756 21474
rect 42700 21420 42756 21422
rect 42140 20300 42196 20356
rect 42140 19794 42196 19796
rect 42140 19742 42142 19794
rect 42142 19742 42194 19794
rect 42194 19742 42196 19794
rect 42140 19740 42196 19742
rect 42140 19404 42196 19460
rect 41692 17724 41748 17780
rect 43148 22258 43204 22260
rect 43148 22206 43150 22258
rect 43150 22206 43202 22258
rect 43202 22206 43204 22258
rect 43148 22204 43204 22206
rect 42476 19740 42532 19796
rect 42700 19122 42756 19124
rect 42700 19070 42702 19122
rect 42702 19070 42754 19122
rect 42754 19070 42756 19122
rect 42700 19068 42756 19070
rect 42924 19404 42980 19460
rect 42364 18226 42420 18228
rect 42364 18174 42366 18226
rect 42366 18174 42418 18226
rect 42418 18174 42420 18226
rect 42364 18172 42420 18174
rect 42476 17948 42532 18004
rect 42364 17106 42420 17108
rect 42364 17054 42366 17106
rect 42366 17054 42418 17106
rect 42418 17054 42420 17106
rect 42364 17052 42420 17054
rect 41580 16940 41636 16996
rect 42028 16882 42084 16884
rect 42028 16830 42030 16882
rect 42030 16830 42082 16882
rect 42082 16830 42084 16882
rect 42028 16828 42084 16830
rect 42140 16716 42196 16772
rect 42252 16492 42308 16548
rect 41916 16380 41972 16436
rect 41356 14530 41412 14532
rect 41356 14478 41358 14530
rect 41358 14478 41410 14530
rect 41410 14478 41412 14530
rect 41356 14476 41412 14478
rect 41468 14418 41524 14420
rect 41468 14366 41470 14418
rect 41470 14366 41522 14418
rect 41522 14366 41524 14418
rect 41468 14364 41524 14366
rect 41468 13020 41524 13076
rect 41244 12236 41300 12292
rect 40460 11788 40516 11844
rect 40348 11394 40404 11396
rect 40348 11342 40350 11394
rect 40350 11342 40402 11394
rect 40402 11342 40404 11394
rect 40348 11340 40404 11342
rect 40348 3388 40404 3444
rect 41020 11116 41076 11172
rect 40796 10444 40852 10500
rect 40908 9772 40964 9828
rect 41468 12178 41524 12180
rect 41468 12126 41470 12178
rect 41470 12126 41522 12178
rect 41522 12126 41524 12178
rect 41468 12124 41524 12126
rect 42028 14642 42084 14644
rect 42028 14590 42030 14642
rect 42030 14590 42082 14642
rect 42082 14590 42084 14642
rect 42028 14588 42084 14590
rect 42588 17052 42644 17108
rect 42588 16658 42644 16660
rect 42588 16606 42590 16658
rect 42590 16606 42642 16658
rect 42642 16606 42644 16658
rect 42588 16604 42644 16606
rect 42812 17948 42868 18004
rect 43148 19346 43204 19348
rect 43148 19294 43150 19346
rect 43150 19294 43202 19346
rect 43202 19294 43204 19346
rect 43148 19292 43204 19294
rect 43036 19180 43092 19236
rect 44940 22930 44996 22932
rect 44940 22878 44942 22930
rect 44942 22878 44994 22930
rect 44994 22878 44996 22930
rect 44940 22876 44996 22878
rect 43596 22258 43652 22260
rect 43596 22206 43598 22258
rect 43598 22206 43650 22258
rect 43650 22206 43652 22258
rect 43596 22204 43652 22206
rect 44044 22146 44100 22148
rect 44044 22094 44046 22146
rect 44046 22094 44098 22146
rect 44098 22094 44100 22146
rect 44044 22092 44100 22094
rect 45052 21980 45108 22036
rect 44268 20802 44324 20804
rect 44268 20750 44270 20802
rect 44270 20750 44322 20802
rect 44322 20750 44324 20802
rect 44268 20748 44324 20750
rect 45276 24162 45332 24164
rect 45276 24110 45278 24162
rect 45278 24110 45330 24162
rect 45330 24110 45332 24162
rect 45276 24108 45332 24110
rect 45276 23154 45332 23156
rect 45276 23102 45278 23154
rect 45278 23102 45330 23154
rect 45330 23102 45332 23154
rect 45276 23100 45332 23102
rect 45500 22876 45556 22932
rect 44828 20300 44884 20356
rect 44940 20188 44996 20244
rect 43484 19234 43540 19236
rect 43484 19182 43486 19234
rect 43486 19182 43538 19234
rect 43538 19182 43540 19234
rect 43484 19180 43540 19182
rect 43372 19068 43428 19124
rect 43260 18396 43316 18452
rect 43708 19852 43764 19908
rect 44044 19404 44100 19460
rect 43484 18338 43540 18340
rect 43484 18286 43486 18338
rect 43486 18286 43538 18338
rect 43538 18286 43540 18338
rect 43484 18284 43540 18286
rect 42812 16716 42868 16772
rect 44604 18620 44660 18676
rect 44156 18562 44212 18564
rect 44156 18510 44158 18562
rect 44158 18510 44210 18562
rect 44210 18510 44212 18562
rect 44156 18508 44212 18510
rect 44044 17778 44100 17780
rect 44044 17726 44046 17778
rect 44046 17726 44098 17778
rect 44098 17726 44100 17778
rect 44044 17724 44100 17726
rect 44268 17612 44324 17668
rect 43820 17388 43876 17444
rect 43036 16716 43092 16772
rect 42924 16492 42980 16548
rect 42700 16380 42756 16436
rect 43260 16940 43316 16996
rect 44044 16994 44100 16996
rect 44044 16942 44046 16994
rect 44046 16942 44098 16994
rect 44098 16942 44100 16994
rect 44044 16940 44100 16942
rect 44716 18562 44772 18564
rect 44716 18510 44718 18562
rect 44718 18510 44770 18562
rect 44770 18510 44772 18562
rect 44716 18508 44772 18510
rect 45164 19740 45220 19796
rect 44940 17724 44996 17780
rect 45052 18396 45108 18452
rect 46396 26684 46452 26740
rect 46284 22370 46340 22372
rect 46284 22318 46286 22370
rect 46286 22318 46338 22370
rect 46338 22318 46340 22370
rect 46284 22316 46340 22318
rect 45836 21026 45892 21028
rect 45836 20974 45838 21026
rect 45838 20974 45890 21026
rect 45890 20974 45892 21026
rect 45836 20972 45892 20974
rect 45612 20748 45668 20804
rect 46284 20802 46340 20804
rect 46284 20750 46286 20802
rect 46286 20750 46338 20802
rect 46338 20750 46340 20802
rect 46284 20748 46340 20750
rect 45500 20690 45556 20692
rect 45500 20638 45502 20690
rect 45502 20638 45554 20690
rect 45554 20638 45556 20690
rect 45500 20636 45556 20638
rect 46396 20524 46452 20580
rect 46844 35196 46900 35252
rect 46956 35084 47012 35140
rect 46956 34636 47012 34692
rect 47180 34636 47236 34692
rect 46956 34076 47012 34132
rect 46732 29148 46788 29204
rect 47292 34524 47348 34580
rect 47180 29538 47236 29540
rect 47180 29486 47182 29538
rect 47182 29486 47234 29538
rect 47234 29486 47236 29538
rect 47180 29484 47236 29486
rect 46844 28252 46900 28308
rect 47180 28252 47236 28308
rect 46732 28140 46788 28196
rect 46844 27804 46900 27860
rect 47404 34130 47460 34132
rect 47404 34078 47406 34130
rect 47406 34078 47458 34130
rect 47458 34078 47460 34130
rect 47404 34076 47460 34078
rect 47964 35474 48020 35476
rect 47964 35422 47966 35474
rect 47966 35422 48018 35474
rect 48018 35422 48020 35474
rect 47964 35420 48020 35422
rect 47964 34242 48020 34244
rect 47964 34190 47966 34242
rect 47966 34190 48018 34242
rect 48018 34190 48020 34242
rect 47964 34188 48020 34190
rect 48636 36258 48692 36260
rect 48636 36206 48638 36258
rect 48638 36206 48690 36258
rect 48690 36206 48692 36258
rect 48636 36204 48692 36206
rect 49532 36652 49588 36708
rect 48748 34242 48804 34244
rect 48748 34190 48750 34242
rect 48750 34190 48802 34242
rect 48802 34190 48804 34242
rect 48748 34188 48804 34190
rect 49084 36370 49140 36372
rect 49084 36318 49086 36370
rect 49086 36318 49138 36370
rect 49138 36318 49140 36370
rect 49084 36316 49140 36318
rect 48972 34130 49028 34132
rect 48972 34078 48974 34130
rect 48974 34078 49026 34130
rect 49026 34078 49028 34130
rect 48972 34076 49028 34078
rect 47740 33516 47796 33572
rect 47964 32562 48020 32564
rect 47964 32510 47966 32562
rect 47966 32510 48018 32562
rect 48018 32510 48020 32562
rect 47964 32508 48020 32510
rect 47516 31836 47572 31892
rect 48188 31836 48244 31892
rect 47516 30828 47572 30884
rect 47852 31052 47908 31108
rect 47404 29426 47460 29428
rect 47404 29374 47406 29426
rect 47406 29374 47458 29426
rect 47458 29374 47460 29426
rect 47404 29372 47460 29374
rect 47852 30380 47908 30436
rect 48860 31052 48916 31108
rect 48860 30882 48916 30884
rect 48860 30830 48862 30882
rect 48862 30830 48914 30882
rect 48914 30830 48916 30882
rect 48860 30828 48916 30830
rect 48188 30098 48244 30100
rect 48188 30046 48190 30098
rect 48190 30046 48242 30098
rect 48242 30046 48244 30098
rect 48188 30044 48244 30046
rect 48748 30044 48804 30100
rect 47852 29538 47908 29540
rect 47852 29486 47854 29538
rect 47854 29486 47906 29538
rect 47906 29486 47908 29538
rect 47852 29484 47908 29486
rect 47404 28642 47460 28644
rect 47404 28590 47406 28642
rect 47406 28590 47458 28642
rect 47458 28590 47460 28642
rect 47404 28588 47460 28590
rect 48076 28252 48132 28308
rect 48860 28082 48916 28084
rect 48860 28030 48862 28082
rect 48862 28030 48914 28082
rect 48914 28030 48916 28082
rect 48860 28028 48916 28030
rect 47852 27916 47908 27972
rect 48636 27916 48692 27972
rect 46620 23436 46676 23492
rect 46956 23772 47012 23828
rect 46620 23100 46676 23156
rect 46620 20748 46676 20804
rect 47292 26236 47348 26292
rect 47516 25004 47572 25060
rect 49084 30156 49140 30212
rect 49084 29314 49140 29316
rect 49084 29262 49086 29314
rect 49086 29262 49138 29314
rect 49138 29262 49140 29314
rect 49084 29260 49140 29262
rect 49980 36594 50036 36596
rect 49980 36542 49982 36594
rect 49982 36542 50034 36594
rect 50034 36542 50036 36594
rect 49980 36540 50036 36542
rect 50428 36594 50484 36596
rect 50428 36542 50430 36594
rect 50430 36542 50482 36594
rect 50482 36542 50484 36594
rect 50428 36540 50484 36542
rect 50988 36540 51044 36596
rect 50092 35810 50148 35812
rect 50092 35758 50094 35810
rect 50094 35758 50146 35810
rect 50146 35758 50148 35810
rect 50092 35756 50148 35758
rect 50316 35420 50372 35476
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50428 35532 50484 35588
rect 49868 34690 49924 34692
rect 49868 34638 49870 34690
rect 49870 34638 49922 34690
rect 49922 34638 49924 34690
rect 49868 34636 49924 34638
rect 50204 34748 50260 34804
rect 49756 34076 49812 34132
rect 50652 35308 50708 35364
rect 50204 33628 50260 33684
rect 49420 31612 49476 31668
rect 50092 31500 50148 31556
rect 49644 30380 49700 30436
rect 49756 29932 49812 29988
rect 49980 29426 50036 29428
rect 49980 29374 49982 29426
rect 49982 29374 50034 29426
rect 50034 29374 50036 29426
rect 49980 29372 50036 29374
rect 49868 28754 49924 28756
rect 49868 28702 49870 28754
rect 49870 28702 49922 28754
rect 49922 28702 49924 28754
rect 49868 28700 49924 28702
rect 49980 27916 50036 27972
rect 50316 32396 50372 32452
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 51100 35644 51156 35700
rect 51772 35420 51828 35476
rect 51548 34972 51604 35028
rect 51660 34914 51716 34916
rect 51660 34862 51662 34914
rect 51662 34862 51714 34914
rect 51714 34862 51716 34914
rect 51660 34860 51716 34862
rect 53340 40460 53396 40516
rect 53452 40402 53508 40404
rect 53452 40350 53454 40402
rect 53454 40350 53506 40402
rect 53506 40350 53508 40402
rect 53452 40348 53508 40350
rect 54908 44380 54964 44436
rect 54572 43148 54628 43204
rect 55020 43036 55076 43092
rect 53676 41244 53732 41300
rect 55132 41916 55188 41972
rect 54796 41132 54852 41188
rect 53564 40124 53620 40180
rect 55580 42252 55636 42308
rect 55356 41692 55412 41748
rect 55244 39788 55300 39844
rect 55356 40236 55412 40292
rect 55804 40348 55860 40404
rect 55020 39004 55076 39060
rect 53004 38946 53060 38948
rect 53004 38894 53006 38946
rect 53006 38894 53058 38946
rect 53058 38894 53060 38946
rect 53004 38892 53060 38894
rect 53452 38834 53508 38836
rect 53452 38782 53454 38834
rect 53454 38782 53506 38834
rect 53506 38782 53508 38834
rect 53452 38780 53508 38782
rect 52220 37378 52276 37380
rect 52220 37326 52222 37378
rect 52222 37326 52274 37378
rect 52274 37326 52276 37378
rect 52220 37324 52276 37326
rect 52668 36988 52724 37044
rect 52556 36540 52612 36596
rect 52108 36370 52164 36372
rect 52108 36318 52110 36370
rect 52110 36318 52162 36370
rect 52162 36318 52164 36370
rect 52108 36316 52164 36318
rect 52220 35980 52276 36036
rect 52108 35644 52164 35700
rect 51996 35420 52052 35476
rect 51996 34972 52052 35028
rect 53116 36988 53172 37044
rect 53116 36316 53172 36372
rect 53004 35980 53060 36036
rect 52892 35810 52948 35812
rect 52892 35758 52894 35810
rect 52894 35758 52946 35810
rect 52946 35758 52948 35810
rect 52892 35756 52948 35758
rect 52220 35308 52276 35364
rect 50988 33964 51044 34020
rect 51436 33458 51492 33460
rect 51436 33406 51438 33458
rect 51438 33406 51490 33458
rect 51490 33406 51492 33458
rect 51436 33404 51492 33406
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50540 32786 50596 32788
rect 50540 32734 50542 32786
rect 50542 32734 50594 32786
rect 50594 32734 50596 32786
rect 50540 32732 50596 32734
rect 51772 33906 51828 33908
rect 51772 33854 51774 33906
rect 51774 33854 51826 33906
rect 51826 33854 51828 33906
rect 51772 33852 51828 33854
rect 52444 35532 52500 35588
rect 53004 35532 53060 35588
rect 52780 34914 52836 34916
rect 52780 34862 52782 34914
rect 52782 34862 52834 34914
rect 52834 34862 52836 34914
rect 52780 34860 52836 34862
rect 53788 37212 53844 37268
rect 53788 36988 53844 37044
rect 54460 36594 54516 36596
rect 54460 36542 54462 36594
rect 54462 36542 54514 36594
rect 54514 36542 54516 36594
rect 54460 36540 54516 36542
rect 53452 35698 53508 35700
rect 53452 35646 53454 35698
rect 53454 35646 53506 35698
rect 53506 35646 53508 35698
rect 53452 35644 53508 35646
rect 56588 40626 56644 40628
rect 56588 40574 56590 40626
rect 56590 40574 56642 40626
rect 56642 40574 56644 40626
rect 56588 40572 56644 40574
rect 57148 40460 57204 40516
rect 56700 40290 56756 40292
rect 56700 40238 56702 40290
rect 56702 40238 56754 40290
rect 56754 40238 56756 40290
rect 56700 40236 56756 40238
rect 56028 39676 56084 39732
rect 56588 39394 56644 39396
rect 56588 39342 56590 39394
rect 56590 39342 56642 39394
rect 56642 39342 56644 39394
rect 56588 39340 56644 39342
rect 56700 38946 56756 38948
rect 56700 38894 56702 38946
rect 56702 38894 56754 38946
rect 56754 38894 56756 38946
rect 56700 38892 56756 38894
rect 57708 42364 57764 42420
rect 57932 43708 57988 43764
rect 57820 40348 57876 40404
rect 57372 38332 57428 38388
rect 57932 37660 57988 37716
rect 55356 36988 55412 37044
rect 58044 36316 58100 36372
rect 55020 35644 55076 35700
rect 55580 35868 55636 35924
rect 55356 34972 55412 35028
rect 51996 33964 52052 34020
rect 51884 33628 51940 33684
rect 52220 33516 52276 33572
rect 52556 33628 52612 33684
rect 52668 33516 52724 33572
rect 51884 32732 51940 32788
rect 51660 32620 51716 32676
rect 50876 31778 50932 31780
rect 50876 31726 50878 31778
rect 50878 31726 50930 31778
rect 50930 31726 50932 31778
rect 50876 31724 50932 31726
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50988 30156 51044 30212
rect 50540 30098 50596 30100
rect 50540 30046 50542 30098
rect 50542 30046 50594 30098
rect 50594 30046 50596 30098
rect 50540 30044 50596 30046
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50428 28642 50484 28644
rect 50428 28590 50430 28642
rect 50430 28590 50482 28642
rect 50482 28590 50484 28642
rect 50428 28588 50484 28590
rect 51212 30044 51268 30100
rect 50876 29426 50932 29428
rect 50876 29374 50878 29426
rect 50878 29374 50930 29426
rect 50930 29374 50932 29426
rect 50876 29372 50932 29374
rect 51884 32562 51940 32564
rect 51884 32510 51886 32562
rect 51886 32510 51938 32562
rect 51938 32510 51940 32562
rect 51884 32508 51940 32510
rect 51436 30380 51492 30436
rect 51548 31724 51604 31780
rect 52220 32562 52276 32564
rect 52220 32510 52222 32562
rect 52222 32510 52274 32562
rect 52274 32510 52276 32562
rect 52220 32508 52276 32510
rect 52556 31778 52612 31780
rect 52556 31726 52558 31778
rect 52558 31726 52610 31778
rect 52610 31726 52612 31778
rect 52556 31724 52612 31726
rect 51996 30882 52052 30884
rect 51996 30830 51998 30882
rect 51998 30830 52050 30882
rect 52050 30830 52052 30882
rect 51996 30828 52052 30830
rect 52108 30268 52164 30324
rect 52220 30492 52276 30548
rect 51996 30098 52052 30100
rect 51996 30046 51998 30098
rect 51998 30046 52050 30098
rect 52050 30046 52052 30098
rect 51996 30044 52052 30046
rect 51436 29986 51492 29988
rect 51436 29934 51438 29986
rect 51438 29934 51490 29986
rect 51490 29934 51492 29986
rect 51436 29932 51492 29934
rect 50316 27916 50372 27972
rect 51436 28530 51492 28532
rect 51436 28478 51438 28530
rect 51438 28478 51490 28530
rect 51490 28478 51492 28530
rect 51436 28476 51492 28478
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 51212 28252 51268 28308
rect 51996 29260 52052 29316
rect 52444 29932 52500 29988
rect 57932 34300 57988 34356
rect 53228 33404 53284 33460
rect 53228 32732 53284 32788
rect 53564 33404 53620 33460
rect 53788 32172 53844 32228
rect 55356 33122 55412 33124
rect 55356 33070 55358 33122
rect 55358 33070 55410 33122
rect 55410 33070 55412 33122
rect 55356 33068 55412 33070
rect 55916 32732 55972 32788
rect 52892 31500 52948 31556
rect 53004 31276 53060 31332
rect 52780 30156 52836 30212
rect 52780 29986 52836 29988
rect 52780 29934 52782 29986
rect 52782 29934 52834 29986
rect 52834 29934 52836 29986
rect 52780 29932 52836 29934
rect 53004 30770 53060 30772
rect 53004 30718 53006 30770
rect 53006 30718 53058 30770
rect 53058 30718 53060 30770
rect 53004 30716 53060 30718
rect 55020 31612 55076 31668
rect 53340 31276 53396 31332
rect 53004 30098 53060 30100
rect 53004 30046 53006 30098
rect 53006 30046 53058 30098
rect 53058 30046 53060 30098
rect 53004 30044 53060 30046
rect 54236 31276 54292 31332
rect 54796 31276 54852 31332
rect 54460 31164 54516 31220
rect 54908 31218 54964 31220
rect 54908 31166 54910 31218
rect 54910 31166 54962 31218
rect 54962 31166 54964 31218
rect 54908 31164 54964 31166
rect 55692 31164 55748 31220
rect 56364 31164 56420 31220
rect 54684 30994 54740 30996
rect 54684 30942 54686 30994
rect 54686 30942 54738 30994
rect 54738 30942 54740 30994
rect 54684 30940 54740 30942
rect 54236 30156 54292 30212
rect 54124 30098 54180 30100
rect 54124 30046 54126 30098
rect 54126 30046 54178 30098
rect 54178 30046 54180 30098
rect 54124 30044 54180 30046
rect 54012 29708 54068 29764
rect 52556 29484 52612 29540
rect 52892 29148 52948 29204
rect 52892 28588 52948 28644
rect 53004 28476 53060 28532
rect 52780 28418 52836 28420
rect 52780 28366 52782 28418
rect 52782 28366 52834 28418
rect 52834 28366 52836 28418
rect 52780 28364 52836 28366
rect 52668 28252 52724 28308
rect 51548 27074 51604 27076
rect 51548 27022 51550 27074
rect 51550 27022 51602 27074
rect 51602 27022 51604 27074
rect 51548 27020 51604 27022
rect 51772 27074 51828 27076
rect 51772 27022 51774 27074
rect 51774 27022 51826 27074
rect 51826 27022 51828 27074
rect 51772 27020 51828 27022
rect 47852 26236 47908 26292
rect 48748 26684 48804 26740
rect 47964 26178 48020 26180
rect 47964 26126 47966 26178
rect 47966 26126 48018 26178
rect 48018 26126 48020 26178
rect 47964 26124 48020 26126
rect 47740 25564 47796 25620
rect 47740 25116 47796 25172
rect 48076 25282 48132 25284
rect 48076 25230 48078 25282
rect 48078 25230 48130 25282
rect 48130 25230 48132 25282
rect 48076 25228 48132 25230
rect 47404 23938 47460 23940
rect 47404 23886 47406 23938
rect 47406 23886 47458 23938
rect 47458 23886 47460 23938
rect 47404 23884 47460 23886
rect 47628 23772 47684 23828
rect 47516 23154 47572 23156
rect 47516 23102 47518 23154
rect 47518 23102 47570 23154
rect 47570 23102 47572 23154
rect 47516 23100 47572 23102
rect 47068 23042 47124 23044
rect 47068 22990 47070 23042
rect 47070 22990 47122 23042
rect 47122 22990 47124 23042
rect 47068 22988 47124 22990
rect 48636 24108 48692 24164
rect 48524 23884 48580 23940
rect 47852 22988 47908 23044
rect 48076 23100 48132 23156
rect 47068 20690 47124 20692
rect 47068 20638 47070 20690
rect 47070 20638 47122 20690
rect 47122 20638 47124 20690
rect 47068 20636 47124 20638
rect 46956 20300 47012 20356
rect 48188 21756 48244 21812
rect 46732 20188 46788 20244
rect 46620 20130 46676 20132
rect 46620 20078 46622 20130
rect 46622 20078 46674 20130
rect 46674 20078 46676 20130
rect 46620 20076 46676 20078
rect 47292 20076 47348 20132
rect 45612 19794 45668 19796
rect 45612 19742 45614 19794
rect 45614 19742 45666 19794
rect 45666 19742 45668 19794
rect 45612 19740 45668 19742
rect 45948 19404 46004 19460
rect 46172 19346 46228 19348
rect 46172 19294 46174 19346
rect 46174 19294 46226 19346
rect 46226 19294 46228 19346
rect 46172 19292 46228 19294
rect 46396 18732 46452 18788
rect 45388 18450 45444 18452
rect 45388 18398 45390 18450
rect 45390 18398 45442 18450
rect 45442 18398 45444 18450
rect 45388 18396 45444 18398
rect 44940 16828 44996 16884
rect 43372 16716 43428 16772
rect 43372 16492 43428 16548
rect 43260 16380 43316 16436
rect 42588 15596 42644 15652
rect 43148 15820 43204 15876
rect 42924 15314 42980 15316
rect 42924 15262 42926 15314
rect 42926 15262 42978 15314
rect 42978 15262 42980 15314
rect 42924 15260 42980 15262
rect 43484 15596 43540 15652
rect 42700 14812 42756 14868
rect 43484 15148 43540 15204
rect 43372 14530 43428 14532
rect 43372 14478 43374 14530
rect 43374 14478 43426 14530
rect 43426 14478 43428 14530
rect 43372 14476 43428 14478
rect 43596 15314 43652 15316
rect 43596 15262 43598 15314
rect 43598 15262 43650 15314
rect 43650 15262 43652 15314
rect 43596 15260 43652 15262
rect 43820 15874 43876 15876
rect 43820 15822 43822 15874
rect 43822 15822 43874 15874
rect 43874 15822 43876 15874
rect 43820 15820 43876 15822
rect 43932 15372 43988 15428
rect 42252 13580 42308 13636
rect 41916 13020 41972 13076
rect 42700 13692 42756 13748
rect 43036 13692 43092 13748
rect 42588 13468 42644 13524
rect 42364 13020 42420 13076
rect 42140 12684 42196 12740
rect 42364 12738 42420 12740
rect 42364 12686 42366 12738
rect 42366 12686 42418 12738
rect 42418 12686 42420 12738
rect 42364 12684 42420 12686
rect 41468 11228 41524 11284
rect 42812 12236 42868 12292
rect 42364 11452 42420 11508
rect 41804 11116 41860 11172
rect 41132 9826 41188 9828
rect 41132 9774 41134 9826
rect 41134 9774 41186 9826
rect 41186 9774 41188 9826
rect 41132 9772 41188 9774
rect 41244 9660 41300 9716
rect 41020 9212 41076 9268
rect 41356 9042 41412 9044
rect 41356 8990 41358 9042
rect 41358 8990 41410 9042
rect 41410 8990 41412 9042
rect 41356 8988 41412 8990
rect 42252 11282 42308 11284
rect 42252 11230 42254 11282
rect 42254 11230 42306 11282
rect 42306 11230 42308 11282
rect 42252 11228 42308 11230
rect 42700 11282 42756 11284
rect 42700 11230 42702 11282
rect 42702 11230 42754 11282
rect 42754 11230 42756 11282
rect 42700 11228 42756 11230
rect 42364 11116 42420 11172
rect 43148 13356 43204 13412
rect 44044 13746 44100 13748
rect 44044 13694 44046 13746
rect 44046 13694 44098 13746
rect 44098 13694 44100 13746
rect 44044 13692 44100 13694
rect 44268 13356 44324 13412
rect 44492 15314 44548 15316
rect 44492 15262 44494 15314
rect 44494 15262 44546 15314
rect 44546 15262 44548 15314
rect 44492 15260 44548 15262
rect 45164 17052 45220 17108
rect 45724 17442 45780 17444
rect 45724 17390 45726 17442
rect 45726 17390 45778 17442
rect 45778 17390 45780 17442
rect 45724 17388 45780 17390
rect 45948 17554 46004 17556
rect 45948 17502 45950 17554
rect 45950 17502 46002 17554
rect 46002 17502 46004 17554
rect 45948 17500 46004 17502
rect 46172 17554 46228 17556
rect 46172 17502 46174 17554
rect 46174 17502 46226 17554
rect 46226 17502 46228 17554
rect 46172 17500 46228 17502
rect 47068 18396 47124 18452
rect 47180 17612 47236 17668
rect 46732 17500 46788 17556
rect 46060 17106 46116 17108
rect 46060 17054 46062 17106
rect 46062 17054 46114 17106
rect 46114 17054 46116 17106
rect 46060 17052 46116 17054
rect 45836 16940 45892 16996
rect 45948 16882 46004 16884
rect 45948 16830 45950 16882
rect 45950 16830 46002 16882
rect 46002 16830 46004 16882
rect 45948 16828 46004 16830
rect 46620 16940 46676 16996
rect 45276 16268 45332 16324
rect 44828 15036 44884 15092
rect 46060 16156 46116 16212
rect 45276 15372 45332 15428
rect 45164 15148 45220 15204
rect 45948 14140 46004 14196
rect 46060 15372 46116 15428
rect 44828 13970 44884 13972
rect 44828 13918 44830 13970
rect 44830 13918 44882 13970
rect 44882 13918 44884 13970
rect 44828 13916 44884 13918
rect 46172 15260 46228 15316
rect 44156 12850 44212 12852
rect 44156 12798 44158 12850
rect 44158 12798 44210 12850
rect 44210 12798 44212 12850
rect 44156 12796 44212 12798
rect 43260 12684 43316 12740
rect 43148 12348 43204 12404
rect 46172 12290 46228 12292
rect 46172 12238 46174 12290
rect 46174 12238 46226 12290
rect 46226 12238 46228 12290
rect 46172 12236 46228 12238
rect 44716 11788 44772 11844
rect 43372 11452 43428 11508
rect 45724 11788 45780 11844
rect 44716 11452 44772 11508
rect 42252 10834 42308 10836
rect 42252 10782 42254 10834
rect 42254 10782 42306 10834
rect 42306 10782 42308 10834
rect 42252 10780 42308 10782
rect 42140 10668 42196 10724
rect 41244 8316 41300 8372
rect 41580 9772 41636 9828
rect 41580 9100 41636 9156
rect 41356 7756 41412 7812
rect 41692 9548 41748 9604
rect 42140 9548 42196 9604
rect 42364 9266 42420 9268
rect 42364 9214 42366 9266
rect 42366 9214 42418 9266
rect 42418 9214 42420 9266
rect 42364 9212 42420 9214
rect 42812 10722 42868 10724
rect 42812 10670 42814 10722
rect 42814 10670 42866 10722
rect 42866 10670 42868 10722
rect 42812 10668 42868 10670
rect 42812 10444 42868 10500
rect 43484 11170 43540 11172
rect 43484 11118 43486 11170
rect 43486 11118 43538 11170
rect 43538 11118 43540 11170
rect 43484 11116 43540 11118
rect 44156 11170 44212 11172
rect 44156 11118 44158 11170
rect 44158 11118 44210 11170
rect 44210 11118 44212 11170
rect 44156 11116 44212 11118
rect 43596 10834 43652 10836
rect 43596 10782 43598 10834
rect 43598 10782 43650 10834
rect 43650 10782 43652 10834
rect 43596 10780 43652 10782
rect 43372 10332 43428 10388
rect 44940 11676 44996 11732
rect 44940 10780 44996 10836
rect 45836 11564 45892 11620
rect 44044 10498 44100 10500
rect 44044 10446 44046 10498
rect 44046 10446 44098 10498
rect 44098 10446 44100 10498
rect 44044 10444 44100 10446
rect 43484 9826 43540 9828
rect 43484 9774 43486 9826
rect 43486 9774 43538 9826
rect 43538 9774 43540 9826
rect 43484 9772 43540 9774
rect 43932 9826 43988 9828
rect 43932 9774 43934 9826
rect 43934 9774 43986 9826
rect 43986 9774 43988 9826
rect 43932 9772 43988 9774
rect 42700 9212 42756 9268
rect 43708 9602 43764 9604
rect 43708 9550 43710 9602
rect 43710 9550 43762 9602
rect 43762 9550 43764 9602
rect 43708 9548 43764 9550
rect 44828 9602 44884 9604
rect 44828 9550 44830 9602
rect 44830 9550 44882 9602
rect 44882 9550 44884 9602
rect 44828 9548 44884 9550
rect 45836 10332 45892 10388
rect 46060 9266 46116 9268
rect 46060 9214 46062 9266
rect 46062 9214 46114 9266
rect 46114 9214 46116 9266
rect 46060 9212 46116 9214
rect 41804 8146 41860 8148
rect 41804 8094 41806 8146
rect 41806 8094 41858 8146
rect 41858 8094 41860 8146
rect 41804 8092 41860 8094
rect 42924 8146 42980 8148
rect 42924 8094 42926 8146
rect 42926 8094 42978 8146
rect 42978 8094 42980 8146
rect 42924 8092 42980 8094
rect 43036 7756 43092 7812
rect 42700 7644 42756 7700
rect 46508 16322 46564 16324
rect 46508 16270 46510 16322
rect 46510 16270 46562 16322
rect 46562 16270 46564 16322
rect 46508 16268 46564 16270
rect 47068 17388 47124 17444
rect 47292 17500 47348 17556
rect 47068 16268 47124 16324
rect 47180 16156 47236 16212
rect 46956 15426 47012 15428
rect 46956 15374 46958 15426
rect 46958 15374 47010 15426
rect 47010 15374 47012 15426
rect 46956 15372 47012 15374
rect 46620 15314 46676 15316
rect 46620 15262 46622 15314
rect 46622 15262 46674 15314
rect 46674 15262 46676 15314
rect 46620 15260 46676 15262
rect 46844 15260 46900 15316
rect 46396 15148 46452 15204
rect 47292 15314 47348 15316
rect 47292 15262 47294 15314
rect 47294 15262 47346 15314
rect 47346 15262 47348 15314
rect 47292 15260 47348 15262
rect 47516 20300 47572 20356
rect 47852 20578 47908 20580
rect 47852 20526 47854 20578
rect 47854 20526 47906 20578
rect 47906 20526 47908 20578
rect 47852 20524 47908 20526
rect 48748 23266 48804 23268
rect 48748 23214 48750 23266
rect 48750 23214 48802 23266
rect 48802 23214 48804 23266
rect 48748 23212 48804 23214
rect 48860 21644 48916 21700
rect 49196 25506 49252 25508
rect 49196 25454 49198 25506
rect 49198 25454 49250 25506
rect 49250 25454 49252 25506
rect 49196 25452 49252 25454
rect 49644 25676 49700 25732
rect 49420 25228 49476 25284
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50988 26348 51044 26404
rect 50316 26124 50372 26180
rect 50316 25394 50372 25396
rect 50316 25342 50318 25394
rect 50318 25342 50370 25394
rect 50370 25342 50372 25394
rect 50316 25340 50372 25342
rect 50204 25004 50260 25060
rect 50204 24780 50260 24836
rect 50092 24108 50148 24164
rect 50652 26290 50708 26292
rect 50652 26238 50654 26290
rect 50654 26238 50706 26290
rect 50706 26238 50708 26290
rect 50652 26236 50708 26238
rect 50876 25564 50932 25620
rect 51660 26402 51716 26404
rect 51660 26350 51662 26402
rect 51662 26350 51714 26402
rect 51714 26350 51716 26402
rect 51660 26348 51716 26350
rect 52220 27468 52276 27524
rect 52220 27132 52276 27188
rect 52108 26236 52164 26292
rect 52220 26908 52276 26964
rect 50988 25452 51044 25508
rect 50540 25394 50596 25396
rect 50540 25342 50542 25394
rect 50542 25342 50594 25394
rect 50594 25342 50596 25394
rect 50540 25340 50596 25342
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50988 25116 51044 25172
rect 51212 25228 51268 25284
rect 51660 25506 51716 25508
rect 51660 25454 51662 25506
rect 51662 25454 51714 25506
rect 51714 25454 51716 25506
rect 51660 25452 51716 25454
rect 52556 27804 52612 27860
rect 52556 27132 52612 27188
rect 53340 28642 53396 28644
rect 53340 28590 53342 28642
rect 53342 28590 53394 28642
rect 53394 28590 53396 28642
rect 53340 28588 53396 28590
rect 53116 28252 53172 28308
rect 53004 27468 53060 27524
rect 52668 27074 52724 27076
rect 52668 27022 52670 27074
rect 52670 27022 52722 27074
rect 52722 27022 52724 27074
rect 52668 27020 52724 27022
rect 52892 26962 52948 26964
rect 52892 26910 52894 26962
rect 52894 26910 52946 26962
rect 52946 26910 52948 26962
rect 52892 26908 52948 26910
rect 53788 29538 53844 29540
rect 53788 29486 53790 29538
rect 53790 29486 53842 29538
rect 53842 29486 53844 29538
rect 53788 29484 53844 29486
rect 54124 29426 54180 29428
rect 54124 29374 54126 29426
rect 54126 29374 54178 29426
rect 54178 29374 54180 29426
rect 54124 29372 54180 29374
rect 53788 28588 53844 28644
rect 53900 28924 53956 28980
rect 53900 28252 53956 28308
rect 54124 28642 54180 28644
rect 54124 28590 54126 28642
rect 54126 28590 54178 28642
rect 54178 28590 54180 28642
rect 54124 28588 54180 28590
rect 54012 27468 54068 27524
rect 54460 30268 54516 30324
rect 55580 30994 55636 30996
rect 55580 30942 55582 30994
rect 55582 30942 55634 30994
rect 55634 30942 55636 30994
rect 55580 30940 55636 30942
rect 54796 30044 54852 30100
rect 54908 30716 54964 30772
rect 54684 29538 54740 29540
rect 54684 29486 54686 29538
rect 54686 29486 54738 29538
rect 54738 29486 54740 29538
rect 54684 29484 54740 29486
rect 54684 29202 54740 29204
rect 54684 29150 54686 29202
rect 54686 29150 54738 29202
rect 54738 29150 54740 29202
rect 54684 29148 54740 29150
rect 54684 28924 54740 28980
rect 55916 30156 55972 30212
rect 55804 29708 55860 29764
rect 55020 29372 55076 29428
rect 55244 29260 55300 29316
rect 56140 28700 56196 28756
rect 54684 28252 54740 28308
rect 54684 27858 54740 27860
rect 54684 27806 54686 27858
rect 54686 27806 54738 27858
rect 54738 27806 54740 27858
rect 54684 27804 54740 27806
rect 54012 27132 54068 27188
rect 52892 26402 52948 26404
rect 52892 26350 52894 26402
rect 52894 26350 52946 26402
rect 52946 26350 52948 26402
rect 52892 26348 52948 26350
rect 53788 26348 53844 26404
rect 52332 26124 52388 26180
rect 53676 26178 53732 26180
rect 53676 26126 53678 26178
rect 53678 26126 53730 26178
rect 53730 26126 53732 26178
rect 53676 26124 53732 26126
rect 51884 25116 51940 25172
rect 51436 25004 51492 25060
rect 50876 24780 50932 24836
rect 51100 24780 51156 24836
rect 50988 24722 51044 24724
rect 50988 24670 50990 24722
rect 50990 24670 51042 24722
rect 51042 24670 51044 24722
rect 50988 24668 51044 24670
rect 49084 23714 49140 23716
rect 49084 23662 49086 23714
rect 49086 23662 49138 23714
rect 49138 23662 49140 23714
rect 49084 23660 49140 23662
rect 49420 23154 49476 23156
rect 49420 23102 49422 23154
rect 49422 23102 49474 23154
rect 49474 23102 49476 23154
rect 49420 23100 49476 23102
rect 50652 24108 50708 24164
rect 50876 23938 50932 23940
rect 50876 23886 50878 23938
rect 50878 23886 50930 23938
rect 50930 23886 50932 23938
rect 50876 23884 50932 23886
rect 51212 23772 51268 23828
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50428 23212 50484 23268
rect 51884 24108 51940 24164
rect 52780 25394 52836 25396
rect 52780 25342 52782 25394
rect 52782 25342 52834 25394
rect 52834 25342 52836 25394
rect 52780 25340 52836 25342
rect 52892 25004 52948 25060
rect 52780 24722 52836 24724
rect 52780 24670 52782 24722
rect 52782 24670 52834 24722
rect 52834 24670 52836 24722
rect 52780 24668 52836 24670
rect 52332 24610 52388 24612
rect 52332 24558 52334 24610
rect 52334 24558 52386 24610
rect 52386 24558 52388 24610
rect 52332 24556 52388 24558
rect 53340 25282 53396 25284
rect 53340 25230 53342 25282
rect 53342 25230 53394 25282
rect 53394 25230 53396 25282
rect 53340 25228 53396 25230
rect 53004 24668 53060 24724
rect 53116 24162 53172 24164
rect 53116 24110 53118 24162
rect 53118 24110 53170 24162
rect 53170 24110 53172 24162
rect 53116 24108 53172 24110
rect 52444 23772 52500 23828
rect 54460 26460 54516 26516
rect 55356 28476 55412 28532
rect 53788 25564 53844 25620
rect 53676 24722 53732 24724
rect 53676 24670 53678 24722
rect 53678 24670 53730 24722
rect 53730 24670 53732 24722
rect 53676 24668 53732 24670
rect 53788 24108 53844 24164
rect 49196 21868 49252 21924
rect 50092 22594 50148 22596
rect 50092 22542 50094 22594
rect 50094 22542 50146 22594
rect 50146 22542 50148 22594
rect 50092 22540 50148 22542
rect 49532 21810 49588 21812
rect 49532 21758 49534 21810
rect 49534 21758 49586 21810
rect 49586 21758 49588 21810
rect 49532 21756 49588 21758
rect 48524 20076 48580 20132
rect 47628 18396 47684 18452
rect 48972 21196 49028 21252
rect 48860 20130 48916 20132
rect 48860 20078 48862 20130
rect 48862 20078 48914 20130
rect 48914 20078 48916 20130
rect 48860 20076 48916 20078
rect 48860 18450 48916 18452
rect 48860 18398 48862 18450
rect 48862 18398 48914 18450
rect 48914 18398 48916 18450
rect 48860 18396 48916 18398
rect 47964 17388 48020 17444
rect 48748 17500 48804 17556
rect 48188 16716 48244 16772
rect 48748 16716 48804 16772
rect 47852 16380 47908 16436
rect 47516 16268 47572 16324
rect 47516 16098 47572 16100
rect 47516 16046 47518 16098
rect 47518 16046 47570 16098
rect 47570 16046 47572 16098
rect 47516 16044 47572 16046
rect 48076 15932 48132 15988
rect 47964 15820 48020 15876
rect 47740 15426 47796 15428
rect 47740 15374 47742 15426
rect 47742 15374 47794 15426
rect 47794 15374 47796 15426
rect 47740 15372 47796 15374
rect 48748 15932 48804 15988
rect 48524 15874 48580 15876
rect 48524 15822 48526 15874
rect 48526 15822 48578 15874
rect 48578 15822 48580 15874
rect 48524 15820 48580 15822
rect 47068 14812 47124 14868
rect 46620 13916 46676 13972
rect 50988 23154 51044 23156
rect 50988 23102 50990 23154
rect 50990 23102 51042 23154
rect 51042 23102 51044 23154
rect 50988 23100 51044 23102
rect 50876 22652 50932 22708
rect 50988 22594 51044 22596
rect 50988 22542 50990 22594
rect 50990 22542 51042 22594
rect 51042 22542 51044 22594
rect 50988 22540 51044 22542
rect 52220 23212 52276 23268
rect 53564 23212 53620 23268
rect 50092 21868 50148 21924
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50204 21644 50260 21700
rect 50204 20914 50260 20916
rect 50204 20862 50206 20914
rect 50206 20862 50258 20914
rect 50258 20862 50260 20914
rect 50204 20860 50260 20862
rect 50540 21644 50596 21700
rect 50428 21586 50484 21588
rect 50428 21534 50430 21586
rect 50430 21534 50482 21586
rect 50482 21534 50484 21586
rect 50428 21532 50484 21534
rect 51100 21810 51156 21812
rect 51100 21758 51102 21810
rect 51102 21758 51154 21810
rect 51154 21758 51156 21810
rect 51100 21756 51156 21758
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 49980 19852 50036 19908
rect 49756 18396 49812 18452
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50428 18396 50484 18452
rect 49196 16770 49252 16772
rect 49196 16718 49198 16770
rect 49198 16718 49250 16770
rect 49250 16718 49252 16770
rect 49196 16716 49252 16718
rect 49420 16716 49476 16772
rect 49084 16380 49140 16436
rect 51772 22258 51828 22260
rect 51772 22206 51774 22258
rect 51774 22206 51826 22258
rect 51826 22206 51828 22258
rect 51772 22204 51828 22206
rect 51660 21756 51716 21812
rect 52780 22652 52836 22708
rect 52892 22258 52948 22260
rect 52892 22206 52894 22258
rect 52894 22206 52946 22258
rect 52946 22206 52948 22258
rect 52892 22204 52948 22206
rect 51548 21586 51604 21588
rect 51548 21534 51550 21586
rect 51550 21534 51602 21586
rect 51602 21534 51604 21586
rect 51548 21532 51604 21534
rect 51548 20972 51604 21028
rect 51996 21644 52052 21700
rect 52108 21420 52164 21476
rect 51548 20802 51604 20804
rect 51548 20750 51550 20802
rect 51550 20750 51602 20802
rect 51602 20750 51604 20802
rect 51548 20748 51604 20750
rect 53788 22146 53844 22148
rect 53788 22094 53790 22146
rect 53790 22094 53842 22146
rect 53842 22094 53844 22146
rect 53788 22092 53844 22094
rect 53452 21980 53508 22036
rect 52892 21810 52948 21812
rect 52892 21758 52894 21810
rect 52894 21758 52946 21810
rect 52946 21758 52948 21810
rect 52892 21756 52948 21758
rect 52444 21698 52500 21700
rect 52444 21646 52446 21698
rect 52446 21646 52498 21698
rect 52498 21646 52500 21698
rect 52444 21644 52500 21646
rect 53116 21644 53172 21700
rect 52668 21026 52724 21028
rect 52668 20974 52670 21026
rect 52670 20974 52722 21026
rect 52722 20974 52724 21026
rect 52668 20972 52724 20974
rect 53676 21756 53732 21812
rect 52108 20748 52164 20804
rect 52220 20860 52276 20916
rect 51996 20524 52052 20580
rect 53228 20914 53284 20916
rect 53228 20862 53230 20914
rect 53230 20862 53282 20914
rect 53282 20862 53284 20914
rect 53228 20860 53284 20862
rect 52444 20748 52500 20804
rect 52444 20018 52500 20020
rect 52444 19966 52446 20018
rect 52446 19966 52498 20018
rect 52498 19966 52500 20018
rect 52444 19964 52500 19966
rect 52780 19068 52836 19124
rect 51996 18450 52052 18452
rect 51996 18398 51998 18450
rect 51998 18398 52050 18450
rect 52050 18398 52052 18450
rect 51996 18396 52052 18398
rect 53004 18396 53060 18452
rect 50764 17666 50820 17668
rect 50764 17614 50766 17666
rect 50766 17614 50818 17666
rect 50818 17614 50820 17666
rect 50764 17612 50820 17614
rect 52332 17612 52388 17668
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50092 16770 50148 16772
rect 50092 16718 50094 16770
rect 50094 16718 50146 16770
rect 50146 16718 50148 16770
rect 50092 16716 50148 16718
rect 50652 16716 50708 16772
rect 49196 16098 49252 16100
rect 49196 16046 49198 16098
rect 49198 16046 49250 16098
rect 49250 16046 49252 16098
rect 49196 16044 49252 16046
rect 51324 17388 51380 17444
rect 51100 16716 51156 16772
rect 50764 16098 50820 16100
rect 50764 16046 50766 16098
rect 50766 16046 50818 16098
rect 50818 16046 50820 16098
rect 50764 16044 50820 16046
rect 50540 15932 50596 15988
rect 50988 15986 51044 15988
rect 50988 15934 50990 15986
rect 50990 15934 51042 15986
rect 51042 15934 51044 15986
rect 50988 15932 51044 15934
rect 49532 15874 49588 15876
rect 49532 15822 49534 15874
rect 49534 15822 49586 15874
rect 49586 15822 49588 15874
rect 49532 15820 49588 15822
rect 49868 15820 49924 15876
rect 49420 15426 49476 15428
rect 49420 15374 49422 15426
rect 49422 15374 49474 15426
rect 49474 15374 49476 15426
rect 49420 15372 49476 15374
rect 48524 14642 48580 14644
rect 48524 14590 48526 14642
rect 48526 14590 48578 14642
rect 48578 14590 48580 14642
rect 48524 14588 48580 14590
rect 49084 14588 49140 14644
rect 48860 14476 48916 14532
rect 47292 13858 47348 13860
rect 47292 13806 47294 13858
rect 47294 13806 47346 13858
rect 47346 13806 47348 13858
rect 47292 13804 47348 13806
rect 47516 13916 47572 13972
rect 49084 13634 49140 13636
rect 49084 13582 49086 13634
rect 49086 13582 49138 13634
rect 49138 13582 49140 13634
rect 49084 13580 49140 13582
rect 49084 11676 49140 11732
rect 47404 11564 47460 11620
rect 49420 14476 49476 14532
rect 46508 9772 46564 9828
rect 46284 3948 46340 4004
rect 50092 15484 50148 15540
rect 49756 14140 49812 14196
rect 51100 15874 51156 15876
rect 51100 15822 51102 15874
rect 51102 15822 51154 15874
rect 51154 15822 51156 15874
rect 51100 15820 51156 15822
rect 50988 15708 51044 15764
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 51660 15874 51716 15876
rect 51660 15822 51662 15874
rect 51662 15822 51714 15874
rect 51714 15822 51716 15874
rect 51660 15820 51716 15822
rect 52556 15820 52612 15876
rect 51548 15708 51604 15764
rect 51100 15484 51156 15540
rect 50428 15372 50484 15428
rect 52780 15874 52836 15876
rect 52780 15822 52782 15874
rect 52782 15822 52834 15874
rect 52834 15822 52836 15874
rect 52780 15820 52836 15822
rect 54796 25564 54852 25620
rect 54684 24946 54740 24948
rect 54684 24894 54686 24946
rect 54686 24894 54738 24946
rect 54738 24894 54740 24946
rect 54684 24892 54740 24894
rect 55692 27858 55748 27860
rect 55692 27806 55694 27858
rect 55694 27806 55746 27858
rect 55746 27806 55748 27858
rect 55692 27804 55748 27806
rect 55692 27132 55748 27188
rect 56700 31218 56756 31220
rect 56700 31166 56702 31218
rect 56702 31166 56754 31218
rect 56754 31166 56756 31218
rect 56700 31164 56756 31166
rect 58156 30322 58212 30324
rect 58156 30270 58158 30322
rect 58158 30270 58210 30322
rect 58210 30270 58212 30322
rect 58156 30268 58212 30270
rect 57148 29650 57204 29652
rect 57148 29598 57150 29650
rect 57150 29598 57202 29650
rect 57202 29598 57204 29650
rect 57148 29596 57204 29598
rect 57596 29596 57652 29652
rect 57484 28924 57540 28980
rect 58156 29650 58212 29652
rect 58156 29598 58158 29650
rect 58158 29598 58210 29650
rect 58210 29598 58212 29650
rect 58156 29596 58212 29598
rect 57820 29148 57876 29204
rect 57820 28700 57876 28756
rect 56364 28588 56420 28644
rect 57148 28642 57204 28644
rect 57148 28590 57150 28642
rect 57150 28590 57202 28642
rect 57202 28590 57204 28642
rect 57148 28588 57204 28590
rect 58156 28642 58212 28644
rect 58156 28590 58158 28642
rect 58158 28590 58210 28642
rect 58210 28590 58212 28642
rect 58156 28588 58212 28590
rect 58156 28252 58212 28308
rect 56140 27356 56196 27412
rect 57596 27580 57652 27636
rect 58156 27580 58212 27636
rect 57820 27244 57876 27300
rect 58156 27186 58212 27188
rect 58156 27134 58158 27186
rect 58158 27134 58210 27186
rect 58210 27134 58212 27186
rect 58156 27132 58212 27134
rect 55244 26514 55300 26516
rect 55244 26462 55246 26514
rect 55246 26462 55298 26514
rect 55298 26462 55300 26514
rect 55244 26460 55300 26462
rect 55356 26178 55412 26180
rect 55356 26126 55358 26178
rect 55358 26126 55410 26178
rect 55410 26126 55412 26178
rect 55356 26124 55412 26126
rect 55468 25564 55524 25620
rect 55356 25116 55412 25172
rect 54796 23212 54852 23268
rect 54124 21980 54180 22036
rect 55244 24610 55300 24612
rect 55244 24558 55246 24610
rect 55246 24558 55298 24610
rect 55298 24558 55300 24610
rect 55244 24556 55300 24558
rect 56700 26178 56756 26180
rect 56700 26126 56702 26178
rect 56702 26126 56754 26178
rect 56754 26126 56756 26178
rect 56700 26124 56756 26126
rect 57820 26796 57876 26852
rect 58044 26796 58100 26852
rect 57484 26290 57540 26292
rect 57484 26238 57486 26290
rect 57486 26238 57538 26290
rect 57538 26238 57540 26290
rect 57484 26236 57540 26238
rect 57148 26012 57204 26068
rect 56924 25900 56980 25956
rect 58044 25900 58100 25956
rect 57036 25788 57092 25844
rect 58156 25618 58212 25620
rect 58156 25566 58158 25618
rect 58158 25566 58210 25618
rect 58210 25566 58212 25618
rect 58156 25564 58212 25566
rect 57036 25004 57092 25060
rect 57596 25116 57652 25172
rect 57484 24946 57540 24948
rect 57484 24894 57486 24946
rect 57486 24894 57538 24946
rect 57538 24894 57540 24946
rect 57484 24892 57540 24894
rect 55244 23996 55300 24052
rect 56028 24610 56084 24612
rect 56028 24558 56030 24610
rect 56030 24558 56082 24610
rect 56082 24558 56084 24610
rect 56028 24556 56084 24558
rect 57148 24444 57204 24500
rect 55580 23266 55636 23268
rect 55580 23214 55582 23266
rect 55582 23214 55634 23266
rect 55634 23214 55636 23266
rect 55580 23212 55636 23214
rect 57484 23436 57540 23492
rect 55468 23042 55524 23044
rect 55468 22990 55470 23042
rect 55470 22990 55522 23042
rect 55522 22990 55524 23042
rect 55468 22988 55524 22990
rect 53676 19234 53732 19236
rect 53676 19182 53678 19234
rect 53678 19182 53730 19234
rect 53730 19182 53732 19234
rect 53676 19180 53732 19182
rect 53452 19122 53508 19124
rect 53452 19070 53454 19122
rect 53454 19070 53506 19122
rect 53506 19070 53508 19122
rect 53452 19068 53508 19070
rect 54012 21532 54068 21588
rect 56700 23042 56756 23044
rect 56700 22990 56702 23042
rect 56702 22990 56754 23042
rect 56754 22990 56756 23042
rect 56700 22988 56756 22990
rect 54908 21756 54964 21812
rect 57148 22764 57204 22820
rect 57036 22428 57092 22484
rect 55244 22092 55300 22148
rect 55356 21756 55412 21812
rect 55132 21586 55188 21588
rect 55132 21534 55134 21586
rect 55134 21534 55186 21586
rect 55186 21534 55188 21586
rect 55132 21532 55188 21534
rect 54012 20914 54068 20916
rect 54012 20862 54014 20914
rect 54014 20862 54066 20914
rect 54066 20862 54068 20914
rect 54012 20860 54068 20862
rect 55020 21474 55076 21476
rect 55020 21422 55022 21474
rect 55022 21422 55074 21474
rect 55074 21422 55076 21474
rect 55020 21420 55076 21422
rect 54572 19180 54628 19236
rect 53564 18284 53620 18340
rect 53340 17388 53396 17444
rect 53116 15874 53172 15876
rect 53116 15822 53118 15874
rect 53118 15822 53170 15874
rect 53170 15822 53172 15874
rect 53116 15820 53172 15822
rect 52780 15148 52836 15204
rect 51660 14588 51716 14644
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 49756 13970 49812 13972
rect 49756 13918 49758 13970
rect 49758 13918 49810 13970
rect 49810 13918 49812 13970
rect 49756 13916 49812 13918
rect 50764 13916 50820 13972
rect 49644 13804 49700 13860
rect 50092 13858 50148 13860
rect 50092 13806 50094 13858
rect 50094 13806 50146 13858
rect 50146 13806 50148 13858
rect 50092 13804 50148 13806
rect 56812 21756 56868 21812
rect 55692 21474 55748 21476
rect 55692 21422 55694 21474
rect 55694 21422 55746 21474
rect 55746 21422 55748 21474
rect 55692 21420 55748 21422
rect 57036 21756 57092 21812
rect 58156 25116 58212 25172
rect 57820 25004 57876 25060
rect 58156 24220 58212 24276
rect 57932 24050 57988 24052
rect 57932 23998 57934 24050
rect 57934 23998 57986 24050
rect 57986 23998 57988 24050
rect 57932 23996 57988 23998
rect 57820 23378 57876 23380
rect 57820 23326 57822 23378
rect 57822 23326 57874 23378
rect 57874 23326 57876 23378
rect 57820 23324 57876 23326
rect 57932 23212 57988 23268
rect 58156 22204 58212 22260
rect 57820 21810 57876 21812
rect 57820 21758 57822 21810
rect 57822 21758 57874 21810
rect 57874 21758 57876 21810
rect 57820 21756 57876 21758
rect 55244 18450 55300 18452
rect 55244 18398 55246 18450
rect 55246 18398 55298 18450
rect 55298 18398 55300 18450
rect 55244 18396 55300 18398
rect 54460 18338 54516 18340
rect 54460 18286 54462 18338
rect 54462 18286 54514 18338
rect 54514 18286 54516 18338
rect 54460 18284 54516 18286
rect 54236 13804 54292 13860
rect 50316 13580 50372 13636
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 49532 3724 49588 3780
rect 40684 3388 40740 3444
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 31602 56252 31612 56308
rect 31668 56252 33180 56308
rect 33236 56252 33246 56308
rect 20178 56028 20188 56084
rect 20244 56028 20860 56084
rect 20916 56028 20926 56084
rect 29474 56028 29484 56084
rect 29540 56028 30604 56084
rect 30660 56028 30670 56084
rect 43250 56028 43260 56084
rect 43316 56028 49532 56084
rect 49588 56028 50428 56084
rect 50484 56028 50494 56084
rect 38322 55916 38332 55972
rect 38388 55916 47628 55972
rect 47684 55916 47694 55972
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 35746 55468 35756 55524
rect 35812 55468 36764 55524
rect 36820 55468 36830 55524
rect 40348 55468 43820 55524
rect 43876 55468 43886 55524
rect 40348 55412 40404 55468
rect 26786 55356 26796 55412
rect 26852 55356 29596 55412
rect 29652 55356 29662 55412
rect 33170 55356 33180 55412
rect 33236 55356 33740 55412
rect 33796 55356 33806 55412
rect 35970 55356 35980 55412
rect 36036 55356 37100 55412
rect 37156 55356 37660 55412
rect 37716 55356 37726 55412
rect 37884 55356 40404 55412
rect 49634 55356 49644 55412
rect 49700 55356 51660 55412
rect 51716 55356 51726 55412
rect 37884 55300 37940 55356
rect 22978 55244 22988 55300
rect 23044 55244 27580 55300
rect 27636 55244 27646 55300
rect 36978 55244 36988 55300
rect 37044 55244 37940 55300
rect 38612 55244 42140 55300
rect 42196 55244 42206 55300
rect 0 55188 800 55216
rect 0 55132 8764 55188
rect 8820 55132 8830 55188
rect 28466 55132 28476 55188
rect 28532 55132 29260 55188
rect 29316 55132 29326 55188
rect 35634 55132 35644 55188
rect 35700 55132 38332 55188
rect 38388 55132 38398 55188
rect 0 55104 800 55132
rect 38612 55076 38668 55244
rect 43922 55132 43932 55188
rect 43988 55132 46396 55188
rect 46452 55132 46462 55188
rect 34626 55020 34636 55076
rect 34692 55020 35084 55076
rect 35140 55020 35150 55076
rect 36418 55020 36428 55076
rect 36484 55020 38668 55076
rect 38770 54908 38780 54964
rect 38836 54908 39116 54964
rect 39172 54908 39182 54964
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 33618 54796 33628 54852
rect 33684 54796 34412 54852
rect 34468 54796 34478 54852
rect 23314 54684 23324 54740
rect 23380 54684 25676 54740
rect 25732 54684 25742 54740
rect 31378 54684 31388 54740
rect 31444 54684 34188 54740
rect 34244 54684 34254 54740
rect 37874 54684 37884 54740
rect 37940 54684 42476 54740
rect 42532 54684 42542 54740
rect 33282 54572 33292 54628
rect 33348 54572 38220 54628
rect 38276 54572 38668 54628
rect 40114 54572 40124 54628
rect 40180 54572 41132 54628
rect 41188 54572 41198 54628
rect 38612 54516 38668 54572
rect 14578 54460 14588 54516
rect 14644 54460 17052 54516
rect 17108 54460 17612 54516
rect 17668 54460 17678 54516
rect 17938 54460 17948 54516
rect 18004 54460 18956 54516
rect 19012 54460 19022 54516
rect 31602 54460 31612 54516
rect 31668 54460 34244 54516
rect 38612 54460 38780 54516
rect 38836 54460 38846 54516
rect 39890 54460 39900 54516
rect 39956 54460 41356 54516
rect 41412 54460 41422 54516
rect 42578 54460 42588 54516
rect 42644 54460 45052 54516
rect 45108 54460 45118 54516
rect 47730 54460 47740 54516
rect 47796 54460 49644 54516
rect 49700 54460 49710 54516
rect 34188 54404 34244 54460
rect 41356 54404 41412 54460
rect 18386 54348 18396 54404
rect 18452 54348 19852 54404
rect 19908 54348 19918 54404
rect 33506 54348 33516 54404
rect 33572 54348 33964 54404
rect 34020 54348 34030 54404
rect 34178 54348 34188 54404
rect 34244 54348 34254 54404
rect 37874 54348 37884 54404
rect 37940 54348 39564 54404
rect 39620 54348 40908 54404
rect 40964 54348 40974 54404
rect 41356 54348 42924 54404
rect 42980 54348 42990 54404
rect 46386 54348 46396 54404
rect 46452 54348 48188 54404
rect 48244 54348 48254 54404
rect 51538 54348 51548 54404
rect 51604 54348 52332 54404
rect 52388 54348 52398 54404
rect 29810 54236 29820 54292
rect 29876 54236 33292 54292
rect 33348 54236 33358 54292
rect 37762 54236 37772 54292
rect 37828 54236 38668 54292
rect 38724 54236 38734 54292
rect 37986 54124 37996 54180
rect 38052 54124 38444 54180
rect 38500 54124 42252 54180
rect 42308 54124 42318 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 37650 54012 37660 54068
rect 37716 54012 38556 54068
rect 38612 54012 38622 54068
rect 42914 54012 42924 54068
rect 42980 54012 43820 54068
rect 43876 54012 46508 54068
rect 46564 54012 46574 54068
rect 15586 53788 15596 53844
rect 15652 53788 17388 53844
rect 17444 53788 17454 53844
rect 18946 53788 18956 53844
rect 19012 53788 20748 53844
rect 20804 53788 20814 53844
rect 33170 53788 33180 53844
rect 33236 53788 34188 53844
rect 34244 53788 34254 53844
rect 36306 53788 36316 53844
rect 36372 53788 37660 53844
rect 37716 53788 37726 53844
rect 38546 53788 38556 53844
rect 38612 53788 39900 53844
rect 39956 53788 39966 53844
rect 40114 53788 40124 53844
rect 40180 53788 41916 53844
rect 41972 53788 41982 53844
rect 42578 53788 42588 53844
rect 42644 53788 42654 53844
rect 44828 53788 45500 53844
rect 45556 53788 45566 53844
rect 45714 53788 45724 53844
rect 45780 53788 47292 53844
rect 47348 53788 47358 53844
rect 42588 53732 42644 53788
rect 44828 53732 44884 53788
rect 17602 53676 17612 53732
rect 17668 53676 18396 53732
rect 18452 53676 18844 53732
rect 18900 53676 19740 53732
rect 19796 53676 19806 53732
rect 19954 53676 19964 53732
rect 20020 53676 20300 53732
rect 20356 53676 21980 53732
rect 22036 53676 22046 53732
rect 22642 53676 22652 53732
rect 22708 53676 24164 53732
rect 27010 53676 27020 53732
rect 27076 53676 28364 53732
rect 28420 53676 29372 53732
rect 29428 53676 30492 53732
rect 30548 53676 30558 53732
rect 33618 53676 33628 53732
rect 33684 53676 36988 53732
rect 37044 53676 37054 53732
rect 39106 53676 39116 53732
rect 39172 53676 41468 53732
rect 41524 53676 42644 53732
rect 43586 53676 43596 53732
rect 43652 53676 44884 53732
rect 45042 53676 45052 53732
rect 45108 53676 48412 53732
rect 48468 53676 49868 53732
rect 49924 53676 49934 53732
rect 24108 53620 24164 53676
rect 14578 53564 14588 53620
rect 14644 53564 15484 53620
rect 15540 53564 15550 53620
rect 17378 53564 17388 53620
rect 17444 53564 17836 53620
rect 17892 53564 17902 53620
rect 18162 53564 18172 53620
rect 18228 53564 18956 53620
rect 19012 53564 19022 53620
rect 19170 53564 19180 53620
rect 19236 53564 20188 53620
rect 20244 53564 22988 53620
rect 23044 53564 23054 53620
rect 24098 53564 24108 53620
rect 24164 53564 25340 53620
rect 25396 53564 27804 53620
rect 27860 53564 29148 53620
rect 29204 53564 29214 53620
rect 29474 53564 29484 53620
rect 29540 53564 35420 53620
rect 35476 53564 35486 53620
rect 38210 53564 38220 53620
rect 38276 53564 40012 53620
rect 40068 53564 40078 53620
rect 44146 53564 44156 53620
rect 44212 53564 46060 53620
rect 46116 53564 46508 53620
rect 46564 53564 46574 53620
rect 47506 53564 47516 53620
rect 47572 53564 49980 53620
rect 50036 53564 50876 53620
rect 50932 53564 50942 53620
rect 47516 53508 47572 53564
rect 16818 53452 16828 53508
rect 16884 53452 17500 53508
rect 17556 53452 17566 53508
rect 19292 53452 19964 53508
rect 20020 53452 20030 53508
rect 22082 53452 22092 53508
rect 22148 53452 23212 53508
rect 23268 53452 23278 53508
rect 25890 53452 25900 53508
rect 25956 53452 26684 53508
rect 26740 53452 27916 53508
rect 27972 53452 29708 53508
rect 29764 53452 29774 53508
rect 32274 53452 32284 53508
rect 32340 53452 34076 53508
rect 34132 53452 34142 53508
rect 42578 53452 42588 53508
rect 42644 53452 43148 53508
rect 43204 53452 45388 53508
rect 45444 53452 45454 53508
rect 45602 53452 45612 53508
rect 45668 53452 46172 53508
rect 46228 53452 47572 53508
rect 49522 53452 49532 53508
rect 49588 53452 50428 53508
rect 50484 53452 50494 53508
rect 50642 53452 50652 53508
rect 50708 53452 50988 53508
rect 51044 53452 51054 53508
rect 19292 53396 19348 53452
rect 18386 53340 18396 53396
rect 18452 53340 19292 53396
rect 19348 53340 19358 53396
rect 21634 53340 21644 53396
rect 21700 53340 22316 53396
rect 22372 53340 22382 53396
rect 26852 53340 36148 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 26852 53284 26908 53340
rect 25218 53228 25228 53284
rect 25284 53228 26908 53284
rect 28130 53228 28140 53284
rect 28196 53228 29596 53284
rect 29652 53228 29662 53284
rect 30706 53228 30716 53284
rect 30772 53228 31276 53284
rect 31332 53228 31342 53284
rect 32722 53228 32732 53284
rect 32788 53228 33516 53284
rect 33572 53228 35868 53284
rect 35924 53228 35934 53284
rect 18946 53116 18956 53172
rect 19012 53116 22204 53172
rect 22260 53116 22270 53172
rect 26898 53116 26908 53172
rect 26964 53116 28028 53172
rect 28084 53116 30156 53172
rect 30212 53116 30940 53172
rect 30996 53116 32508 53172
rect 32564 53116 33292 53172
rect 33348 53116 34636 53172
rect 34692 53116 34702 53172
rect 36092 53060 36148 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 38658 53116 38668 53172
rect 38724 53116 41020 53172
rect 41076 53116 41086 53172
rect 50082 53116 50092 53172
rect 50148 53116 50988 53172
rect 51044 53116 51054 53172
rect 17714 53004 17724 53060
rect 17780 53004 18172 53060
rect 18228 53004 22092 53060
rect 22148 53004 22158 53060
rect 22978 53004 22988 53060
rect 23044 53004 24444 53060
rect 24500 53004 25676 53060
rect 25732 53004 25742 53060
rect 30482 53004 30492 53060
rect 30548 53004 31836 53060
rect 31892 53004 31902 53060
rect 36092 53004 37324 53060
rect 37380 53004 40236 53060
rect 40292 53004 40302 53060
rect 42018 53004 42028 53060
rect 42084 53004 43708 53060
rect 43764 53004 44044 53060
rect 44100 53004 44110 53060
rect 31490 52892 31500 52948
rect 31556 52892 34412 52948
rect 34468 52892 34478 52948
rect 34850 52892 34860 52948
rect 34916 52892 35980 52948
rect 36036 52892 36046 52948
rect 49746 52892 49756 52948
rect 49812 52892 50540 52948
rect 50596 52892 50876 52948
rect 50932 52892 50942 52948
rect 51314 52892 51324 52948
rect 51380 52892 52444 52948
rect 52500 52892 52510 52948
rect 50876 52836 50932 52892
rect 16930 52780 16940 52836
rect 16996 52780 18172 52836
rect 18228 52780 18620 52836
rect 18676 52780 21644 52836
rect 21700 52780 21710 52836
rect 29586 52780 29596 52836
rect 29652 52780 37996 52836
rect 38052 52780 38062 52836
rect 47170 52780 47180 52836
rect 47236 52780 48188 52836
rect 48244 52780 48748 52836
rect 48804 52780 48814 52836
rect 50876 52780 51660 52836
rect 51716 52780 51726 52836
rect 24658 52668 24668 52724
rect 24724 52668 25452 52724
rect 25508 52668 26572 52724
rect 26628 52668 29260 52724
rect 29316 52668 29326 52724
rect 20402 52556 20412 52612
rect 20468 52556 24220 52612
rect 24276 52556 25116 52612
rect 25172 52556 26348 52612
rect 26404 52556 29484 52612
rect 29540 52556 29550 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 21858 52444 21868 52500
rect 21924 52444 28812 52500
rect 28868 52444 29372 52500
rect 29428 52444 29438 52500
rect 17714 52332 17724 52388
rect 17780 52332 17790 52388
rect 18050 52332 18060 52388
rect 18116 52332 24220 52388
rect 24276 52332 25228 52388
rect 25284 52332 25294 52388
rect 25778 52332 25788 52388
rect 25844 52332 26796 52388
rect 26852 52332 26862 52388
rect 30258 52332 30268 52388
rect 30324 52332 31388 52388
rect 31444 52332 31454 52388
rect 17724 52276 17780 52332
rect 17724 52220 18228 52276
rect 20626 52220 20636 52276
rect 20692 52220 21420 52276
rect 21476 52220 21486 52276
rect 24658 52220 24668 52276
rect 24724 52220 25340 52276
rect 25396 52220 25406 52276
rect 29698 52220 29708 52276
rect 29764 52220 30492 52276
rect 30548 52220 30558 52276
rect 40226 52220 40236 52276
rect 40292 52220 46620 52276
rect 46676 52220 47180 52276
rect 47236 52220 47246 52276
rect 18172 52164 18228 52220
rect 16268 52108 17388 52164
rect 17444 52108 17454 52164
rect 17826 52108 17836 52164
rect 17892 52108 17902 52164
rect 18162 52108 18172 52164
rect 18228 52108 18238 52164
rect 19170 52108 19180 52164
rect 19236 52108 19740 52164
rect 19796 52108 20412 52164
rect 20468 52108 20478 52164
rect 20738 52108 20748 52164
rect 20804 52108 21980 52164
rect 22036 52108 22046 52164
rect 22418 52108 22428 52164
rect 22484 52108 23548 52164
rect 23604 52108 25452 52164
rect 25508 52108 25518 52164
rect 26226 52108 26236 52164
rect 26292 52108 27020 52164
rect 27076 52108 27086 52164
rect 50306 52108 50316 52164
rect 50372 52108 50652 52164
rect 50708 52108 51324 52164
rect 51380 52108 51390 52164
rect 53554 52108 53564 52164
rect 53620 52108 54572 52164
rect 54628 52108 54638 52164
rect 16268 52052 16324 52108
rect 17836 52052 17892 52108
rect 16258 51996 16268 52052
rect 16324 51996 16334 52052
rect 16482 51996 16492 52052
rect 16548 51996 18788 52052
rect 25666 51996 25676 52052
rect 25732 51996 26908 52052
rect 26964 51996 26974 52052
rect 30034 51996 30044 52052
rect 30100 51996 31724 52052
rect 31780 51996 33068 52052
rect 33124 51996 33134 52052
rect 34402 51996 34412 52052
rect 34468 51996 39228 52052
rect 39284 51996 39452 52052
rect 39508 51996 39518 52052
rect 46050 51996 46060 52052
rect 46116 51996 46956 52052
rect 47012 51996 47022 52052
rect 49298 51996 49308 52052
rect 49364 51996 49756 52052
rect 49812 51996 49822 52052
rect 50204 51996 50764 52052
rect 50820 51996 50830 52052
rect 18732 51828 18788 51996
rect 50204 51828 50260 51996
rect 18722 51772 18732 51828
rect 18788 51772 18798 51828
rect 37202 51772 37212 51828
rect 37268 51772 44156 51828
rect 44212 51772 49420 51828
rect 49476 51772 49980 51828
rect 50036 51772 50046 51828
rect 50194 51772 50204 51828
rect 50260 51772 50270 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 17042 51660 17052 51716
rect 17108 51660 17948 51716
rect 18004 51660 19516 51716
rect 19572 51660 19582 51716
rect 49980 51604 50036 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 17602 51548 17612 51604
rect 17668 51548 23324 51604
rect 23380 51548 23390 51604
rect 29138 51548 29148 51604
rect 29204 51548 29708 51604
rect 29764 51548 29774 51604
rect 33954 51548 33964 51604
rect 34020 51548 34636 51604
rect 34692 51548 34702 51604
rect 49980 51548 50988 51604
rect 51044 51548 51054 51604
rect 23650 51436 23660 51492
rect 23716 51436 28364 51492
rect 28420 51436 28430 51492
rect 28588 51436 34972 51492
rect 35028 51436 36988 51492
rect 37044 51436 37054 51492
rect 46050 51436 46060 51492
rect 46116 51436 47852 51492
rect 47908 51436 47918 51492
rect 52434 51436 52444 51492
rect 52500 51436 54684 51492
rect 54740 51436 55580 51492
rect 55636 51436 55646 51492
rect 28588 51268 28644 51436
rect 34514 51324 34524 51380
rect 34580 51324 35980 51380
rect 36036 51324 36046 51380
rect 38770 51324 38780 51380
rect 38836 51324 41356 51380
rect 41412 51324 41422 51380
rect 42578 51324 42588 51380
rect 42644 51324 43820 51380
rect 43876 51324 43886 51380
rect 45378 51324 45388 51380
rect 45444 51324 46620 51380
rect 46676 51324 48748 51380
rect 48804 51324 53116 51380
rect 53172 51324 53900 51380
rect 53956 51324 53966 51380
rect 14578 51212 14588 51268
rect 14644 51212 16156 51268
rect 16212 51212 16222 51268
rect 19394 51212 19404 51268
rect 19460 51212 22988 51268
rect 23044 51212 23436 51268
rect 23492 51212 23502 51268
rect 26786 51212 26796 51268
rect 26852 51212 28588 51268
rect 28644 51212 28654 51268
rect 34738 51212 34748 51268
rect 34804 51212 37212 51268
rect 37268 51212 37278 51268
rect 39554 51212 39564 51268
rect 39620 51212 41132 51268
rect 41188 51212 41198 51268
rect 49186 51212 49196 51268
rect 49252 51212 50204 51268
rect 50260 51212 50270 51268
rect 38994 51100 39004 51156
rect 39060 51100 40796 51156
rect 40852 51100 40862 51156
rect 51986 51100 51996 51156
rect 52052 51100 52668 51156
rect 52724 51100 52734 51156
rect 50866 50988 50876 51044
rect 50932 50988 51436 51044
rect 51492 50988 52556 51044
rect 52612 50988 52622 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 14690 50764 14700 50820
rect 14756 50764 17052 50820
rect 17108 50764 17118 50820
rect 38882 50764 38892 50820
rect 38948 50764 40908 50820
rect 40964 50764 40974 50820
rect 13682 50652 13692 50708
rect 13748 50652 15820 50708
rect 15876 50652 15886 50708
rect 27570 50652 27580 50708
rect 27636 50652 37100 50708
rect 37156 50652 37166 50708
rect 37538 50652 37548 50708
rect 37604 50652 38332 50708
rect 38388 50652 40852 50708
rect 50082 50652 50092 50708
rect 50148 50652 51996 50708
rect 52052 50652 52062 50708
rect 53452 50652 53564 50708
rect 53620 50652 53630 50708
rect 40796 50596 40852 50652
rect 53452 50596 53508 50652
rect 15698 50540 15708 50596
rect 15764 50540 16380 50596
rect 16436 50540 16446 50596
rect 19058 50540 19068 50596
rect 19124 50540 20188 50596
rect 20244 50540 20254 50596
rect 23762 50540 23772 50596
rect 23828 50540 24556 50596
rect 24612 50540 24622 50596
rect 28354 50540 28364 50596
rect 28420 50540 30716 50596
rect 30772 50540 30782 50596
rect 35970 50540 35980 50596
rect 36036 50540 36540 50596
rect 36596 50540 39116 50596
rect 39172 50540 39182 50596
rect 40786 50540 40796 50596
rect 40852 50540 41916 50596
rect 41972 50540 49308 50596
rect 49364 50540 50876 50596
rect 50932 50540 50942 50596
rect 51202 50540 51212 50596
rect 51268 50540 51884 50596
rect 51940 50540 53508 50596
rect 12898 50428 12908 50484
rect 12964 50428 13580 50484
rect 13636 50428 13646 50484
rect 21756 50428 22092 50484
rect 22148 50428 22158 50484
rect 28466 50428 28476 50484
rect 28532 50428 29932 50484
rect 29988 50428 29998 50484
rect 33618 50428 33628 50484
rect 33684 50428 34076 50484
rect 34132 50428 35308 50484
rect 35364 50428 35374 50484
rect 38210 50428 38220 50484
rect 38276 50428 41244 50484
rect 41300 50428 41310 50484
rect 43362 50428 43372 50484
rect 43428 50428 44940 50484
rect 44996 50428 45006 50484
rect 50306 50428 50316 50484
rect 50372 50428 51996 50484
rect 52052 50428 52062 50484
rect 19730 50316 19740 50372
rect 19796 50316 20636 50372
rect 20692 50316 20702 50372
rect 21756 50260 21812 50428
rect 32162 50316 32172 50372
rect 32228 50316 32732 50372
rect 32788 50316 32798 50372
rect 41458 50316 41468 50372
rect 41524 50316 45052 50372
rect 45108 50316 45118 50372
rect 21746 50204 21756 50260
rect 21812 50204 21822 50260
rect 25442 50204 25452 50260
rect 25508 50204 27244 50260
rect 27300 50204 34300 50260
rect 34356 50204 34366 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 26786 50092 26796 50148
rect 26852 50092 27356 50148
rect 27412 50092 27422 50148
rect 30482 50092 30492 50148
rect 30548 50092 30940 50148
rect 30996 50092 34748 50148
rect 34804 50092 44716 50148
rect 44772 50092 44782 50148
rect 16482 49980 16492 50036
rect 16548 49980 17836 50036
rect 17892 49980 18396 50036
rect 18452 49980 18462 50036
rect 20626 49980 20636 50036
rect 20692 49980 21756 50036
rect 21812 49980 21822 50036
rect 29250 49980 29260 50036
rect 29316 49980 30044 50036
rect 30100 49980 30110 50036
rect 34290 49980 34300 50036
rect 34356 49980 35980 50036
rect 36036 49980 36046 50036
rect 36306 49980 36316 50036
rect 36372 49980 37212 50036
rect 37268 49980 37278 50036
rect 44594 49980 44604 50036
rect 44660 49980 45276 50036
rect 45332 49980 45342 50036
rect 48066 49980 48076 50036
rect 48132 49980 48860 50036
rect 48916 49980 48926 50036
rect 54114 49980 54124 50036
rect 54180 49980 54796 50036
rect 54852 49980 54862 50036
rect 2034 49868 2044 49924
rect 2100 49868 3948 49924
rect 4004 49868 4014 49924
rect 10098 49868 10108 49924
rect 10164 49868 12236 49924
rect 12292 49868 13468 49924
rect 13524 49868 14028 49924
rect 14084 49868 14094 49924
rect 15708 49868 24668 49924
rect 24724 49868 26572 49924
rect 26628 49868 27580 49924
rect 27636 49868 27646 49924
rect 29474 49868 29484 49924
rect 29540 49868 32508 49924
rect 32564 49868 32574 49924
rect 49074 49868 49084 49924
rect 49140 49868 49756 49924
rect 49812 49868 49822 49924
rect 52882 49868 52892 49924
rect 52948 49868 53900 49924
rect 53956 49868 53966 49924
rect 0 49812 800 49840
rect 15708 49812 15764 49868
rect 0 49756 1932 49812
rect 1988 49756 1998 49812
rect 13346 49756 13356 49812
rect 13412 49756 15708 49812
rect 15764 49756 15774 49812
rect 15922 49756 15932 49812
rect 15988 49756 17500 49812
rect 17556 49756 17566 49812
rect 18498 49756 18508 49812
rect 18564 49756 19516 49812
rect 19572 49756 21308 49812
rect 21364 49756 21374 49812
rect 25442 49756 25452 49812
rect 25508 49756 26124 49812
rect 26180 49756 26190 49812
rect 28802 49756 28812 49812
rect 28868 49756 30156 49812
rect 30212 49756 30222 49812
rect 31490 49756 31500 49812
rect 31556 49756 32172 49812
rect 32228 49756 32238 49812
rect 36082 49756 36092 49812
rect 36148 49756 37548 49812
rect 37604 49756 37614 49812
rect 41682 49756 41692 49812
rect 41748 49756 44940 49812
rect 44996 49756 45388 49812
rect 45444 49756 47068 49812
rect 47124 49756 47134 49812
rect 0 49728 800 49756
rect 17052 49700 17108 49756
rect 18508 49700 18564 49756
rect 1698 49644 1708 49700
rect 1764 49644 2492 49700
rect 2548 49644 2558 49700
rect 17042 49644 17052 49700
rect 17108 49644 17118 49700
rect 17378 49644 17388 49700
rect 17444 49644 18564 49700
rect 19618 49644 19628 49700
rect 19684 49644 20412 49700
rect 20468 49644 20478 49700
rect 25218 49644 25228 49700
rect 25284 49644 27468 49700
rect 27524 49644 27534 49700
rect 36194 49644 36204 49700
rect 36260 49644 36988 49700
rect 37044 49644 37054 49700
rect 40338 49644 40348 49700
rect 40404 49644 41020 49700
rect 41076 49644 41086 49700
rect 15026 49532 15036 49588
rect 15092 49532 15820 49588
rect 15876 49532 17276 49588
rect 17332 49532 17724 49588
rect 17780 49532 17790 49588
rect 38322 49532 38332 49588
rect 38388 49532 43260 49588
rect 43316 49532 43326 49588
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 0 49140 800 49168
rect 0 49084 1708 49140
rect 1764 49084 1774 49140
rect 25778 49084 25788 49140
rect 25844 49084 27020 49140
rect 27076 49084 27086 49140
rect 28578 49084 28588 49140
rect 28644 49084 33964 49140
rect 34020 49084 34030 49140
rect 39890 49084 39900 49140
rect 39956 49084 50764 49140
rect 50820 49084 50830 49140
rect 0 49056 800 49084
rect 15138 48972 15148 49028
rect 15204 48972 15820 49028
rect 15876 48972 38108 49028
rect 38164 48972 38174 49028
rect 49186 48972 49196 49028
rect 49252 48972 50204 49028
rect 50260 48972 50270 49028
rect 12226 48860 12236 48916
rect 12292 48860 13356 48916
rect 13412 48860 13422 48916
rect 15026 48860 15036 48916
rect 15092 48860 16156 48916
rect 16212 48860 16222 48916
rect 20066 48860 20076 48916
rect 20132 48860 22204 48916
rect 22260 48860 22540 48916
rect 22596 48860 22606 48916
rect 28914 48860 28924 48916
rect 28980 48860 29932 48916
rect 29988 48860 29998 48916
rect 33058 48860 33068 48916
rect 33124 48860 33404 48916
rect 33460 48860 33470 48916
rect 42018 48860 42028 48916
rect 42084 48860 42924 48916
rect 42980 48860 42990 48916
rect 43586 48860 43596 48916
rect 43652 48860 44492 48916
rect 44548 48860 44558 48916
rect 50866 48860 50876 48916
rect 50932 48860 51884 48916
rect 51940 48860 52668 48916
rect 52724 48860 54124 48916
rect 54180 48860 54190 48916
rect 13458 48748 13468 48804
rect 13524 48748 15148 48804
rect 15204 48748 15214 48804
rect 16706 48748 16716 48804
rect 16772 48748 17164 48804
rect 17220 48748 17230 48804
rect 23538 48748 23548 48804
rect 23604 48748 24332 48804
rect 24388 48748 24398 48804
rect 30034 48748 30044 48804
rect 30100 48748 31388 48804
rect 31444 48748 31836 48804
rect 31892 48748 31902 48804
rect 35084 48748 36316 48804
rect 36372 48748 37436 48804
rect 37492 48748 38444 48804
rect 38500 48748 38510 48804
rect 41794 48748 41804 48804
rect 41860 48748 42476 48804
rect 42532 48748 42542 48804
rect 43026 48748 43036 48804
rect 43092 48748 45164 48804
rect 45220 48748 46396 48804
rect 46452 48748 46462 48804
rect 53330 48748 53340 48804
rect 53396 48748 55468 48804
rect 55524 48748 55534 48804
rect 31836 48692 31892 48748
rect 35084 48692 35140 48748
rect 31836 48636 33180 48692
rect 33236 48636 33740 48692
rect 33796 48636 35084 48692
rect 35140 48636 35150 48692
rect 36754 48636 36764 48692
rect 36820 48636 37996 48692
rect 38052 48636 38062 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 36082 48524 36092 48580
rect 36148 48524 39004 48580
rect 39060 48524 39070 48580
rect 0 48468 800 48496
rect 0 48412 1708 48468
rect 1764 48412 2492 48468
rect 2548 48412 2558 48468
rect 25442 48412 25452 48468
rect 25508 48412 26796 48468
rect 26852 48412 26862 48468
rect 42130 48412 42140 48468
rect 42196 48412 42812 48468
rect 42868 48412 42878 48468
rect 50418 48412 50428 48468
rect 50484 48412 51324 48468
rect 51380 48412 51390 48468
rect 0 48384 800 48412
rect 2034 48300 2044 48356
rect 2100 48300 5964 48356
rect 6020 48300 6030 48356
rect 16482 48300 16492 48356
rect 16548 48300 17836 48356
rect 17892 48300 18060 48356
rect 18116 48300 30940 48356
rect 30996 48300 31006 48356
rect 36866 48300 36876 48356
rect 36932 48300 37660 48356
rect 37716 48300 37726 48356
rect 12002 48188 12012 48244
rect 12068 48188 12908 48244
rect 12964 48188 12974 48244
rect 19506 48188 19516 48244
rect 19572 48188 21868 48244
rect 21924 48188 24108 48244
rect 24164 48188 24174 48244
rect 25106 48188 25116 48244
rect 25172 48188 26908 48244
rect 26964 48188 26974 48244
rect 29250 48188 29260 48244
rect 29316 48188 30380 48244
rect 30436 48188 30446 48244
rect 35634 48188 35644 48244
rect 35700 48188 48748 48244
rect 48804 48188 49532 48244
rect 49588 48188 50204 48244
rect 50260 48188 50270 48244
rect 14690 48076 14700 48132
rect 14756 48076 16380 48132
rect 16436 48076 16446 48132
rect 25554 48076 25564 48132
rect 25620 48076 27580 48132
rect 27636 48076 27646 48132
rect 27794 48076 27804 48132
rect 27860 48076 29372 48132
rect 29428 48076 29438 48132
rect 36418 48076 36428 48132
rect 36484 48076 36988 48132
rect 37044 48076 37054 48132
rect 40450 48076 40460 48132
rect 40516 48076 41356 48132
rect 41412 48076 47404 48132
rect 47460 48076 48188 48132
rect 48244 48076 48254 48132
rect 49858 48076 49868 48132
rect 49924 48076 51772 48132
rect 51828 48076 53116 48132
rect 53172 48076 53182 48132
rect 48188 48020 48244 48076
rect 24882 47964 24892 48020
rect 24948 47964 26908 48020
rect 26964 47964 26974 48020
rect 34850 47964 34860 48020
rect 34916 47964 40124 48020
rect 40180 47964 40190 48020
rect 48188 47964 50428 48020
rect 50484 47964 50494 48020
rect 25330 47852 25340 47908
rect 25396 47852 26572 47908
rect 26628 47852 26638 47908
rect 0 47796 800 47824
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 0 47740 1708 47796
rect 1764 47740 2492 47796
rect 2548 47740 2558 47796
rect 12898 47740 12908 47796
rect 12964 47740 13132 47796
rect 13188 47740 24668 47796
rect 24724 47740 25564 47796
rect 25620 47740 25630 47796
rect 31938 47740 31948 47796
rect 32004 47740 32844 47796
rect 32900 47740 32910 47796
rect 36876 47740 51212 47796
rect 51268 47740 51278 47796
rect 0 47712 800 47740
rect 36876 47684 36932 47740
rect 35522 47628 35532 47684
rect 35588 47628 36876 47684
rect 36932 47628 36942 47684
rect 37426 47628 37436 47684
rect 37492 47628 38780 47684
rect 38836 47628 39900 47684
rect 39956 47628 39966 47684
rect 35746 47516 35756 47572
rect 35812 47516 40460 47572
rect 40516 47516 40526 47572
rect 51762 47516 51772 47572
rect 51828 47516 52332 47572
rect 52388 47516 52398 47572
rect 17154 47404 17164 47460
rect 17220 47404 17612 47460
rect 17668 47404 19516 47460
rect 19572 47404 19582 47460
rect 24882 47404 24892 47460
rect 24948 47404 25676 47460
rect 25732 47404 25742 47460
rect 26450 47404 26460 47460
rect 26516 47404 27020 47460
rect 27076 47404 34972 47460
rect 35028 47404 36092 47460
rect 36148 47404 36428 47460
rect 36484 47404 36494 47460
rect 37426 47404 37436 47460
rect 37492 47404 38892 47460
rect 38948 47404 38958 47460
rect 40114 47404 40124 47460
rect 40180 47404 41244 47460
rect 41300 47404 41310 47460
rect 36306 47292 36316 47348
rect 36372 47292 37772 47348
rect 37828 47292 37838 47348
rect 2034 47180 2044 47236
rect 2100 47180 3612 47236
rect 3668 47180 3678 47236
rect 26226 47180 26236 47236
rect 26292 47180 27692 47236
rect 27748 47180 27758 47236
rect 27906 47180 27916 47236
rect 27972 47180 34300 47236
rect 34356 47180 34366 47236
rect 34514 47180 34524 47236
rect 34580 47180 36092 47236
rect 36148 47180 36158 47236
rect 36754 47180 36764 47236
rect 36820 47180 37884 47236
rect 37940 47180 37950 47236
rect 40002 47180 40012 47236
rect 40068 47180 40460 47236
rect 40516 47180 40526 47236
rect 41458 47180 41468 47236
rect 41524 47180 44940 47236
rect 44996 47180 47292 47236
rect 47348 47180 49196 47236
rect 49252 47180 49644 47236
rect 49700 47180 49710 47236
rect 0 47124 800 47152
rect 0 47068 1708 47124
rect 1764 47068 2492 47124
rect 2548 47068 2558 47124
rect 27794 47068 27804 47124
rect 27860 47068 29148 47124
rect 29204 47068 29214 47124
rect 30146 47068 30156 47124
rect 30212 47068 35196 47124
rect 35252 47068 35756 47124
rect 35812 47068 35822 47124
rect 46050 47068 46060 47124
rect 46116 47068 47740 47124
rect 47796 47068 49756 47124
rect 49812 47068 49822 47124
rect 0 47040 800 47068
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 8418 46956 8428 47012
rect 8484 46956 9660 47012
rect 9716 46956 9726 47012
rect 13234 46956 13244 47012
rect 13300 46956 14028 47012
rect 14084 46956 14094 47012
rect 26338 46956 26348 47012
rect 26404 46956 31836 47012
rect 31892 46956 32172 47012
rect 32228 46956 37996 47012
rect 38052 46956 38062 47012
rect 15250 46844 15260 46900
rect 15316 46844 16044 46900
rect 16100 46844 17948 46900
rect 18004 46844 18620 46900
rect 18676 46844 18686 46900
rect 21074 46844 21084 46900
rect 21140 46844 22540 46900
rect 22596 46844 25340 46900
rect 25396 46844 25406 46900
rect 47058 46844 47068 46900
rect 47124 46844 48748 46900
rect 48804 46844 48814 46900
rect 10994 46732 11004 46788
rect 11060 46732 11788 46788
rect 11844 46732 11854 46788
rect 16706 46732 16716 46788
rect 16772 46732 30156 46788
rect 30212 46732 30222 46788
rect 30818 46732 30828 46788
rect 30884 46732 32284 46788
rect 32340 46732 34076 46788
rect 34132 46732 40908 46788
rect 40964 46732 40974 46788
rect 46610 46732 46620 46788
rect 46676 46732 49420 46788
rect 49476 46732 49486 46788
rect 51986 46732 51996 46788
rect 52052 46732 52668 46788
rect 52724 46732 52734 46788
rect 11666 46620 11676 46676
rect 11732 46620 12460 46676
rect 12516 46620 12526 46676
rect 16342 46620 16380 46676
rect 16436 46620 16446 46676
rect 17938 46620 17948 46676
rect 18004 46620 20188 46676
rect 20244 46620 20254 46676
rect 20514 46620 20524 46676
rect 20580 46620 22092 46676
rect 22148 46620 22158 46676
rect 27570 46620 27580 46676
rect 27636 46620 29148 46676
rect 29204 46620 30940 46676
rect 30996 46620 31006 46676
rect 36642 46620 36652 46676
rect 36708 46620 37884 46676
rect 37940 46620 37950 46676
rect 40450 46620 40460 46676
rect 40516 46620 41132 46676
rect 41188 46620 41198 46676
rect 20188 46564 20244 46620
rect 9874 46508 9884 46564
rect 9940 46508 11788 46564
rect 11844 46508 11854 46564
rect 20188 46508 20636 46564
rect 20692 46508 20702 46564
rect 36194 46508 36204 46564
rect 36260 46508 37100 46564
rect 37156 46508 37166 46564
rect 38322 46508 38332 46564
rect 38388 46508 39004 46564
rect 39060 46508 40012 46564
rect 40068 46508 40078 46564
rect 50530 46508 50540 46564
rect 50596 46508 50988 46564
rect 51044 46508 51054 46564
rect 0 46452 800 46480
rect 0 46396 1708 46452
rect 1764 46396 2940 46452
rect 2996 46396 3006 46452
rect 32834 46396 32844 46452
rect 32900 46396 33964 46452
rect 34020 46396 37324 46452
rect 37380 46396 37390 46452
rect 41906 46396 41916 46452
rect 41972 46396 43708 46452
rect 43764 46396 43774 46452
rect 0 46368 800 46396
rect 41010 46284 41020 46340
rect 41076 46284 42140 46340
rect 42196 46284 42206 46340
rect 44370 46284 44380 46340
rect 44436 46284 45052 46340
rect 45108 46284 45118 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 45826 46172 45836 46228
rect 45892 46172 55244 46228
rect 55300 46172 55310 46228
rect 13122 46060 13132 46116
rect 13188 46060 13580 46116
rect 13636 46060 13646 46116
rect 17938 46060 17948 46116
rect 18004 46060 18284 46116
rect 18340 46060 18350 46116
rect 19618 46060 19628 46116
rect 19684 46060 20804 46116
rect 31714 46060 31724 46116
rect 31780 46060 32060 46116
rect 32116 46060 36484 46116
rect 37986 46060 37996 46116
rect 38052 46060 38668 46116
rect 38724 46060 40460 46116
rect 40516 46060 42140 46116
rect 42196 46060 42206 46116
rect 46834 46060 46844 46116
rect 46900 46060 48300 46116
rect 48356 46060 48972 46116
rect 49028 46060 49038 46116
rect 20748 46004 20804 46060
rect 11218 45948 11228 46004
rect 11284 45948 11294 46004
rect 14690 45948 14700 46004
rect 14756 45948 15148 46004
rect 15204 45948 15214 46004
rect 19842 45948 19852 46004
rect 19908 45948 20524 46004
rect 20580 45948 20590 46004
rect 20738 45948 20748 46004
rect 20804 45948 23604 46004
rect 23874 45948 23884 46004
rect 23940 45948 26460 46004
rect 26516 45948 26526 46004
rect 33954 45948 33964 46004
rect 34020 45948 36204 46004
rect 36260 45948 36270 46004
rect 0 45780 800 45808
rect 11228 45780 11284 45948
rect 15698 45836 15708 45892
rect 15764 45836 17612 45892
rect 17668 45836 17678 45892
rect 20402 45836 20412 45892
rect 20468 45836 21868 45892
rect 21924 45836 21934 45892
rect 23548 45780 23604 45948
rect 36428 45892 36484 46060
rect 40226 45948 40236 46004
rect 40292 45948 40796 46004
rect 40852 45948 40862 46004
rect 50418 45948 50428 46004
rect 50484 45948 50988 46004
rect 51044 45948 51054 46004
rect 33394 45836 33404 45892
rect 33460 45836 35868 45892
rect 35924 45836 35934 45892
rect 36428 45836 39956 45892
rect 40114 45836 40124 45892
rect 40180 45836 41580 45892
rect 41636 45836 42364 45892
rect 42420 45836 42430 45892
rect 43698 45836 43708 45892
rect 43764 45836 45164 45892
rect 45220 45836 45230 45892
rect 46162 45836 46172 45892
rect 46228 45836 47292 45892
rect 47348 45836 47358 45892
rect 49634 45836 49644 45892
rect 49700 45836 52668 45892
rect 52724 45836 52734 45892
rect 0 45724 2380 45780
rect 2436 45724 3164 45780
rect 3220 45724 3230 45780
rect 11228 45724 11788 45780
rect 11844 45724 12572 45780
rect 12628 45724 13916 45780
rect 13972 45724 13982 45780
rect 22754 45724 22764 45780
rect 22820 45724 22830 45780
rect 23548 45724 24332 45780
rect 24388 45724 35532 45780
rect 35588 45724 35598 45780
rect 0 45696 800 45724
rect 22764 45668 22820 45724
rect 39900 45668 39956 45836
rect 45378 45724 45388 45780
rect 45444 45724 47964 45780
rect 48020 45724 48030 45780
rect 10780 45612 12236 45668
rect 12292 45612 14476 45668
rect 14532 45612 14542 45668
rect 16818 45612 16828 45668
rect 16884 45612 19964 45668
rect 20020 45612 20300 45668
rect 20356 45612 21868 45668
rect 21924 45612 21934 45668
rect 22764 45612 28028 45668
rect 28084 45612 28094 45668
rect 28802 45612 28812 45668
rect 28868 45612 29260 45668
rect 29316 45612 29326 45668
rect 32284 45612 34860 45668
rect 34916 45612 34926 45668
rect 39890 45612 39900 45668
rect 39956 45612 43372 45668
rect 43428 45612 43438 45668
rect 45826 45612 45836 45668
rect 45892 45612 51996 45668
rect 52052 45612 53004 45668
rect 53060 45612 53070 45668
rect 10780 45556 10836 45612
rect 32284 45556 32340 45612
rect 10770 45500 10780 45556
rect 10836 45500 10846 45556
rect 11666 45500 11676 45556
rect 11732 45500 13692 45556
rect 13748 45500 14252 45556
rect 14308 45500 14318 45556
rect 21410 45500 21420 45556
rect 21476 45500 23044 45556
rect 23762 45500 23772 45556
rect 23828 45500 25340 45556
rect 25396 45500 25406 45556
rect 26852 45500 32340 45556
rect 33394 45500 33404 45556
rect 33460 45500 33470 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 22988 45444 23044 45500
rect 26852 45444 26908 45500
rect 33404 45444 33460 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 12226 45388 12236 45444
rect 12292 45388 13244 45444
rect 13300 45388 13310 45444
rect 21634 45388 21644 45444
rect 21700 45388 22764 45444
rect 22820 45388 22830 45444
rect 22988 45388 26908 45444
rect 30156 45388 33460 45444
rect 51650 45388 51660 45444
rect 51716 45388 52220 45444
rect 52276 45388 52286 45444
rect 30156 45332 30212 45388
rect 12114 45276 12124 45332
rect 12180 45276 14140 45332
rect 14196 45276 22092 45332
rect 22148 45276 23660 45332
rect 23716 45276 25340 45332
rect 25396 45276 30212 45332
rect 31378 45276 31388 45332
rect 31444 45276 32284 45332
rect 32340 45276 33404 45332
rect 33460 45276 33470 45332
rect 33842 45276 33852 45332
rect 33908 45276 34748 45332
rect 34804 45276 34814 45332
rect 50754 45276 50764 45332
rect 50820 45276 54684 45332
rect 54740 45276 54750 45332
rect 2034 45164 2044 45220
rect 2100 45164 6748 45220
rect 6804 45164 6814 45220
rect 11218 45164 11228 45220
rect 11284 45164 15372 45220
rect 15428 45164 15438 45220
rect 23212 45164 25228 45220
rect 25284 45164 27132 45220
rect 27188 45164 27198 45220
rect 31938 45164 31948 45220
rect 32004 45164 32508 45220
rect 32564 45164 34412 45220
rect 34468 45164 34478 45220
rect 43474 45164 43484 45220
rect 43540 45164 43932 45220
rect 43988 45164 45164 45220
rect 45220 45164 45230 45220
rect 0 45108 800 45136
rect 23212 45108 23268 45164
rect 0 45052 1820 45108
rect 1876 45052 1886 45108
rect 14690 45052 14700 45108
rect 14756 45052 15260 45108
rect 15316 45052 15326 45108
rect 17490 45052 17500 45108
rect 17556 45052 20748 45108
rect 20804 45052 23212 45108
rect 23268 45052 23278 45108
rect 26226 45052 26236 45108
rect 26292 45052 27020 45108
rect 27076 45052 27086 45108
rect 29474 45052 29484 45108
rect 29540 45052 30380 45108
rect 30436 45052 30446 45108
rect 31714 45052 31724 45108
rect 31780 45052 33180 45108
rect 33236 45052 33246 45108
rect 34514 45052 34524 45108
rect 34580 45052 35084 45108
rect 35140 45052 35150 45108
rect 42130 45052 42140 45108
rect 42196 45052 42812 45108
rect 42868 45052 42878 45108
rect 43138 45052 43148 45108
rect 43204 45052 43708 45108
rect 43764 45052 43774 45108
rect 0 45024 800 45052
rect 1698 44940 1708 44996
rect 1764 44940 2492 44996
rect 2548 44940 2558 44996
rect 9762 44940 9772 44996
rect 9828 44940 10892 44996
rect 10948 44940 10958 44996
rect 23538 44940 23548 44996
rect 23604 44940 23884 44996
rect 23940 44940 23950 44996
rect 31490 44940 31500 44996
rect 31556 44940 33628 44996
rect 33684 44940 33694 44996
rect 33842 44940 33852 44996
rect 33908 44940 34748 44996
rect 34804 44940 34814 44996
rect 43250 44940 43260 44996
rect 43316 44940 43820 44996
rect 43876 44940 43886 44996
rect 46274 44940 46284 44996
rect 46340 44940 47068 44996
rect 47124 44940 47134 44996
rect 51202 44940 51212 44996
rect 51268 44940 52108 44996
rect 52164 44940 52174 44996
rect 15092 44828 21756 44884
rect 21812 44828 26460 44884
rect 26516 44828 26526 44884
rect 45154 44828 45164 44884
rect 45220 44828 46508 44884
rect 46564 44828 47852 44884
rect 47908 44828 47918 44884
rect 15092 44772 15148 44828
rect 13906 44716 13916 44772
rect 13972 44716 15148 44772
rect 15474 44716 15484 44772
rect 15540 44716 17276 44772
rect 17332 44716 17342 44772
rect 29922 44716 29932 44772
rect 29988 44716 33292 44772
rect 33348 44716 34132 44772
rect 35746 44716 35756 44772
rect 35812 44716 45388 44772
rect 45444 44716 45454 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 34076 44660 34132 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 10098 44604 10108 44660
rect 10164 44604 14924 44660
rect 14980 44604 15820 44660
rect 15876 44604 15886 44660
rect 24966 44604 25004 44660
rect 25060 44604 25070 44660
rect 34066 44604 34076 44660
rect 34132 44604 34412 44660
rect 34468 44604 34478 44660
rect 38668 44604 38892 44660
rect 38948 44604 38958 44660
rect 38668 44548 38724 44604
rect 2146 44492 2156 44548
rect 2212 44492 5292 44548
rect 5348 44492 5358 44548
rect 15138 44492 15148 44548
rect 15204 44492 15484 44548
rect 15540 44492 15550 44548
rect 25554 44492 25564 44548
rect 25620 44492 25900 44548
rect 25956 44492 25966 44548
rect 26114 44492 26124 44548
rect 26180 44492 26796 44548
rect 26852 44492 38108 44548
rect 38164 44492 38174 44548
rect 38658 44492 38668 44548
rect 38724 44492 38734 44548
rect 51090 44492 51100 44548
rect 51156 44492 52556 44548
rect 52612 44492 52622 44548
rect 0 44436 800 44464
rect 59200 44436 60000 44464
rect 0 44380 1708 44436
rect 1764 44380 1774 44436
rect 24210 44380 24220 44436
rect 24276 44380 25004 44436
rect 25060 44380 31836 44436
rect 31892 44380 31902 44436
rect 43250 44380 43260 44436
rect 43316 44380 43820 44436
rect 43876 44380 43886 44436
rect 50978 44380 50988 44436
rect 51044 44380 51884 44436
rect 51940 44380 51950 44436
rect 54898 44380 54908 44436
rect 54964 44380 60000 44436
rect 0 44352 800 44380
rect 59200 44352 60000 44380
rect 13010 44268 13020 44324
rect 13076 44268 13916 44324
rect 13972 44268 13982 44324
rect 15586 44268 15596 44324
rect 15652 44268 16380 44324
rect 16436 44268 16446 44324
rect 25890 44268 25900 44324
rect 25956 44268 27132 44324
rect 27188 44268 27198 44324
rect 29138 44268 29148 44324
rect 29204 44268 32508 44324
rect 32564 44268 33964 44324
rect 34020 44268 34524 44324
rect 34580 44268 34590 44324
rect 38546 44268 38556 44324
rect 38612 44212 38668 44324
rect 42130 44268 42140 44324
rect 42196 44268 43036 44324
rect 43092 44268 43102 44324
rect 13570 44156 13580 44212
rect 13636 44156 14140 44212
rect 14196 44156 14206 44212
rect 18386 44156 18396 44212
rect 18452 44156 19404 44212
rect 19460 44156 21980 44212
rect 22036 44156 22652 44212
rect 22708 44156 22718 44212
rect 33842 44156 33852 44212
rect 33908 44156 34860 44212
rect 34916 44156 34926 44212
rect 38612 44156 39340 44212
rect 39396 44156 40236 44212
rect 40292 44156 51212 44212
rect 51268 44156 51278 44212
rect 11442 44044 11452 44100
rect 11508 44044 12012 44100
rect 12068 44044 13132 44100
rect 13188 44044 13198 44100
rect 33618 44044 33628 44100
rect 33684 44044 34748 44100
rect 34804 44044 34814 44100
rect 42802 44044 42812 44100
rect 42868 44044 43932 44100
rect 43988 44044 43998 44100
rect 50754 44044 50764 44100
rect 50820 44044 51436 44100
rect 51492 44044 51502 44100
rect 50978 43932 50988 43988
rect 51044 43932 51082 43988
rect 51650 43932 51660 43988
rect 51716 43932 51726 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 2706 43820 2716 43876
rect 2772 43820 3724 43876
rect 3780 43820 3790 43876
rect 22306 43820 22316 43876
rect 22372 43820 22382 43876
rect 28354 43820 28364 43876
rect 28420 43820 28924 43876
rect 28980 43820 28990 43876
rect 0 43764 800 43792
rect 22316 43764 22372 43820
rect 0 43708 1932 43764
rect 1988 43708 1998 43764
rect 13468 43708 15484 43764
rect 15540 43708 15550 43764
rect 19954 43708 19964 43764
rect 20020 43708 21420 43764
rect 21476 43708 21486 43764
rect 22316 43708 25284 43764
rect 27458 43708 27468 43764
rect 27524 43708 30380 43764
rect 30436 43708 30446 43764
rect 33058 43708 33068 43764
rect 33124 43708 33404 43764
rect 33460 43708 34412 43764
rect 34468 43708 34478 43764
rect 34636 43708 35308 43764
rect 35364 43708 35374 43764
rect 37762 43708 37772 43764
rect 37828 43708 38668 43764
rect 38724 43708 42140 43764
rect 42196 43708 42206 43764
rect 0 43680 800 43708
rect 13468 43652 13524 43708
rect 2034 43596 2044 43652
rect 2100 43596 6860 43652
rect 6916 43596 6926 43652
rect 12002 43596 12012 43652
rect 12068 43596 13524 43652
rect 14466 43596 14476 43652
rect 14532 43596 17500 43652
rect 17556 43596 17566 43652
rect 18946 43596 18956 43652
rect 19012 43596 19852 43652
rect 19908 43596 20524 43652
rect 20580 43596 20972 43652
rect 21028 43596 21038 43652
rect 24546 43596 24556 43652
rect 24612 43596 24622 43652
rect 4274 43484 4284 43540
rect 4340 43484 8092 43540
rect 8148 43484 8158 43540
rect 8642 43484 8652 43540
rect 8708 43484 10556 43540
rect 10612 43484 12236 43540
rect 12292 43484 13916 43540
rect 13972 43484 13982 43540
rect 17500 43428 17556 43596
rect 24556 43540 24612 43596
rect 20178 43484 20188 43540
rect 20244 43484 20748 43540
rect 20804 43484 20814 43540
rect 23986 43484 23996 43540
rect 24052 43484 24612 43540
rect 25228 43540 25284 43708
rect 34636 43652 34692 43708
rect 51660 43652 51716 43932
rect 59200 43764 60000 43792
rect 57922 43708 57932 43764
rect 57988 43708 60000 43764
rect 59200 43680 60000 43708
rect 25666 43596 25676 43652
rect 25732 43596 26572 43652
rect 26628 43596 27020 43652
rect 27076 43596 27086 43652
rect 27906 43596 27916 43652
rect 27972 43596 29036 43652
rect 29092 43596 29102 43652
rect 33506 43596 33516 43652
rect 33572 43596 34188 43652
rect 34244 43596 34254 43652
rect 34412 43596 34692 43652
rect 40114 43596 40124 43652
rect 40180 43596 41020 43652
rect 41076 43596 41086 43652
rect 47842 43596 47852 43652
rect 47908 43596 48860 43652
rect 48916 43596 48926 43652
rect 49970 43596 49980 43652
rect 50036 43596 50988 43652
rect 51044 43596 51716 43652
rect 53106 43596 53116 43652
rect 53172 43596 54460 43652
rect 54516 43596 54526 43652
rect 34412 43540 34468 43596
rect 25228 43484 29596 43540
rect 29652 43484 29662 43540
rect 34402 43484 34412 43540
rect 34468 43484 34478 43540
rect 36306 43484 36316 43540
rect 36372 43484 37660 43540
rect 37716 43484 37726 43540
rect 46050 43484 46060 43540
rect 46116 43484 47628 43540
rect 47684 43484 47694 43540
rect 50372 43484 51772 43540
rect 51828 43484 51838 43540
rect 3826 43372 3836 43428
rect 3892 43372 5740 43428
rect 5796 43372 8204 43428
rect 8260 43372 8270 43428
rect 11330 43372 11340 43428
rect 11396 43372 13580 43428
rect 13636 43372 13646 43428
rect 17500 43372 24556 43428
rect 24612 43372 24622 43428
rect 26450 43372 26460 43428
rect 26516 43372 27132 43428
rect 27188 43372 27198 43428
rect 50372 43316 50428 43484
rect 16818 43260 16828 43316
rect 16884 43260 17836 43316
rect 17892 43260 17902 43316
rect 22502 43260 22540 43316
rect 22596 43260 22606 43316
rect 26562 43260 26572 43316
rect 26628 43260 28140 43316
rect 28196 43260 28206 43316
rect 42018 43260 42028 43316
rect 42084 43260 43820 43316
rect 43876 43260 43886 43316
rect 49858 43260 49868 43316
rect 49924 43260 50428 43316
rect 12450 43148 12460 43204
rect 12516 43148 13468 43204
rect 13524 43148 15148 43204
rect 17714 43148 17724 43204
rect 17780 43148 19068 43204
rect 19124 43148 19134 43204
rect 52994 43148 53004 43204
rect 53060 43148 54572 43204
rect 54628 43148 54638 43204
rect 0 43092 800 43120
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 0 43036 1708 43092
rect 1764 43036 2492 43092
rect 2548 43036 2558 43092
rect 0 43008 800 43036
rect 15092 42980 15148 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 59200 43092 60000 43120
rect 20066 43036 20076 43092
rect 20132 43036 23996 43092
rect 24052 43036 24062 43092
rect 51398 43036 51436 43092
rect 51492 43036 51502 43092
rect 55010 43036 55020 43092
rect 55076 43036 60000 43092
rect 59200 43008 60000 43036
rect 7858 42924 7868 42980
rect 7924 42924 11228 42980
rect 11284 42924 11294 42980
rect 12786 42924 12796 42980
rect 12852 42924 13468 42980
rect 13524 42924 13534 42980
rect 14018 42924 14028 42980
rect 14084 42924 14364 42980
rect 14420 42924 14430 42980
rect 15092 42924 18172 42980
rect 18228 42924 25788 42980
rect 25844 42924 25854 42980
rect 41570 42924 41580 42980
rect 41636 42924 45724 42980
rect 45780 42924 49756 42980
rect 49812 42924 50652 42980
rect 50708 42924 50718 42980
rect 9986 42812 9996 42868
rect 10052 42812 10444 42868
rect 10500 42812 11004 42868
rect 11060 42812 11070 42868
rect 18274 42812 18284 42868
rect 18340 42812 24332 42868
rect 24388 42812 25676 42868
rect 25732 42812 25742 42868
rect 29810 42812 29820 42868
rect 29876 42812 30268 42868
rect 30324 42812 33740 42868
rect 33796 42812 35532 42868
rect 35588 42812 38668 42868
rect 50950 42812 50988 42868
rect 51044 42812 51054 42868
rect 2146 42700 2156 42756
rect 2212 42700 5852 42756
rect 5908 42700 5918 42756
rect 11330 42700 11340 42756
rect 11396 42700 12012 42756
rect 12068 42700 12078 42756
rect 13682 42700 13692 42756
rect 13748 42700 14812 42756
rect 14868 42700 14878 42756
rect 22754 42700 22764 42756
rect 22820 42700 23100 42756
rect 23156 42700 23166 42756
rect 23426 42700 23436 42756
rect 23492 42700 23884 42756
rect 23940 42700 23950 42756
rect 24546 42700 24556 42756
rect 24612 42700 25116 42756
rect 25172 42700 27244 42756
rect 27300 42700 27310 42756
rect 34738 42700 34748 42756
rect 34804 42700 35420 42756
rect 35476 42700 35486 42756
rect 38612 42644 38668 42812
rect 42242 42700 42252 42756
rect 42308 42700 42476 42756
rect 42532 42700 42542 42756
rect 46498 42700 46508 42756
rect 46564 42700 47404 42756
rect 47460 42700 47470 42756
rect 50754 42700 50764 42756
rect 50820 42700 53116 42756
rect 53172 42700 53182 42756
rect 2034 42588 2044 42644
rect 2100 42588 4844 42644
rect 4900 42588 4910 42644
rect 7522 42588 7532 42644
rect 7588 42588 8764 42644
rect 8820 42588 8830 42644
rect 11554 42588 11564 42644
rect 11620 42588 12572 42644
rect 12628 42588 12638 42644
rect 17826 42588 17836 42644
rect 17892 42588 19404 42644
rect 19460 42588 19470 42644
rect 23762 42588 23772 42644
rect 23828 42588 25340 42644
rect 25396 42588 26572 42644
rect 26628 42588 26638 42644
rect 28242 42588 28252 42644
rect 28308 42588 28700 42644
rect 28756 42588 29260 42644
rect 29316 42588 32732 42644
rect 32788 42588 38500 42644
rect 38612 42588 42364 42644
rect 42420 42588 42430 42644
rect 38444 42532 38500 42588
rect 13682 42476 13692 42532
rect 13748 42476 14700 42532
rect 14756 42476 15148 42532
rect 15204 42476 16044 42532
rect 16100 42476 16110 42532
rect 21298 42476 21308 42532
rect 21364 42476 22316 42532
rect 22372 42476 22382 42532
rect 22978 42476 22988 42532
rect 23044 42476 24220 42532
rect 24276 42476 24780 42532
rect 24836 42476 25900 42532
rect 25956 42476 25966 42532
rect 26226 42476 26236 42532
rect 26292 42476 32788 42532
rect 34178 42476 34188 42532
rect 34244 42476 34748 42532
rect 34804 42476 34814 42532
rect 38434 42476 38444 42532
rect 38500 42476 38892 42532
rect 38948 42476 48860 42532
rect 48916 42476 49308 42532
rect 49364 42476 49374 42532
rect 0 42420 800 42448
rect 32732 42420 32788 42476
rect 59200 42420 60000 42448
rect 0 42364 1708 42420
rect 1764 42364 2492 42420
rect 2548 42364 2558 42420
rect 26562 42364 26572 42420
rect 26628 42364 29372 42420
rect 29428 42364 29438 42420
rect 32732 42364 38668 42420
rect 57698 42364 57708 42420
rect 57764 42364 60000 42420
rect 0 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 35830 42252 35868 42308
rect 35924 42252 35934 42308
rect 5842 42140 5852 42196
rect 5908 42140 7084 42196
rect 7140 42140 7150 42196
rect 26646 42140 26684 42196
rect 26740 42140 26750 42196
rect 33730 42140 33740 42196
rect 33796 42140 34524 42196
rect 34580 42140 35084 42196
rect 35140 42140 35150 42196
rect 38612 42084 38668 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 59200 42336 60000 42364
rect 50978 42252 50988 42308
rect 51044 42252 55580 42308
rect 55636 42252 55646 42308
rect 40114 42140 40124 42196
rect 40180 42140 41580 42196
rect 41636 42140 47852 42196
rect 47908 42140 47918 42196
rect 51426 42140 51436 42196
rect 51492 42140 51884 42196
rect 51940 42140 51950 42196
rect 12562 42028 12572 42084
rect 12628 42028 13580 42084
rect 13636 42028 13646 42084
rect 21410 42028 21420 42084
rect 21476 42028 26908 42084
rect 30034 42028 30044 42084
rect 30100 42028 30716 42084
rect 30772 42028 30782 42084
rect 31266 42028 31276 42084
rect 31332 42028 32844 42084
rect 32900 42028 32910 42084
rect 38612 42028 42252 42084
rect 42308 42028 42318 42084
rect 51324 42028 52668 42084
rect 52724 42028 52734 42084
rect 26852 41972 26908 42028
rect 51324 41972 51380 42028
rect 2594 41916 2604 41972
rect 2660 41916 4284 41972
rect 4340 41916 4350 41972
rect 4946 41916 4956 41972
rect 5012 41916 6300 41972
rect 6356 41916 6366 41972
rect 12338 41916 12348 41972
rect 12404 41916 13468 41972
rect 13524 41916 13534 41972
rect 13794 41916 13804 41972
rect 13860 41916 15036 41972
rect 15092 41916 15102 41972
rect 19058 41916 19068 41972
rect 19124 41916 20748 41972
rect 20804 41916 20814 41972
rect 23650 41916 23660 41972
rect 23716 41916 24108 41972
rect 24164 41916 24174 41972
rect 26852 41916 30492 41972
rect 30548 41916 30558 41972
rect 30930 41916 30940 41972
rect 30996 41916 32396 41972
rect 32452 41916 32462 41972
rect 35074 41916 35084 41972
rect 35140 41916 36428 41972
rect 36484 41916 36494 41972
rect 45042 41916 45052 41972
rect 45108 41916 47516 41972
rect 47572 41916 47964 41972
rect 48020 41916 48030 41972
rect 51314 41916 51324 41972
rect 51380 41916 51390 41972
rect 51874 41916 51884 41972
rect 51940 41916 55132 41972
rect 55188 41916 55198 41972
rect 51884 41860 51940 41916
rect 2706 41804 2716 41860
rect 2772 41804 11116 41860
rect 11172 41804 12796 41860
rect 12852 41804 12862 41860
rect 22978 41804 22988 41860
rect 23044 41804 24668 41860
rect 24724 41804 26908 41860
rect 27346 41804 27356 41860
rect 27412 41804 31388 41860
rect 31444 41804 31454 41860
rect 38210 41804 38220 41860
rect 38276 41804 38780 41860
rect 38836 41804 38846 41860
rect 41570 41804 41580 41860
rect 41636 41804 42364 41860
rect 42420 41804 42430 41860
rect 45266 41804 45276 41860
rect 45332 41804 45342 41860
rect 45490 41804 45500 41860
rect 45556 41804 46508 41860
rect 46564 41804 46574 41860
rect 46722 41804 46732 41860
rect 46788 41804 50876 41860
rect 50932 41804 51940 41860
rect 0 41748 800 41776
rect 0 41692 1708 41748
rect 1764 41692 2940 41748
rect 2996 41692 3006 41748
rect 0 41664 800 41692
rect 26852 41636 26908 41804
rect 45276 41748 45332 41804
rect 59200 41748 60000 41776
rect 29026 41692 29036 41748
rect 29092 41692 30268 41748
rect 30324 41692 30334 41748
rect 30706 41692 30716 41748
rect 30772 41692 33740 41748
rect 33796 41692 33806 41748
rect 45276 41692 49644 41748
rect 49700 41692 49710 41748
rect 55346 41692 55356 41748
rect 55412 41692 60000 41748
rect 59200 41664 60000 41692
rect 26852 41580 30100 41636
rect 38434 41580 38444 41636
rect 38500 41580 39676 41636
rect 39732 41580 45836 41636
rect 45892 41580 45902 41636
rect 47618 41580 47628 41636
rect 47684 41580 49308 41636
rect 49364 41580 49374 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 30044 41524 30100 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 19618 41468 19628 41524
rect 19684 41468 20188 41524
rect 20244 41468 26908 41524
rect 30034 41468 30044 41524
rect 30100 41468 30110 41524
rect 41682 41468 41692 41524
rect 41748 41468 45612 41524
rect 45668 41468 45678 41524
rect 26852 41412 26908 41468
rect 2034 41356 2044 41412
rect 2100 41356 8092 41412
rect 8148 41356 8158 41412
rect 24882 41356 24892 41412
rect 24948 41356 25676 41412
rect 25732 41356 25742 41412
rect 26852 41356 37436 41412
rect 37492 41356 41020 41412
rect 41076 41356 41468 41412
rect 41524 41356 41534 41412
rect 47058 41356 47068 41412
rect 47124 41356 53452 41412
rect 53508 41356 53518 41412
rect 14018 41244 14028 41300
rect 14084 41244 14924 41300
rect 14980 41244 14990 41300
rect 21410 41244 21420 41300
rect 21476 41244 22092 41300
rect 22148 41244 23996 41300
rect 24052 41244 24062 41300
rect 53666 41244 53676 41300
rect 53732 41244 56868 41300
rect 1810 41132 1820 41188
rect 1876 41132 2492 41188
rect 2548 41132 2558 41188
rect 10882 41132 10892 41188
rect 10948 41132 14252 41188
rect 14308 41132 14318 41188
rect 15026 41132 15036 41188
rect 15092 41132 15820 41188
rect 15876 41132 15886 41188
rect 22418 41132 22428 41188
rect 22484 41132 22494 41188
rect 23090 41132 23100 41188
rect 23156 41132 24332 41188
rect 24388 41132 24398 41188
rect 27906 41132 27916 41188
rect 27972 41132 28812 41188
rect 28868 41132 30716 41188
rect 30772 41132 30782 41188
rect 45826 41132 45836 41188
rect 45892 41132 47628 41188
rect 47684 41132 47694 41188
rect 48738 41132 48748 41188
rect 48804 41132 52668 41188
rect 52724 41132 52734 41188
rect 53218 41132 53228 41188
rect 53284 41132 54796 41188
rect 54852 41132 54862 41188
rect 0 41076 800 41104
rect 22428 41076 22484 41132
rect 56812 41076 56868 41244
rect 59200 41076 60000 41104
rect 0 41020 2380 41076
rect 2436 41020 3164 41076
rect 3220 41020 3230 41076
rect 13234 41020 13244 41076
rect 13300 41020 13692 41076
rect 13748 41020 13758 41076
rect 14578 41020 14588 41076
rect 14644 41020 16380 41076
rect 16436 41020 16446 41076
rect 19394 41020 19404 41076
rect 19460 41020 19852 41076
rect 19908 41020 19918 41076
rect 22428 41020 23212 41076
rect 23268 41020 23278 41076
rect 24098 41020 24108 41076
rect 24164 41020 24444 41076
rect 24500 41020 25004 41076
rect 25060 41020 27020 41076
rect 27076 41020 27086 41076
rect 32498 41020 32508 41076
rect 32564 41020 45052 41076
rect 45108 41020 45276 41076
rect 45332 41020 45342 41076
rect 47506 41020 47516 41076
rect 47572 41020 49084 41076
rect 49140 41020 49150 41076
rect 56812 41020 60000 41076
rect 0 40992 800 41020
rect 59200 40992 60000 41020
rect 9090 40908 9100 40964
rect 9156 40908 13804 40964
rect 13860 40908 13870 40964
rect 14690 40908 14700 40964
rect 14756 40908 15932 40964
rect 15988 40908 15998 40964
rect 16594 40908 16604 40964
rect 16660 40908 20244 40964
rect 22754 40908 22764 40964
rect 22820 40908 24556 40964
rect 24612 40908 24622 40964
rect 35634 40908 35644 40964
rect 35700 40908 35868 40964
rect 35924 40908 35934 40964
rect 36194 40908 36204 40964
rect 36260 40908 36988 40964
rect 37044 40908 37660 40964
rect 37716 40908 37726 40964
rect 44370 40908 44380 40964
rect 44436 40908 45612 40964
rect 45668 40908 45948 40964
rect 46004 40908 46014 40964
rect 51650 40908 51660 40964
rect 51716 40908 52108 40964
rect 52164 40908 52174 40964
rect 16604 40628 16660 40908
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 20188 40740 20244 40908
rect 21858 40796 21868 40852
rect 21924 40796 30044 40852
rect 30100 40796 30940 40852
rect 30996 40796 31612 40852
rect 31668 40796 31678 40852
rect 36642 40796 36652 40852
rect 36708 40796 37100 40852
rect 37156 40796 37166 40852
rect 41458 40796 41468 40852
rect 41524 40796 42028 40852
rect 42084 40796 42094 40852
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 19366 40684 19404 40740
rect 19460 40684 19470 40740
rect 20188 40684 22764 40740
rect 22820 40684 22830 40740
rect 25778 40684 25788 40740
rect 25844 40684 27916 40740
rect 27972 40684 27982 40740
rect 28466 40684 28476 40740
rect 28532 40684 29148 40740
rect 29204 40684 29484 40740
rect 29540 40684 29550 40740
rect 38098 40684 38108 40740
rect 38164 40684 38668 40740
rect 38724 40684 43932 40740
rect 43988 40684 46396 40740
rect 46452 40684 46462 40740
rect 12898 40572 12908 40628
rect 12964 40572 14084 40628
rect 14914 40572 14924 40628
rect 14980 40572 16660 40628
rect 21298 40572 21308 40628
rect 21364 40572 22204 40628
rect 22260 40572 24444 40628
rect 24500 40572 25228 40628
rect 25284 40572 25294 40628
rect 26646 40572 26684 40628
rect 26740 40572 26750 40628
rect 35634 40572 35644 40628
rect 35700 40572 36092 40628
rect 36148 40572 36158 40628
rect 41682 40572 41692 40628
rect 41748 40572 42252 40628
rect 42308 40572 42318 40628
rect 53106 40572 53116 40628
rect 53172 40572 56588 40628
rect 56644 40572 56654 40628
rect 14028 40516 14084 40572
rect 8306 40460 8316 40516
rect 8372 40460 10668 40516
rect 10724 40460 11452 40516
rect 11508 40460 11518 40516
rect 14018 40460 14028 40516
rect 14084 40460 16940 40516
rect 16996 40460 17006 40516
rect 18722 40460 18732 40516
rect 18788 40460 20580 40516
rect 22530 40460 22540 40516
rect 22596 40460 23436 40516
rect 23492 40460 23502 40516
rect 24770 40460 24780 40516
rect 24836 40460 25004 40516
rect 25060 40460 25070 40516
rect 41346 40460 41356 40516
rect 41412 40460 42588 40516
rect 42644 40460 43484 40516
rect 43540 40460 43550 40516
rect 44940 40460 46508 40516
rect 46564 40460 46574 40516
rect 53330 40460 53340 40516
rect 53396 40460 57148 40516
rect 57204 40460 57214 40516
rect 0 40404 800 40432
rect 0 40348 1820 40404
rect 1876 40348 1886 40404
rect 4610 40348 4620 40404
rect 4676 40348 7700 40404
rect 16370 40348 16380 40404
rect 16436 40348 18844 40404
rect 18900 40348 18910 40404
rect 0 40320 800 40348
rect 7644 40292 7700 40348
rect 1698 40236 1708 40292
rect 1764 40236 2492 40292
rect 2548 40236 2558 40292
rect 7634 40236 7644 40292
rect 7700 40236 9548 40292
rect 9604 40236 9614 40292
rect 13458 40236 13468 40292
rect 13524 40236 14252 40292
rect 14308 40236 14318 40292
rect 15474 40236 15484 40292
rect 15540 40236 16828 40292
rect 16884 40236 16894 40292
rect 20524 40180 20580 40460
rect 44940 40404 44996 40460
rect 59200 40404 60000 40432
rect 21186 40348 21196 40404
rect 21252 40348 21644 40404
rect 21700 40348 21868 40404
rect 21924 40348 21934 40404
rect 23986 40348 23996 40404
rect 24052 40348 25228 40404
rect 25284 40348 26292 40404
rect 26236 40292 26292 40348
rect 31892 40348 32508 40404
rect 32564 40348 32574 40404
rect 33180 40348 33852 40404
rect 33908 40348 33918 40404
rect 37090 40348 37100 40404
rect 37156 40348 38780 40404
rect 38836 40348 38846 40404
rect 41570 40348 41580 40404
rect 41636 40348 44940 40404
rect 44996 40348 45006 40404
rect 45266 40348 45276 40404
rect 45332 40348 48412 40404
rect 48468 40348 48860 40404
rect 48916 40348 49308 40404
rect 49364 40348 51212 40404
rect 51268 40348 51278 40404
rect 51650 40348 51660 40404
rect 51716 40348 53452 40404
rect 53508 40348 53518 40404
rect 53900 40348 55804 40404
rect 55860 40348 55870 40404
rect 57810 40348 57820 40404
rect 57876 40348 60000 40404
rect 31892 40292 31948 40348
rect 33180 40292 33236 40348
rect 53900 40292 53956 40348
rect 59200 40320 60000 40348
rect 23202 40236 23212 40292
rect 23268 40236 25340 40292
rect 25396 40236 25406 40292
rect 26226 40236 26236 40292
rect 26292 40236 26302 40292
rect 29250 40236 29260 40292
rect 29316 40236 29932 40292
rect 29988 40236 31948 40292
rect 33170 40236 33180 40292
rect 33236 40236 33246 40292
rect 43362 40236 43372 40292
rect 43428 40236 43932 40292
rect 43988 40236 43998 40292
rect 44258 40236 44268 40292
rect 44324 40236 47068 40292
rect 47124 40236 47134 40292
rect 52210 40236 52220 40292
rect 52276 40236 53956 40292
rect 55346 40236 55356 40292
rect 55412 40236 56700 40292
rect 56756 40236 56766 40292
rect 2034 40124 2044 40180
rect 2100 40124 8764 40180
rect 8820 40124 8830 40180
rect 20524 40124 24108 40180
rect 24164 40124 24174 40180
rect 31042 40124 31052 40180
rect 31108 40124 32284 40180
rect 32340 40124 32350 40180
rect 42802 40124 42812 40180
rect 42868 40124 43820 40180
rect 43876 40124 43886 40180
rect 44594 40124 44604 40180
rect 44660 40124 44670 40180
rect 48066 40124 48076 40180
rect 48132 40124 53564 40180
rect 53620 40124 53630 40180
rect 44604 40068 44660 40124
rect 8530 40012 8540 40068
rect 8596 40012 8988 40068
rect 9044 40012 24332 40068
rect 24388 40012 24398 40068
rect 36642 40012 36652 40068
rect 36708 40012 44660 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 23762 39900 23772 39956
rect 23828 39900 26236 39956
rect 26292 39900 26302 39956
rect 30146 39900 30156 39956
rect 30212 39900 33516 39956
rect 33572 39900 33582 39956
rect 40338 39900 40348 39956
rect 40404 39900 48748 39956
rect 48804 39900 48814 39956
rect 30790 39788 30828 39844
rect 30884 39788 30894 39844
rect 38612 39788 41020 39844
rect 41076 39788 43148 39844
rect 43204 39788 43214 39844
rect 55234 39788 55244 39844
rect 55300 39788 56868 39844
rect 0 39732 800 39760
rect 38612 39732 38668 39788
rect 56812 39732 56868 39788
rect 59200 39732 60000 39760
rect 0 39676 1932 39732
rect 1988 39676 1998 39732
rect 8372 39676 10892 39732
rect 10948 39676 10958 39732
rect 11106 39676 11116 39732
rect 11172 39676 11564 39732
rect 11620 39676 12964 39732
rect 26114 39676 26124 39732
rect 26180 39676 27580 39732
rect 27636 39676 27646 39732
rect 28242 39676 28252 39732
rect 28308 39676 29260 39732
rect 29316 39676 29326 39732
rect 30258 39676 30268 39732
rect 30324 39676 31164 39732
rect 31220 39676 31230 39732
rect 32834 39676 32844 39732
rect 32900 39676 37548 39732
rect 37604 39676 38668 39732
rect 51202 39676 51212 39732
rect 51268 39676 52780 39732
rect 52836 39676 56028 39732
rect 56084 39676 56094 39732
rect 56812 39676 60000 39732
rect 0 39648 800 39676
rect 8372 39620 8428 39676
rect 10892 39620 10948 39676
rect 12908 39620 12964 39676
rect 59200 39648 60000 39676
rect 4274 39564 4284 39620
rect 4340 39564 7084 39620
rect 7140 39564 8428 39620
rect 9538 39564 9548 39620
rect 9604 39564 9996 39620
rect 10052 39564 10062 39620
rect 10892 39564 11900 39620
rect 11956 39564 11966 39620
rect 12898 39564 12908 39620
rect 12964 39564 13580 39620
rect 13636 39564 13646 39620
rect 16818 39564 16828 39620
rect 16884 39564 18396 39620
rect 18452 39564 18462 39620
rect 26450 39564 26460 39620
rect 26516 39564 27692 39620
rect 27748 39564 27758 39620
rect 32498 39564 32508 39620
rect 32564 39564 35868 39620
rect 35924 39564 37212 39620
rect 37268 39564 37772 39620
rect 37828 39564 38444 39620
rect 38500 39564 38510 39620
rect 44818 39564 44828 39620
rect 44884 39564 45836 39620
rect 45892 39564 45902 39620
rect 19058 39452 19068 39508
rect 19124 39452 33964 39508
rect 34020 39452 34030 39508
rect 37212 39452 41244 39508
rect 41300 39452 41310 39508
rect 24322 39340 24332 39396
rect 24388 39340 28028 39396
rect 28084 39340 28094 39396
rect 32386 39340 32396 39396
rect 32452 39340 34860 39396
rect 34916 39340 34926 39396
rect 35298 39340 35308 39396
rect 35364 39340 36540 39396
rect 36596 39340 36606 39396
rect 37212 39284 37268 39452
rect 38434 39340 38444 39396
rect 38500 39340 38892 39396
rect 38948 39340 38958 39396
rect 42354 39340 42364 39396
rect 42420 39340 50316 39396
rect 50372 39340 51772 39396
rect 51828 39340 56588 39396
rect 56644 39340 56654 39396
rect 21942 39228 21980 39284
rect 22036 39228 22046 39284
rect 25106 39228 25116 39284
rect 25172 39228 32508 39284
rect 32564 39228 32574 39284
rect 32732 39228 37268 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 5282 39116 5292 39172
rect 5348 39116 6188 39172
rect 6244 39116 6254 39172
rect 0 39060 800 39088
rect 0 39004 1708 39060
rect 1764 39004 1774 39060
rect 9986 39004 9996 39060
rect 10052 39004 10220 39060
rect 10276 39004 11116 39060
rect 11172 39004 11182 39060
rect 12450 39004 12460 39060
rect 12516 39004 13580 39060
rect 13636 39004 13646 39060
rect 27122 39004 27132 39060
rect 27188 39004 28140 39060
rect 28196 39004 28206 39060
rect 30230 39004 30268 39060
rect 30324 39004 30334 39060
rect 0 38976 800 39004
rect 32732 38948 32788 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 34178 39116 34188 39172
rect 34244 39116 41580 39172
rect 41636 39116 41646 39172
rect 59200 39060 60000 39088
rect 33954 39004 33964 39060
rect 34020 39004 34300 39060
rect 34356 39004 37044 39060
rect 55010 39004 55020 39060
rect 55076 39004 60000 39060
rect 36988 38948 37044 39004
rect 59200 38976 60000 39004
rect 2034 38892 2044 38948
rect 2100 38892 4620 38948
rect 4676 38892 4686 38948
rect 16034 38892 16044 38948
rect 16100 38892 17724 38948
rect 17780 38892 17790 38948
rect 22418 38892 22428 38948
rect 22484 38892 22764 38948
rect 22820 38892 32788 38948
rect 35410 38892 35420 38948
rect 35476 38892 35980 38948
rect 36036 38892 36046 38948
rect 36614 38892 36652 38948
rect 36708 38892 36718 38948
rect 36978 38892 36988 38948
rect 37044 38892 37324 38948
rect 37380 38892 45500 38948
rect 45556 38892 50876 38948
rect 50932 38892 52444 38948
rect 52500 38892 53004 38948
rect 53060 38892 56700 38948
rect 56756 38892 56766 38948
rect 4722 38780 4732 38836
rect 4788 38780 5740 38836
rect 5796 38780 5806 38836
rect 5954 38780 5964 38836
rect 6020 38780 6860 38836
rect 6916 38780 6926 38836
rect 25778 38780 25788 38836
rect 25844 38780 26908 38836
rect 26964 38780 26974 38836
rect 35420 38780 35700 38836
rect 44258 38780 44268 38836
rect 44324 38780 53452 38836
rect 53508 38780 53518 38836
rect 5740 38724 5796 38780
rect 35420 38724 35476 38780
rect 35644 38724 35700 38780
rect 5740 38668 6748 38724
rect 6804 38668 6814 38724
rect 27682 38668 27692 38724
rect 27748 38668 29596 38724
rect 29652 38668 29662 38724
rect 35410 38668 35420 38724
rect 35476 38668 35486 38724
rect 35634 38668 35644 38724
rect 35700 38668 35710 38724
rect 42242 38668 42252 38724
rect 42308 38668 42420 38724
rect 43250 38668 43260 38724
rect 43316 38668 44156 38724
rect 44212 38668 45500 38724
rect 45556 38668 45566 38724
rect 47170 38668 47180 38724
rect 47236 38668 49532 38724
rect 49588 38668 49598 38724
rect 42364 38612 42420 38668
rect 5170 38556 5180 38612
rect 5236 38556 6188 38612
rect 6244 38556 6254 38612
rect 21410 38556 21420 38612
rect 21476 38556 21756 38612
rect 21812 38556 21822 38612
rect 42354 38556 42364 38612
rect 42420 38556 42430 38612
rect 46610 38556 46620 38612
rect 46676 38556 46956 38612
rect 47012 38556 47022 38612
rect 5058 38444 5068 38500
rect 5124 38444 5628 38500
rect 5684 38444 6244 38500
rect 18722 38444 18732 38500
rect 18788 38444 25116 38500
rect 25172 38444 25182 38500
rect 28886 38444 28924 38500
rect 28980 38444 28990 38500
rect 38612 38444 39228 38500
rect 39284 38444 39564 38500
rect 39620 38444 39630 38500
rect 0 38388 800 38416
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 6188 38388 6244 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 0 38332 1708 38388
rect 1764 38332 2492 38388
rect 2548 38332 2558 38388
rect 6178 38332 6188 38388
rect 6244 38332 6254 38388
rect 12562 38332 12572 38388
rect 12628 38332 31388 38388
rect 31444 38332 31836 38388
rect 31892 38332 31902 38388
rect 35634 38332 35644 38388
rect 35700 38332 36204 38388
rect 36260 38332 36270 38388
rect 0 38304 800 38332
rect 38612 38276 38668 38444
rect 59200 38388 60000 38416
rect 57362 38332 57372 38388
rect 57428 38332 60000 38388
rect 59200 38304 60000 38332
rect 5842 38220 5852 38276
rect 5908 38220 6076 38276
rect 6132 38220 6142 38276
rect 31052 38220 38668 38276
rect 46834 38220 46844 38276
rect 46900 38220 47292 38276
rect 47348 38220 47358 38276
rect 14130 38108 14140 38164
rect 14196 38108 14812 38164
rect 14868 38108 15148 38164
rect 23762 38108 23772 38164
rect 23828 38108 25676 38164
rect 25732 38108 26124 38164
rect 26180 38108 26190 38164
rect 30146 38108 30156 38164
rect 30212 38108 30828 38164
rect 30884 38108 30894 38164
rect 15092 38052 15148 38108
rect 31052 38052 31108 38220
rect 34962 38108 34972 38164
rect 35028 38108 35980 38164
rect 36036 38108 37772 38164
rect 37828 38108 37838 38164
rect 40338 38108 40348 38164
rect 40404 38108 40908 38164
rect 40964 38108 50876 38164
rect 50932 38108 50942 38164
rect 37772 38052 37828 38108
rect 10882 37996 10892 38052
rect 10948 37996 11564 38052
rect 11620 37996 12012 38052
rect 12068 37996 12078 38052
rect 13010 37996 13020 38052
rect 13076 37996 13804 38052
rect 13860 37996 13870 38052
rect 15092 37996 15820 38052
rect 15876 37996 15886 38052
rect 19954 37996 19964 38052
rect 20020 37996 21196 38052
rect 21252 37996 21262 38052
rect 30706 37996 30716 38052
rect 30772 37996 31108 38052
rect 33506 37996 33516 38052
rect 33572 37996 37100 38052
rect 37156 37996 37166 38052
rect 37772 37996 42812 38052
rect 42868 37996 42878 38052
rect 46610 37996 46620 38052
rect 46676 37996 47068 38052
rect 47124 37996 47134 38052
rect 2034 37884 2044 37940
rect 2100 37884 5404 37940
rect 5460 37884 6076 37940
rect 6132 37884 6412 37940
rect 6468 37884 6478 37940
rect 7634 37884 7644 37940
rect 7700 37884 8764 37940
rect 8820 37884 8830 37940
rect 11330 37884 11340 37940
rect 11396 37884 12236 37940
rect 12292 37884 12302 37940
rect 15474 37884 15484 37940
rect 15540 37884 16604 37940
rect 16660 37884 16670 37940
rect 20850 37884 20860 37940
rect 20916 37884 21756 37940
rect 21812 37884 22316 37940
rect 22372 37884 30492 37940
rect 30548 37884 31388 37940
rect 31444 37884 31454 37940
rect 34290 37884 34300 37940
rect 34356 37884 35084 37940
rect 35140 37884 35150 37940
rect 40562 37884 40572 37940
rect 40628 37884 42028 37940
rect 42084 37884 42094 37940
rect 47842 37884 47852 37940
rect 47908 37884 49532 37940
rect 49588 37884 49598 37940
rect 14242 37772 14252 37828
rect 14308 37772 21308 37828
rect 21364 37772 21374 37828
rect 26002 37772 26012 37828
rect 26068 37772 26908 37828
rect 27794 37772 27804 37828
rect 27860 37772 28588 37828
rect 28644 37772 29036 37828
rect 29092 37772 29102 37828
rect 33954 37772 33964 37828
rect 34020 37772 34636 37828
rect 34692 37772 34702 37828
rect 0 37716 800 37744
rect 0 37660 1708 37716
rect 1764 37660 2492 37716
rect 2548 37660 2558 37716
rect 0 37632 800 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 26852 37604 26908 37772
rect 59200 37716 60000 37744
rect 36194 37660 36204 37716
rect 36260 37660 36988 37716
rect 37044 37660 37054 37716
rect 57922 37660 57932 37716
rect 57988 37660 60000 37716
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 59200 37632 60000 37660
rect 6402 37548 6412 37604
rect 6468 37548 7308 37604
rect 7364 37548 7374 37604
rect 7522 37548 7532 37604
rect 7588 37548 18060 37604
rect 18116 37548 18126 37604
rect 26852 37548 33068 37604
rect 33124 37548 33404 37604
rect 33460 37548 33470 37604
rect 33842 37548 33852 37604
rect 33908 37548 40012 37604
rect 40068 37548 40078 37604
rect 33404 37492 33460 37548
rect 2034 37436 2044 37492
rect 2100 37436 5068 37492
rect 5124 37436 5134 37492
rect 11442 37436 11452 37492
rect 11508 37436 33180 37492
rect 33236 37436 33246 37492
rect 33404 37436 34412 37492
rect 34468 37436 34478 37492
rect 35186 37436 35196 37492
rect 35252 37436 41356 37492
rect 41412 37436 45836 37492
rect 45892 37436 45902 37492
rect 48402 37436 48412 37492
rect 48468 37436 50428 37492
rect 50484 37436 50494 37492
rect 6514 37324 6524 37380
rect 6580 37324 6972 37380
rect 7028 37324 7038 37380
rect 12674 37324 12684 37380
rect 12740 37324 14812 37380
rect 14868 37324 14878 37380
rect 20178 37324 20188 37380
rect 20244 37324 21644 37380
rect 21700 37324 21710 37380
rect 29138 37324 29148 37380
rect 29204 37324 35308 37380
rect 35364 37324 35374 37380
rect 35970 37324 35980 37380
rect 36036 37324 36540 37380
rect 36596 37324 36652 37380
rect 36708 37324 37436 37380
rect 37492 37324 37502 37380
rect 40338 37324 40348 37380
rect 40404 37324 41132 37380
rect 41188 37324 41198 37380
rect 46274 37324 46284 37380
rect 46340 37324 46508 37380
rect 46564 37324 46574 37380
rect 51202 37324 51212 37380
rect 51268 37324 52220 37380
rect 52276 37324 52286 37380
rect 14354 37212 14364 37268
rect 14420 37212 14700 37268
rect 14756 37212 16156 37268
rect 16212 37212 16222 37268
rect 20514 37212 20524 37268
rect 20580 37212 21420 37268
rect 21476 37212 21486 37268
rect 21830 37212 21868 37268
rect 21924 37212 22316 37268
rect 22372 37212 23380 37268
rect 23538 37212 23548 37268
rect 23604 37212 25676 37268
rect 25732 37212 25742 37268
rect 28018 37212 28028 37268
rect 28084 37212 28812 37268
rect 28868 37212 28878 37268
rect 33180 37212 37772 37268
rect 37828 37212 38556 37268
rect 38612 37212 38622 37268
rect 39778 37212 39788 37268
rect 39844 37212 40908 37268
rect 40964 37212 40974 37268
rect 46050 37212 46060 37268
rect 46116 37212 46396 37268
rect 46452 37212 46462 37268
rect 46610 37212 46620 37268
rect 46676 37212 47068 37268
rect 47124 37212 48076 37268
rect 48132 37212 48860 37268
rect 48916 37212 48926 37268
rect 51538 37212 51548 37268
rect 51604 37212 53788 37268
rect 53844 37212 53854 37268
rect 23324 37156 23380 37212
rect 33180 37156 33236 37212
rect 12562 37100 12572 37156
rect 12628 37100 13356 37156
rect 13412 37100 13422 37156
rect 16268 37100 16940 37156
rect 16996 37100 17006 37156
rect 21298 37100 21308 37156
rect 21364 37100 23100 37156
rect 23156 37100 23166 37156
rect 23324 37100 33236 37156
rect 33292 37100 38220 37156
rect 38276 37100 38286 37156
rect 39330 37100 39340 37156
rect 39396 37100 41020 37156
rect 41076 37100 41086 37156
rect 0 37044 800 37072
rect 16268 37044 16324 37100
rect 33292 37044 33348 37100
rect 38220 37044 38276 37100
rect 59200 37044 60000 37072
rect 0 36988 1708 37044
rect 1764 36988 2940 37044
rect 2996 36988 3006 37044
rect 15698 36988 15708 37044
rect 15764 36988 16324 37044
rect 16482 36988 16492 37044
rect 16548 36988 17500 37044
rect 17556 36988 24836 37044
rect 28466 36988 28476 37044
rect 28532 36988 29260 37044
rect 29316 36988 29326 37044
rect 32498 36988 32508 37044
rect 32564 36988 33292 37044
rect 33348 36988 33358 37044
rect 34402 36988 34412 37044
rect 34468 36988 35308 37044
rect 35364 36988 35374 37044
rect 35634 36988 35644 37044
rect 35700 36988 36316 37044
rect 36372 36988 36382 37044
rect 38220 36988 41804 37044
rect 41860 36988 41870 37044
rect 51314 36988 51324 37044
rect 51380 36988 52668 37044
rect 52724 36988 52734 37044
rect 53106 36988 53116 37044
rect 53172 36988 53788 37044
rect 53844 36988 53854 37044
rect 55346 36988 55356 37044
rect 55412 36988 60000 37044
rect 0 36960 800 36988
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 24780 36820 24836 36988
rect 59200 36960 60000 36988
rect 27010 36876 27020 36932
rect 27076 36876 27916 36932
rect 27972 36876 27982 36932
rect 30034 36876 30044 36932
rect 30100 36876 30716 36932
rect 30772 36876 30782 36932
rect 40898 36876 40908 36932
rect 40964 36876 41916 36932
rect 41972 36876 41982 36932
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 24770 36764 24780 36820
rect 24836 36764 26908 36820
rect 27570 36764 27580 36820
rect 27636 36764 28140 36820
rect 28196 36764 28206 36820
rect 26852 36708 26908 36764
rect 17154 36652 17164 36708
rect 17220 36652 26348 36708
rect 26404 36652 26414 36708
rect 26852 36652 32732 36708
rect 32788 36652 32798 36708
rect 34514 36652 34524 36708
rect 34580 36652 36092 36708
rect 36148 36652 36158 36708
rect 36876 36652 36988 36708
rect 37044 36652 37054 36708
rect 42578 36652 42588 36708
rect 42644 36652 43260 36708
rect 43316 36652 43326 36708
rect 46722 36652 46732 36708
rect 46788 36652 49532 36708
rect 49588 36652 49598 36708
rect 36876 36596 36932 36652
rect 2706 36540 2716 36596
rect 2772 36540 6636 36596
rect 6692 36540 6702 36596
rect 7298 36540 7308 36596
rect 7364 36540 8428 36596
rect 8484 36540 8494 36596
rect 19506 36540 19516 36596
rect 19572 36540 20636 36596
rect 20692 36540 33404 36596
rect 33460 36540 33470 36596
rect 34066 36540 34076 36596
rect 34132 36540 36932 36596
rect 37090 36540 37100 36596
rect 37156 36540 49980 36596
rect 50036 36540 50428 36596
rect 50484 36540 50988 36596
rect 51044 36540 51054 36596
rect 52546 36540 52556 36596
rect 52612 36540 54460 36596
rect 54516 36540 54526 36596
rect 34076 36484 34132 36540
rect 1698 36428 1708 36484
rect 1764 36428 2492 36484
rect 2548 36428 2558 36484
rect 11778 36428 11788 36484
rect 11844 36428 13356 36484
rect 13412 36428 13804 36484
rect 13860 36428 14476 36484
rect 14532 36428 14542 36484
rect 16706 36428 16716 36484
rect 16772 36428 17836 36484
rect 17892 36428 18508 36484
rect 18564 36428 18574 36484
rect 26786 36428 26796 36484
rect 26852 36428 27580 36484
rect 27636 36428 27646 36484
rect 31602 36428 31612 36484
rect 31668 36428 32172 36484
rect 32228 36428 34132 36484
rect 34626 36428 34636 36484
rect 34692 36428 38668 36484
rect 39554 36428 39564 36484
rect 39620 36428 40236 36484
rect 40292 36428 40302 36484
rect 41692 36428 42812 36484
rect 42868 36428 47516 36484
rect 47572 36428 47582 36484
rect 0 36372 800 36400
rect 38612 36372 38668 36428
rect 41692 36372 41748 36428
rect 59200 36372 60000 36400
rect 0 36316 2380 36372
rect 2436 36316 3164 36372
rect 3220 36316 3230 36372
rect 17378 36316 17388 36372
rect 17444 36316 17948 36372
rect 18004 36316 24780 36372
rect 24836 36316 24846 36372
rect 27794 36316 27804 36372
rect 27860 36316 28028 36372
rect 28084 36316 28094 36372
rect 34290 36316 34300 36372
rect 34356 36316 35532 36372
rect 35588 36316 35598 36372
rect 35746 36316 35756 36372
rect 35812 36316 35868 36372
rect 35924 36316 35934 36372
rect 38612 36316 41748 36372
rect 41906 36316 41916 36372
rect 41972 36316 49084 36372
rect 49140 36316 52108 36372
rect 52164 36316 53116 36372
rect 53172 36316 53182 36372
rect 58034 36316 58044 36372
rect 58100 36316 60000 36372
rect 0 36288 800 36316
rect 59200 36288 60000 36316
rect 2034 36204 2044 36260
rect 2100 36204 5292 36260
rect 5348 36204 5358 36260
rect 16034 36204 16044 36260
rect 16100 36204 17164 36260
rect 17220 36204 17230 36260
rect 22978 36204 22988 36260
rect 23044 36204 23380 36260
rect 25554 36204 25564 36260
rect 25620 36204 26572 36260
rect 26628 36204 26638 36260
rect 26898 36204 26908 36260
rect 26964 36204 28700 36260
rect 28756 36204 28766 36260
rect 29698 36204 29708 36260
rect 29764 36204 31052 36260
rect 31108 36204 31836 36260
rect 31892 36204 31902 36260
rect 35074 36204 35084 36260
rect 35140 36204 35644 36260
rect 35700 36204 35710 36260
rect 41794 36204 41804 36260
rect 41860 36204 42476 36260
rect 42532 36204 42542 36260
rect 43698 36204 43708 36260
rect 43764 36204 44940 36260
rect 44996 36204 45836 36260
rect 45892 36204 45902 36260
rect 46162 36204 46172 36260
rect 46228 36204 47180 36260
rect 47236 36204 47246 36260
rect 48066 36204 48076 36260
rect 48132 36204 48636 36260
rect 48692 36204 48702 36260
rect 23324 36148 23380 36204
rect 23314 36092 23324 36148
rect 23380 36092 24332 36148
rect 24388 36092 25116 36148
rect 25172 36092 30044 36148
rect 30100 36092 30110 36148
rect 30258 36092 30268 36148
rect 30324 36092 30362 36148
rect 30706 36092 30716 36148
rect 30772 36092 39004 36148
rect 39060 36092 40572 36148
rect 40628 36092 41132 36148
rect 41188 36092 41198 36148
rect 41906 36092 41916 36148
rect 41972 36092 42252 36148
rect 42308 36092 42318 36148
rect 46050 36092 46060 36148
rect 46116 36092 46956 36148
rect 47012 36092 47022 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 30454 35980 30492 36036
rect 30548 35980 30558 36036
rect 30716 35924 30772 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 39666 35980 39676 36036
rect 39732 35980 40236 36036
rect 40292 35980 40302 36036
rect 52210 35980 52220 36036
rect 52276 35980 53004 36036
rect 53060 35980 53070 36036
rect 14578 35868 14588 35924
rect 14644 35868 15596 35924
rect 15652 35868 15662 35924
rect 24098 35868 24108 35924
rect 24164 35868 24668 35924
rect 24724 35868 30772 35924
rect 36978 35868 36988 35924
rect 37044 35868 41244 35924
rect 41300 35868 41310 35924
rect 45490 35868 45500 35924
rect 45556 35868 55580 35924
rect 55636 35868 55646 35924
rect 7970 35756 7980 35812
rect 8036 35756 8316 35812
rect 8372 35756 12012 35812
rect 12068 35756 12078 35812
rect 12450 35756 12460 35812
rect 12516 35756 14364 35812
rect 14420 35756 15036 35812
rect 15092 35756 15102 35812
rect 27794 35756 27804 35812
rect 27860 35756 31164 35812
rect 31220 35756 31612 35812
rect 31668 35756 38668 35812
rect 45266 35756 45276 35812
rect 45332 35756 46508 35812
rect 46564 35756 46574 35812
rect 47170 35756 47180 35812
rect 47236 35756 47852 35812
rect 47908 35756 47918 35812
rect 48066 35756 48076 35812
rect 48132 35756 50092 35812
rect 50148 35756 52892 35812
rect 52948 35756 52958 35812
rect 0 35700 800 35728
rect 38612 35700 38668 35756
rect 51100 35700 51156 35756
rect 59200 35700 60000 35728
rect 0 35644 1708 35700
rect 1764 35644 1774 35700
rect 4274 35644 4284 35700
rect 4340 35644 7532 35700
rect 7588 35644 7598 35700
rect 14130 35644 14140 35700
rect 14196 35644 15148 35700
rect 23650 35644 23660 35700
rect 23716 35644 23726 35700
rect 30818 35644 30828 35700
rect 30884 35644 31276 35700
rect 31332 35644 31342 35700
rect 32722 35644 32732 35700
rect 32788 35644 34188 35700
rect 34244 35644 38388 35700
rect 38612 35644 40908 35700
rect 40964 35644 40974 35700
rect 42018 35644 42028 35700
rect 42084 35644 43484 35700
rect 43540 35644 43550 35700
rect 51090 35644 51100 35700
rect 51156 35644 51166 35700
rect 52098 35644 52108 35700
rect 52164 35644 53452 35700
rect 53508 35644 53518 35700
rect 55010 35644 55020 35700
rect 55076 35644 60000 35700
rect 0 35616 800 35644
rect 5170 35532 5180 35588
rect 5236 35532 8428 35588
rect 8484 35532 9548 35588
rect 9604 35532 11004 35588
rect 11060 35532 12908 35588
rect 12964 35532 12974 35588
rect 15092 35532 15148 35644
rect 23660 35588 23716 35644
rect 15204 35532 15214 35588
rect 23426 35532 23436 35588
rect 23492 35532 25452 35588
rect 25508 35532 29036 35588
rect 29092 35532 29102 35588
rect 30258 35532 30268 35588
rect 30324 35532 30604 35588
rect 30660 35532 30670 35588
rect 32946 35532 32956 35588
rect 33012 35532 34076 35588
rect 34132 35532 34142 35588
rect 35186 35532 35196 35588
rect 35252 35532 37548 35588
rect 37604 35532 38108 35588
rect 38164 35532 38174 35588
rect 12562 35420 12572 35476
rect 12628 35420 13692 35476
rect 13748 35420 13758 35476
rect 30454 35420 30492 35476
rect 30548 35420 30558 35476
rect 10994 35308 11004 35364
rect 11060 35308 14252 35364
rect 14308 35308 14318 35364
rect 22642 35308 22652 35364
rect 22708 35308 22718 35364
rect 28914 35308 28924 35364
rect 28980 35308 29708 35364
rect 29764 35308 30828 35364
rect 30884 35308 30894 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 22652 35252 22708 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 38332 35252 38388 35644
rect 59200 35616 60000 35644
rect 42802 35532 42812 35588
rect 42868 35532 45948 35588
rect 46004 35532 46014 35588
rect 50418 35532 50428 35588
rect 50484 35532 52444 35588
rect 52500 35532 53004 35588
rect 53060 35532 53070 35588
rect 46498 35420 46508 35476
rect 46564 35420 47964 35476
rect 48020 35420 48030 35476
rect 50306 35420 50316 35476
rect 50372 35420 51772 35476
rect 51828 35420 51996 35476
rect 52052 35420 52062 35476
rect 50316 35364 50372 35420
rect 42690 35308 42700 35364
rect 42756 35308 43260 35364
rect 43316 35308 50372 35364
rect 50642 35308 50652 35364
rect 50708 35308 52220 35364
rect 52276 35308 52286 35364
rect 22652 35196 23548 35252
rect 23604 35196 23614 35252
rect 31490 35196 31500 35252
rect 31556 35196 32508 35252
rect 32564 35196 33740 35252
rect 33796 35196 33806 35252
rect 38332 35196 40908 35252
rect 40964 35196 41468 35252
rect 41524 35196 46844 35252
rect 46900 35196 46910 35252
rect 31686 35084 31724 35140
rect 31780 35084 31790 35140
rect 37650 35084 37660 35140
rect 37716 35084 40012 35140
rect 40068 35084 40078 35140
rect 43474 35084 43484 35140
rect 43540 35084 44940 35140
rect 44996 35084 45006 35140
rect 46610 35084 46620 35140
rect 46676 35084 46956 35140
rect 47012 35084 47022 35140
rect 0 35028 800 35056
rect 59200 35028 60000 35056
rect 0 34972 1932 35028
rect 1988 34972 1998 35028
rect 34514 34972 34524 35028
rect 34580 34972 35868 35028
rect 35924 34972 37100 35028
rect 37156 34972 37166 35028
rect 51538 34972 51548 35028
rect 51604 34972 51996 35028
rect 52052 34972 52062 35028
rect 55346 34972 55356 35028
rect 55412 34972 60000 35028
rect 0 34944 800 34972
rect 59200 34944 60000 34972
rect 23202 34860 23212 34916
rect 23268 34860 24108 34916
rect 24164 34860 24174 34916
rect 27542 34860 27580 34916
rect 27636 34860 28140 34916
rect 28196 34860 28206 34916
rect 39442 34860 39452 34916
rect 39508 34860 40124 34916
rect 40180 34860 40190 34916
rect 41990 34860 42028 34916
rect 42084 34860 42094 34916
rect 42354 34860 42364 34916
rect 42420 34860 42924 34916
rect 42980 34860 42990 34916
rect 51650 34860 51660 34916
rect 51716 34860 52780 34916
rect 52836 34860 52846 34916
rect 21634 34748 21644 34804
rect 21700 34748 22876 34804
rect 22932 34748 22942 34804
rect 23874 34748 23884 34804
rect 23940 34748 31388 34804
rect 31444 34748 31454 34804
rect 31836 34748 38668 34804
rect 39218 34748 39228 34804
rect 39284 34748 39788 34804
rect 39844 34748 50204 34804
rect 50260 34748 50270 34804
rect 31836 34692 31892 34748
rect 38612 34692 38668 34748
rect 13346 34636 13356 34692
rect 13412 34636 14140 34692
rect 14196 34636 14206 34692
rect 22418 34636 22428 34692
rect 22484 34636 23212 34692
rect 23268 34636 23278 34692
rect 23762 34636 23772 34692
rect 23828 34636 24444 34692
rect 24500 34636 24510 34692
rect 26450 34636 26460 34692
rect 26516 34636 27244 34692
rect 27300 34636 27310 34692
rect 28802 34636 28812 34692
rect 28868 34636 29484 34692
rect 29540 34636 30268 34692
rect 30324 34636 31892 34692
rect 33730 34636 33740 34692
rect 33796 34636 34300 34692
rect 34356 34636 35532 34692
rect 35588 34636 35598 34692
rect 38612 34636 38780 34692
rect 38836 34636 38846 34692
rect 39666 34636 39676 34692
rect 39732 34636 40348 34692
rect 40404 34636 40414 34692
rect 41682 34636 41692 34692
rect 41748 34636 44044 34692
rect 44100 34636 44110 34692
rect 45938 34636 45948 34692
rect 46004 34636 46956 34692
rect 47012 34636 47022 34692
rect 47170 34636 47180 34692
rect 47236 34636 49868 34692
rect 49924 34636 49934 34692
rect 33954 34524 33964 34580
rect 34020 34524 34748 34580
rect 34804 34524 36428 34580
rect 36484 34524 36494 34580
rect 45826 34524 45836 34580
rect 45892 34524 47292 34580
rect 47348 34524 47358 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 34962 34412 34972 34468
rect 35028 34412 36540 34468
rect 36596 34412 36606 34468
rect 59200 34356 60000 34384
rect 10994 34300 11004 34356
rect 11060 34300 12236 34356
rect 12292 34300 12684 34356
rect 12740 34300 15148 34356
rect 15204 34300 17052 34356
rect 17108 34300 17118 34356
rect 17602 34300 17612 34356
rect 17668 34300 18396 34356
rect 18452 34300 18462 34356
rect 27906 34300 27916 34356
rect 27972 34300 29988 34356
rect 34374 34300 34412 34356
rect 34468 34300 34478 34356
rect 37090 34300 37100 34356
rect 37156 34300 41132 34356
rect 41188 34300 42028 34356
rect 42084 34300 42094 34356
rect 57922 34300 57932 34356
rect 57988 34300 60000 34356
rect 17612 34244 17668 34300
rect 29932 34244 29988 34300
rect 59200 34272 60000 34300
rect 16146 34188 16156 34244
rect 16212 34188 17668 34244
rect 20962 34188 20972 34244
rect 21028 34188 28028 34244
rect 28084 34188 28094 34244
rect 29922 34188 29932 34244
rect 29988 34188 30492 34244
rect 30548 34188 30558 34244
rect 47954 34188 47964 34244
rect 48020 34188 48748 34244
rect 48804 34188 48814 34244
rect 1922 34076 1932 34132
rect 1988 34076 5068 34132
rect 5124 34076 5628 34132
rect 5684 34076 5694 34132
rect 16370 34076 16380 34132
rect 16436 34076 17948 34132
rect 18004 34076 18014 34132
rect 34402 34076 34412 34132
rect 34468 34076 36204 34132
rect 36260 34076 36270 34132
rect 46946 34076 46956 34132
rect 47012 34076 47404 34132
rect 47460 34076 47470 34132
rect 48962 34076 48972 34132
rect 49028 34076 49756 34132
rect 49812 34076 49822 34132
rect 4284 33964 10220 34020
rect 10276 33964 11004 34020
rect 11060 33964 11070 34020
rect 17714 33964 17724 34020
rect 17780 33964 18508 34020
rect 18564 33964 18574 34020
rect 23538 33964 23548 34020
rect 23604 33964 31612 34020
rect 31668 33964 32284 34020
rect 32340 33964 32350 34020
rect 34178 33964 34188 34020
rect 34244 33964 34748 34020
rect 34804 33964 36652 34020
rect 36708 33964 36718 34020
rect 42018 33964 42028 34020
rect 42084 33964 43708 34020
rect 43764 33964 43774 34020
rect 50978 33964 50988 34020
rect 51044 33964 51996 34020
rect 52052 33964 52062 34020
rect 4284 33908 4340 33964
rect 4274 33852 4284 33908
rect 4340 33852 4350 33908
rect 5842 33852 5852 33908
rect 5908 33852 7196 33908
rect 7252 33852 8652 33908
rect 8708 33852 10556 33908
rect 10612 33852 11564 33908
rect 11620 33852 11630 33908
rect 33618 33852 33628 33908
rect 33684 33852 34972 33908
rect 35028 33852 35038 33908
rect 36754 33852 36764 33908
rect 36820 33852 37772 33908
rect 37828 33852 37838 33908
rect 50372 33852 51772 33908
rect 51828 33852 51838 33908
rect 18498 33740 18508 33796
rect 18564 33740 21756 33796
rect 21812 33740 22764 33796
rect 22820 33740 22830 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 50372 33684 50428 33852
rect 18274 33628 18284 33684
rect 18340 33628 19068 33684
rect 19124 33628 19134 33684
rect 35634 33628 35644 33684
rect 35700 33628 36540 33684
rect 36596 33628 37436 33684
rect 37492 33628 37502 33684
rect 38994 33628 39004 33684
rect 39060 33628 40348 33684
rect 40404 33628 40414 33684
rect 46610 33628 46620 33684
rect 46676 33628 48748 33684
rect 48804 33628 48814 33684
rect 50194 33628 50204 33684
rect 50260 33628 50428 33684
rect 51874 33628 51884 33684
rect 51940 33628 52556 33684
rect 52612 33628 52622 33684
rect 18834 33516 18844 33572
rect 18900 33516 25900 33572
rect 25956 33516 25966 33572
rect 31014 33516 31052 33572
rect 31108 33516 31118 33572
rect 45826 33516 45836 33572
rect 45892 33516 47740 33572
rect 47796 33516 52220 33572
rect 52276 33516 52668 33572
rect 52724 33516 52734 33572
rect 4722 33404 4732 33460
rect 4788 33404 5292 33460
rect 5348 33404 5740 33460
rect 5796 33404 5806 33460
rect 7074 33404 7084 33460
rect 7140 33404 8540 33460
rect 8596 33404 10444 33460
rect 10500 33404 11452 33460
rect 11508 33404 11518 33460
rect 14242 33404 14252 33460
rect 14308 33404 15484 33460
rect 15540 33404 15550 33460
rect 20290 33404 20300 33460
rect 20356 33404 21084 33460
rect 21140 33404 21868 33460
rect 21924 33404 21934 33460
rect 30930 33404 30940 33460
rect 30996 33404 31276 33460
rect 31332 33404 31342 33460
rect 51426 33404 51436 33460
rect 51492 33404 53228 33460
rect 53284 33404 53564 33460
rect 53620 33404 53630 33460
rect 12898 33292 12908 33348
rect 12964 33292 13580 33348
rect 13636 33292 14028 33348
rect 14084 33292 14094 33348
rect 19506 33292 19516 33348
rect 19572 33292 22988 33348
rect 23044 33292 24220 33348
rect 24276 33292 24892 33348
rect 24948 33292 25340 33348
rect 25396 33292 25406 33348
rect 15474 33180 15484 33236
rect 15540 33180 16492 33236
rect 16548 33180 16558 33236
rect 22502 33180 22540 33236
rect 22596 33180 22606 33236
rect 24546 33180 24556 33236
rect 24612 33180 25676 33236
rect 25732 33180 25742 33236
rect 28578 33180 28588 33236
rect 28644 33180 31276 33236
rect 31332 33180 31342 33236
rect 31714 33180 31724 33236
rect 31780 33180 32508 33236
rect 32564 33180 32574 33236
rect 39442 33180 39452 33236
rect 39508 33180 39676 33236
rect 39732 33180 39742 33236
rect 44258 33180 44268 33236
rect 44324 33180 45612 33236
rect 45668 33180 45678 33236
rect 5842 33068 5852 33124
rect 5908 33068 6300 33124
rect 6356 33068 6366 33124
rect 11666 33068 11676 33124
rect 11732 33068 13468 33124
rect 13524 33068 14364 33124
rect 14420 33068 14924 33124
rect 14980 33068 14990 33124
rect 15138 33068 15148 33124
rect 15204 33068 16156 33124
rect 16212 33068 16222 33124
rect 16818 33068 16828 33124
rect 16884 33068 17612 33124
rect 17668 33068 23548 33124
rect 23604 33068 23614 33124
rect 32050 33068 32060 33124
rect 32116 33068 32956 33124
rect 33012 33068 33022 33124
rect 33842 33068 33852 33124
rect 33908 33068 34300 33124
rect 34356 33068 34366 33124
rect 35298 33068 35308 33124
rect 35364 33068 35980 33124
rect 36036 33068 37100 33124
rect 37156 33068 37166 33124
rect 40002 33068 40012 33124
rect 40068 33068 55356 33124
rect 55412 33068 55422 33124
rect 14242 32956 14252 33012
rect 14308 32956 17276 33012
rect 17332 32956 17342 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 14466 32844 14476 32900
rect 14532 32844 15148 32900
rect 15204 32844 15214 32900
rect 25666 32844 25676 32900
rect 25732 32844 27804 32900
rect 27860 32844 29484 32900
rect 29540 32844 29550 32900
rect 14550 32732 14588 32788
rect 14644 32732 14654 32788
rect 18610 32732 18620 32788
rect 18676 32732 19740 32788
rect 19796 32732 20860 32788
rect 20916 32732 22540 32788
rect 22596 32732 23548 32788
rect 24434 32732 24444 32788
rect 24500 32732 25564 32788
rect 25620 32732 25630 32788
rect 28466 32732 28476 32788
rect 28532 32732 29820 32788
rect 29876 32732 29886 32788
rect 38882 32732 38892 32788
rect 38948 32732 39340 32788
rect 39396 32732 39406 32788
rect 50530 32732 50540 32788
rect 50596 32732 51884 32788
rect 51940 32732 53228 32788
rect 53284 32732 55916 32788
rect 55972 32732 55982 32788
rect 23492 32676 23548 32732
rect 4610 32620 4620 32676
rect 4676 32620 5404 32676
rect 5460 32620 5470 32676
rect 6962 32620 6972 32676
rect 7028 32620 7532 32676
rect 7588 32620 9772 32676
rect 9828 32620 9838 32676
rect 23492 32620 25228 32676
rect 25284 32620 25294 32676
rect 25890 32620 25900 32676
rect 25956 32620 30044 32676
rect 30100 32620 31388 32676
rect 31444 32620 31454 32676
rect 35410 32620 35420 32676
rect 35476 32620 36316 32676
rect 36372 32620 36382 32676
rect 50372 32620 51660 32676
rect 51716 32620 51726 32676
rect 8530 32508 8540 32564
rect 8596 32508 9996 32564
rect 10052 32508 10062 32564
rect 15362 32508 15372 32564
rect 15428 32508 15932 32564
rect 15988 32508 15998 32564
rect 25442 32508 25452 32564
rect 25508 32508 26908 32564
rect 32946 32508 32956 32564
rect 33012 32508 33740 32564
rect 33796 32508 41692 32564
rect 41748 32508 42812 32564
rect 42868 32508 45052 32564
rect 45108 32508 47964 32564
rect 48020 32508 48030 32564
rect 6290 32396 6300 32452
rect 6356 32396 7644 32452
rect 7700 32396 8316 32452
rect 8372 32396 12348 32452
rect 12404 32396 12414 32452
rect 15092 32396 16828 32452
rect 16884 32396 16894 32452
rect 0 32340 800 32368
rect 15092 32340 15148 32396
rect 0 32284 1708 32340
rect 1764 32284 1774 32340
rect 13906 32284 13916 32340
rect 13972 32284 14140 32340
rect 14196 32284 14364 32340
rect 14420 32284 15148 32340
rect 26852 32340 26908 32508
rect 29250 32396 29260 32452
rect 29316 32396 33852 32452
rect 33908 32396 33918 32452
rect 35970 32396 35980 32452
rect 36036 32396 37212 32452
rect 37268 32396 38332 32452
rect 38388 32396 38398 32452
rect 50306 32396 50316 32452
rect 50372 32396 50428 32620
rect 51874 32508 51884 32564
rect 51940 32508 52220 32564
rect 52276 32508 52286 32564
rect 26852 32284 27244 32340
rect 27300 32284 29148 32340
rect 29204 32284 29708 32340
rect 29764 32284 31052 32340
rect 31108 32284 31836 32340
rect 31892 32284 40684 32340
rect 40740 32284 41244 32340
rect 41300 32284 41310 32340
rect 42130 32284 42140 32340
rect 42196 32284 42252 32340
rect 42308 32284 42318 32340
rect 0 32256 800 32284
rect 39442 32172 39452 32228
rect 39508 32172 41468 32228
rect 41524 32172 44604 32228
rect 44660 32172 53788 32228
rect 53844 32172 53854 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 13346 32060 13356 32116
rect 13412 32060 13804 32116
rect 13860 32060 14140 32116
rect 14196 32060 14206 32116
rect 23202 32060 23212 32116
rect 23268 32060 23660 32116
rect 23716 32060 23726 32116
rect 36754 32060 36764 32116
rect 36820 32060 40348 32116
rect 40404 32060 40414 32116
rect 4060 31948 5180 32004
rect 5236 31948 5246 32004
rect 5394 31948 5404 32004
rect 5460 31948 6188 32004
rect 6244 31948 6254 32004
rect 7634 31948 7644 32004
rect 7700 31948 9548 32004
rect 9604 31948 9614 32004
rect 26674 31948 26684 32004
rect 26740 31948 45836 32004
rect 45892 31948 45902 32004
rect 4060 31892 4116 31948
rect 3042 31836 3052 31892
rect 3108 31836 3388 31892
rect 3444 31836 3454 31892
rect 4050 31836 4060 31892
rect 4116 31836 4126 31892
rect 6300 31836 10220 31892
rect 10276 31836 11564 31892
rect 11620 31836 11630 31892
rect 14914 31836 14924 31892
rect 14980 31836 15820 31892
rect 15876 31836 15886 31892
rect 23986 31836 23996 31892
rect 24052 31836 24668 31892
rect 24724 31836 24734 31892
rect 28578 31836 28588 31892
rect 28644 31836 29148 31892
rect 29204 31836 30380 31892
rect 30436 31836 30446 31892
rect 38546 31836 38556 31892
rect 38612 31836 39452 31892
rect 39508 31836 39518 31892
rect 43586 31836 43596 31892
rect 43652 31836 45388 31892
rect 45444 31836 45454 31892
rect 47506 31836 47516 31892
rect 47572 31836 48188 31892
rect 48244 31836 48254 31892
rect 3714 31724 3724 31780
rect 3780 31724 4620 31780
rect 4676 31724 4686 31780
rect 0 31668 800 31696
rect 6300 31668 6356 31836
rect 6514 31724 6524 31780
rect 6580 31724 9436 31780
rect 9492 31724 9502 31780
rect 9650 31724 9660 31780
rect 9716 31724 29484 31780
rect 29540 31724 30156 31780
rect 30212 31724 30222 31780
rect 36866 31724 36876 31780
rect 36932 31724 38444 31780
rect 38500 31724 38510 31780
rect 50866 31724 50876 31780
rect 50932 31724 51548 31780
rect 51604 31724 52556 31780
rect 52612 31724 52622 31780
rect 0 31612 1876 31668
rect 2930 31612 2940 31668
rect 2996 31612 3836 31668
rect 3892 31612 3902 31668
rect 4498 31612 4508 31668
rect 4564 31612 5516 31668
rect 5572 31612 5964 31668
rect 6020 31612 6356 31668
rect 8978 31612 8988 31668
rect 9044 31612 10108 31668
rect 10164 31612 10174 31668
rect 10322 31612 10332 31668
rect 10388 31612 10668 31668
rect 10724 31612 10734 31668
rect 11330 31612 11340 31668
rect 11396 31612 12124 31668
rect 12180 31612 12190 31668
rect 14690 31612 14700 31668
rect 14756 31612 14766 31668
rect 14914 31612 14924 31668
rect 14980 31612 15260 31668
rect 15316 31612 15326 31668
rect 15586 31612 15596 31668
rect 15652 31612 17164 31668
rect 17220 31612 17230 31668
rect 17378 31612 17388 31668
rect 17444 31612 18732 31668
rect 18788 31612 18798 31668
rect 20514 31612 20524 31668
rect 20580 31612 22876 31668
rect 22932 31612 22942 31668
rect 23874 31612 23884 31668
rect 23940 31612 24556 31668
rect 24612 31612 24622 31668
rect 26002 31612 26012 31668
rect 26068 31612 32172 31668
rect 32228 31612 35868 31668
rect 35924 31612 45948 31668
rect 46004 31612 46508 31668
rect 46564 31612 49420 31668
rect 49476 31612 49486 31668
rect 52892 31612 55020 31668
rect 55076 31612 55086 31668
rect 0 31584 800 31612
rect 1820 31220 1876 31612
rect 2034 31500 2044 31556
rect 2100 31500 2110 31556
rect 3154 31500 3164 31556
rect 3220 31500 4732 31556
rect 4788 31500 4798 31556
rect 5058 31500 5068 31556
rect 5124 31500 10220 31556
rect 10276 31500 10286 31556
rect 2044 31332 2100 31500
rect 10444 31444 10500 31612
rect 14700 31556 14756 31612
rect 52892 31556 52948 31612
rect 11106 31500 11116 31556
rect 11172 31500 12572 31556
rect 12628 31500 12638 31556
rect 14700 31500 16380 31556
rect 16436 31500 16446 31556
rect 22530 31500 22540 31556
rect 22596 31500 24780 31556
rect 24836 31500 24846 31556
rect 29810 31500 29820 31556
rect 29876 31500 30268 31556
rect 30324 31500 30334 31556
rect 31714 31500 31724 31556
rect 31780 31500 43148 31556
rect 43204 31500 44156 31556
rect 44212 31500 44222 31556
rect 50082 31500 50092 31556
rect 50148 31500 52892 31556
rect 52948 31500 52958 31556
rect 7522 31388 7532 31444
rect 7588 31388 9100 31444
rect 9156 31388 9548 31444
rect 9604 31388 10500 31444
rect 13906 31388 13916 31444
rect 13972 31388 16940 31444
rect 16996 31388 17006 31444
rect 21522 31388 21532 31444
rect 21588 31388 33964 31444
rect 34020 31388 34300 31444
rect 34356 31388 36988 31444
rect 37044 31388 37054 31444
rect 39638 31388 39676 31444
rect 39732 31388 43596 31444
rect 43652 31388 43662 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 2044 31276 8540 31332
rect 8596 31276 8606 31332
rect 15698 31276 15708 31332
rect 15764 31276 17724 31332
rect 17780 31276 17790 31332
rect 22530 31276 22540 31332
rect 22596 31276 24444 31332
rect 24500 31276 24510 31332
rect 52994 31276 53004 31332
rect 53060 31276 53340 31332
rect 53396 31276 54236 31332
rect 54292 31276 54796 31332
rect 54852 31276 54862 31332
rect 1810 31164 1820 31220
rect 1876 31164 5964 31220
rect 6020 31164 6030 31220
rect 17154 31164 17164 31220
rect 17220 31164 18844 31220
rect 18900 31164 18910 31220
rect 20290 31164 20300 31220
rect 20356 31164 22316 31220
rect 22372 31164 22988 31220
rect 23044 31164 23054 31220
rect 24658 31164 24668 31220
rect 24724 31164 25452 31220
rect 25508 31164 25518 31220
rect 29922 31164 29932 31220
rect 29988 31164 30716 31220
rect 30772 31164 31948 31220
rect 32004 31164 33180 31220
rect 33236 31164 33246 31220
rect 36642 31164 36652 31220
rect 36708 31164 37100 31220
rect 37156 31164 38108 31220
rect 38164 31164 38174 31220
rect 41682 31164 41692 31220
rect 41748 31164 42700 31220
rect 42756 31164 54460 31220
rect 54516 31164 54908 31220
rect 54964 31164 55692 31220
rect 55748 31164 56364 31220
rect 56420 31164 56700 31220
rect 56756 31164 56766 31220
rect 2034 31052 2044 31108
rect 2100 31052 8428 31108
rect 8484 31052 9100 31108
rect 9156 31052 9166 31108
rect 30258 31052 30268 31108
rect 30324 31052 31724 31108
rect 31780 31052 31790 31108
rect 38612 31052 40124 31108
rect 40180 31052 41020 31108
rect 41076 31052 41086 31108
rect 44594 31052 44604 31108
rect 44660 31052 45724 31108
rect 45780 31052 45790 31108
rect 46022 31052 46060 31108
rect 46116 31052 46126 31108
rect 47842 31052 47852 31108
rect 47908 31052 48860 31108
rect 48916 31052 48926 31108
rect 0 30996 800 31024
rect 38612 30996 38668 31052
rect 0 30940 2380 30996
rect 2436 30940 3164 30996
rect 3220 30940 3230 30996
rect 10770 30940 10780 30996
rect 10836 30940 12460 30996
rect 12516 30940 12526 30996
rect 16370 30940 16380 30996
rect 16436 30940 17724 30996
rect 17780 30940 17790 30996
rect 18610 30940 18620 30996
rect 18676 30940 19068 30996
rect 19124 30940 19628 30996
rect 19684 30940 19852 30996
rect 19908 30940 21868 30996
rect 21924 30940 21934 30996
rect 23090 30940 23100 30996
rect 23156 30940 23772 30996
rect 23828 30940 23838 30996
rect 24434 30940 24444 30996
rect 24500 30940 29484 30996
rect 29540 30940 29550 30996
rect 29810 30940 29820 30996
rect 29876 30940 31836 30996
rect 31892 30940 31902 30996
rect 34150 30940 34188 30996
rect 34244 30940 34254 30996
rect 36726 30940 36764 30996
rect 36820 30940 36830 30996
rect 38098 30940 38108 30996
rect 38164 30940 38668 30996
rect 54674 30940 54684 30996
rect 54740 30940 55580 30996
rect 55636 30940 55646 30996
rect 0 30912 800 30940
rect 3042 30828 3052 30884
rect 3108 30828 6412 30884
rect 6468 30828 6478 30884
rect 12786 30828 12796 30884
rect 12852 30828 13244 30884
rect 13300 30828 14364 30884
rect 14420 30828 14430 30884
rect 15138 30828 15148 30884
rect 15204 30828 15596 30884
rect 15652 30828 15662 30884
rect 23650 30828 23660 30884
rect 23716 30828 25340 30884
rect 25396 30828 25406 30884
rect 31154 30828 31164 30884
rect 31220 30828 33852 30884
rect 33908 30828 33918 30884
rect 35858 30828 35868 30884
rect 35924 30828 37212 30884
rect 37268 30828 37278 30884
rect 38546 30828 38556 30884
rect 38612 30828 39676 30884
rect 39732 30828 40796 30884
rect 40852 30828 40862 30884
rect 41010 30828 41020 30884
rect 41076 30828 43036 30884
rect 43092 30828 43102 30884
rect 44034 30828 44044 30884
rect 44100 30828 45052 30884
rect 45108 30828 47516 30884
rect 47572 30828 48860 30884
rect 48916 30828 51996 30884
rect 52052 30828 54964 30884
rect 54908 30772 54964 30828
rect 2706 30716 2716 30772
rect 2772 30716 9324 30772
rect 9380 30716 9996 30772
rect 10052 30716 11004 30772
rect 11060 30716 11070 30772
rect 19170 30716 19180 30772
rect 19236 30716 24332 30772
rect 24388 30716 24398 30772
rect 31938 30716 31948 30772
rect 32004 30716 33516 30772
rect 33572 30716 33582 30772
rect 34972 30716 35644 30772
rect 35700 30716 35710 30772
rect 36502 30716 36540 30772
rect 36596 30716 36606 30772
rect 37874 30716 37884 30772
rect 37940 30716 39340 30772
rect 39396 30716 39406 30772
rect 50372 30716 53004 30772
rect 53060 30716 53070 30772
rect 54898 30716 54908 30772
rect 54964 30716 54974 30772
rect 27794 30604 27804 30660
rect 27860 30604 30492 30660
rect 30548 30604 31500 30660
rect 31556 30604 31566 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 34972 30548 35028 30716
rect 50372 30660 50428 30716
rect 36306 30604 36316 30660
rect 36372 30604 50428 30660
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 16482 30492 16492 30548
rect 16548 30492 17164 30548
rect 17220 30492 18060 30548
rect 18116 30492 18732 30548
rect 18788 30492 18798 30548
rect 21746 30492 21756 30548
rect 21812 30492 34636 30548
rect 34692 30492 35028 30548
rect 36978 30492 36988 30548
rect 37044 30492 37548 30548
rect 37604 30492 37614 30548
rect 43698 30492 43708 30548
rect 43764 30492 52220 30548
rect 52276 30492 52286 30548
rect 3378 30380 3388 30436
rect 3444 30380 7980 30436
rect 8036 30380 8876 30436
rect 8932 30380 8942 30436
rect 11554 30380 11564 30436
rect 11620 30380 17388 30436
rect 17444 30380 21532 30436
rect 21588 30380 22316 30436
rect 22372 30380 22382 30436
rect 22530 30380 22540 30436
rect 22596 30380 22876 30436
rect 22932 30380 22942 30436
rect 31602 30380 31612 30436
rect 31668 30380 31678 30436
rect 34412 30380 38108 30436
rect 38164 30380 38174 30436
rect 46050 30380 46060 30436
rect 46116 30380 47852 30436
rect 47908 30380 49644 30436
rect 49700 30380 51436 30436
rect 51492 30380 51502 30436
rect 0 30324 800 30352
rect 31612 30324 31668 30380
rect 34412 30324 34468 30380
rect 0 30268 3052 30324
rect 3108 30268 3118 30324
rect 9538 30268 9548 30324
rect 9604 30268 10220 30324
rect 10276 30268 10286 30324
rect 13010 30268 13020 30324
rect 13076 30268 15372 30324
rect 15428 30268 15438 30324
rect 22418 30268 22428 30324
rect 22484 30268 23548 30324
rect 23604 30268 23614 30324
rect 29698 30268 29708 30324
rect 29764 30268 30156 30324
rect 30212 30268 30222 30324
rect 31612 30268 34412 30324
rect 34468 30268 34478 30324
rect 35074 30268 35084 30324
rect 35140 30268 37212 30324
rect 37268 30268 37278 30324
rect 52098 30268 52108 30324
rect 52164 30268 54460 30324
rect 54516 30268 58156 30324
rect 58212 30268 58222 30324
rect 0 30240 800 30268
rect 2818 30156 2828 30212
rect 2884 30156 5740 30212
rect 5796 30156 5806 30212
rect 8194 30156 8204 30212
rect 8260 30156 10556 30212
rect 10612 30156 10622 30212
rect 16930 30156 16940 30212
rect 16996 30156 17836 30212
rect 17892 30156 18956 30212
rect 19012 30156 19022 30212
rect 24210 30156 24220 30212
rect 24276 30156 26908 30212
rect 31602 30156 31612 30212
rect 31668 30156 33740 30212
rect 33796 30156 34524 30212
rect 34580 30156 34590 30212
rect 34822 30156 34860 30212
rect 34916 30156 34926 30212
rect 35522 30156 35532 30212
rect 35588 30156 36316 30212
rect 36372 30156 37772 30212
rect 37828 30156 37838 30212
rect 38210 30156 38220 30212
rect 38276 30156 38668 30212
rect 38724 30156 38734 30212
rect 40226 30156 40236 30212
rect 40292 30156 40684 30212
rect 40740 30156 40750 30212
rect 49074 30156 49084 30212
rect 49140 30156 50988 30212
rect 51044 30156 51054 30212
rect 52770 30156 52780 30212
rect 52836 30156 54236 30212
rect 54292 30156 55916 30212
rect 55972 30156 55982 30212
rect 2482 30044 2492 30100
rect 2548 30044 3612 30100
rect 3668 30044 3678 30100
rect 4498 30044 4508 30100
rect 4564 30044 5964 30100
rect 6020 30044 6030 30100
rect 8642 30044 8652 30100
rect 8708 30044 9660 30100
rect 9716 30044 10444 30100
rect 10500 30044 10510 30100
rect 13794 30044 13804 30100
rect 13860 30044 17724 30100
rect 17780 30044 17790 30100
rect 19282 30044 19292 30100
rect 19348 30044 24052 30100
rect 23996 29988 24052 30044
rect 26852 29988 26908 30156
rect 30818 30044 30828 30100
rect 30884 30044 31836 30100
rect 31892 30044 33068 30100
rect 33124 30044 33134 30100
rect 34150 30044 34188 30100
rect 34244 30044 34254 30100
rect 37426 30044 37436 30100
rect 37492 30044 38108 30100
rect 38164 30044 38174 30100
rect 44370 30044 44380 30100
rect 44436 30044 48188 30100
rect 48244 30044 48254 30100
rect 48738 30044 48748 30100
rect 48804 30044 50540 30100
rect 50596 30044 50606 30100
rect 51202 30044 51212 30100
rect 51268 30044 51996 30100
rect 52052 30044 53004 30100
rect 53060 30044 53070 30100
rect 54114 30044 54124 30100
rect 54180 30044 54796 30100
rect 54852 30044 54862 30100
rect 54124 29988 54180 30044
rect 7970 29932 7980 29988
rect 8036 29932 9772 29988
rect 9828 29932 9838 29988
rect 12002 29932 12012 29988
rect 12068 29932 12572 29988
rect 12628 29932 17612 29988
rect 17668 29932 19516 29988
rect 19572 29932 19582 29988
rect 23986 29932 23996 29988
rect 24052 29932 24892 29988
rect 24948 29932 24958 29988
rect 26852 29932 34860 29988
rect 34916 29932 34926 29988
rect 37986 29932 37996 29988
rect 38052 29932 39452 29988
rect 39508 29932 40012 29988
rect 40068 29932 40078 29988
rect 49746 29932 49756 29988
rect 49812 29932 51436 29988
rect 51492 29932 51502 29988
rect 52434 29932 52444 29988
rect 52500 29932 52780 29988
rect 52836 29932 54180 29988
rect 35410 29820 35420 29876
rect 35476 29820 36092 29876
rect 36148 29820 36158 29876
rect 36390 29820 36428 29876
rect 36484 29820 36494 29876
rect 38098 29820 38108 29876
rect 38164 29820 39004 29876
rect 39060 29820 39070 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 14578 29708 14588 29764
rect 14644 29708 14700 29764
rect 14756 29708 14766 29764
rect 32162 29708 32172 29764
rect 32228 29708 35644 29764
rect 35700 29708 35710 29764
rect 36614 29708 36652 29764
rect 36708 29708 36718 29764
rect 37538 29708 37548 29764
rect 37604 29708 37884 29764
rect 37940 29708 37950 29764
rect 38434 29708 38444 29764
rect 38500 29708 39228 29764
rect 39284 29708 39294 29764
rect 54002 29708 54012 29764
rect 54068 29708 55804 29764
rect 55860 29708 55870 29764
rect 0 29652 800 29680
rect 35644 29652 35700 29708
rect 59200 29652 60000 29680
rect 0 29596 1764 29652
rect 2034 29596 2044 29652
rect 2100 29596 6972 29652
rect 7028 29596 7038 29652
rect 8530 29596 8540 29652
rect 8596 29596 8876 29652
rect 8932 29596 10108 29652
rect 10164 29596 10780 29652
rect 10836 29596 10846 29652
rect 21634 29596 21644 29652
rect 21700 29596 22428 29652
rect 22484 29596 22494 29652
rect 23426 29596 23436 29652
rect 23492 29596 27916 29652
rect 27972 29596 27982 29652
rect 33516 29596 33852 29652
rect 33908 29596 34300 29652
rect 34356 29596 34366 29652
rect 35644 29596 38556 29652
rect 38612 29596 38622 29652
rect 41906 29596 41916 29652
rect 41972 29596 57148 29652
rect 57204 29596 57214 29652
rect 57586 29596 57596 29652
rect 57652 29596 58156 29652
rect 58212 29596 60000 29652
rect 0 29568 800 29596
rect 1708 29428 1764 29596
rect 2706 29484 2716 29540
rect 2772 29484 15148 29540
rect 22306 29484 22316 29540
rect 22372 29484 23324 29540
rect 23380 29484 23390 29540
rect 27234 29484 27244 29540
rect 27300 29484 33292 29540
rect 33348 29484 33358 29540
rect 1698 29372 1708 29428
rect 1764 29372 3164 29428
rect 3220 29372 3230 29428
rect 7858 29372 7868 29428
rect 7924 29372 8092 29428
rect 8148 29372 8988 29428
rect 9044 29372 9054 29428
rect 15092 29316 15148 29484
rect 29474 29372 29484 29428
rect 29540 29372 29932 29428
rect 29988 29372 30940 29428
rect 30996 29372 31006 29428
rect 33516 29316 33572 29596
rect 59200 29568 60000 29596
rect 34402 29484 34412 29540
rect 34468 29484 34524 29540
rect 34580 29484 34590 29540
rect 37100 29484 43708 29540
rect 43764 29484 44156 29540
rect 44212 29484 44222 29540
rect 45938 29484 45948 29540
rect 46004 29484 47180 29540
rect 47236 29484 47246 29540
rect 47842 29484 47852 29540
rect 47908 29484 52556 29540
rect 52612 29484 52622 29540
rect 53778 29484 53788 29540
rect 53844 29484 54684 29540
rect 54740 29484 54750 29540
rect 34402 29372 34412 29428
rect 34468 29372 35196 29428
rect 35252 29372 35262 29428
rect 36278 29372 36316 29428
rect 36372 29372 36382 29428
rect 2370 29260 2380 29316
rect 2436 29260 5068 29316
rect 5124 29260 5134 29316
rect 15092 29260 22036 29316
rect 24882 29260 24892 29316
rect 24948 29260 26908 29316
rect 31042 29260 31052 29316
rect 31108 29260 31836 29316
rect 31892 29260 31902 29316
rect 33282 29260 33292 29316
rect 33348 29260 33572 29316
rect 36418 29260 36428 29316
rect 36484 29260 36876 29316
rect 36932 29260 36942 29316
rect 21980 29204 22036 29260
rect 26852 29204 26908 29260
rect 37100 29204 37156 29484
rect 37538 29372 37548 29428
rect 37604 29372 38780 29428
rect 38836 29372 39452 29428
rect 39508 29372 39518 29428
rect 40674 29372 40684 29428
rect 40740 29372 42700 29428
rect 42756 29372 42766 29428
rect 43362 29372 43372 29428
rect 43428 29372 47404 29428
rect 47460 29372 47470 29428
rect 49970 29372 49980 29428
rect 50036 29372 50876 29428
rect 50932 29372 50942 29428
rect 54114 29372 54124 29428
rect 54180 29372 55020 29428
rect 55076 29372 55086 29428
rect 38546 29260 38556 29316
rect 38612 29260 39004 29316
rect 39060 29260 39070 29316
rect 42466 29260 42476 29316
rect 42532 29260 43260 29316
rect 43316 29260 43326 29316
rect 43810 29260 43820 29316
rect 43876 29260 49084 29316
rect 49140 29260 49150 29316
rect 51986 29260 51996 29316
rect 52052 29260 55244 29316
rect 55300 29260 55310 29316
rect 4498 29148 4508 29204
rect 4564 29148 5740 29204
rect 5796 29148 5806 29204
rect 17826 29148 17836 29204
rect 17892 29148 18620 29204
rect 18676 29148 18686 29204
rect 21970 29148 21980 29204
rect 22036 29148 22046 29204
rect 26852 29148 33404 29204
rect 33460 29148 33852 29204
rect 33908 29148 33918 29204
rect 34076 29148 37156 29204
rect 42578 29148 42588 29204
rect 42644 29148 44940 29204
rect 44996 29148 45006 29204
rect 46694 29148 46732 29204
rect 46788 29148 46798 29204
rect 52882 29148 52892 29204
rect 52948 29148 54684 29204
rect 54740 29148 54750 29204
rect 57810 29148 57820 29204
rect 57876 29148 57886 29204
rect 34076 29092 34132 29148
rect 57820 29092 57876 29148
rect 32946 29036 32956 29092
rect 33012 29036 34132 29092
rect 35746 29036 35756 29092
rect 35812 29036 36652 29092
rect 36708 29036 36718 29092
rect 40786 29036 40796 29092
rect 40852 29036 41468 29092
rect 41524 29036 43092 29092
rect 0 28980 800 29008
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 43036 28980 43092 29036
rect 50372 29036 57876 29092
rect 50372 28980 50428 29036
rect 59200 28980 60000 29008
rect 0 28924 2380 28980
rect 2436 28924 2446 28980
rect 25666 28924 25676 28980
rect 25732 28924 26796 28980
rect 0 28896 800 28924
rect 26852 28868 26908 28980
rect 35970 28924 35980 28980
rect 36036 28924 36428 28980
rect 36484 28924 37324 28980
rect 37380 28924 37390 28980
rect 38612 28924 42476 28980
rect 42532 28924 42542 28980
rect 43026 28924 43036 28980
rect 43092 28924 44268 28980
rect 44324 28924 50428 28980
rect 53890 28924 53900 28980
rect 53956 28924 54684 28980
rect 54740 28924 54750 28980
rect 57474 28924 57484 28980
rect 57540 28924 60000 28980
rect 38612 28868 38668 28924
rect 59200 28896 60000 28924
rect 25218 28812 25228 28868
rect 25284 28812 26684 28868
rect 26740 28812 26750 28868
rect 26852 28812 38668 28868
rect 43922 28812 43932 28868
rect 43988 28812 46172 28868
rect 46228 28812 46238 28868
rect 7746 28700 7756 28756
rect 7812 28700 8092 28756
rect 8148 28700 8158 28756
rect 18498 28700 18508 28756
rect 18564 28700 19292 28756
rect 19348 28700 20188 28756
rect 20244 28700 20254 28756
rect 22194 28700 22204 28756
rect 22260 28700 24668 28756
rect 24724 28700 26348 28756
rect 26404 28700 26414 28756
rect 26562 28700 26572 28756
rect 26628 28700 30828 28756
rect 30884 28700 30894 28756
rect 31826 28700 31836 28756
rect 31892 28700 32396 28756
rect 32452 28700 32462 28756
rect 33394 28700 33404 28756
rect 33460 28700 34412 28756
rect 34468 28700 34478 28756
rect 34822 28700 34860 28756
rect 34916 28700 34926 28756
rect 35308 28700 36428 28756
rect 36484 28700 36494 28756
rect 36726 28700 36764 28756
rect 36820 28700 36830 28756
rect 37426 28700 37436 28756
rect 37492 28700 38668 28756
rect 44370 28700 44380 28756
rect 44436 28700 49868 28756
rect 49924 28700 49934 28756
rect 56130 28700 56140 28756
rect 56196 28700 57820 28756
rect 57876 28700 57886 28756
rect 35308 28644 35364 28700
rect 38612 28644 38668 28700
rect 6962 28588 6972 28644
rect 7028 28588 7420 28644
rect 7476 28588 8204 28644
rect 8260 28588 8270 28644
rect 25890 28588 25900 28644
rect 25956 28588 26460 28644
rect 26516 28588 26526 28644
rect 28354 28588 28364 28644
rect 28420 28588 29596 28644
rect 29652 28588 29662 28644
rect 32050 28588 32060 28644
rect 32116 28588 33292 28644
rect 33348 28588 33358 28644
rect 34066 28588 34076 28644
rect 34132 28588 35364 28644
rect 35522 28588 35532 28644
rect 35588 28588 36316 28644
rect 36372 28588 36382 28644
rect 36530 28588 36540 28644
rect 36596 28588 37548 28644
rect 37604 28588 37614 28644
rect 38612 28588 43260 28644
rect 43316 28588 43596 28644
rect 43652 28588 43662 28644
rect 44146 28588 44156 28644
rect 44212 28588 47404 28644
rect 47460 28588 47470 28644
rect 50418 28588 50428 28644
rect 50484 28588 52892 28644
rect 52948 28588 52958 28644
rect 53330 28588 53340 28644
rect 53396 28588 53788 28644
rect 53844 28588 54124 28644
rect 54180 28588 54190 28644
rect 54684 28588 56364 28644
rect 56420 28588 56430 28644
rect 57138 28588 57148 28644
rect 57204 28588 58156 28644
rect 58212 28588 58222 28644
rect 2482 28476 2492 28532
rect 2548 28476 3612 28532
rect 3668 28476 3678 28532
rect 3938 28476 3948 28532
rect 4004 28476 4844 28532
rect 4900 28476 5628 28532
rect 5684 28476 5694 28532
rect 12786 28476 12796 28532
rect 12852 28476 13580 28532
rect 13636 28476 13646 28532
rect 24210 28476 24220 28532
rect 24276 28476 26012 28532
rect 26068 28476 26078 28532
rect 33618 28476 33628 28532
rect 33684 28476 35084 28532
rect 35140 28476 35150 28532
rect 35746 28476 35756 28532
rect 35812 28476 36204 28532
rect 36260 28476 36540 28532
rect 36596 28476 36606 28532
rect 43698 28476 43708 28532
rect 43764 28476 44604 28532
rect 44660 28476 44670 28532
rect 51426 28476 51436 28532
rect 51492 28476 53004 28532
rect 53060 28476 53070 28532
rect 1698 28364 1708 28420
rect 1764 28364 5068 28420
rect 5124 28364 5134 28420
rect 8642 28364 8652 28420
rect 8708 28364 9996 28420
rect 10052 28364 10062 28420
rect 12562 28364 12572 28420
rect 12628 28364 14028 28420
rect 14084 28364 14094 28420
rect 21970 28364 21980 28420
rect 22036 28364 23996 28420
rect 24052 28364 24062 28420
rect 35858 28364 35868 28420
rect 35924 28364 36316 28420
rect 36372 28364 36382 28420
rect 36614 28364 36652 28420
rect 36708 28364 36718 28420
rect 38434 28364 38444 28420
rect 38500 28364 39004 28420
rect 39060 28364 39070 28420
rect 45266 28364 45276 28420
rect 45332 28364 46396 28420
rect 46452 28364 52780 28420
rect 52836 28364 52846 28420
rect 0 28308 800 28336
rect 1708 28308 1764 28364
rect 54684 28308 54740 28588
rect 55356 28532 55412 28588
rect 55346 28476 55356 28532
rect 55412 28476 55422 28532
rect 59200 28308 60000 28336
rect 0 28252 1764 28308
rect 3490 28252 3500 28308
rect 3556 28252 4620 28308
rect 4676 28252 4686 28308
rect 10994 28252 11004 28308
rect 11060 28252 11564 28308
rect 11620 28252 12684 28308
rect 12740 28252 12750 28308
rect 41234 28252 41244 28308
rect 41300 28252 43484 28308
rect 43540 28252 43550 28308
rect 46834 28252 46844 28308
rect 46900 28252 47180 28308
rect 47236 28252 48076 28308
rect 48132 28252 48142 28308
rect 51202 28252 51212 28308
rect 51268 28252 52668 28308
rect 52724 28252 52734 28308
rect 53106 28252 53116 28308
rect 53172 28252 53900 28308
rect 53956 28252 53966 28308
rect 54674 28252 54684 28308
rect 54740 28252 54750 28308
rect 58146 28252 58156 28308
rect 58212 28252 60000 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 59200 28224 60000 28252
rect 46162 28140 46172 28196
rect 46228 28140 46732 28196
rect 46788 28140 46798 28196
rect 2706 28028 2716 28084
rect 2772 28028 19068 28084
rect 19124 28028 19628 28084
rect 19684 28028 19694 28084
rect 28354 28028 28364 28084
rect 28420 28028 29260 28084
rect 29316 28028 29326 28084
rect 29698 28028 29708 28084
rect 29764 28028 30268 28084
rect 30324 28028 31052 28084
rect 31108 28028 31118 28084
rect 41458 28028 41468 28084
rect 41524 28028 41804 28084
rect 41860 28028 42364 28084
rect 42420 28028 43036 28084
rect 43092 28028 43102 28084
rect 45388 28028 48860 28084
rect 48916 28028 48926 28084
rect 45388 27972 45444 28028
rect 3266 27916 3276 27972
rect 3332 27916 3724 27972
rect 3780 27916 3790 27972
rect 5058 27916 5068 27972
rect 5124 27916 5964 27972
rect 6020 27916 6030 27972
rect 12786 27916 12796 27972
rect 12852 27916 13916 27972
rect 13972 27916 13982 27972
rect 28578 27916 28588 27972
rect 28644 27916 29372 27972
rect 29428 27916 29438 27972
rect 35980 27916 42588 27972
rect 42644 27916 42654 27972
rect 45378 27916 45388 27972
rect 45444 27916 45454 27972
rect 47842 27916 47852 27972
rect 47908 27916 47918 27972
rect 48626 27916 48636 27972
rect 48692 27916 49980 27972
rect 50036 27916 50046 27972
rect 50306 27916 50316 27972
rect 4162 27804 4172 27860
rect 4228 27804 5292 27860
rect 5348 27804 5358 27860
rect 8866 27804 8876 27860
rect 8932 27804 9772 27860
rect 9828 27804 10444 27860
rect 10500 27804 10510 27860
rect 11778 27804 11788 27860
rect 11844 27804 13132 27860
rect 13188 27804 13198 27860
rect 17826 27804 17836 27860
rect 17892 27804 18284 27860
rect 18340 27804 18350 27860
rect 21634 27804 21644 27860
rect 21700 27804 22428 27860
rect 22484 27804 22494 27860
rect 25890 27804 25900 27860
rect 25956 27804 26684 27860
rect 26740 27804 26750 27860
rect 27570 27804 27580 27860
rect 27636 27804 31948 27860
rect 32004 27804 32014 27860
rect 35980 27748 36036 27916
rect 47852 27860 47908 27916
rect 50372 27860 50428 27972
rect 38658 27804 38668 27860
rect 38724 27804 39228 27860
rect 39284 27804 39294 27860
rect 40114 27804 40124 27860
rect 40180 27804 41356 27860
rect 41412 27804 42140 27860
rect 42196 27804 42206 27860
rect 42802 27804 42812 27860
rect 42868 27804 43820 27860
rect 43876 27804 43886 27860
rect 46386 27804 46396 27860
rect 46452 27804 46844 27860
rect 46900 27804 46910 27860
rect 47852 27804 52556 27860
rect 52612 27804 52622 27860
rect 54674 27804 54684 27860
rect 54740 27804 55692 27860
rect 55748 27804 55758 27860
rect 2034 27692 2044 27748
rect 2100 27692 3388 27748
rect 4834 27692 4844 27748
rect 4900 27692 5404 27748
rect 5460 27692 5470 27748
rect 17602 27692 17612 27748
rect 17668 27692 18172 27748
rect 18228 27692 18238 27748
rect 20066 27692 20076 27748
rect 20132 27692 21420 27748
rect 21476 27692 21486 27748
rect 35970 27692 35980 27748
rect 36036 27692 36046 27748
rect 38210 27692 38220 27748
rect 38276 27692 38780 27748
rect 38836 27692 38846 27748
rect 44034 27692 44044 27748
rect 44100 27692 44716 27748
rect 44772 27692 44782 27748
rect 0 27636 800 27664
rect 3332 27636 3388 27692
rect 59200 27636 60000 27664
rect 0 27580 2604 27636
rect 2660 27580 2670 27636
rect 3332 27580 7420 27636
rect 7476 27580 7486 27636
rect 7970 27580 7980 27636
rect 8036 27580 8540 27636
rect 8596 27580 8606 27636
rect 8978 27580 8988 27636
rect 9044 27580 9548 27636
rect 9604 27580 9614 27636
rect 30482 27580 30492 27636
rect 30548 27580 35588 27636
rect 37202 27580 37212 27636
rect 37268 27580 40908 27636
rect 40964 27580 40974 27636
rect 46358 27580 46396 27636
rect 46452 27580 46462 27636
rect 57586 27580 57596 27636
rect 57652 27580 58156 27636
rect 58212 27580 60000 27636
rect 0 27552 800 27580
rect 35532 27524 35588 27580
rect 59200 27552 60000 27580
rect 9212 27468 12740 27524
rect 18274 27468 18284 27524
rect 18340 27468 32060 27524
rect 32116 27468 34748 27524
rect 34804 27468 34814 27524
rect 35532 27468 40236 27524
rect 40292 27468 42588 27524
rect 42644 27468 45388 27524
rect 45444 27468 45454 27524
rect 52210 27468 52220 27524
rect 52276 27468 53004 27524
rect 53060 27468 54012 27524
rect 54068 27468 54078 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 1698 27356 1708 27412
rect 1764 27356 3388 27412
rect 3444 27356 3454 27412
rect 9212 27300 9268 27468
rect 10210 27356 10220 27412
rect 10276 27356 11788 27412
rect 11844 27356 11854 27412
rect 12450 27356 12460 27412
rect 12516 27356 12526 27412
rect 2034 27244 2044 27300
rect 2100 27244 9268 27300
rect 12460 27188 12516 27356
rect 12684 27300 12740 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 14578 27356 14588 27412
rect 14644 27356 15932 27412
rect 15988 27356 22764 27412
rect 22820 27356 30492 27412
rect 30548 27356 30558 27412
rect 35532 27356 56140 27412
rect 56196 27356 56206 27412
rect 35532 27300 35588 27356
rect 12684 27244 19852 27300
rect 19908 27244 19918 27300
rect 26852 27244 33180 27300
rect 33236 27244 33246 27300
rect 33954 27244 33964 27300
rect 34020 27244 34188 27300
rect 34244 27244 35308 27300
rect 35364 27244 35588 27300
rect 36306 27244 36316 27300
rect 36372 27244 37324 27300
rect 37380 27244 37390 27300
rect 38098 27244 38108 27300
rect 38164 27244 57820 27300
rect 57876 27244 57886 27300
rect 26852 27188 26908 27244
rect 2706 27132 2716 27188
rect 2772 27132 3556 27188
rect 3714 27132 3724 27188
rect 3780 27132 4508 27188
rect 4564 27132 4574 27188
rect 4844 27132 12516 27188
rect 13682 27132 13692 27188
rect 13748 27132 14028 27188
rect 14084 27132 18732 27188
rect 18788 27132 18798 27188
rect 18946 27132 18956 27188
rect 19012 27132 26908 27188
rect 31164 27132 32620 27188
rect 32676 27132 33628 27188
rect 33684 27132 33694 27188
rect 34738 27132 34748 27188
rect 34804 27132 38668 27188
rect 39890 27132 39900 27188
rect 39956 27132 44828 27188
rect 44884 27132 44894 27188
rect 45826 27132 45836 27188
rect 45892 27132 52220 27188
rect 52276 27132 52286 27188
rect 52546 27132 52556 27188
rect 52612 27132 54012 27188
rect 54068 27132 54078 27188
rect 55682 27132 55692 27188
rect 55748 27132 58156 27188
rect 58212 27132 58222 27188
rect 3500 27076 3556 27132
rect 4844 27076 4900 27132
rect 3500 27020 4900 27076
rect 5058 27020 5068 27076
rect 5124 27020 6188 27076
rect 6244 27020 6254 27076
rect 0 26964 800 26992
rect 12124 26964 12180 27132
rect 31164 27076 31220 27132
rect 12898 27020 12908 27076
rect 12964 27020 13244 27076
rect 13300 27020 14700 27076
rect 14756 27020 19628 27076
rect 19684 27020 19694 27076
rect 20402 27020 20412 27076
rect 20468 27020 21308 27076
rect 21364 27020 23100 27076
rect 23156 27020 23436 27076
rect 23492 27020 23502 27076
rect 23874 27020 23884 27076
rect 23940 27020 25228 27076
rect 25284 27020 31164 27076
rect 31220 27020 31230 27076
rect 31602 27020 31612 27076
rect 31668 27020 32060 27076
rect 32116 27020 32126 27076
rect 32274 27020 32284 27076
rect 32340 27020 35756 27076
rect 35812 27020 35822 27076
rect 36418 27020 36428 27076
rect 36484 27020 37212 27076
rect 37268 27020 37278 27076
rect 37762 27020 37772 27076
rect 37828 27020 37838 27076
rect 31612 26964 31668 27020
rect 37772 26964 37828 27020
rect 0 26908 1708 26964
rect 1764 26908 1774 26964
rect 2482 26908 2492 26964
rect 2548 26908 5740 26964
rect 5796 26908 5806 26964
rect 7970 26908 7980 26964
rect 8036 26908 8988 26964
rect 9044 26908 9054 26964
rect 12114 26908 12124 26964
rect 12180 26908 12190 26964
rect 20178 26908 20188 26964
rect 20244 26908 21084 26964
rect 21140 26908 21532 26964
rect 21588 26908 21598 26964
rect 28252 26908 30940 26964
rect 30996 26908 31668 26964
rect 31826 26908 31836 26964
rect 31892 26908 32956 26964
rect 33012 26908 33022 26964
rect 33954 26908 33964 26964
rect 34020 26908 34748 26964
rect 34804 26908 36876 26964
rect 36932 26908 36942 26964
rect 37212 26908 37828 26964
rect 38612 26964 38668 27132
rect 40786 27020 40796 27076
rect 40852 27020 41468 27076
rect 41524 27020 41534 27076
rect 43036 27020 44156 27076
rect 44212 27020 44222 27076
rect 51538 27020 51548 27076
rect 51604 27020 51614 27076
rect 51762 27020 51772 27076
rect 51828 27020 52668 27076
rect 52724 27020 52734 27076
rect 43036 26964 43092 27020
rect 51548 26964 51604 27020
rect 59200 26964 60000 26992
rect 38612 26908 43036 26964
rect 43092 26908 43102 26964
rect 43250 26908 43260 26964
rect 43316 26908 44044 26964
rect 44100 26908 44110 26964
rect 51548 26908 52220 26964
rect 52276 26908 52892 26964
rect 52948 26908 52958 26964
rect 58156 26908 60000 26964
rect 0 26880 800 26908
rect 4050 26796 4060 26852
rect 4116 26796 4732 26852
rect 4788 26796 4798 26852
rect 28252 26740 28308 26908
rect 37212 26852 37268 26908
rect 58156 26852 58212 26908
rect 59200 26880 60000 26908
rect 36418 26796 36428 26852
rect 36484 26796 37212 26852
rect 37268 26796 37278 26852
rect 37762 26796 37772 26852
rect 37828 26796 38444 26852
rect 38500 26796 57820 26852
rect 57876 26796 57886 26852
rect 58034 26796 58044 26852
rect 58100 26796 58212 26852
rect 14018 26684 14028 26740
rect 14084 26684 14588 26740
rect 14644 26684 14654 26740
rect 18498 26684 18508 26740
rect 18564 26684 18956 26740
rect 19012 26684 19022 26740
rect 25442 26684 25452 26740
rect 25508 26684 28308 26740
rect 28466 26684 28476 26740
rect 28532 26684 28924 26740
rect 28980 26684 30604 26740
rect 30660 26684 30670 26740
rect 31686 26684 31724 26740
rect 31780 26684 31790 26740
rect 42018 26684 42028 26740
rect 42084 26684 42700 26740
rect 42756 26684 43820 26740
rect 43876 26684 43886 26740
rect 46022 26684 46060 26740
rect 46116 26684 46126 26740
rect 46386 26684 46396 26740
rect 46452 26684 46732 26740
rect 46788 26684 46798 26740
rect 48710 26684 48748 26740
rect 48804 26684 48814 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 3490 26572 3500 26628
rect 3556 26572 3948 26628
rect 4004 26572 4014 26628
rect 14252 26572 15036 26628
rect 15092 26572 15102 26628
rect 2034 26460 2044 26516
rect 2100 26460 9996 26516
rect 10052 26460 11004 26516
rect 11060 26460 11070 26516
rect 924 26348 2492 26404
rect 2548 26348 2558 26404
rect 4498 26348 4508 26404
rect 4564 26348 4844 26404
rect 4900 26348 5964 26404
rect 6020 26348 6030 26404
rect 0 26292 800 26320
rect 924 26292 980 26348
rect 14252 26292 14308 26572
rect 14466 26460 14476 26516
rect 14532 26460 14542 26516
rect 17490 26460 17500 26516
rect 17556 26460 18060 26516
rect 18116 26460 18126 26516
rect 21186 26460 21196 26516
rect 21252 26460 22764 26516
rect 22820 26460 22830 26516
rect 24546 26460 24556 26516
rect 24612 26460 25340 26516
rect 25396 26460 25406 26516
rect 27570 26460 27580 26516
rect 27636 26460 28140 26516
rect 28196 26460 28206 26516
rect 34626 26460 34636 26516
rect 34692 26460 35532 26516
rect 35588 26460 36428 26516
rect 36484 26460 40012 26516
rect 40068 26460 40078 26516
rect 41990 26460 42028 26516
rect 42084 26460 42094 26516
rect 43362 26460 43372 26516
rect 43428 26460 43932 26516
rect 43988 26460 43998 26516
rect 54450 26460 54460 26516
rect 54516 26460 55244 26516
rect 55300 26460 55310 26516
rect 0 26236 980 26292
rect 4050 26236 4060 26292
rect 4116 26236 8428 26292
rect 8484 26236 8494 26292
rect 14242 26236 14252 26292
rect 14308 26236 14318 26292
rect 0 26208 800 26236
rect 2482 26124 2492 26180
rect 2548 26124 3836 26180
rect 3892 26124 3902 26180
rect 4610 26124 4620 26180
rect 4676 26124 5404 26180
rect 5460 26124 5470 26180
rect 7298 26124 7308 26180
rect 7364 26124 9548 26180
rect 9604 26124 9614 26180
rect 14476 26068 14532 26460
rect 18060 26404 18116 26460
rect 18060 26348 22428 26404
rect 22484 26348 24668 26404
rect 24724 26348 24734 26404
rect 37986 26348 37996 26404
rect 38052 26348 38556 26404
rect 38612 26348 38622 26404
rect 42578 26348 42588 26404
rect 42644 26348 43148 26404
rect 43204 26348 44044 26404
rect 44100 26348 44604 26404
rect 44660 26348 44670 26404
rect 50978 26348 50988 26404
rect 51044 26348 51660 26404
rect 51716 26348 51726 26404
rect 52882 26348 52892 26404
rect 52948 26348 53788 26404
rect 53844 26348 53854 26404
rect 59200 26292 60000 26320
rect 16706 26236 16716 26292
rect 16772 26236 17500 26292
rect 17556 26236 17566 26292
rect 21746 26236 21756 26292
rect 21812 26236 25900 26292
rect 25956 26236 25966 26292
rect 27682 26236 27692 26292
rect 27748 26236 29148 26292
rect 29204 26236 31500 26292
rect 31556 26236 31566 26292
rect 40002 26236 40012 26292
rect 40068 26236 42476 26292
rect 42532 26236 42542 26292
rect 47282 26236 47292 26292
rect 47348 26236 47852 26292
rect 47908 26236 47918 26292
rect 50642 26236 50652 26292
rect 50708 26236 50988 26292
rect 51044 26236 52108 26292
rect 52164 26236 52174 26292
rect 57474 26236 57484 26292
rect 57540 26236 60000 26292
rect 59200 26208 60000 26236
rect 23314 26124 23324 26180
rect 23380 26124 24108 26180
rect 24164 26124 24780 26180
rect 24836 26124 24846 26180
rect 30370 26124 30380 26180
rect 30436 26124 33964 26180
rect 34020 26124 34030 26180
rect 47954 26124 47964 26180
rect 48020 26124 50316 26180
rect 50372 26124 50382 26180
rect 52322 26124 52332 26180
rect 52388 26124 53676 26180
rect 53732 26124 53742 26180
rect 55346 26124 55356 26180
rect 55412 26124 56700 26180
rect 56756 26124 56766 26180
rect 3714 26012 3724 26068
rect 3780 26012 6188 26068
rect 6244 26012 6254 26068
rect 10434 26012 10444 26068
rect 10500 26012 11676 26068
rect 11732 26012 11742 26068
rect 14466 26012 14476 26068
rect 14532 26012 14542 26068
rect 22978 26012 22988 26068
rect 23044 26012 23548 26068
rect 23604 26012 35084 26068
rect 35140 26012 35980 26068
rect 36036 26012 36046 26068
rect 50372 26012 57148 26068
rect 57204 26012 57214 26068
rect 50372 25956 50428 26012
rect 20626 25900 20636 25956
rect 20692 25900 21980 25956
rect 22036 25900 33740 25956
rect 33796 25900 34412 25956
rect 34468 25900 34478 25956
rect 39218 25900 39228 25956
rect 39284 25900 40348 25956
rect 40404 25900 41468 25956
rect 41524 25900 50428 25956
rect 56914 25900 56924 25956
rect 56980 25900 58044 25956
rect 58100 25900 58110 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 1586 25788 1596 25844
rect 1652 25788 4340 25844
rect 24546 25788 24556 25844
rect 24612 25788 24892 25844
rect 24948 25788 25452 25844
rect 25508 25788 25518 25844
rect 25890 25788 25900 25844
rect 25956 25788 26236 25844
rect 26292 25788 34188 25844
rect 34244 25788 34254 25844
rect 39106 25788 39116 25844
rect 39172 25788 39340 25844
rect 39396 25788 41132 25844
rect 41188 25788 57036 25844
rect 57092 25788 57102 25844
rect 4284 25732 4340 25788
rect 2258 25676 2268 25732
rect 2324 25676 4060 25732
rect 4116 25676 4126 25732
rect 4284 25676 5852 25732
rect 5908 25676 5918 25732
rect 6178 25676 6188 25732
rect 6244 25676 13916 25732
rect 13972 25676 13982 25732
rect 21746 25676 21756 25732
rect 21812 25676 29708 25732
rect 29764 25676 29774 25732
rect 35746 25676 35756 25732
rect 35812 25676 38780 25732
rect 38836 25676 38846 25732
rect 49634 25676 49644 25732
rect 49700 25676 49710 25732
rect 0 25620 800 25648
rect 49644 25620 49700 25676
rect 59200 25620 60000 25648
rect 0 25564 1708 25620
rect 1764 25564 1774 25620
rect 2594 25564 2604 25620
rect 2660 25564 7980 25620
rect 8036 25564 8046 25620
rect 15026 25564 15036 25620
rect 15092 25564 15484 25620
rect 15540 25564 18396 25620
rect 18452 25564 18462 25620
rect 26236 25564 28476 25620
rect 28532 25564 28542 25620
rect 38612 25564 42252 25620
rect 42308 25564 42318 25620
rect 47730 25564 47740 25620
rect 47796 25564 50876 25620
rect 50932 25564 51716 25620
rect 53778 25564 53788 25620
rect 53844 25564 54796 25620
rect 54852 25564 55468 25620
rect 55524 25564 58156 25620
rect 58212 25564 58222 25620
rect 0 25536 800 25564
rect 1708 25508 1764 25564
rect 26236 25508 26292 25564
rect 38612 25508 38668 25564
rect 51660 25508 51716 25564
rect 59164 25536 60000 25620
rect 1708 25452 7756 25508
rect 7812 25452 7822 25508
rect 9202 25452 9212 25508
rect 9268 25452 17612 25508
rect 17668 25452 17678 25508
rect 19394 25452 19404 25508
rect 19460 25452 20300 25508
rect 20356 25452 20366 25508
rect 22866 25452 22876 25508
rect 22932 25452 26236 25508
rect 26292 25452 26302 25508
rect 26786 25452 26796 25508
rect 26852 25452 28140 25508
rect 28196 25452 28206 25508
rect 35252 25452 38668 25508
rect 39778 25452 39788 25508
rect 39844 25452 40572 25508
rect 40628 25452 40638 25508
rect 49186 25452 49196 25508
rect 49252 25452 50988 25508
rect 51044 25452 51054 25508
rect 51650 25452 51660 25508
rect 51716 25452 51726 25508
rect 35252 25396 35308 25452
rect 59164 25396 59220 25536
rect 2706 25340 2716 25396
rect 2772 25340 3164 25396
rect 3220 25340 4060 25396
rect 4116 25340 4126 25396
rect 19506 25340 19516 25396
rect 19572 25340 21308 25396
rect 21364 25340 21374 25396
rect 26898 25340 26908 25396
rect 26964 25340 27244 25396
rect 27300 25340 27310 25396
rect 27458 25340 27468 25396
rect 27524 25340 27804 25396
rect 27860 25340 35308 25396
rect 38546 25340 38556 25396
rect 38612 25340 40236 25396
rect 40292 25340 40302 25396
rect 50306 25340 50316 25396
rect 50372 25284 50428 25396
rect 50530 25340 50540 25396
rect 50596 25340 52780 25396
rect 52836 25340 52846 25396
rect 59164 25340 59332 25396
rect 1810 25228 1820 25284
rect 1876 25228 4844 25284
rect 4900 25228 5964 25284
rect 6020 25228 8428 25284
rect 13458 25228 13468 25284
rect 13524 25228 14700 25284
rect 14756 25228 14766 25284
rect 15138 25228 15148 25284
rect 15204 25228 17948 25284
rect 18004 25228 19292 25284
rect 19348 25228 19358 25284
rect 19842 25228 19852 25284
rect 19908 25228 22428 25284
rect 22484 25228 22494 25284
rect 26114 25228 26124 25284
rect 26180 25228 27356 25284
rect 27412 25228 27422 25284
rect 29810 25228 29820 25284
rect 29876 25228 34076 25284
rect 34132 25228 34142 25284
rect 37762 25228 37772 25284
rect 37828 25228 38332 25284
rect 38388 25228 39116 25284
rect 39172 25228 39182 25284
rect 48066 25228 48076 25284
rect 48132 25228 49420 25284
rect 49476 25228 49486 25284
rect 50372 25228 51212 25284
rect 51268 25228 53340 25284
rect 53396 25228 53406 25284
rect 8372 25172 8428 25228
rect 59276 25172 59332 25340
rect 3490 25116 3500 25172
rect 3556 25116 3948 25172
rect 4004 25116 5516 25172
rect 5572 25116 5582 25172
rect 5842 25116 5852 25172
rect 5908 25116 6412 25172
rect 6468 25116 6478 25172
rect 8372 25116 9660 25172
rect 9716 25116 10108 25172
rect 10164 25116 11116 25172
rect 11172 25116 11900 25172
rect 11956 25116 11966 25172
rect 14914 25116 14924 25172
rect 14980 25116 15596 25172
rect 15652 25116 15662 25172
rect 26852 25116 34636 25172
rect 34692 25116 34702 25172
rect 45938 25116 45948 25172
rect 46004 25116 47740 25172
rect 47796 25116 47806 25172
rect 50978 25116 50988 25172
rect 51044 25116 51884 25172
rect 51940 25116 55356 25172
rect 55412 25116 55422 25172
rect 57586 25116 57596 25172
rect 57652 25116 58156 25172
rect 58212 25116 59332 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 26852 25060 26908 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 3332 25004 18732 25060
rect 18788 25004 19404 25060
rect 19460 25004 19470 25060
rect 22418 25004 22428 25060
rect 22484 25004 26908 25060
rect 27010 25004 27020 25060
rect 27076 25004 27804 25060
rect 27860 25004 27870 25060
rect 29474 25004 29484 25060
rect 29540 25004 29550 25060
rect 36418 25004 36428 25060
rect 36484 25004 47516 25060
rect 47572 25004 47582 25060
rect 50194 25004 50204 25060
rect 50260 25004 50428 25060
rect 51426 25004 51436 25060
rect 51492 25004 52892 25060
rect 52948 25004 52958 25060
rect 57026 25004 57036 25060
rect 57092 25004 57820 25060
rect 57876 25004 57886 25060
rect 0 24948 800 24976
rect 3332 24948 3388 25004
rect 0 24892 1708 24948
rect 1764 24892 1774 24948
rect 2706 24892 2716 24948
rect 2772 24892 3388 24948
rect 3602 24892 3612 24948
rect 3668 24892 4172 24948
rect 4228 24892 4238 24948
rect 27570 24892 27580 24948
rect 27636 24892 28028 24948
rect 28084 24892 28094 24948
rect 0 24864 800 24892
rect 29484 24836 29540 25004
rect 50372 24948 50428 25004
rect 59200 24948 60000 24976
rect 35074 24892 35084 24948
rect 35140 24892 36092 24948
rect 36148 24892 36158 24948
rect 50372 24892 51156 24948
rect 54674 24892 54684 24948
rect 54740 24892 57484 24948
rect 57540 24892 60000 24948
rect 51100 24836 51156 24892
rect 59200 24864 60000 24892
rect 4722 24780 4732 24836
rect 4788 24780 6188 24836
rect 6244 24780 6254 24836
rect 16594 24780 16604 24836
rect 16660 24780 19068 24836
rect 19124 24780 19134 24836
rect 23986 24780 23996 24836
rect 24052 24780 29540 24836
rect 34738 24780 34748 24836
rect 34804 24780 35420 24836
rect 35476 24780 35486 24836
rect 36418 24780 36428 24836
rect 36484 24780 37660 24836
rect 37716 24780 37726 24836
rect 40348 24780 41020 24836
rect 41076 24780 41086 24836
rect 50194 24780 50204 24836
rect 50260 24780 50876 24836
rect 50932 24780 50942 24836
rect 51090 24780 51100 24836
rect 51156 24780 51166 24836
rect 40348 24724 40404 24780
rect 2370 24668 2380 24724
rect 2436 24668 7308 24724
rect 7364 24668 7374 24724
rect 10546 24668 10556 24724
rect 10612 24668 13692 24724
rect 13748 24668 14364 24724
rect 14420 24668 14430 24724
rect 30258 24668 30268 24724
rect 30324 24668 33068 24724
rect 33124 24668 33134 24724
rect 33506 24668 33516 24724
rect 33572 24668 33964 24724
rect 34020 24668 34030 24724
rect 35746 24668 35756 24724
rect 35812 24668 37884 24724
rect 37940 24668 40348 24724
rect 40404 24668 40414 24724
rect 40898 24668 40908 24724
rect 40964 24668 42924 24724
rect 42980 24668 42990 24724
rect 44482 24668 44492 24724
rect 44548 24668 50988 24724
rect 51044 24668 51054 24724
rect 52770 24668 52780 24724
rect 52836 24668 53004 24724
rect 53060 24668 53676 24724
rect 53732 24668 53742 24724
rect 5394 24556 5404 24612
rect 5460 24556 7084 24612
rect 7140 24556 7150 24612
rect 12226 24556 12236 24612
rect 12292 24556 14812 24612
rect 14868 24556 14878 24612
rect 24770 24556 24780 24612
rect 24836 24556 25452 24612
rect 25508 24556 25518 24612
rect 28690 24556 28700 24612
rect 28756 24556 29820 24612
rect 29876 24556 29886 24612
rect 32620 24556 40684 24612
rect 40740 24556 40750 24612
rect 44594 24556 44604 24612
rect 44660 24556 52332 24612
rect 52388 24556 52398 24612
rect 55234 24556 55244 24612
rect 55300 24556 56028 24612
rect 56084 24556 56094 24612
rect 5730 24444 5740 24500
rect 5796 24444 6300 24500
rect 6356 24444 6366 24500
rect 12450 24332 12460 24388
rect 12516 24332 13132 24388
rect 13188 24332 13198 24388
rect 13906 24332 13916 24388
rect 13972 24332 14700 24388
rect 14756 24332 14766 24388
rect 20290 24332 20300 24388
rect 20356 24332 20860 24388
rect 20916 24332 20926 24388
rect 26226 24332 26236 24388
rect 26292 24332 29372 24388
rect 29428 24332 29438 24388
rect 0 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 0 24220 2380 24276
rect 2436 24220 2446 24276
rect 25890 24220 25900 24276
rect 25956 24220 32284 24276
rect 32340 24220 32350 24276
rect 0 24192 800 24220
rect 32620 24164 32676 24556
rect 38434 24444 38444 24500
rect 38500 24444 39788 24500
rect 39844 24444 39854 24500
rect 40562 24444 40572 24500
rect 40628 24444 41916 24500
rect 41972 24444 43148 24500
rect 43204 24444 57148 24500
rect 57204 24444 57214 24500
rect 36978 24332 36988 24388
rect 37044 24332 39564 24388
rect 39620 24332 39630 24388
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 59200 24276 60000 24304
rect 58146 24220 58156 24276
rect 58212 24220 60000 24276
rect 59200 24192 60000 24220
rect 18946 24108 18956 24164
rect 19012 24108 19516 24164
rect 19572 24108 32676 24164
rect 44370 24108 44380 24164
rect 44436 24108 45276 24164
rect 45332 24108 45342 24164
rect 48626 24108 48636 24164
rect 48692 24108 50092 24164
rect 50148 24108 50158 24164
rect 50642 24108 50652 24164
rect 50708 24108 51884 24164
rect 51940 24108 53116 24164
rect 53172 24108 53788 24164
rect 53844 24108 53854 24164
rect 1698 23996 1708 24052
rect 1764 23996 5068 24052
rect 5124 23996 5134 24052
rect 6626 23996 6636 24052
rect 6692 23996 9548 24052
rect 9604 23996 12908 24052
rect 12964 23996 12974 24052
rect 16482 23996 16492 24052
rect 16548 23996 17724 24052
rect 17780 23996 17790 24052
rect 19954 23996 19964 24052
rect 20020 23996 20188 24052
rect 20244 23996 30604 24052
rect 30660 23996 31276 24052
rect 31332 23996 31342 24052
rect 40338 23996 40348 24052
rect 40404 23996 42140 24052
rect 42196 23996 42206 24052
rect 55234 23996 55244 24052
rect 55300 23996 57932 24052
rect 57988 23996 57998 24052
rect 21522 23884 21532 23940
rect 21588 23884 22204 23940
rect 22260 23884 22270 23940
rect 25666 23884 25676 23940
rect 25732 23884 26460 23940
rect 26516 23884 27356 23940
rect 27412 23884 27422 23940
rect 27570 23884 27580 23940
rect 27636 23884 27674 23940
rect 37986 23884 37996 23940
rect 38052 23884 39116 23940
rect 39172 23884 41468 23940
rect 41524 23884 41534 23940
rect 46498 23884 46508 23940
rect 46564 23884 47404 23940
rect 47460 23884 48524 23940
rect 48580 23884 49140 23940
rect 50866 23884 50876 23940
rect 50932 23884 50988 23940
rect 51044 23884 51054 23940
rect 3714 23772 3724 23828
rect 3780 23772 5292 23828
rect 5348 23772 5358 23828
rect 5730 23772 5740 23828
rect 5796 23772 6636 23828
rect 6692 23772 7028 23828
rect 19058 23772 19068 23828
rect 19124 23772 21308 23828
rect 21364 23772 21374 23828
rect 39554 23772 39564 23828
rect 39620 23772 41804 23828
rect 41860 23772 41870 23828
rect 46946 23772 46956 23828
rect 47012 23772 47628 23828
rect 47684 23772 47694 23828
rect 6972 23716 7028 23772
rect 49084 23716 49140 23884
rect 51202 23772 51212 23828
rect 51268 23772 52444 23828
rect 52500 23772 52510 23828
rect 3938 23660 3948 23716
rect 4004 23660 4844 23716
rect 4900 23660 5964 23716
rect 6020 23660 6030 23716
rect 6962 23660 6972 23716
rect 7028 23660 9884 23716
rect 9940 23660 9950 23716
rect 32834 23660 32844 23716
rect 32900 23660 34748 23716
rect 34804 23660 34814 23716
rect 38770 23660 38780 23716
rect 38836 23660 43484 23716
rect 43540 23660 43550 23716
rect 49074 23660 49084 23716
rect 49140 23660 49150 23716
rect 59200 23604 60000 23632
rect 5730 23548 5740 23604
rect 5796 23548 6300 23604
rect 6356 23548 9212 23604
rect 9268 23548 12572 23604
rect 12628 23548 12638 23604
rect 36978 23548 36988 23604
rect 37044 23548 37996 23604
rect 38052 23548 38062 23604
rect 42242 23548 42252 23604
rect 42308 23548 42318 23604
rect 43148 23548 43820 23604
rect 43876 23548 43886 23604
rect 57484 23548 60000 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 42252 23492 42308 23548
rect 43148 23492 43204 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 57484 23492 57540 23548
rect 59200 23520 60000 23548
rect 9426 23436 9436 23492
rect 9492 23436 9884 23492
rect 9940 23436 9950 23492
rect 11526 23436 11564 23492
rect 11620 23436 11630 23492
rect 32050 23436 32060 23492
rect 32116 23436 33180 23492
rect 33236 23436 35476 23492
rect 37314 23436 37324 23492
rect 37380 23436 38220 23492
rect 38276 23436 38556 23492
rect 38612 23436 38622 23492
rect 42252 23436 42812 23492
rect 42868 23436 42878 23492
rect 43138 23436 43148 23492
rect 43204 23436 43214 23492
rect 45042 23436 45052 23492
rect 45108 23436 46620 23492
rect 46676 23436 46686 23492
rect 57474 23436 57484 23492
rect 57540 23436 57550 23492
rect 35420 23380 35476 23436
rect 4834 23324 4844 23380
rect 4900 23324 8764 23380
rect 8820 23324 8830 23380
rect 9874 23324 9884 23380
rect 9940 23324 9950 23380
rect 11778 23324 11788 23380
rect 11844 23324 11882 23380
rect 12002 23324 12012 23380
rect 12068 23324 13804 23380
rect 13860 23324 14812 23380
rect 14868 23324 14878 23380
rect 16818 23324 16828 23380
rect 16884 23324 17388 23380
rect 17444 23324 18060 23380
rect 18116 23324 18126 23380
rect 33618 23324 33628 23380
rect 33684 23324 34972 23380
rect 35028 23324 35038 23380
rect 35420 23324 37772 23380
rect 37828 23324 37838 23380
rect 38098 23324 38108 23380
rect 38164 23324 38668 23380
rect 42354 23324 42364 23380
rect 42420 23324 43484 23380
rect 43540 23324 57820 23380
rect 57876 23324 57886 23380
rect 9884 23268 9940 23324
rect 7410 23212 7420 23268
rect 7476 23212 9660 23268
rect 9716 23212 9726 23268
rect 9884 23212 16492 23268
rect 16548 23212 16558 23268
rect 21970 23212 21980 23268
rect 22036 23212 26908 23268
rect 26964 23212 27580 23268
rect 27636 23212 27646 23268
rect 29026 23212 29036 23268
rect 29092 23212 30492 23268
rect 30548 23212 30940 23268
rect 30996 23212 31006 23268
rect 31350 23212 31388 23268
rect 31444 23212 31454 23268
rect 32498 23212 32508 23268
rect 32564 23212 33348 23268
rect 33842 23212 33852 23268
rect 33908 23212 35196 23268
rect 35252 23212 35262 23268
rect 33292 23156 33348 23212
rect 38612 23156 38668 23324
rect 43698 23212 43708 23268
rect 43764 23212 48748 23268
rect 48804 23212 48814 23268
rect 50418 23212 50428 23268
rect 50484 23212 52220 23268
rect 52276 23212 52286 23268
rect 53554 23212 53564 23268
rect 53620 23212 54796 23268
rect 54852 23212 55580 23268
rect 55636 23212 57932 23268
rect 57988 23212 57998 23268
rect 2930 23100 2940 23156
rect 2996 23100 6300 23156
rect 6356 23100 6366 23156
rect 8866 23100 8876 23156
rect 8932 23100 9996 23156
rect 10052 23100 10062 23156
rect 12348 23100 12796 23156
rect 12852 23100 12862 23156
rect 27682 23100 27692 23156
rect 27748 23100 30044 23156
rect 30100 23100 31052 23156
rect 31108 23100 31118 23156
rect 31490 23100 31500 23156
rect 31556 23100 33068 23156
rect 33124 23100 33134 23156
rect 33292 23100 34076 23156
rect 34132 23100 34636 23156
rect 34692 23100 34702 23156
rect 38612 23100 38892 23156
rect 38948 23100 38958 23156
rect 39330 23100 39340 23156
rect 39396 23100 40236 23156
rect 40292 23100 40908 23156
rect 40964 23100 40974 23156
rect 43362 23100 43372 23156
rect 43428 23100 45276 23156
rect 45332 23100 45342 23156
rect 46610 23100 46620 23156
rect 46676 23100 47516 23156
rect 47572 23100 47582 23156
rect 48066 23100 48076 23156
rect 48132 23100 49420 23156
rect 49476 23100 50988 23156
rect 51044 23100 51054 23156
rect 12348 23044 12404 23100
rect 3602 22988 3612 23044
rect 3668 22988 4620 23044
rect 4676 22988 5292 23044
rect 5348 22988 6636 23044
rect 6692 22988 6702 23044
rect 11890 22988 11900 23044
rect 11956 22988 12404 23044
rect 12674 22988 12684 23044
rect 12740 22988 13132 23044
rect 13188 22988 18956 23044
rect 19012 22988 19022 23044
rect 19842 22988 19852 23044
rect 19908 22988 20636 23044
rect 20692 22988 20702 23044
rect 21858 22988 21868 23044
rect 21924 22988 22428 23044
rect 22484 22988 22494 23044
rect 23874 22988 23884 23044
rect 23940 22988 24780 23044
rect 24836 22988 24846 23044
rect 28802 22988 28812 23044
rect 28868 22988 29148 23044
rect 29204 22988 29596 23044
rect 29652 22988 29662 23044
rect 31686 22988 31724 23044
rect 31780 22988 31790 23044
rect 33954 22988 33964 23044
rect 34020 22988 34524 23044
rect 34580 22988 34590 23044
rect 34962 22988 34972 23044
rect 35028 22988 35756 23044
rect 35812 22988 35822 23044
rect 39106 22988 39116 23044
rect 39172 22988 42756 23044
rect 42914 22988 42924 23044
rect 42980 22988 43932 23044
rect 43988 22988 44380 23044
rect 44436 22988 44446 23044
rect 44716 22988 47068 23044
rect 47124 22988 47852 23044
rect 47908 22988 47918 23044
rect 55458 22988 55468 23044
rect 55524 22988 56700 23044
rect 56756 22988 56766 23044
rect 0 22932 800 22960
rect 23884 22932 23940 22988
rect 42700 22932 42756 22988
rect 44716 22932 44772 22988
rect 59200 22932 60000 22960
rect 0 22876 1708 22932
rect 1764 22876 1774 22932
rect 10546 22876 10556 22932
rect 10612 22876 23940 22932
rect 29026 22876 29036 22932
rect 29092 22876 29820 22932
rect 29876 22876 29886 22932
rect 32050 22876 32060 22932
rect 32116 22876 32956 22932
rect 33012 22876 33022 22932
rect 34374 22876 34412 22932
rect 34468 22876 34478 22932
rect 34962 22876 34972 22932
rect 35028 22876 37100 22932
rect 37156 22876 37166 22932
rect 37538 22876 37548 22932
rect 37604 22876 38668 22932
rect 39218 22876 39228 22932
rect 39284 22876 42476 22932
rect 42532 22876 42542 22932
rect 42700 22876 44772 22932
rect 44930 22876 44940 22932
rect 44996 22876 45500 22932
rect 45556 22876 45566 22932
rect 59052 22876 60000 22932
rect 0 22848 800 22876
rect 11526 22764 11564 22820
rect 11620 22764 11630 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 38612 22708 38668 22876
rect 40450 22764 40460 22820
rect 40516 22764 41468 22820
rect 41524 22764 57148 22820
rect 57204 22764 57214 22820
rect 59052 22708 59108 22876
rect 59200 22848 60000 22876
rect 26852 22652 28364 22708
rect 28420 22652 29372 22708
rect 29428 22652 30884 22708
rect 34066 22652 34076 22708
rect 34132 22652 34524 22708
rect 34580 22652 34590 22708
rect 38612 22652 41748 22708
rect 50866 22652 50876 22708
rect 50932 22652 52780 22708
rect 52836 22652 52846 22708
rect 59052 22652 59332 22708
rect 11554 22540 11564 22596
rect 11620 22540 13468 22596
rect 13524 22540 13534 22596
rect 1698 22428 1708 22484
rect 1764 22428 6188 22484
rect 6244 22428 6254 22484
rect 9426 22428 9436 22484
rect 9492 22428 9996 22484
rect 10052 22428 10556 22484
rect 10612 22428 10622 22484
rect 11330 22428 11340 22484
rect 11396 22428 12012 22484
rect 12068 22428 12078 22484
rect 17938 22428 17948 22484
rect 18004 22428 19180 22484
rect 19236 22428 21868 22484
rect 21924 22428 21934 22484
rect 7522 22316 7532 22372
rect 7588 22316 13468 22372
rect 13524 22316 13534 22372
rect 0 22260 800 22288
rect 0 22204 1708 22260
rect 1764 22204 1774 22260
rect 6626 22204 6636 22260
rect 6692 22204 7868 22260
rect 7924 22204 7934 22260
rect 9212 22204 15260 22260
rect 15316 22204 15326 22260
rect 0 22176 800 22204
rect 9212 22036 9268 22204
rect 14690 22092 14700 22148
rect 14756 22092 15148 22148
rect 15204 22092 15214 22148
rect 18284 22036 18340 22428
rect 26852 22260 26908 22652
rect 28130 22540 28140 22596
rect 28196 22540 29708 22596
rect 29764 22540 30044 22596
rect 30100 22540 30110 22596
rect 30828 22484 30884 22652
rect 41692 22596 41748 22652
rect 33394 22540 33404 22596
rect 33460 22540 33852 22596
rect 33908 22540 33918 22596
rect 34738 22540 34748 22596
rect 34804 22540 35868 22596
rect 35924 22540 35934 22596
rect 38098 22540 38108 22596
rect 38164 22540 39116 22596
rect 39172 22540 39182 22596
rect 39442 22540 39452 22596
rect 39508 22540 39518 22596
rect 41682 22540 41692 22596
rect 41748 22540 41758 22596
rect 50082 22540 50092 22596
rect 50148 22540 50988 22596
rect 51044 22540 51054 22596
rect 39452 22484 39508 22540
rect 30828 22428 38668 22484
rect 38612 22372 38668 22428
rect 39452 22428 40236 22484
rect 40292 22428 40684 22484
rect 40740 22428 40750 22484
rect 41234 22428 41244 22484
rect 41300 22428 41916 22484
rect 41972 22428 57036 22484
rect 57092 22428 57102 22484
rect 39452 22372 39508 22428
rect 30930 22316 30940 22372
rect 30996 22316 31500 22372
rect 31556 22316 31566 22372
rect 31826 22316 31836 22372
rect 31892 22316 32396 22372
rect 32452 22316 32462 22372
rect 33618 22316 33628 22372
rect 33684 22316 36204 22372
rect 36260 22316 36270 22372
rect 38612 22316 39508 22372
rect 42018 22316 42028 22372
rect 42084 22316 43036 22372
rect 43092 22316 46284 22372
rect 46340 22316 46350 22372
rect 59276 22260 59332 22652
rect 18722 22204 18732 22260
rect 18788 22204 26908 22260
rect 28578 22204 28588 22260
rect 28644 22204 30492 22260
rect 30548 22204 30558 22260
rect 32274 22204 32284 22260
rect 32340 22204 32956 22260
rect 33012 22204 33022 22260
rect 34290 22204 34300 22260
rect 34356 22204 35756 22260
rect 35812 22204 35822 22260
rect 36428 22204 38892 22260
rect 38948 22204 39564 22260
rect 39620 22204 39630 22260
rect 39778 22204 39788 22260
rect 39844 22204 40236 22260
rect 40292 22204 40302 22260
rect 41794 22204 41804 22260
rect 41860 22204 43148 22260
rect 43204 22204 43596 22260
rect 43652 22204 43662 22260
rect 51762 22204 51772 22260
rect 51828 22204 52892 22260
rect 52948 22204 52958 22260
rect 58146 22204 58156 22260
rect 58212 22204 59332 22260
rect 28018 22092 28028 22148
rect 28084 22092 29148 22148
rect 29204 22092 29214 22148
rect 29586 22092 29596 22148
rect 29652 22092 30716 22148
rect 30772 22092 30782 22148
rect 31826 22092 31836 22148
rect 31892 22092 32620 22148
rect 32676 22092 32686 22148
rect 33618 22092 33628 22148
rect 33684 22092 34076 22148
rect 34132 22092 34142 22148
rect 34402 22092 34412 22148
rect 34468 22092 34860 22148
rect 34916 22092 35532 22148
rect 35588 22092 35598 22148
rect 36428 22036 36484 22204
rect 37314 22092 37324 22148
rect 37380 22092 38220 22148
rect 38276 22092 38286 22148
rect 42130 22092 42140 22148
rect 42196 22092 42364 22148
rect 42420 22092 44044 22148
rect 44100 22092 44110 22148
rect 53778 22092 53788 22148
rect 53844 22092 55244 22148
rect 55300 22092 55310 22148
rect 2930 21980 2940 22036
rect 2996 21980 9268 22036
rect 9426 21980 9436 22036
rect 9492 21980 9502 22036
rect 18274 21980 18284 22036
rect 18340 21980 18350 22036
rect 20962 21980 20972 22036
rect 21028 21980 21980 22036
rect 22036 21980 22046 22036
rect 32386 21980 32396 22036
rect 32452 21980 35868 22036
rect 35924 21980 36484 22036
rect 37874 21980 37884 22036
rect 37940 21980 38556 22036
rect 38612 21980 38622 22036
rect 42578 21980 42588 22036
rect 42644 21980 45052 22036
rect 45108 21980 45118 22036
rect 53442 21980 53452 22036
rect 53508 21980 54124 22036
rect 54180 21980 54190 22036
rect 9436 21924 9492 21980
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 7298 21868 7308 21924
rect 7364 21868 8316 21924
rect 8372 21868 9492 21924
rect 12338 21868 12348 21924
rect 12404 21868 13020 21924
rect 13076 21868 13086 21924
rect 13458 21868 13468 21924
rect 13524 21868 14252 21924
rect 14308 21868 16156 21924
rect 16212 21868 17500 21924
rect 17556 21868 17566 21924
rect 23436 21868 25340 21924
rect 25396 21868 28252 21924
rect 28308 21868 31052 21924
rect 31108 21868 31118 21924
rect 33170 21868 33180 21924
rect 33236 21868 33964 21924
rect 34020 21868 34412 21924
rect 34468 21868 34478 21924
rect 34860 21868 36316 21924
rect 36372 21868 36382 21924
rect 40674 21868 40684 21924
rect 40740 21868 42924 21924
rect 42980 21868 42990 21924
rect 49186 21868 49196 21924
rect 49252 21868 50092 21924
rect 50148 21868 50158 21924
rect 1698 21756 1708 21812
rect 1764 21756 1774 21812
rect 2482 21756 2492 21812
rect 2548 21756 3836 21812
rect 3892 21756 3902 21812
rect 12674 21756 12684 21812
rect 12740 21756 13356 21812
rect 13412 21756 13692 21812
rect 13748 21756 13758 21812
rect 14252 21756 16604 21812
rect 16660 21756 16670 21812
rect 17602 21756 17612 21812
rect 17668 21756 19180 21812
rect 19236 21756 19246 21812
rect 21186 21756 21196 21812
rect 21252 21756 21756 21812
rect 21812 21756 21822 21812
rect 1708 21700 1764 21756
rect 1708 21644 5740 21700
rect 5796 21644 5806 21700
rect 0 21588 800 21616
rect 14252 21588 14308 21756
rect 23436 21700 23492 21868
rect 34860 21812 34916 21868
rect 26002 21756 26012 21812
rect 26068 21756 26572 21812
rect 26628 21756 26638 21812
rect 29138 21756 29148 21812
rect 29204 21756 31500 21812
rect 31556 21756 31566 21812
rect 31714 21756 31724 21812
rect 31780 21756 32172 21812
rect 32228 21756 32238 21812
rect 34850 21756 34860 21812
rect 34916 21756 34926 21812
rect 40002 21756 40012 21812
rect 40068 21756 41020 21812
rect 41076 21756 41086 21812
rect 48178 21756 48188 21812
rect 48244 21756 49532 21812
rect 49588 21756 51100 21812
rect 51156 21756 51166 21812
rect 51650 21756 51660 21812
rect 51716 21756 52892 21812
rect 52948 21756 52958 21812
rect 53666 21756 53676 21812
rect 53732 21756 54908 21812
rect 54964 21756 55356 21812
rect 55412 21756 56812 21812
rect 56868 21756 56878 21812
rect 57026 21756 57036 21812
rect 57092 21756 57820 21812
rect 57876 21756 57886 21812
rect 16706 21644 16716 21700
rect 16772 21644 17500 21700
rect 17556 21644 17566 21700
rect 21410 21644 21420 21700
rect 21476 21644 22092 21700
rect 22148 21644 23492 21700
rect 26898 21644 26908 21700
rect 26964 21644 28476 21700
rect 28532 21644 30828 21700
rect 30884 21644 30894 21700
rect 33730 21644 33740 21700
rect 33796 21644 34300 21700
rect 34356 21644 34366 21700
rect 39890 21644 39900 21700
rect 39956 21644 41468 21700
rect 41524 21644 41534 21700
rect 48850 21644 48860 21700
rect 48916 21644 50036 21700
rect 50194 21644 50204 21700
rect 50260 21644 50540 21700
rect 50596 21644 50606 21700
rect 51986 21644 51996 21700
rect 52052 21644 52444 21700
rect 52500 21644 53116 21700
rect 53172 21644 53182 21700
rect 0 21532 2604 21588
rect 2660 21532 5292 21588
rect 5348 21532 5358 21588
rect 8530 21532 8540 21588
rect 8596 21532 9436 21588
rect 9492 21532 9502 21588
rect 14242 21532 14252 21588
rect 14308 21532 14318 21588
rect 14914 21532 14924 21588
rect 14980 21532 17388 21588
rect 17444 21532 17454 21588
rect 18834 21532 18844 21588
rect 18900 21532 28028 21588
rect 28084 21532 28094 21588
rect 28354 21532 28364 21588
rect 28420 21532 29484 21588
rect 29540 21532 29550 21588
rect 38098 21532 38108 21588
rect 38164 21532 38892 21588
rect 38948 21532 39788 21588
rect 39844 21532 39854 21588
rect 0 21504 800 21532
rect 49980 21476 50036 21644
rect 50418 21532 50428 21588
rect 50484 21532 51548 21588
rect 51604 21532 51614 21588
rect 54002 21532 54012 21588
rect 54068 21532 55132 21588
rect 55188 21532 55198 21588
rect 2258 21420 2268 21476
rect 2324 21420 8092 21476
rect 8148 21420 10780 21476
rect 10836 21420 10846 21476
rect 13682 21420 13692 21476
rect 13748 21420 14588 21476
rect 14644 21420 14654 21476
rect 15138 21420 15148 21476
rect 15204 21420 24500 21476
rect 24658 21420 24668 21476
rect 24724 21420 26012 21476
rect 26068 21420 26078 21476
rect 26226 21420 26236 21476
rect 26292 21420 26684 21476
rect 26740 21420 28476 21476
rect 28532 21420 28542 21476
rect 31378 21420 31388 21476
rect 31444 21420 31500 21476
rect 31556 21420 31566 21476
rect 35858 21420 35868 21476
rect 35924 21420 36764 21476
rect 36820 21420 36830 21476
rect 37650 21420 37660 21476
rect 37716 21420 38668 21476
rect 38724 21420 39004 21476
rect 39060 21420 39070 21476
rect 41906 21420 41916 21476
rect 41972 21420 42700 21476
rect 42756 21420 42766 21476
rect 49980 21420 52108 21476
rect 52164 21420 52174 21476
rect 55010 21420 55020 21476
rect 55076 21420 55692 21476
rect 55748 21420 55758 21476
rect 24444 21364 24500 21420
rect 3266 21308 3276 21364
rect 3332 21308 6300 21364
rect 6356 21308 6366 21364
rect 9398 21308 9436 21364
rect 9492 21308 9502 21364
rect 15922 21308 15932 21364
rect 15988 21308 18172 21364
rect 18228 21308 18238 21364
rect 24444 21308 25564 21364
rect 25620 21308 25630 21364
rect 30482 21308 30492 21364
rect 30548 21308 32284 21364
rect 32340 21308 32350 21364
rect 35298 21308 35308 21364
rect 35364 21308 36204 21364
rect 36260 21308 38668 21364
rect 38612 21252 38668 21308
rect 3714 21196 3724 21252
rect 3780 21196 4172 21252
rect 4228 21196 4238 21252
rect 16594 21196 16604 21252
rect 16660 21196 18508 21252
rect 18564 21196 18574 21252
rect 28018 21196 28028 21252
rect 28084 21196 30716 21252
rect 30772 21196 34412 21252
rect 34468 21196 34478 21252
rect 38612 21196 48972 21252
rect 49028 21196 49038 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 26982 21084 27020 21140
rect 27076 21084 27086 21140
rect 2370 20972 2380 21028
rect 2436 20972 7980 21028
rect 8036 20972 8204 21028
rect 8260 20972 8876 21028
rect 8932 20972 8942 21028
rect 37650 20972 37660 21028
rect 37716 20972 38332 21028
rect 38388 20972 38398 21028
rect 41346 20972 41356 21028
rect 41412 20972 45836 21028
rect 45892 20972 45902 21028
rect 51538 20972 51548 21028
rect 51604 20972 52668 21028
rect 52724 20972 52734 21028
rect 0 20916 800 20944
rect 0 20860 1708 20916
rect 1764 20860 1774 20916
rect 2258 20860 2268 20916
rect 2324 20860 7308 20916
rect 7364 20860 7374 20916
rect 21858 20860 21868 20916
rect 21924 20860 23436 20916
rect 23492 20860 23884 20916
rect 23940 20860 24668 20916
rect 24724 20860 25340 20916
rect 25396 20860 25406 20916
rect 28466 20860 28476 20916
rect 28532 20860 31052 20916
rect 31108 20860 31118 20916
rect 31378 20860 31388 20916
rect 31444 20860 33180 20916
rect 33236 20860 33246 20916
rect 40338 20860 40348 20916
rect 40404 20860 50204 20916
rect 50260 20860 50270 20916
rect 52210 20860 52220 20916
rect 52276 20860 53228 20916
rect 53284 20860 54012 20916
rect 54068 20860 54078 20916
rect 0 20832 800 20860
rect 2930 20748 2940 20804
rect 2996 20748 3388 20804
rect 3826 20748 3836 20804
rect 3892 20748 4172 20804
rect 4228 20748 4238 20804
rect 4834 20748 4844 20804
rect 4900 20748 5964 20804
rect 6020 20748 6030 20804
rect 7410 20748 7420 20804
rect 7476 20748 8652 20804
rect 8708 20748 8718 20804
rect 17714 20748 17724 20804
rect 17780 20748 18508 20804
rect 18564 20748 18574 20804
rect 18834 20748 18844 20804
rect 18900 20748 19404 20804
rect 19460 20748 19964 20804
rect 20020 20748 20030 20804
rect 20850 20748 20860 20804
rect 20916 20748 21980 20804
rect 22036 20748 22428 20804
rect 22484 20748 22494 20804
rect 28130 20748 28140 20804
rect 28196 20748 30044 20804
rect 30100 20748 30110 20804
rect 33954 20748 33964 20804
rect 34020 20748 34412 20804
rect 34468 20748 34478 20804
rect 36082 20748 36092 20804
rect 36148 20748 37436 20804
rect 37492 20748 37502 20804
rect 40450 20748 40460 20804
rect 40516 20748 41804 20804
rect 41860 20748 41870 20804
rect 44258 20748 44268 20804
rect 44324 20748 45612 20804
rect 45668 20748 46284 20804
rect 46340 20748 46350 20804
rect 46582 20748 46620 20804
rect 46676 20748 46686 20804
rect 51538 20748 51548 20804
rect 51604 20748 52108 20804
rect 52164 20748 52444 20804
rect 52500 20748 52510 20804
rect 3332 20692 3388 20748
rect 3332 20636 8876 20692
rect 8932 20636 10108 20692
rect 10164 20636 10174 20692
rect 2482 20524 2492 20580
rect 2548 20524 3500 20580
rect 3556 20524 3566 20580
rect 7298 20524 7308 20580
rect 7364 20524 8540 20580
rect 8596 20524 12012 20580
rect 12068 20524 12078 20580
rect 19628 20468 19684 20748
rect 20738 20636 20748 20692
rect 20804 20636 21756 20692
rect 21812 20636 22316 20692
rect 22372 20636 22382 20692
rect 24546 20636 24556 20692
rect 24612 20636 29932 20692
rect 29988 20636 29998 20692
rect 39330 20636 39340 20692
rect 39396 20636 40908 20692
rect 40964 20636 40974 20692
rect 45490 20636 45500 20692
rect 45556 20636 47068 20692
rect 47124 20636 47134 20692
rect 26674 20524 26684 20580
rect 26740 20524 28364 20580
rect 28420 20524 28430 20580
rect 28578 20524 28588 20580
rect 28644 20524 29484 20580
rect 29540 20524 29550 20580
rect 29810 20524 29820 20580
rect 29876 20524 31164 20580
rect 31220 20524 31230 20580
rect 33058 20524 33068 20580
rect 33124 20524 34748 20580
rect 34804 20524 34814 20580
rect 35186 20524 35196 20580
rect 35252 20524 35868 20580
rect 35924 20524 35934 20580
rect 38612 20524 39116 20580
rect 39172 20524 39182 20580
rect 40562 20524 40572 20580
rect 40628 20524 41020 20580
rect 41076 20524 41086 20580
rect 46386 20524 46396 20580
rect 46452 20524 47852 20580
rect 47908 20524 51996 20580
rect 52052 20524 52062 20580
rect 38612 20468 38668 20524
rect 19618 20412 19628 20468
rect 19684 20412 19694 20468
rect 26852 20412 31500 20468
rect 31556 20412 31566 20468
rect 36530 20412 36540 20468
rect 36596 20412 38668 20468
rect 38994 20412 39004 20468
rect 39060 20412 39340 20468
rect 39396 20412 39406 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 26852 20356 26908 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 1484 20300 2716 20356
rect 2772 20300 2782 20356
rect 6290 20300 6300 20356
rect 6356 20300 6366 20356
rect 7522 20300 7532 20356
rect 7588 20300 7644 20356
rect 7700 20300 9660 20356
rect 9716 20300 9726 20356
rect 16118 20300 16156 20356
rect 16212 20300 16222 20356
rect 20514 20300 20524 20356
rect 20580 20300 26908 20356
rect 30370 20300 30380 20356
rect 30436 20300 32956 20356
rect 33012 20300 33022 20356
rect 39442 20300 39452 20356
rect 39508 20300 39900 20356
rect 39956 20300 41020 20356
rect 41076 20300 41468 20356
rect 41524 20300 41534 20356
rect 42130 20300 42140 20356
rect 42196 20300 42206 20356
rect 44818 20300 44828 20356
rect 44884 20300 46956 20356
rect 47012 20300 47516 20356
rect 47572 20300 47582 20356
rect 0 20244 800 20272
rect 1484 20244 1540 20300
rect 0 20188 1540 20244
rect 1698 20188 1708 20244
rect 1764 20188 2604 20244
rect 2660 20188 2670 20244
rect 0 20160 800 20188
rect 6300 20132 6356 20300
rect 20524 20244 20580 20300
rect 42140 20244 42196 20300
rect 6738 20188 6748 20244
rect 6804 20188 20580 20244
rect 6300 20076 7700 20132
rect 8866 20076 8876 20132
rect 8932 20076 10556 20132
rect 10612 20076 10622 20132
rect 11778 20076 11788 20132
rect 11844 20076 12012 20132
rect 12068 20076 12078 20132
rect 14018 20076 14028 20132
rect 14084 20076 15036 20132
rect 15092 20076 15102 20132
rect 27122 20076 27132 20132
rect 27188 20076 27916 20132
rect 27972 20076 27982 20132
rect 33618 20076 33628 20132
rect 33684 20076 34972 20132
rect 35028 20076 35038 20132
rect 7644 20020 7700 20076
rect 35252 20020 35308 20244
rect 35364 20188 36092 20244
rect 36148 20188 36158 20244
rect 42140 20188 44940 20244
rect 44996 20188 46732 20244
rect 46788 20188 46798 20244
rect 46610 20076 46620 20132
rect 46676 20076 47292 20132
rect 47348 20076 48524 20132
rect 48580 20076 48860 20132
rect 48916 20076 48926 20132
rect 7644 19964 9548 20020
rect 9604 19964 9614 20020
rect 9874 19964 9884 20020
rect 9940 19964 9950 20020
rect 14802 19964 14812 20020
rect 14868 19964 15372 20020
rect 15428 19964 15438 20020
rect 21186 19964 21196 20020
rect 21252 19964 24108 20020
rect 24164 19964 24174 20020
rect 34178 19964 34188 20020
rect 34244 19964 34860 20020
rect 34916 19964 35308 20020
rect 36306 19964 36316 20020
rect 36372 19964 37212 20020
rect 37268 19964 37278 20020
rect 50372 19964 52444 20020
rect 52500 19964 52510 20020
rect 9884 19908 9940 19964
rect 50372 19908 50428 19964
rect 1708 19852 5628 19908
rect 5684 19852 5694 19908
rect 7410 19852 7420 19908
rect 7476 19852 7486 19908
rect 9202 19852 9212 19908
rect 9268 19852 9940 19908
rect 22194 19852 22204 19908
rect 22260 19852 23660 19908
rect 23716 19852 23726 19908
rect 37090 19852 37100 19908
rect 37156 19852 38108 19908
rect 38164 19852 38174 19908
rect 39666 19852 39676 19908
rect 39732 19852 43708 19908
rect 43764 19852 43774 19908
rect 49970 19852 49980 19908
rect 50036 19852 50428 19908
rect 0 19572 800 19600
rect 1708 19572 1764 19852
rect 7420 19796 7476 19852
rect 4162 19740 4172 19796
rect 4228 19740 4900 19796
rect 6962 19740 6972 19796
rect 7028 19740 7476 19796
rect 10210 19740 10220 19796
rect 10276 19740 11452 19796
rect 11508 19740 13244 19796
rect 13300 19740 14364 19796
rect 14420 19740 14430 19796
rect 22306 19740 22316 19796
rect 22372 19740 23548 19796
rect 23604 19740 23614 19796
rect 23874 19740 23884 19796
rect 23940 19740 26908 19796
rect 33282 19740 33292 19796
rect 33348 19740 38668 19796
rect 38724 19740 39564 19796
rect 39620 19740 39630 19796
rect 39778 19740 39788 19796
rect 39844 19740 40236 19796
rect 40292 19740 40302 19796
rect 42130 19740 42140 19796
rect 42196 19740 42476 19796
rect 42532 19740 42542 19796
rect 45154 19740 45164 19796
rect 45220 19740 45612 19796
rect 45668 19740 45678 19796
rect 4844 19684 4900 19740
rect 4834 19628 4844 19684
rect 4900 19628 4910 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 0 19516 1708 19572
rect 1764 19516 1774 19572
rect 0 19488 800 19516
rect 26852 19460 26908 19740
rect 39788 19684 39844 19740
rect 39106 19628 39116 19684
rect 39172 19628 39844 19684
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 3378 19404 3388 19460
rect 3444 19404 6412 19460
rect 6468 19404 6478 19460
rect 26852 19404 41020 19460
rect 41076 19404 42140 19460
rect 42196 19404 42924 19460
rect 42980 19404 42990 19460
rect 44034 19404 44044 19460
rect 44100 19404 45948 19460
rect 46004 19404 46014 19460
rect 6178 19292 6188 19348
rect 6244 19292 8428 19348
rect 8484 19292 8494 19348
rect 12898 19292 12908 19348
rect 12964 19292 13580 19348
rect 13636 19292 13646 19348
rect 24434 19292 24444 19348
rect 24500 19292 25676 19348
rect 25732 19292 25742 19348
rect 31266 19292 31276 19348
rect 31332 19292 31612 19348
rect 31668 19292 31724 19348
rect 31780 19292 35868 19348
rect 35924 19292 35934 19348
rect 37762 19292 37772 19348
rect 37828 19292 38556 19348
rect 38612 19236 38668 19348
rect 43138 19292 43148 19348
rect 43204 19292 46172 19348
rect 46228 19292 46238 19348
rect 3798 19180 3836 19236
rect 3892 19180 3902 19236
rect 8306 19180 8316 19236
rect 8372 19180 9884 19236
rect 9940 19180 9950 19236
rect 12002 19180 12012 19236
rect 12068 19180 16044 19236
rect 16100 19180 16110 19236
rect 18610 19180 18620 19236
rect 18676 19180 19628 19236
rect 19684 19180 19694 19236
rect 21074 19180 21084 19236
rect 21140 19180 21644 19236
rect 21700 19180 21710 19236
rect 22316 19180 22540 19236
rect 22596 19180 25228 19236
rect 25284 19180 28028 19236
rect 28084 19180 28094 19236
rect 28578 19180 28588 19236
rect 28644 19180 29708 19236
rect 29764 19180 29774 19236
rect 32834 19180 32844 19236
rect 32900 19180 33516 19236
rect 33572 19180 33582 19236
rect 36754 19180 36764 19236
rect 36820 19180 38108 19236
rect 38164 19180 38174 19236
rect 38612 19180 43036 19236
rect 43092 19180 43484 19236
rect 43540 19180 43550 19236
rect 53666 19180 53676 19236
rect 53732 19180 54572 19236
rect 54628 19180 54638 19236
rect 22316 19124 22372 19180
rect 2706 19068 2716 19124
rect 2772 19068 6076 19124
rect 6132 19068 8092 19124
rect 8148 19068 8158 19124
rect 13682 19068 13692 19124
rect 13748 19068 14476 19124
rect 14532 19068 14542 19124
rect 15670 19068 15708 19124
rect 15764 19068 15774 19124
rect 16482 19068 16492 19124
rect 16548 19068 17276 19124
rect 17332 19068 17342 19124
rect 19516 19068 21196 19124
rect 21252 19068 21262 19124
rect 22306 19068 22316 19124
rect 22372 19068 22382 19124
rect 26114 19068 26124 19124
rect 26180 19068 26908 19124
rect 26964 19068 27132 19124
rect 27188 19068 27198 19124
rect 33180 19068 42700 19124
rect 42756 19068 43372 19124
rect 43428 19068 43438 19124
rect 52770 19068 52780 19124
rect 52836 19068 53452 19124
rect 53508 19068 53518 19124
rect 19516 19012 19572 19068
rect 2034 18956 2044 19012
rect 2100 18956 3388 19012
rect 7522 18956 7532 19012
rect 7588 18956 8652 19012
rect 8708 18956 9660 19012
rect 9716 18956 11116 19012
rect 11172 18956 19572 19012
rect 19628 18956 20412 19012
rect 20468 18956 20860 19012
rect 20916 18956 21084 19012
rect 21140 18956 21150 19012
rect 26786 18956 26796 19012
rect 26852 18956 32956 19012
rect 33012 18956 33022 19012
rect 0 18900 800 18928
rect 3332 18900 3388 18956
rect 0 18844 2380 18900
rect 2436 18844 3164 18900
rect 3220 18844 3230 18900
rect 3332 18844 15484 18900
rect 15540 18844 15550 18900
rect 15698 18844 15708 18900
rect 15764 18844 16156 18900
rect 16212 18844 16222 18900
rect 0 18816 800 18844
rect 19628 18788 19684 18956
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 8978 18732 8988 18788
rect 9044 18732 9324 18788
rect 9380 18732 10332 18788
rect 10388 18732 10398 18788
rect 11228 18732 12460 18788
rect 12516 18732 12526 18788
rect 15586 18732 15596 18788
rect 15652 18732 19404 18788
rect 19460 18732 19684 18788
rect 26562 18732 26572 18788
rect 26628 18732 27132 18788
rect 27188 18732 29036 18788
rect 29092 18732 29102 18788
rect 8866 18620 8876 18676
rect 8932 18620 9212 18676
rect 9268 18620 10220 18676
rect 10276 18620 11004 18676
rect 11060 18620 11070 18676
rect 11228 18564 11284 18732
rect 33180 18676 33236 19068
rect 35746 18956 35756 19012
rect 35812 18956 36652 19012
rect 36708 18956 36718 19012
rect 38518 18956 38556 19012
rect 38612 18956 38622 19012
rect 11638 18620 11676 18676
rect 11732 18620 11742 18676
rect 15026 18620 15036 18676
rect 15092 18620 16604 18676
rect 16660 18620 33236 18676
rect 33292 18844 39564 18900
rect 39620 18844 39630 18900
rect 33292 18564 33348 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 36194 18732 36204 18788
rect 36260 18732 36652 18788
rect 36708 18732 36718 18788
rect 37762 18732 37772 18788
rect 37828 18732 46396 18788
rect 46452 18732 46462 18788
rect 35858 18620 35868 18676
rect 35924 18620 36428 18676
rect 36484 18620 36494 18676
rect 40114 18620 40124 18676
rect 40180 18620 44604 18676
rect 44660 18620 44670 18676
rect 3612 18508 4620 18564
rect 4676 18508 4686 18564
rect 4834 18508 4844 18564
rect 4900 18508 7308 18564
rect 7364 18508 11284 18564
rect 12450 18508 12460 18564
rect 12516 18508 13804 18564
rect 13860 18508 13870 18564
rect 15474 18508 15484 18564
rect 15540 18508 15820 18564
rect 15876 18508 15886 18564
rect 16930 18508 16940 18564
rect 16996 18508 18844 18564
rect 18900 18508 18910 18564
rect 30146 18508 30156 18564
rect 30212 18508 33348 18564
rect 36726 18508 36764 18564
rect 36820 18508 36830 18564
rect 41346 18508 41356 18564
rect 41412 18508 44156 18564
rect 44212 18508 44716 18564
rect 44772 18508 44782 18564
rect 3612 18452 3668 18508
rect 3602 18396 3612 18452
rect 3668 18396 3678 18452
rect 3938 18396 3948 18452
rect 4004 18396 4284 18452
rect 4340 18396 4350 18452
rect 4498 18396 4508 18452
rect 4564 18396 5740 18452
rect 5796 18396 5806 18452
rect 7858 18396 7868 18452
rect 7924 18396 7934 18452
rect 8530 18396 8540 18452
rect 8596 18396 11340 18452
rect 11396 18396 11676 18452
rect 11732 18396 11742 18452
rect 15250 18396 15260 18452
rect 15316 18396 15932 18452
rect 15988 18396 17948 18452
rect 18004 18396 18014 18452
rect 19282 18396 19292 18452
rect 19348 18396 24724 18452
rect 25218 18396 25228 18452
rect 25284 18396 26684 18452
rect 26740 18396 26750 18452
rect 30930 18396 30940 18452
rect 30996 18396 32060 18452
rect 32116 18396 32126 18452
rect 33058 18396 33068 18452
rect 33124 18396 33516 18452
rect 33572 18396 33582 18452
rect 38546 18396 38556 18452
rect 38612 18396 39228 18452
rect 39284 18396 39294 18452
rect 39666 18396 39676 18452
rect 39732 18396 40348 18452
rect 40404 18396 43260 18452
rect 43316 18396 45052 18452
rect 45108 18396 45118 18452
rect 45378 18396 45388 18452
rect 45444 18396 47068 18452
rect 47124 18396 47628 18452
rect 47684 18396 48860 18452
rect 48916 18396 49756 18452
rect 49812 18396 50428 18452
rect 50484 18396 51996 18452
rect 52052 18396 53004 18452
rect 53060 18396 55244 18452
rect 55300 18396 55310 18452
rect 7868 18340 7924 18396
rect 24668 18340 24724 18396
rect 4386 18284 4396 18340
rect 4452 18284 5068 18340
rect 5124 18284 5134 18340
rect 7868 18284 8764 18340
rect 8820 18284 8830 18340
rect 22866 18284 22876 18340
rect 22932 18284 23884 18340
rect 23940 18284 24444 18340
rect 24500 18284 24510 18340
rect 24668 18284 26908 18340
rect 27010 18284 27020 18340
rect 27076 18284 31948 18340
rect 32004 18284 32014 18340
rect 32610 18284 32620 18340
rect 32676 18284 33180 18340
rect 33236 18284 33246 18340
rect 37996 18284 43484 18340
rect 43540 18284 43550 18340
rect 53554 18284 53564 18340
rect 53620 18284 54460 18340
rect 54516 18284 54526 18340
rect 0 18228 800 18256
rect 26852 18228 26908 18284
rect 37996 18228 38052 18284
rect 0 18172 1708 18228
rect 1764 18172 1774 18228
rect 3332 18172 6972 18228
rect 7028 18172 7038 18228
rect 7634 18172 7644 18228
rect 7700 18172 10332 18228
rect 10388 18172 10398 18228
rect 13906 18172 13916 18228
rect 13972 18172 15036 18228
rect 15092 18172 15102 18228
rect 19730 18172 19740 18228
rect 19796 18172 26348 18228
rect 26404 18172 26414 18228
rect 26852 18172 28028 18228
rect 28084 18172 28094 18228
rect 31602 18172 31612 18228
rect 31668 18172 35924 18228
rect 36418 18172 36428 18228
rect 36484 18172 37548 18228
rect 37604 18172 38052 18228
rect 38108 18172 42364 18228
rect 42420 18172 42430 18228
rect 0 18144 800 18172
rect 3332 17892 3388 18172
rect 10332 18116 10388 18172
rect 35868 18116 35924 18172
rect 38108 18116 38164 18172
rect 10332 18060 13020 18116
rect 13076 18060 13086 18116
rect 20290 18060 20300 18116
rect 20356 18060 30940 18116
rect 30996 18060 31006 18116
rect 35868 18060 36652 18116
rect 36708 18060 36718 18116
rect 37314 18060 37324 18116
rect 37380 18060 38164 18116
rect 38612 18060 41468 18116
rect 41524 18060 41534 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 8866 17948 8876 18004
rect 8932 17948 9324 18004
rect 9380 17948 9390 18004
rect 16146 17948 16156 18004
rect 16212 17948 17164 18004
rect 17220 17948 17230 18004
rect 24210 17948 24220 18004
rect 24276 17948 25228 18004
rect 25284 17948 25294 18004
rect 28242 17948 28252 18004
rect 28308 17948 29372 18004
rect 29428 17948 30156 18004
rect 30212 17948 30222 18004
rect 31042 17948 31052 18004
rect 31108 17948 34300 18004
rect 34356 17948 34366 18004
rect 25228 17892 25284 17948
rect 38612 17892 38668 18060
rect 39778 17948 39788 18004
rect 39844 17948 40348 18004
rect 40404 17948 40414 18004
rect 42466 17948 42476 18004
rect 42532 17948 42812 18004
rect 42868 17948 42878 18004
rect 2034 17836 2044 17892
rect 2100 17836 3388 17892
rect 22082 17836 22092 17892
rect 22148 17836 25004 17892
rect 25060 17836 25070 17892
rect 25228 17836 38668 17892
rect 1698 17724 1708 17780
rect 1764 17724 5068 17780
rect 5124 17724 5134 17780
rect 7298 17724 7308 17780
rect 7364 17724 8316 17780
rect 8372 17724 8382 17780
rect 13346 17724 13356 17780
rect 13412 17724 13692 17780
rect 13748 17724 13758 17780
rect 17378 17724 17388 17780
rect 17444 17724 18284 17780
rect 18340 17724 18350 17780
rect 30930 17724 30940 17780
rect 30996 17724 31388 17780
rect 31444 17724 31454 17780
rect 32050 17724 32060 17780
rect 32116 17724 41244 17780
rect 41300 17724 41310 17780
rect 41682 17724 41692 17780
rect 41748 17724 44044 17780
rect 44100 17724 44940 17780
rect 44996 17724 45006 17780
rect 41692 17668 41748 17724
rect 2930 17612 2940 17668
rect 2996 17612 6188 17668
rect 6244 17612 6254 17668
rect 7532 17612 8876 17668
rect 8932 17612 8942 17668
rect 20514 17612 20524 17668
rect 20580 17612 21420 17668
rect 21476 17612 22876 17668
rect 22932 17612 22942 17668
rect 26898 17612 26908 17668
rect 26964 17612 27580 17668
rect 27636 17612 27646 17668
rect 27794 17612 27804 17668
rect 27860 17612 28364 17668
rect 28420 17612 30268 17668
rect 30324 17612 30334 17668
rect 32386 17612 32396 17668
rect 32452 17612 33292 17668
rect 33348 17612 33404 17668
rect 33460 17612 33470 17668
rect 36754 17612 36764 17668
rect 36820 17612 37884 17668
rect 37940 17612 37950 17668
rect 39666 17612 39676 17668
rect 39732 17612 41748 17668
rect 44258 17612 44268 17668
rect 44324 17612 47180 17668
rect 47236 17612 47246 17668
rect 50754 17612 50764 17668
rect 50820 17612 52332 17668
rect 52388 17612 52398 17668
rect 0 17556 800 17584
rect 7532 17556 7588 17612
rect 41244 17556 41300 17612
rect 0 17500 1708 17556
rect 1764 17500 1774 17556
rect 7522 17500 7532 17556
rect 7588 17500 7598 17556
rect 7746 17500 7756 17556
rect 7812 17500 8092 17556
rect 8148 17500 8158 17556
rect 13906 17500 13916 17556
rect 13972 17500 14476 17556
rect 14532 17500 14542 17556
rect 24770 17500 24780 17556
rect 24836 17500 25340 17556
rect 25396 17500 25406 17556
rect 26898 17500 26908 17556
rect 26964 17500 28588 17556
rect 28644 17500 28654 17556
rect 29138 17500 29148 17556
rect 29204 17500 31724 17556
rect 31780 17500 31790 17556
rect 41234 17500 41244 17556
rect 41300 17500 41310 17556
rect 45938 17500 45948 17556
rect 46004 17500 46014 17556
rect 46162 17500 46172 17556
rect 46228 17500 46732 17556
rect 46788 17500 47292 17556
rect 47348 17500 48748 17556
rect 48804 17500 48814 17556
rect 0 17472 800 17500
rect 45948 17444 46004 17500
rect 10882 17388 10892 17444
rect 10948 17388 15596 17444
rect 15652 17388 16716 17444
rect 16772 17388 16782 17444
rect 26002 17388 26012 17444
rect 26068 17388 27468 17444
rect 27524 17388 27534 17444
rect 28466 17388 28476 17444
rect 28532 17388 30492 17444
rect 30548 17388 30558 17444
rect 33170 17388 33180 17444
rect 33236 17388 33964 17444
rect 34020 17388 34030 17444
rect 34290 17388 34300 17444
rect 34356 17388 34748 17444
rect 34804 17388 34814 17444
rect 43810 17388 43820 17444
rect 43876 17388 45724 17444
rect 45780 17388 45790 17444
rect 45948 17388 47068 17444
rect 47124 17388 47964 17444
rect 48020 17388 48030 17444
rect 51202 17388 51212 17444
rect 51268 17388 51324 17444
rect 51380 17388 53340 17444
rect 53396 17388 53406 17444
rect 1586 17276 1596 17332
rect 1652 17276 4340 17332
rect 6850 17276 6860 17332
rect 6916 17276 7868 17332
rect 7924 17276 7934 17332
rect 11302 17276 11340 17332
rect 11396 17276 11406 17332
rect 28578 17276 28588 17332
rect 28644 17276 30044 17332
rect 30100 17276 30110 17332
rect 34514 17276 34524 17332
rect 34580 17276 34972 17332
rect 35028 17276 36428 17332
rect 36484 17276 37436 17332
rect 37492 17276 37502 17332
rect 4284 17108 4340 17276
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 29474 17164 29484 17220
rect 29540 17164 31052 17220
rect 31108 17164 31118 17220
rect 3154 17052 3164 17108
rect 3220 17052 4060 17108
rect 4116 17052 4126 17108
rect 4274 17052 4284 17108
rect 4340 17052 4350 17108
rect 10210 17052 10220 17108
rect 10276 17052 11340 17108
rect 11396 17052 11676 17108
rect 11732 17052 11742 17108
rect 18946 17052 18956 17108
rect 19012 17052 19404 17108
rect 19460 17052 20076 17108
rect 20132 17052 20412 17108
rect 20468 17052 20478 17108
rect 20738 17052 20748 17108
rect 20804 17052 21756 17108
rect 21812 17052 22428 17108
rect 22484 17052 22494 17108
rect 25778 17052 25788 17108
rect 25844 17052 26908 17108
rect 26964 17052 26974 17108
rect 34402 17052 34412 17108
rect 34468 17052 37772 17108
rect 37828 17052 37838 17108
rect 42354 17052 42364 17108
rect 42420 17052 42588 17108
rect 42644 17052 42654 17108
rect 45154 17052 45164 17108
rect 45220 17052 46060 17108
rect 46116 17052 46126 17108
rect 13122 16940 13132 16996
rect 13188 16940 14700 16996
rect 14756 16940 15036 16996
rect 15092 16940 15102 16996
rect 27682 16940 27692 16996
rect 27748 16940 28476 16996
rect 28532 16940 29484 16996
rect 29540 16940 30268 16996
rect 30324 16940 30334 16996
rect 0 16884 800 16912
rect 37772 16884 37828 17052
rect 38994 16940 39004 16996
rect 39060 16940 39452 16996
rect 39508 16940 41580 16996
rect 41636 16940 43260 16996
rect 43316 16940 44044 16996
rect 44100 16940 44110 16996
rect 45826 16940 45836 16996
rect 45892 16940 46620 16996
rect 46676 16940 46686 16996
rect 0 16828 2380 16884
rect 2436 16828 5180 16884
rect 5236 16828 5246 16884
rect 21970 16828 21980 16884
rect 22036 16828 25228 16884
rect 25284 16828 25676 16884
rect 25732 16828 25742 16884
rect 32498 16828 32508 16884
rect 32564 16828 33180 16884
rect 33236 16828 33246 16884
rect 37772 16828 39116 16884
rect 39172 16828 39676 16884
rect 39732 16828 39742 16884
rect 41916 16828 42028 16884
rect 42084 16828 42094 16884
rect 44930 16828 44940 16884
rect 44996 16828 45948 16884
rect 46004 16828 46014 16884
rect 0 16800 800 16828
rect 22764 16772 22820 16828
rect 2482 16716 2492 16772
rect 2548 16716 3276 16772
rect 3332 16716 3342 16772
rect 4274 16716 4284 16772
rect 4340 16716 5068 16772
rect 5124 16716 5134 16772
rect 5506 16716 5516 16772
rect 5572 16716 6636 16772
rect 6692 16716 6702 16772
rect 22754 16716 22764 16772
rect 22820 16716 22830 16772
rect 24658 16716 24668 16772
rect 24724 16716 25564 16772
rect 25620 16716 25630 16772
rect 26786 16716 26796 16772
rect 26852 16716 27356 16772
rect 27412 16716 28364 16772
rect 28420 16716 28430 16772
rect 33618 16716 33628 16772
rect 33684 16716 33964 16772
rect 34020 16716 34030 16772
rect 34850 16716 34860 16772
rect 34916 16716 36876 16772
rect 36932 16716 36942 16772
rect 37986 16716 37996 16772
rect 38052 16716 39228 16772
rect 39284 16716 39294 16772
rect 41916 16660 41972 16828
rect 42130 16716 42140 16772
rect 42196 16716 42812 16772
rect 42868 16716 42878 16772
rect 43026 16716 43036 16772
rect 43092 16716 43372 16772
rect 43428 16716 43438 16772
rect 48178 16716 48188 16772
rect 48244 16716 48748 16772
rect 48804 16716 49196 16772
rect 49252 16716 49262 16772
rect 49410 16716 49420 16772
rect 49476 16716 50092 16772
rect 50148 16716 50652 16772
rect 50708 16716 51100 16772
rect 51156 16716 51166 16772
rect 2034 16604 2044 16660
rect 2100 16604 14028 16660
rect 14084 16604 14812 16660
rect 14868 16604 14878 16660
rect 15698 16604 15708 16660
rect 15764 16604 17276 16660
rect 17332 16604 17342 16660
rect 23986 16604 23996 16660
rect 24052 16604 28588 16660
rect 28644 16604 28654 16660
rect 41916 16604 42588 16660
rect 42644 16604 42654 16660
rect 6962 16492 6972 16548
rect 7028 16492 8204 16548
rect 8260 16492 9884 16548
rect 9940 16492 16156 16548
rect 16212 16492 16716 16548
rect 16772 16492 16782 16548
rect 27346 16492 27356 16548
rect 27412 16492 33292 16548
rect 33348 16492 33358 16548
rect 37538 16492 37548 16548
rect 37604 16492 42252 16548
rect 42308 16492 42318 16548
rect 42914 16492 42924 16548
rect 42980 16492 43372 16548
rect 43428 16492 43438 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 25442 16380 25452 16436
rect 25508 16380 26908 16436
rect 35746 16380 35756 16436
rect 35812 16380 36316 16436
rect 36372 16380 38220 16436
rect 38276 16380 38286 16436
rect 41906 16380 41916 16436
rect 41972 16380 42700 16436
rect 42756 16380 43260 16436
rect 43316 16380 43326 16436
rect 47842 16380 47852 16436
rect 47908 16380 49084 16436
rect 49140 16380 49150 16436
rect 2706 16268 2716 16324
rect 2772 16268 6972 16324
rect 7028 16268 8092 16324
rect 8148 16268 8764 16324
rect 8820 16268 8830 16324
rect 11666 16268 11676 16324
rect 11732 16268 11742 16324
rect 17042 16268 17052 16324
rect 17108 16268 18396 16324
rect 18452 16268 18462 16324
rect 0 16212 800 16240
rect 11676 16212 11732 16268
rect 26852 16212 26908 16380
rect 31266 16268 31276 16324
rect 31332 16268 33068 16324
rect 33124 16268 33134 16324
rect 37090 16268 37100 16324
rect 37156 16268 37548 16324
rect 37604 16268 37614 16324
rect 45266 16268 45276 16324
rect 45332 16268 46508 16324
rect 46564 16268 47068 16324
rect 47124 16268 47134 16324
rect 47292 16268 47516 16324
rect 47572 16268 47582 16324
rect 47292 16212 47348 16268
rect 0 16156 1708 16212
rect 1764 16156 1774 16212
rect 4050 16156 4060 16212
rect 4116 16156 4620 16212
rect 4676 16156 4686 16212
rect 11676 16156 12124 16212
rect 12180 16156 14364 16212
rect 14420 16156 14430 16212
rect 26852 16156 46060 16212
rect 46116 16156 46126 16212
rect 47170 16156 47180 16212
rect 47236 16156 47348 16212
rect 0 16128 800 16156
rect 11778 16044 11788 16100
rect 11844 16044 12348 16100
rect 12404 16044 12414 16100
rect 21522 16044 21532 16100
rect 21588 16044 22204 16100
rect 22260 16044 22270 16100
rect 22978 16044 22988 16100
rect 23044 16044 23660 16100
rect 23716 16044 23726 16100
rect 25554 16044 25564 16100
rect 25620 16044 26572 16100
rect 26628 16044 26638 16100
rect 26982 16044 27020 16100
rect 27076 16044 27086 16100
rect 33842 16044 33852 16100
rect 33908 16044 34748 16100
rect 34804 16044 34814 16100
rect 35522 16044 35532 16100
rect 35588 16044 38108 16100
rect 38164 16044 38174 16100
rect 47506 16044 47516 16100
rect 47572 16044 49196 16100
rect 49252 16044 49262 16100
rect 50372 16044 50764 16100
rect 50820 16044 50830 16100
rect 22204 15988 22260 16044
rect 11330 15932 11340 15988
rect 11396 15932 11406 15988
rect 12786 15932 12796 15988
rect 12852 15932 13692 15988
rect 13748 15932 13758 15988
rect 22204 15932 23772 15988
rect 23828 15932 23838 15988
rect 24546 15932 24556 15988
rect 24612 15932 27692 15988
rect 27748 15932 27758 15988
rect 32722 15932 32732 15988
rect 32788 15932 32798 15988
rect 33030 15932 33068 15988
rect 33124 15932 33134 15988
rect 35634 15932 35644 15988
rect 35700 15932 36988 15988
rect 37044 15932 37054 15988
rect 37426 15932 37436 15988
rect 37492 15932 37884 15988
rect 37940 15932 37950 15988
rect 48066 15932 48076 15988
rect 48132 15932 48748 15988
rect 48804 15932 48814 15988
rect 11340 15876 11396 15932
rect 32732 15876 32788 15932
rect 50372 15876 50428 16044
rect 50530 15932 50540 15988
rect 50596 15932 50988 15988
rect 51044 15932 51054 15988
rect 7074 15820 7084 15876
rect 7140 15820 8988 15876
rect 9044 15820 9054 15876
rect 11340 15820 23100 15876
rect 23156 15820 23166 15876
rect 32732 15820 33292 15876
rect 33348 15820 34300 15876
rect 34356 15820 34366 15876
rect 35970 15820 35980 15876
rect 36036 15820 37324 15876
rect 37380 15820 37390 15876
rect 43138 15820 43148 15876
rect 43204 15820 43820 15876
rect 43876 15820 43886 15876
rect 47954 15820 47964 15876
rect 48020 15820 48524 15876
rect 48580 15820 49532 15876
rect 49588 15820 49598 15876
rect 49858 15820 49868 15876
rect 49924 15820 50428 15876
rect 51090 15820 51100 15876
rect 51156 15820 51212 15876
rect 51268 15820 51278 15876
rect 51650 15820 51660 15876
rect 51716 15820 52556 15876
rect 52612 15820 52622 15876
rect 52770 15820 52780 15876
rect 52836 15820 53116 15876
rect 53172 15820 53182 15876
rect 3714 15708 3724 15764
rect 3780 15708 4732 15764
rect 4788 15708 4798 15764
rect 50978 15708 50988 15764
rect 51044 15708 51548 15764
rect 51604 15708 51614 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 1698 15596 1708 15652
rect 1764 15596 4844 15652
rect 4900 15596 4910 15652
rect 8306 15596 8316 15652
rect 8372 15596 9436 15652
rect 9492 15596 9660 15652
rect 9716 15596 9726 15652
rect 9874 15596 9884 15652
rect 9940 15596 11004 15652
rect 11060 15596 13132 15652
rect 13188 15596 14028 15652
rect 14084 15596 14094 15652
rect 15092 15596 15260 15652
rect 15316 15596 15326 15652
rect 33842 15596 33852 15652
rect 33908 15596 33918 15652
rect 38098 15596 38108 15652
rect 38164 15596 38892 15652
rect 38948 15596 38958 15652
rect 42578 15596 42588 15652
rect 42644 15596 43484 15652
rect 43540 15596 43550 15652
rect 0 15540 800 15568
rect 0 15484 2380 15540
rect 2436 15484 2446 15540
rect 2706 15484 2716 15540
rect 2772 15484 4004 15540
rect 5954 15484 5964 15540
rect 6020 15484 6188 15540
rect 6244 15484 10444 15540
rect 10500 15484 10510 15540
rect 0 15456 800 15484
rect 2380 15428 2436 15484
rect 3948 15428 4004 15484
rect 15092 15428 15148 15596
rect 33852 15540 33908 15596
rect 31826 15484 31836 15540
rect 31892 15484 32620 15540
rect 32676 15484 33908 15540
rect 35186 15484 35196 15540
rect 35252 15484 35980 15540
rect 36036 15484 36046 15540
rect 37090 15484 37100 15540
rect 37156 15484 39228 15540
rect 39284 15484 39294 15540
rect 46060 15484 48244 15540
rect 50082 15484 50092 15540
rect 50148 15484 51100 15540
rect 51156 15484 51166 15540
rect 35980 15428 36036 15484
rect 46060 15428 46116 15484
rect 2034 15372 2044 15428
rect 2100 15372 2110 15428
rect 2380 15372 3612 15428
rect 3668 15372 3678 15428
rect 3948 15372 14700 15428
rect 14756 15372 15148 15428
rect 28018 15372 28028 15428
rect 28084 15372 28812 15428
rect 28868 15372 28878 15428
rect 31042 15372 31052 15428
rect 31108 15372 31276 15428
rect 31332 15372 31948 15428
rect 32004 15372 32284 15428
rect 32340 15372 33068 15428
rect 33124 15372 33134 15428
rect 35980 15372 38668 15428
rect 43922 15372 43932 15428
rect 43988 15372 45276 15428
rect 45332 15372 45342 15428
rect 46050 15372 46060 15428
rect 46116 15372 46126 15428
rect 46946 15372 46956 15428
rect 47012 15372 47740 15428
rect 47796 15372 47806 15428
rect 2044 15204 2100 15372
rect 3042 15260 3052 15316
rect 3108 15260 4060 15316
rect 4116 15260 4126 15316
rect 4498 15260 4508 15316
rect 4564 15260 6076 15316
rect 6132 15260 6142 15316
rect 6738 15260 6748 15316
rect 6804 15260 8092 15316
rect 8148 15260 8652 15316
rect 8708 15260 9884 15316
rect 9940 15260 9950 15316
rect 13010 15260 13020 15316
rect 13076 15260 13804 15316
rect 13860 15260 13870 15316
rect 14354 15260 14364 15316
rect 14420 15260 16156 15316
rect 16212 15260 16222 15316
rect 16594 15260 16604 15316
rect 16660 15260 17948 15316
rect 18004 15260 18014 15316
rect 22418 15260 22428 15316
rect 22484 15260 25228 15316
rect 25284 15260 25900 15316
rect 25956 15260 25966 15316
rect 25900 15204 25956 15260
rect 26852 15204 26908 15316
rect 26964 15260 26974 15316
rect 38210 15260 38220 15316
rect 38276 15260 38444 15316
rect 38500 15260 38510 15316
rect 38612 15204 38668 15372
rect 42914 15260 42924 15316
rect 42980 15260 43596 15316
rect 43652 15260 43662 15316
rect 44482 15260 44492 15316
rect 44548 15260 44558 15316
rect 44828 15260 46172 15316
rect 46228 15260 46620 15316
rect 46676 15260 46686 15316
rect 46834 15260 46844 15316
rect 46900 15260 47292 15316
rect 47348 15260 47358 15316
rect 44492 15204 44548 15260
rect 2044 15148 7084 15204
rect 7140 15148 7150 15204
rect 8418 15148 8428 15204
rect 8484 15148 10108 15204
rect 10164 15148 10174 15204
rect 16706 15148 16716 15204
rect 16772 15148 17612 15204
rect 17668 15148 17678 15204
rect 18386 15148 18396 15204
rect 18452 15148 18956 15204
rect 19012 15148 19740 15204
rect 19796 15148 19806 15204
rect 22978 15148 22988 15204
rect 23044 15148 23324 15204
rect 23380 15148 23390 15204
rect 25900 15148 26908 15204
rect 31602 15148 31612 15204
rect 31668 15148 32396 15204
rect 32452 15148 32462 15204
rect 33516 15148 33852 15204
rect 33908 15148 33918 15204
rect 35410 15148 35420 15204
rect 35476 15148 35756 15204
rect 35812 15148 35822 15204
rect 38612 15148 38780 15204
rect 38836 15148 40012 15204
rect 40068 15148 40078 15204
rect 43474 15148 43484 15204
rect 43540 15148 44548 15204
rect 33516 15092 33572 15148
rect 44828 15092 44884 15260
rect 48188 15204 48244 15484
rect 49410 15372 49420 15428
rect 49476 15372 50428 15428
rect 50484 15372 50494 15428
rect 45154 15148 45164 15204
rect 45220 15148 46396 15204
rect 46452 15148 46462 15204
rect 48188 15148 52780 15204
rect 52836 15148 52846 15204
rect 1698 15036 1708 15092
rect 1764 15036 5964 15092
rect 6020 15036 6030 15092
rect 6962 15036 6972 15092
rect 7028 15036 7420 15092
rect 7476 15036 7486 15092
rect 15586 15036 15596 15092
rect 15652 15036 16380 15092
rect 16436 15036 16446 15092
rect 27234 15036 27244 15092
rect 27300 15036 30604 15092
rect 30660 15036 30670 15092
rect 32050 15036 32060 15092
rect 32116 15036 33292 15092
rect 33348 15036 33358 15092
rect 33506 15036 33516 15092
rect 33572 15036 33582 15092
rect 34150 15036 34188 15092
rect 34244 15036 34254 15092
rect 44818 15036 44828 15092
rect 44884 15036 44894 15092
rect 0 14868 800 14896
rect 1708 14868 1764 15036
rect 16118 14924 16156 14980
rect 16212 14924 16222 14980
rect 34066 14924 34076 14980
rect 34132 14924 34142 14980
rect 37538 14924 37548 14980
rect 37604 14924 37996 14980
rect 38052 14924 38062 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 0 14812 1764 14868
rect 25330 14812 25340 14868
rect 25396 14812 26348 14868
rect 26404 14812 26908 14868
rect 26964 14812 27916 14868
rect 27972 14812 27982 14868
rect 0 14784 800 14812
rect 2034 14700 2044 14756
rect 2100 14700 11676 14756
rect 11732 14700 11742 14756
rect 2706 14588 2716 14644
rect 2772 14588 11900 14644
rect 11956 14588 12572 14644
rect 12628 14588 12638 14644
rect 18834 14588 18844 14644
rect 18900 14588 19628 14644
rect 19684 14588 19694 14644
rect 34076 14532 34132 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 35858 14812 35868 14868
rect 35924 14812 36148 14868
rect 36278 14812 36316 14868
rect 36372 14812 36382 14868
rect 42690 14812 42700 14868
rect 42756 14812 47068 14868
rect 47124 14812 47134 14868
rect 36092 14756 36148 14812
rect 36082 14700 36092 14756
rect 36148 14700 36158 14756
rect 42018 14588 42028 14644
rect 42084 14588 46620 14644
rect 46676 14588 46686 14644
rect 48514 14588 48524 14644
rect 48580 14588 49084 14644
rect 49140 14588 51660 14644
rect 51716 14588 51726 14644
rect 2482 14476 2492 14532
rect 2548 14476 5068 14532
rect 5124 14476 5134 14532
rect 7746 14476 7756 14532
rect 7812 14476 8204 14532
rect 8260 14476 8270 14532
rect 10434 14476 10444 14532
rect 10500 14476 13916 14532
rect 13972 14476 14812 14532
rect 14868 14476 14878 14532
rect 18498 14476 18508 14532
rect 18564 14476 18732 14532
rect 18788 14476 18798 14532
rect 19506 14476 19516 14532
rect 19572 14476 20300 14532
rect 20356 14476 20366 14532
rect 26674 14476 26684 14532
rect 26740 14476 27580 14532
rect 27636 14476 27646 14532
rect 33282 14476 33292 14532
rect 33348 14476 34076 14532
rect 34132 14476 34142 14532
rect 34962 14476 34972 14532
rect 35028 14476 37212 14532
rect 37268 14476 38444 14532
rect 38500 14476 38510 14532
rect 39554 14476 39564 14532
rect 39620 14476 41356 14532
rect 41412 14476 41422 14532
rect 43362 14476 43372 14532
rect 43428 14476 48860 14532
rect 48916 14476 49420 14532
rect 49476 14476 49486 14532
rect 2492 14308 2548 14476
rect 7298 14364 7308 14420
rect 7364 14364 8316 14420
rect 8372 14364 8382 14420
rect 17042 14364 17052 14420
rect 17108 14364 18060 14420
rect 18116 14364 18126 14420
rect 18386 14364 18396 14420
rect 18452 14364 19404 14420
rect 19460 14364 19470 14420
rect 26002 14364 26012 14420
rect 26068 14364 26796 14420
rect 26852 14364 27468 14420
rect 27524 14364 27534 14420
rect 29698 14364 29708 14420
rect 29764 14364 39452 14420
rect 39508 14364 41468 14420
rect 41524 14364 41534 14420
rect 924 14252 2548 14308
rect 7970 14252 7980 14308
rect 8036 14252 8046 14308
rect 34962 14252 34972 14308
rect 35028 14252 36988 14308
rect 37044 14252 37548 14308
rect 37604 14252 37614 14308
rect 0 14196 800 14224
rect 924 14196 980 14252
rect 7980 14196 8036 14252
rect 0 14140 980 14196
rect 7746 14140 7756 14196
rect 7812 14140 8036 14196
rect 20178 14140 20188 14196
rect 20244 14140 26012 14196
rect 26068 14140 26078 14196
rect 35970 14140 35980 14196
rect 36036 14140 36652 14196
rect 36708 14140 36718 14196
rect 45938 14140 45948 14196
rect 46004 14140 47572 14196
rect 49746 14140 49756 14196
rect 49812 14140 50428 14196
rect 0 14112 800 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 7186 14028 7196 14084
rect 7252 14028 7980 14084
rect 8036 14028 8046 14084
rect 23090 14028 23100 14084
rect 23156 14028 37884 14084
rect 37940 14028 37950 14084
rect 47516 13972 47572 14140
rect 50372 13972 50428 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 11106 13916 11116 13972
rect 11172 13916 13020 13972
rect 13076 13916 13086 13972
rect 16818 13916 16828 13972
rect 16884 13916 17836 13972
rect 17892 13916 17902 13972
rect 22866 13916 22876 13972
rect 22932 13916 24668 13972
rect 24724 13916 25004 13972
rect 25060 13916 25070 13972
rect 25554 13916 25564 13972
rect 25620 13916 27020 13972
rect 27076 13916 27086 13972
rect 31154 13916 31164 13972
rect 31220 13916 31612 13972
rect 31668 13916 31678 13972
rect 37762 13916 37772 13972
rect 37828 13916 39340 13972
rect 39396 13916 39406 13972
rect 44818 13916 44828 13972
rect 44884 13916 46620 13972
rect 46676 13916 46686 13972
rect 47506 13916 47516 13972
rect 47572 13916 49756 13972
rect 49812 13916 49822 13972
rect 50372 13916 50764 13972
rect 50820 13916 50830 13972
rect 7606 13804 7644 13860
rect 7700 13804 7710 13860
rect 27122 13804 27132 13860
rect 27188 13804 29372 13860
rect 29428 13804 31052 13860
rect 31108 13804 31118 13860
rect 33282 13804 33292 13860
rect 33348 13804 34524 13860
rect 34580 13804 34590 13860
rect 36764 13804 41132 13860
rect 41188 13804 41198 13860
rect 47282 13804 47292 13860
rect 47348 13804 49644 13860
rect 49700 13804 50092 13860
rect 50148 13804 50158 13860
rect 50372 13804 54236 13860
rect 54292 13804 54302 13860
rect 36764 13748 36820 13804
rect 2706 13692 2716 13748
rect 2772 13692 9996 13748
rect 10052 13692 10062 13748
rect 11442 13692 11452 13748
rect 11508 13692 13804 13748
rect 13860 13692 15036 13748
rect 15092 13692 15102 13748
rect 25330 13692 25340 13748
rect 25396 13692 26012 13748
rect 26068 13692 26078 13748
rect 34066 13692 34076 13748
rect 34132 13692 35420 13748
rect 35476 13692 35486 13748
rect 36754 13692 36764 13748
rect 36820 13692 36830 13748
rect 38770 13692 38780 13748
rect 38836 13692 39452 13748
rect 39508 13692 42700 13748
rect 42756 13692 42766 13748
rect 43026 13692 43036 13748
rect 43092 13692 44044 13748
rect 44100 13692 44110 13748
rect 3332 13580 5068 13636
rect 5124 13580 5134 13636
rect 16370 13580 16380 13636
rect 16436 13580 17276 13636
rect 17332 13580 17342 13636
rect 18050 13580 18060 13636
rect 18116 13580 18396 13636
rect 18452 13580 18462 13636
rect 20178 13580 20188 13636
rect 20244 13580 21532 13636
rect 21588 13580 21598 13636
rect 29922 13580 29932 13636
rect 29988 13580 39564 13636
rect 39620 13580 39630 13636
rect 41122 13580 41132 13636
rect 41188 13580 42252 13636
rect 42308 13580 42318 13636
rect 49074 13580 49084 13636
rect 49140 13580 50316 13636
rect 50372 13580 50428 13804
rect 0 13524 800 13552
rect 0 13468 1764 13524
rect 3266 13468 3276 13524
rect 3332 13468 3388 13580
rect 4284 13468 5292 13524
rect 5348 13468 5358 13524
rect 16482 13468 16492 13524
rect 16548 13468 17612 13524
rect 17668 13468 17678 13524
rect 27794 13468 27804 13524
rect 27860 13468 28924 13524
rect 28980 13468 28990 13524
rect 34738 13468 34748 13524
rect 34804 13468 36204 13524
rect 36260 13468 36652 13524
rect 36708 13468 36718 13524
rect 41010 13468 41020 13524
rect 41076 13468 42588 13524
rect 42644 13468 42654 13524
rect 0 13440 800 13468
rect 1708 13412 1764 13468
rect 4284 13412 4340 13468
rect 1698 13356 1708 13412
rect 1764 13356 1774 13412
rect 4274 13356 4284 13412
rect 4340 13356 4350 13412
rect 6962 13356 6972 13412
rect 7028 13356 8092 13412
rect 8148 13356 8158 13412
rect 26226 13356 26236 13412
rect 26292 13356 26572 13412
rect 26628 13356 28252 13412
rect 28308 13356 28318 13412
rect 30930 13356 30940 13412
rect 30996 13356 31836 13412
rect 31892 13356 31902 13412
rect 43138 13356 43148 13412
rect 43204 13356 44268 13412
rect 44324 13356 44334 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 13570 13244 13580 13300
rect 13636 13244 13916 13300
rect 13972 13244 13982 13300
rect 24994 13244 25004 13300
rect 25060 13244 26908 13300
rect 26852 13188 26908 13244
rect 12562 13132 12572 13188
rect 12628 13132 13468 13188
rect 13524 13132 13534 13188
rect 26852 13132 40404 13188
rect 2482 13020 2492 13076
rect 2548 13020 3388 13076
rect 3444 13020 3454 13076
rect 4918 13020 4956 13076
rect 5012 13020 5022 13076
rect 26450 13020 26460 13076
rect 26516 13020 26796 13076
rect 26852 13020 26862 13076
rect 2370 12908 2380 12964
rect 2436 12908 5740 12964
rect 5796 12908 5806 12964
rect 24108 12908 26908 12964
rect 26964 12908 26974 12964
rect 28354 12908 28364 12964
rect 28420 12908 29148 12964
rect 29204 12908 29214 12964
rect 30706 12908 30716 12964
rect 30772 12908 31612 12964
rect 31668 12908 31678 12964
rect 0 12852 800 12880
rect 2380 12852 2436 12908
rect 24108 12852 24164 12908
rect 0 12796 2436 12852
rect 24098 12796 24108 12852
rect 24164 12796 24174 12852
rect 24658 12796 24668 12852
rect 24724 12796 25116 12852
rect 25172 12796 25182 12852
rect 31378 12796 31388 12852
rect 31444 12796 33404 12852
rect 33460 12796 33470 12852
rect 0 12768 800 12796
rect 40348 12740 40404 13132
rect 40674 13020 40684 13076
rect 40740 13020 41468 13076
rect 41524 13020 41534 13076
rect 41906 13020 41916 13076
rect 41972 13020 42364 13076
rect 42420 13020 42430 13076
rect 41122 12796 41132 12852
rect 41188 12796 44156 12852
rect 44212 12796 44222 12852
rect 2034 12684 2044 12740
rect 2100 12684 10444 12740
rect 10500 12684 10510 12740
rect 10658 12684 10668 12740
rect 10724 12684 13692 12740
rect 13748 12684 14700 12740
rect 14756 12684 14766 12740
rect 22530 12684 22540 12740
rect 22596 12684 24220 12740
rect 24276 12684 24286 12740
rect 26002 12684 26012 12740
rect 26068 12684 26908 12740
rect 26964 12684 27356 12740
rect 27412 12684 27422 12740
rect 32498 12684 32508 12740
rect 32564 12684 34300 12740
rect 34356 12684 35196 12740
rect 35252 12684 35262 12740
rect 37762 12684 37772 12740
rect 37828 12684 38556 12740
rect 38612 12684 38622 12740
rect 40338 12684 40348 12740
rect 40404 12684 42140 12740
rect 42196 12684 42206 12740
rect 42354 12684 42364 12740
rect 42420 12684 43260 12740
rect 43316 12684 43326 12740
rect 1698 12572 1708 12628
rect 1764 12572 4172 12628
rect 4228 12572 4238 12628
rect 19058 12572 19068 12628
rect 19124 12572 19134 12628
rect 31490 12572 31500 12628
rect 31556 12572 31948 12628
rect 32004 12572 32014 12628
rect 33366 12572 33404 12628
rect 33460 12572 33470 12628
rect 2034 12460 2044 12516
rect 2100 12460 6412 12516
rect 6468 12460 7756 12516
rect 7812 12460 7822 12516
rect 13542 12460 13580 12516
rect 13636 12460 13646 12516
rect 19068 12404 19124 12572
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 38518 12460 38556 12516
rect 38612 12460 38622 12516
rect 3602 12348 3612 12404
rect 3668 12348 4508 12404
rect 4564 12348 5852 12404
rect 5908 12348 5918 12404
rect 13122 12348 13132 12404
rect 13188 12348 14140 12404
rect 14196 12348 14206 12404
rect 14690 12348 14700 12404
rect 14756 12348 15484 12404
rect 15540 12348 15550 12404
rect 19068 12348 19740 12404
rect 19796 12348 19806 12404
rect 28130 12348 28140 12404
rect 28196 12348 28924 12404
rect 28980 12348 29820 12404
rect 29876 12348 29886 12404
rect 30930 12348 30940 12404
rect 30996 12348 31612 12404
rect 31668 12348 31836 12404
rect 31892 12348 31902 12404
rect 32050 12348 32060 12404
rect 32116 12348 33180 12404
rect 33236 12348 33246 12404
rect 38770 12348 38780 12404
rect 38836 12348 43148 12404
rect 43204 12348 43214 12404
rect 31836 12292 31892 12348
rect 4834 12236 4844 12292
rect 4900 12236 4956 12292
rect 5012 12236 5022 12292
rect 6066 12236 6076 12292
rect 6132 12236 6860 12292
rect 6916 12236 6926 12292
rect 13010 12236 13020 12292
rect 13076 12236 13692 12292
rect 13748 12236 13758 12292
rect 18610 12236 18620 12292
rect 18676 12236 19180 12292
rect 19236 12236 20636 12292
rect 20692 12236 20702 12292
rect 28242 12236 28252 12292
rect 28308 12236 29148 12292
rect 29204 12236 29214 12292
rect 29586 12236 29596 12292
rect 29652 12236 30492 12292
rect 30548 12236 30558 12292
rect 31836 12236 32508 12292
rect 32564 12236 32574 12292
rect 33954 12236 33964 12292
rect 34020 12236 34972 12292
rect 35028 12236 37772 12292
rect 37828 12236 37838 12292
rect 38658 12236 38668 12292
rect 38724 12236 39452 12292
rect 39508 12236 39518 12292
rect 41234 12236 41244 12292
rect 41300 12236 42812 12292
rect 42868 12236 46172 12292
rect 46228 12236 46238 12292
rect 0 12180 800 12208
rect 34636 12180 34692 12236
rect 0 12124 1708 12180
rect 1764 12124 5292 12180
rect 5348 12124 5358 12180
rect 11778 12124 11788 12180
rect 11844 12124 13244 12180
rect 13300 12124 13310 12180
rect 27346 12124 27356 12180
rect 27412 12124 29484 12180
rect 29540 12124 29550 12180
rect 34626 12124 34636 12180
rect 34692 12124 34702 12180
rect 37538 12124 37548 12180
rect 37604 12124 38444 12180
rect 38500 12124 38510 12180
rect 40898 12124 40908 12180
rect 40964 12124 41468 12180
rect 41524 12124 41534 12180
rect 0 12096 800 12124
rect 2594 12012 2604 12068
rect 2660 12012 3276 12068
rect 3332 12012 3342 12068
rect 9986 12012 9996 12068
rect 10052 12012 32060 12068
rect 32116 12012 32126 12068
rect 34178 12012 34188 12068
rect 34244 12012 34748 12068
rect 34804 12012 34972 12068
rect 35028 12012 35038 12068
rect 38098 12012 38108 12068
rect 38164 12012 39116 12068
rect 39172 12012 39182 12068
rect 9996 11956 10052 12012
rect 32060 11956 32116 12012
rect 3378 11900 3388 11956
rect 3444 11900 6860 11956
rect 6916 11900 6926 11956
rect 8642 11900 8652 11956
rect 8708 11900 9100 11956
rect 9156 11900 10052 11956
rect 13010 11900 13020 11956
rect 13076 11900 13580 11956
rect 13636 11900 13646 11956
rect 32060 11900 40572 11956
rect 40628 11900 40638 11956
rect 8978 11788 8988 11844
rect 9044 11788 10108 11844
rect 10164 11788 10174 11844
rect 12338 11788 12348 11844
rect 12404 11788 13580 11844
rect 13636 11788 16604 11844
rect 16660 11788 17388 11844
rect 17444 11788 17454 11844
rect 34066 11788 34076 11844
rect 34132 11788 34524 11844
rect 34580 11788 34590 11844
rect 39890 11788 39900 11844
rect 39956 11788 40460 11844
rect 40516 11788 40526 11844
rect 44706 11788 44716 11844
rect 44772 11788 45724 11844
rect 45780 11788 45790 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 2482 11676 2492 11732
rect 2548 11676 3948 11732
rect 4004 11676 4014 11732
rect 13906 11676 13916 11732
rect 13972 11676 15372 11732
rect 15428 11676 15438 11732
rect 17714 11676 17724 11732
rect 17780 11676 20860 11732
rect 20916 11676 20926 11732
rect 25890 11676 25900 11732
rect 25956 11676 26796 11732
rect 26852 11676 27580 11732
rect 27636 11676 28364 11732
rect 28420 11676 28430 11732
rect 38294 11676 38332 11732
rect 38388 11676 38398 11732
rect 44930 11676 44940 11732
rect 44996 11676 49084 11732
rect 49140 11676 49150 11732
rect 2034 11564 2044 11620
rect 2100 11564 7644 11620
rect 7700 11564 7710 11620
rect 12898 11564 12908 11620
rect 12964 11564 17052 11620
rect 17108 11564 17118 11620
rect 38182 11564 38220 11620
rect 38276 11564 38286 11620
rect 45826 11564 45836 11620
rect 45892 11564 47404 11620
rect 47460 11564 47470 11620
rect 0 11508 800 11536
rect 0 11452 1708 11508
rect 1764 11452 1774 11508
rect 3154 11452 3164 11508
rect 3220 11452 5740 11508
rect 5796 11452 5806 11508
rect 11330 11452 11340 11508
rect 11396 11452 12796 11508
rect 12852 11452 12862 11508
rect 24658 11452 24668 11508
rect 24724 11452 25340 11508
rect 25396 11452 27132 11508
rect 27188 11452 27198 11508
rect 34290 11452 34300 11508
rect 34356 11452 35196 11508
rect 35252 11452 35262 11508
rect 38668 11452 38780 11508
rect 38836 11452 39004 11508
rect 39060 11452 39070 11508
rect 42354 11452 42364 11508
rect 42420 11452 43372 11508
rect 43428 11452 44716 11508
rect 44772 11452 44782 11508
rect 0 11424 800 11452
rect 38668 11396 38724 11452
rect 2706 11340 2716 11396
rect 2772 11340 11452 11396
rect 11508 11340 11518 11396
rect 12226 11340 12236 11396
rect 12292 11340 14028 11396
rect 14084 11340 14094 11396
rect 16594 11340 16604 11396
rect 16660 11340 16940 11396
rect 16996 11340 17006 11396
rect 26002 11340 26012 11396
rect 26068 11340 30268 11396
rect 30324 11340 30334 11396
rect 31266 11340 31276 11396
rect 31332 11340 32172 11396
rect 32228 11340 32238 11396
rect 33618 11340 33628 11396
rect 33684 11340 34860 11396
rect 34916 11340 34926 11396
rect 37090 11340 37100 11396
rect 37156 11340 38332 11396
rect 38388 11340 38398 11396
rect 38546 11340 38556 11396
rect 38612 11340 38724 11396
rect 39778 11340 39788 11396
rect 39844 11340 40348 11396
rect 40404 11340 40414 11396
rect 4946 11228 4956 11284
rect 5012 11228 5628 11284
rect 5684 11228 5694 11284
rect 29138 11228 29148 11284
rect 29204 11228 29932 11284
rect 29988 11228 31500 11284
rect 31556 11228 31566 11284
rect 37762 11228 37772 11284
rect 37828 11228 38332 11284
rect 38388 11228 38668 11284
rect 39666 11228 39676 11284
rect 39732 11228 41468 11284
rect 41524 11228 41534 11284
rect 42242 11228 42252 11284
rect 42308 11228 42700 11284
rect 42756 11228 42766 11284
rect 38612 11172 38668 11228
rect 10658 11116 10668 11172
rect 10724 11116 11900 11172
rect 11956 11116 11966 11172
rect 14690 11116 14700 11172
rect 14756 11116 17164 11172
rect 17220 11116 17230 11172
rect 38406 11116 38444 11172
rect 38500 11116 38510 11172
rect 38612 11116 39900 11172
rect 39956 11116 41020 11172
rect 41076 11116 41804 11172
rect 41860 11116 41870 11172
rect 42354 11116 42364 11172
rect 42420 11116 43484 11172
rect 43540 11116 44156 11172
rect 44212 11116 44222 11172
rect 12450 11004 12460 11060
rect 12516 11004 15148 11060
rect 15092 10948 15148 11004
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 12114 10892 12124 10948
rect 12180 10892 12572 10948
rect 12628 10892 13804 10948
rect 13860 10892 13870 10948
rect 15092 10892 16324 10948
rect 35858 10892 35868 10948
rect 35924 10892 38220 10948
rect 38276 10892 38286 10948
rect 0 10836 800 10864
rect 16268 10836 16324 10892
rect 0 10780 2380 10836
rect 2436 10780 2446 10836
rect 3938 10780 3948 10836
rect 4004 10780 5516 10836
rect 5572 10780 7308 10836
rect 7364 10780 7374 10836
rect 7858 10780 7868 10836
rect 7924 10780 8540 10836
rect 8596 10780 8606 10836
rect 9538 10780 9548 10836
rect 9604 10780 10220 10836
rect 10276 10780 11564 10836
rect 11620 10780 11630 10836
rect 13234 10780 13244 10836
rect 13300 10780 15708 10836
rect 15764 10780 15774 10836
rect 16268 10780 18396 10836
rect 18452 10780 18462 10836
rect 36194 10780 36204 10836
rect 36260 10780 36540 10836
rect 36596 10780 36988 10836
rect 37044 10780 37054 10836
rect 38770 10780 38780 10836
rect 38836 10780 42252 10836
rect 42308 10780 42318 10836
rect 43586 10780 43596 10836
rect 43652 10780 44940 10836
rect 44996 10780 45006 10836
rect 0 10752 800 10780
rect 1698 10668 1708 10724
rect 1764 10668 2492 10724
rect 2548 10668 2558 10724
rect 4386 10668 4396 10724
rect 4452 10668 4956 10724
rect 5012 10668 5964 10724
rect 6020 10668 9660 10724
rect 9716 10668 9726 10724
rect 12786 10668 12796 10724
rect 12852 10668 13916 10724
rect 13972 10668 13982 10724
rect 6514 10556 6524 10612
rect 6580 10556 7084 10612
rect 7140 10556 7868 10612
rect 7924 10556 9548 10612
rect 9604 10556 9614 10612
rect 5618 10444 5628 10500
rect 5684 10444 6188 10500
rect 6244 10444 8428 10500
rect 8484 10444 8494 10500
rect 16268 10388 16324 10780
rect 26114 10668 26124 10724
rect 26180 10668 27244 10724
rect 27300 10668 27310 10724
rect 35410 10668 35420 10724
rect 35476 10668 38220 10724
rect 38276 10668 38668 10724
rect 42130 10668 42140 10724
rect 42196 10668 42812 10724
rect 42868 10668 42878 10724
rect 16594 10556 16604 10612
rect 16660 10556 17388 10612
rect 17444 10556 18396 10612
rect 18452 10556 18462 10612
rect 20738 10444 20748 10500
rect 20804 10444 22092 10500
rect 22148 10444 22158 10500
rect 26786 10444 26796 10500
rect 26852 10444 26908 10668
rect 38612 10612 38668 10668
rect 32386 10556 32396 10612
rect 32452 10556 33180 10612
rect 33236 10556 34524 10612
rect 34580 10556 35756 10612
rect 35812 10556 35822 10612
rect 36082 10556 36092 10612
rect 36148 10556 37324 10612
rect 37380 10556 38108 10612
rect 38164 10556 38174 10612
rect 38612 10556 39004 10612
rect 39060 10556 39070 10612
rect 35970 10444 35980 10500
rect 36036 10444 37100 10500
rect 37156 10444 37884 10500
rect 37940 10444 37950 10500
rect 39778 10444 39788 10500
rect 39844 10444 40796 10500
rect 40852 10444 42812 10500
rect 42868 10444 44044 10500
rect 44100 10444 44110 10500
rect 5170 10332 5180 10388
rect 5236 10332 10444 10388
rect 10500 10332 12460 10388
rect 12516 10332 12526 10388
rect 16258 10332 16268 10388
rect 16324 10332 16334 10388
rect 34066 10332 34076 10388
rect 34132 10332 38444 10388
rect 38500 10332 38668 10388
rect 43362 10332 43372 10388
rect 43428 10332 45836 10388
rect 45892 10332 45902 10388
rect 38612 10276 38668 10332
rect 38612 10220 39228 10276
rect 39284 10220 39294 10276
rect 0 10164 800 10192
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 0 10108 3052 10164
rect 3108 10108 3836 10164
rect 3892 10108 3902 10164
rect 13794 10108 13804 10164
rect 13860 10108 14812 10164
rect 14868 10108 14878 10164
rect 16034 10108 16044 10164
rect 16100 10108 17052 10164
rect 17108 10108 17118 10164
rect 23650 10108 23660 10164
rect 23716 10108 25116 10164
rect 25172 10108 25182 10164
rect 37874 10108 37884 10164
rect 37940 10108 38668 10164
rect 38724 10108 40012 10164
rect 40068 10108 40078 10164
rect 0 10080 800 10108
rect 27234 9996 27244 10052
rect 27300 9996 27804 10052
rect 27860 9996 28812 10052
rect 28868 9996 28878 10052
rect 30034 9996 30044 10052
rect 30100 9996 33068 10052
rect 33124 9996 33134 10052
rect 4274 9884 4284 9940
rect 4340 9884 5516 9940
rect 5572 9884 5582 9940
rect 16370 9884 16380 9940
rect 16436 9884 16828 9940
rect 16884 9884 16894 9940
rect 2034 9772 2044 9828
rect 2100 9772 5068 9828
rect 5124 9772 5134 9828
rect 8754 9772 8764 9828
rect 8820 9772 11788 9828
rect 11844 9772 11854 9828
rect 16706 9772 16716 9828
rect 16772 9772 17724 9828
rect 17780 9772 17790 9828
rect 19058 9772 19068 9828
rect 19124 9772 19852 9828
rect 19908 9772 22652 9828
rect 22708 9772 22718 9828
rect 23874 9772 23884 9828
rect 23940 9772 27020 9828
rect 27076 9772 28028 9828
rect 28084 9772 28094 9828
rect 39442 9772 39452 9828
rect 39508 9772 40908 9828
rect 40964 9772 41132 9828
rect 41188 9772 41198 9828
rect 41570 9772 41580 9828
rect 41636 9772 43484 9828
rect 43540 9772 43550 9828
rect 43922 9772 43932 9828
rect 43988 9772 46508 9828
rect 46564 9772 46574 9828
rect 43932 9716 43988 9772
rect 2706 9660 2716 9716
rect 2772 9660 6076 9716
rect 6132 9660 6142 9716
rect 13682 9660 13692 9716
rect 13748 9660 15148 9716
rect 15204 9660 15214 9716
rect 17490 9660 17500 9716
rect 17556 9660 18172 9716
rect 18228 9660 19404 9716
rect 19460 9660 20076 9716
rect 20132 9660 20142 9716
rect 31378 9660 31388 9716
rect 31444 9660 31836 9716
rect 31892 9660 31902 9716
rect 34514 9660 34524 9716
rect 34580 9660 35756 9716
rect 35812 9660 35822 9716
rect 40114 9660 40124 9716
rect 40180 9660 41244 9716
rect 41300 9660 43988 9716
rect 20738 9548 20748 9604
rect 20804 9548 21868 9604
rect 21924 9548 24668 9604
rect 24724 9548 25228 9604
rect 25284 9548 25294 9604
rect 27906 9548 27916 9604
rect 27972 9548 28588 9604
rect 28644 9548 28654 9604
rect 41682 9548 41692 9604
rect 41748 9548 42140 9604
rect 42196 9548 43708 9604
rect 43764 9548 44828 9604
rect 44884 9548 44894 9604
rect 13010 9436 13020 9492
rect 13076 9436 14476 9492
rect 14532 9436 14542 9492
rect 28242 9436 28252 9492
rect 28308 9436 35084 9492
rect 35140 9436 35150 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 7522 9324 7532 9380
rect 7588 9324 8428 9380
rect 8484 9324 16380 9380
rect 16436 9324 16446 9380
rect 21074 9324 21084 9380
rect 21140 9324 33740 9380
rect 33796 9324 33806 9380
rect 5954 9212 5964 9268
rect 6020 9212 9772 9268
rect 9828 9212 9838 9268
rect 16258 9212 16268 9268
rect 16324 9212 17052 9268
rect 17108 9212 17118 9268
rect 22978 9212 22988 9268
rect 23044 9212 23436 9268
rect 23492 9212 26684 9268
rect 26740 9212 27692 9268
rect 27748 9212 34972 9268
rect 35028 9212 35038 9268
rect 35186 9212 35196 9268
rect 35252 9212 35868 9268
rect 35924 9212 35934 9268
rect 41010 9212 41020 9268
rect 41076 9212 42364 9268
rect 42420 9212 42430 9268
rect 42690 9212 42700 9268
rect 42756 9212 46060 9268
rect 46116 9212 46126 9268
rect 18050 9100 18060 9156
rect 18116 9100 19516 9156
rect 19572 9100 19582 9156
rect 24098 9100 24108 9156
rect 24164 9100 26796 9156
rect 26852 9100 26862 9156
rect 35298 9100 35308 9156
rect 35364 9100 39788 9156
rect 39844 9100 41580 9156
rect 41636 9100 41646 9156
rect 25218 8988 25228 9044
rect 25284 8988 27020 9044
rect 27076 8988 27086 9044
rect 29474 8988 29484 9044
rect 29540 8988 30268 9044
rect 30324 8988 30334 9044
rect 38210 8988 38220 9044
rect 38276 8988 38892 9044
rect 38948 8988 38958 9044
rect 39666 8988 39676 9044
rect 39732 8988 41356 9044
rect 41412 8988 41422 9044
rect 8082 8876 8092 8932
rect 8148 8876 9660 8932
rect 9716 8876 9726 8932
rect 38322 8876 38332 8932
rect 38388 8876 39900 8932
rect 39956 8876 39966 8932
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 5058 8428 5068 8484
rect 5124 8428 7364 8484
rect 9762 8428 9772 8484
rect 9828 8428 11228 8484
rect 11284 8428 11294 8484
rect 12674 8428 12684 8484
rect 12740 8428 15932 8484
rect 15988 8428 15998 8484
rect 33954 8428 33964 8484
rect 34020 8428 35420 8484
rect 35476 8428 35486 8484
rect 39554 8428 39564 8484
rect 39620 8428 39630 8484
rect 7308 8372 7364 8428
rect 12684 8372 12740 8428
rect 14588 8372 14644 8428
rect 39564 8372 39620 8428
rect 7298 8316 7308 8372
rect 7364 8316 7980 8372
rect 8036 8316 8764 8372
rect 8820 8316 8830 8372
rect 10770 8316 10780 8372
rect 10836 8316 12740 8372
rect 14578 8316 14588 8372
rect 14644 8316 14654 8372
rect 39564 8316 41244 8372
rect 41300 8316 41310 8372
rect 9874 8204 9884 8260
rect 9940 8204 12236 8260
rect 12292 8204 13692 8260
rect 13748 8204 13758 8260
rect 18946 8204 18956 8260
rect 19012 8204 19292 8260
rect 19348 8204 20076 8260
rect 20132 8204 20142 8260
rect 31490 8204 31500 8260
rect 31556 8204 33180 8260
rect 33236 8204 33246 8260
rect 10210 8092 10220 8148
rect 10276 8092 10668 8148
rect 10724 8092 10734 8148
rect 41794 8092 41804 8148
rect 41860 8092 42924 8148
rect 42980 8092 42990 8148
rect 10546 7980 10556 8036
rect 10612 7980 12124 8036
rect 12180 7980 12190 8036
rect 12562 7980 12572 8036
rect 12628 7980 13580 8036
rect 13636 7980 13646 8036
rect 37538 7980 37548 8036
rect 37604 7980 38220 8036
rect 38276 7980 38286 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 41346 7756 41356 7812
rect 41412 7756 43036 7812
rect 43092 7756 43102 7812
rect 8978 7644 8988 7700
rect 9044 7644 9772 7700
rect 9828 7644 9838 7700
rect 33170 7644 33180 7700
rect 33236 7644 35532 7700
rect 35588 7644 36428 7700
rect 36484 7644 36876 7700
rect 36932 7644 40124 7700
rect 40180 7644 42700 7700
rect 42756 7644 42766 7700
rect 16370 7420 16380 7476
rect 16436 7420 18508 7476
rect 18564 7420 18574 7476
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 18050 6524 18060 6580
rect 18116 6524 18284 6580
rect 18340 6524 18350 6580
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 35074 4956 35084 5012
rect 35140 4956 36652 5012
rect 36708 4956 36718 5012
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 17826 3948 17836 4004
rect 17892 3948 18396 4004
rect 18452 3948 18462 4004
rect 38658 3948 38668 4004
rect 38724 3948 46284 4004
rect 46340 3948 46350 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 18022 3724 18060 3780
rect 18116 3724 18126 3780
rect 34738 3724 34748 3780
rect 34804 3724 49532 3780
rect 49588 3724 49598 3780
rect 35410 3612 35420 3668
rect 35476 3612 36092 3668
rect 36148 3612 36158 3668
rect 32946 3500 32956 3556
rect 33012 3500 33516 3556
rect 33572 3500 33582 3556
rect 36306 3500 36316 3556
rect 36372 3500 37100 3556
rect 37156 3500 37548 3556
rect 37604 3500 37614 3556
rect 37874 3500 37884 3556
rect 37940 3500 39004 3556
rect 39060 3500 39070 3556
rect 18162 3388 18172 3444
rect 18228 3388 18620 3444
rect 18676 3388 18686 3444
rect 29596 3388 30268 3444
rect 30324 3388 30334 3444
rect 35186 3388 35196 3444
rect 35252 3388 35756 3444
rect 35812 3388 36204 3444
rect 36260 3388 36270 3444
rect 39890 3388 39900 3444
rect 39956 3388 40348 3444
rect 40404 3388 40684 3444
rect 40740 3388 40750 3444
rect 29596 3332 29652 3388
rect 29586 3276 29596 3332
rect 29652 3276 29662 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 22540 46844 22596 46900
rect 16380 46620 16436 46676
rect 50988 46508 51044 46564
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 25004 44604 25060 44660
rect 50988 44380 51044 44436
rect 16380 44268 16436 44324
rect 21980 44156 22036 44212
rect 51436 44044 51492 44100
rect 50988 43932 51044 43988
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 28924 43820 28980 43876
rect 50988 43596 51044 43652
rect 22540 43260 22596 43316
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 51436 43036 51492 43092
rect 50988 42812 51044 42868
rect 42252 42700 42308 42756
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 35868 42252 35924 42308
rect 26684 42140 26740 42196
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 42252 42028 42308 42084
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19404 41020 19460 41076
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 19404 40684 19460 40740
rect 26684 40572 26740 40628
rect 35644 40572 35700 40628
rect 25004 40460 25060 40516
rect 21868 40348 21924 40404
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 30828 39788 30884 39844
rect 21980 39228 22036 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 30268 39004 30324 39060
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 36652 38892 36708 38948
rect 35644 38668 35700 38724
rect 42252 38668 42308 38724
rect 28924 38444 28980 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 36652 37324 36708 37380
rect 21868 37212 21924 37268
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 35868 36316 35924 36372
rect 30268 36092 30324 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 30492 35980 30548 36036
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 46508 35756 46564 35812
rect 30828 35644 30884 35700
rect 30268 35532 30324 35588
rect 30492 35420 30548 35476
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 31724 35084 31780 35140
rect 27580 34860 27636 34916
rect 42028 34860 42084 34916
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 34412 34300 34468 34356
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 48748 33628 48804 33684
rect 31052 33516 31108 33572
rect 22540 33180 22596 33236
rect 39676 33180 39732 33236
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 14588 32732 14644 32788
rect 42252 32284 42308 32340
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 22540 31500 22596 31556
rect 31724 31500 31780 31556
rect 39676 31388 39732 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 46060 31052 46116 31108
rect 34188 30940 34244 30996
rect 36764 30940 36820 30996
rect 36540 30716 36596 30772
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 22540 30380 22596 30436
rect 34860 30156 34916 30212
rect 34188 30044 34244 30100
rect 19516 29932 19572 29988
rect 36428 29820 36484 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 14588 29708 14644 29764
rect 36652 29708 36708 29764
rect 34412 29484 34468 29540
rect 36316 29372 36372 29428
rect 46732 29148 46788 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 20188 28700 20244 28756
rect 34860 28700 34916 28756
rect 36764 28700 36820 28756
rect 36540 28476 36596 28532
rect 36316 28364 36372 28420
rect 36652 28364 36708 28420
rect 46396 28364 46452 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 31052 28028 31108 28084
rect 46396 27580 46452 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 31724 26684 31780 26740
rect 46060 26684 46116 26740
rect 46732 26684 46788 26740
rect 48748 26684 48804 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 42028 26460 42084 26516
rect 50988 26236 51044 26292
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 36428 25004 36484 25060
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19516 24108 19572 24164
rect 20188 23996 20244 24052
rect 27580 23884 27636 23940
rect 46508 23884 46564 23940
rect 50988 23884 51044 23940
rect 42252 23548 42308 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 9884 23436 9940 23492
rect 11564 23436 11620 23492
rect 11788 23324 11844 23380
rect 34972 23324 35028 23380
rect 31388 23212 31444 23268
rect 31724 22988 31780 23044
rect 34412 22876 34468 22932
rect 34972 22876 35028 22932
rect 11564 22764 11620 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 9436 22428 9492 22484
rect 34412 22092 34468 22148
rect 38220 22092 38276 22148
rect 42140 22092 42196 22148
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 31388 21420 31444 21476
rect 9436 21308 9492 21364
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 27020 21084 27076 21140
rect 3836 20748 3892 20804
rect 46620 20748 46676 20804
rect 33068 20524 33124 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 7644 20300 7700 20356
rect 16156 20300 16212 20356
rect 11788 20076 11844 20132
rect 34188 19964 34244 20020
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 31724 19292 31780 19348
rect 3836 19180 3892 19236
rect 9884 19180 9940 19236
rect 15708 19068 15764 19124
rect 26908 19068 26964 19124
rect 15708 18844 15764 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 38556 18956 38612 19012
rect 11676 18620 11732 18676
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 36764 18508 36820 18564
rect 7644 18172 7700 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 26908 17612 26964 17668
rect 33404 17612 33460 17668
rect 36764 17612 36820 17668
rect 51212 17388 51268 17444
rect 11340 17276 11396 17332
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 11676 17052 11732 17108
rect 26908 17052 26964 17108
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 36316 16380 36372 16436
rect 37548 16268 37604 16324
rect 27020 16044 27076 16100
rect 11340 15932 11396 15988
rect 33068 15932 33124 15988
rect 51212 15820 51268 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 34188 15036 34244 15092
rect 16156 14924 16212 14980
rect 37548 14924 37604 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 36316 14812 36372 14868
rect 46620 14588 46676 14644
rect 38444 14476 38500 14532
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 7644 13804 7700 13860
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 4956 13020 5012 13076
rect 42140 12684 42196 12740
rect 33404 12572 33460 12628
rect 13580 12460 13636 12516
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 38556 12460 38612 12516
rect 4956 12236 5012 12292
rect 13580 11900 13636 11956
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 38332 11676 38388 11732
rect 38220 11564 38276 11620
rect 38332 11228 38388 11284
rect 38444 11116 38500 11172
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 18060 6524 18116 6580
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 18060 3724 18116 3780
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 16380 46676 16436 46686
rect 16380 44324 16436 46620
rect 16380 44258 16436 44268
rect 19808 45500 20128 47012
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 19808 43932 20128 45444
rect 22540 46900 22596 46910
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19404 41076 19460 41086
rect 19404 40740 19460 41020
rect 19404 40674 19460 40684
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 19808 39228 20128 40740
rect 21980 44212 22036 44222
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 21868 40404 21924 40414
rect 21868 37268 21924 40348
rect 21980 39284 22036 44156
rect 22540 43316 22596 46844
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 22540 43250 22596 43260
rect 25004 44660 25060 44670
rect 25004 40516 25060 44604
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 28924 43876 28980 43886
rect 26684 42196 26740 42206
rect 26684 40628 26740 42140
rect 26684 40562 26740 40572
rect 25004 40450 25060 40460
rect 21980 39218 22036 39228
rect 28924 38500 28980 43820
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50988 46564 51044 46574
rect 50988 44436 51044 46508
rect 50988 43988 51044 44380
rect 50988 43922 51044 43932
rect 51436 44100 51492 44110
rect 42252 42756 42308 42766
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35868 42308 35924 42318
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 30828 39844 30884 39854
rect 28924 38434 28980 38444
rect 30268 39060 30324 39070
rect 21868 37202 21924 37212
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 30268 36148 30324 39004
rect 30268 35588 30324 36092
rect 30268 35522 30324 35532
rect 30492 36036 30548 36046
rect 30492 35476 30548 35980
rect 30828 35700 30884 39788
rect 30828 35634 30884 35644
rect 35168 38444 35488 39956
rect 35644 40628 35700 40638
rect 35644 38724 35700 40572
rect 35644 38658 35700 38668
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 30492 35410 30548 35420
rect 35168 35308 35488 36820
rect 35868 36372 35924 42252
rect 42252 42084 42308 42700
rect 36652 38948 36708 38958
rect 36652 37380 36708 38892
rect 42252 38724 42308 42028
rect 42252 38658 42308 38668
rect 50528 42364 50848 43876
rect 50988 43652 51044 43662
rect 50988 42868 51044 43596
rect 51436 43092 51492 44044
rect 51436 43026 51492 43036
rect 50988 42802 51044 42812
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 36652 37314 36708 37324
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 35868 36306 35924 36316
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 31724 35140 31780 35150
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 27580 34916 27636 34926
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 14588 32788 14644 32798
rect 14588 29764 14644 32732
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 14588 29698 14644 29708
rect 19516 29988 19572 29998
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 19516 24164 19572 29932
rect 19516 24098 19572 24108
rect 19808 29820 20128 31332
rect 22540 33236 22596 33246
rect 22540 31556 22596 33180
rect 22540 30436 22596 31500
rect 22540 30370 22596 30380
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 20188 28756 20244 28766
rect 20188 24052 20244 28700
rect 20188 23986 20244 23996
rect 27580 23940 27636 34860
rect 31052 33572 31108 33582
rect 31052 28084 31108 33516
rect 31052 28018 31108 28028
rect 31724 31556 31780 35084
rect 31724 26740 31780 31500
rect 34412 34356 34468 34366
rect 34188 30996 34244 31006
rect 34188 30100 34244 30940
rect 34188 30034 34244 30044
rect 34412 29540 34468 34300
rect 35168 33740 35488 35252
rect 46508 35812 46564 35822
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 42028 34916 42084 34926
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 39676 33236 39732 33246
rect 39676 31444 39732 33180
rect 39676 31378 39732 31388
rect 36764 30996 36820 31006
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 34412 29474 34468 29484
rect 34860 30212 34916 30222
rect 34860 28756 34916 30156
rect 34860 28690 34916 28700
rect 35168 29036 35488 30548
rect 36540 30772 36596 30782
rect 36428 29876 36484 29886
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 31724 26674 31780 26684
rect 35168 27468 35488 28980
rect 36316 29428 36372 29438
rect 36316 28420 36372 29372
rect 36316 28354 36372 28364
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 27580 23874 27636 23884
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 36428 25060 36484 29820
rect 36540 28532 36596 30716
rect 36540 28466 36596 28476
rect 36652 29764 36708 29774
rect 36652 28420 36708 29708
rect 36764 28756 36820 30940
rect 36764 28690 36820 28700
rect 36652 28354 36708 28364
rect 42028 26516 42084 34860
rect 42028 26450 42084 26460
rect 42252 32340 42308 32350
rect 36428 24994 36484 25004
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 9884 23492 9940 23502
rect 9436 22484 9492 22494
rect 9436 21364 9492 22428
rect 9436 21298 9492 21308
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 3836 20804 3892 20814
rect 3836 19236 3892 20748
rect 3836 19170 3892 19180
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 7644 20356 7700 20366
rect 7644 18228 7700 20300
rect 9884 19236 9940 23436
rect 11564 23492 11620 23502
rect 11564 22820 11620 23436
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 11564 22754 11620 22764
rect 11788 23380 11844 23390
rect 11788 20132 11844 23324
rect 19808 21980 20128 23492
rect 34972 23380 35028 23390
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 31388 23268 31444 23278
rect 31388 21476 31444 23212
rect 31388 21410 31444 21420
rect 31724 23044 31780 23054
rect 11788 20066 11844 20076
rect 16156 20356 16212 20366
rect 9884 19170 9940 19180
rect 15708 19124 15764 19134
rect 15708 18900 15764 19068
rect 15708 18834 15764 18844
rect 7644 13860 7700 18172
rect 11676 18676 11732 18686
rect 11340 17332 11396 17342
rect 11340 15988 11396 17276
rect 11676 17108 11732 18620
rect 11676 17042 11732 17052
rect 11340 15922 11396 15932
rect 16156 14980 16212 20300
rect 16156 14914 16212 14924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 27020 21140 27076 21150
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 26908 19124 26964 19134
rect 26908 17668 26964 19068
rect 26908 17108 26964 17612
rect 26908 17042 26964 17052
rect 27020 16100 27076 21084
rect 31724 19348 31780 22988
rect 34412 22932 34468 22942
rect 34412 22148 34468 22876
rect 34972 22932 35028 23324
rect 34972 22866 35028 22876
rect 34412 22082 34468 22092
rect 35168 22764 35488 24276
rect 42252 23604 42308 32284
rect 46060 31108 46116 31118
rect 46060 26740 46116 31052
rect 46396 28420 46452 28430
rect 46396 27636 46452 28364
rect 46396 27570 46452 27580
rect 46060 26674 46116 26684
rect 46508 23940 46564 35756
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 48748 33684 48804 33694
rect 46732 29204 46788 29214
rect 46732 26740 46788 29148
rect 46732 26674 46788 26684
rect 48748 26740 48804 33628
rect 48748 26674 48804 26684
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 46508 23874 46564 23884
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 42252 23538 42308 23548
rect 50528 23548 50848 25060
rect 50988 26292 51044 26302
rect 50988 23940 51044 26236
rect 50988 23874 51044 23884
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 31724 19282 31780 19292
rect 33068 20580 33124 20590
rect 27020 16034 27076 16044
rect 33068 15988 33124 20524
rect 34188 20020 34244 20030
rect 33068 15922 33124 15932
rect 33404 17668 33460 17678
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 7644 13794 7700 13804
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4956 13076 5012 13086
rect 4956 12292 5012 13020
rect 19808 12572 20128 14084
rect 4956 12226 5012 12236
rect 13580 12516 13636 12526
rect 13580 11956 13636 12460
rect 13580 11890 13636 11900
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 33404 12628 33460 17612
rect 34188 15092 34244 19964
rect 34188 15026 34244 15036
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 38220 22148 38276 22158
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 36764 18564 36820 18574
rect 36764 17668 36820 18508
rect 36764 17602 36820 17612
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 33404 12562 33460 12572
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 36316 16436 36372 16446
rect 36316 14868 36372 16380
rect 37548 16324 37604 16334
rect 37548 14980 37604 16268
rect 37548 14914 37604 14924
rect 36316 14802 36372 14812
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 18060 6580 18116 6590
rect 18060 3780 18116 6524
rect 18060 3714 18116 3724
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 38220 11620 38276 22092
rect 42140 22148 42196 22158
rect 38556 19012 38612 19022
rect 38444 14532 38500 14542
rect 38220 11554 38276 11564
rect 38332 11732 38388 11742
rect 38332 11284 38388 11676
rect 38332 11218 38388 11228
rect 38444 11172 38500 14476
rect 38556 12516 38612 18956
rect 42140 12740 42196 22092
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 46620 20804 46676 20814
rect 46620 14644 46676 20748
rect 46620 14578 46676 14588
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 51212 17444 51268 17454
rect 51212 15876 51268 17388
rect 51212 15810 51268 15820
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 42140 12674 42196 12684
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 38556 12450 38612 12460
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 38444 11106 38500 11116
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1424_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11872 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1425_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31472 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1426_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32144 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1427_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10976 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1428_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7616 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1429_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8512 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1430_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11088 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1431_
timestamp 1698431365
transform -1 0 10864 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1432_
timestamp 1698431365
transform 1 0 28000 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1433_
timestamp 1698431365
transform 1 0 30128 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1434_
timestamp 1698431365
transform 1 0 20496 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1435_
timestamp 1698431365
transform 1 0 32032 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1436_
timestamp 1698431365
transform -1 0 38528 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1437_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20496 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1438_
timestamp 1698431365
transform -1 0 19264 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1439_
timestamp 1698431365
transform 1 0 37072 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1440_
timestamp 1698431365
transform -1 0 30912 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1441_
timestamp 1698431365
transform 1 0 30128 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1442_
timestamp 1698431365
transform 1 0 28896 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1443_
timestamp 1698431365
transform 1 0 27216 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1444_
timestamp 1698431365
transform -1 0 31808 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1445_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29680 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1446_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11200 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1447_
timestamp 1698431365
transform 1 0 33824 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1448_
timestamp 1698431365
transform -1 0 35392 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1449_
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1450_
timestamp 1698431365
transform -1 0 32704 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1451_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31360 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1452_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32144 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1453_
timestamp 1698431365
transform 1 0 20160 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1454_
timestamp 1698431365
transform 1 0 35728 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1455_
timestamp 1698431365
transform -1 0 36512 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1456_
timestamp 1698431365
transform 1 0 20272 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1457_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20272 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1458_
timestamp 1698431365
transform -1 0 34272 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1459_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30128 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1460_
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1461_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20272 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1462_
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1463_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1464_
timestamp 1698431365
transform -1 0 29680 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1465_
timestamp 1698431365
transform 1 0 41104 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1466_
timestamp 1698431365
transform -1 0 40096 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1467_
timestamp 1698431365
transform -1 0 30688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1468_
timestamp 1698431365
transform 1 0 41664 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1469_
timestamp 1698431365
transform 1 0 30464 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1470_
timestamp 1698431365
transform 1 0 30688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1471_
timestamp 1698431365
transform 1 0 29456 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1472_
timestamp 1698431365
transform -1 0 34944 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1473_
timestamp 1698431365
transform -1 0 20944 0 1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1474_
timestamp 1698431365
transform 1 0 21616 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1475_
timestamp 1698431365
transform 1 0 26880 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1476_
timestamp 1698431365
transform 1 0 27664 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1477_
timestamp 1698431365
transform 1 0 29232 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1478_
timestamp 1698431365
transform -1 0 29904 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1479_
timestamp 1698431365
transform 1 0 29008 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1480_
timestamp 1698431365
transform -1 0 29008 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1481_
timestamp 1698431365
transform 1 0 27888 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1482_
timestamp 1698431365
transform 1 0 29344 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1483_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19712 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1484_
timestamp 1698431365
transform -1 0 23072 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1485_
timestamp 1698431365
transform 1 0 22512 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1486_
timestamp 1698431365
transform 1 0 23856 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1487_
timestamp 1698431365
transform 1 0 22400 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1488_
timestamp 1698431365
transform 1 0 24192 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1489_
timestamp 1698431365
transform 1 0 24192 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1490_
timestamp 1698431365
transform 1 0 25312 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1491_
timestamp 1698431365
transform -1 0 35840 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1492_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25872 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1493_
timestamp 1698431365
transform -1 0 26992 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1494_
timestamp 1698431365
transform -1 0 26432 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1495_
timestamp 1698431365
transform 1 0 20944 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1496_
timestamp 1698431365
transform 1 0 21952 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1497_
timestamp 1698431365
transform 1 0 22176 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1498_
timestamp 1698431365
transform -1 0 23744 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1499_
timestamp 1698431365
transform 1 0 23296 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1500_
timestamp 1698431365
transform 1 0 23072 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1501_
timestamp 1698431365
transform 1 0 23408 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1502_
timestamp 1698431365
transform 1 0 27776 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1503_
timestamp 1698431365
transform 1 0 26096 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1504_
timestamp 1698431365
transform -1 0 27216 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1505_
timestamp 1698431365
transform -1 0 27440 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1506_
timestamp 1698431365
transform -1 0 24192 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1507_
timestamp 1698431365
transform 1 0 37632 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1508_
timestamp 1698431365
transform -1 0 44240 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1509_
timestamp 1698431365
transform 1 0 23408 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1510_
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1511_
timestamp 1698431365
transform 1 0 25088 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1512_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1513_
timestamp 1698431365
transform 1 0 27776 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1514_
timestamp 1698431365
transform -1 0 28784 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1515_
timestamp 1698431365
transform 1 0 28672 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1516_
timestamp 1698431365
transform 1 0 27552 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1517_
timestamp 1698431365
transform 1 0 34496 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1518_
timestamp 1698431365
transform 1 0 37520 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1519_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26656 0 1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1520_
timestamp 1698431365
transform -1 0 39088 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1521_
timestamp 1698431365
transform 1 0 36848 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1522_
timestamp 1698431365
transform 1 0 25984 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1523_
timestamp 1698431365
transform 1 0 32928 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1524_
timestamp 1698431365
transform -1 0 37632 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1525_
timestamp 1698431365
transform -1 0 46032 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1526_
timestamp 1698431365
transform 1 0 35840 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1527_
timestamp 1698431365
transform 1 0 36736 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1528_
timestamp 1698431365
transform 1 0 37184 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1529_
timestamp 1698431365
transform 1 0 35616 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1530_
timestamp 1698431365
transform -1 0 35616 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1531_
timestamp 1698431365
transform 1 0 24080 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1532_
timestamp 1698431365
transform 1 0 34608 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1533_
timestamp 1698431365
transform 1 0 35952 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1534_
timestamp 1698431365
transform 1 0 33824 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1535_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34720 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1536_
timestamp 1698431365
transform 1 0 33824 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1537_
timestamp 1698431365
transform -1 0 33600 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1538_
timestamp 1698431365
transform 1 0 35392 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1539_
timestamp 1698431365
transform 1 0 32032 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1540_
timestamp 1698431365
transform 1 0 33824 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1541_
timestamp 1698431365
transform 1 0 32032 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1542_
timestamp 1698431365
transform 1 0 34272 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1543_
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1544_
timestamp 1698431365
transform 1 0 34272 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1545_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34384 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1546_
timestamp 1698431365
transform -1 0 33600 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1547_
timestamp 1698431365
transform -1 0 32704 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1548_
timestamp 1698431365
transform 1 0 32704 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1549_
timestamp 1698431365
transform 1 0 36960 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1550_
timestamp 1698431365
transform -1 0 36960 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1551_
timestamp 1698431365
transform -1 0 34944 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1552_
timestamp 1698431365
transform 1 0 34944 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1553_
timestamp 1698431365
transform -1 0 36288 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1554_
timestamp 1698431365
transform 1 0 34944 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1555_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36064 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1556_
timestamp 1698431365
transform -1 0 34608 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1557_
timestamp 1698431365
transform 1 0 34608 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1558_
timestamp 1698431365
transform -1 0 32704 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1559_
timestamp 1698431365
transform 1 0 31024 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1560_
timestamp 1698431365
transform -1 0 33824 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1561_
timestamp 1698431365
transform -1 0 34944 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1562_
timestamp 1698431365
transform -1 0 36064 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1563_
timestamp 1698431365
transform 1 0 31360 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1564_
timestamp 1698431365
transform 1 0 33040 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1565_
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1566_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43232 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1567_
timestamp 1698431365
transform -1 0 36400 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1568_
timestamp 1698431365
transform -1 0 36512 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1569_
timestamp 1698431365
transform -1 0 35728 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1570_
timestamp 1698431365
transform 1 0 33936 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1571_
timestamp 1698431365
transform 1 0 42896 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1572_
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1573_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1574_
timestamp 1698431365
transform 1 0 36400 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1575_
timestamp 1698431365
transform 1 0 41104 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1576_
timestamp 1698431365
transform 1 0 40992 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1577_
timestamp 1698431365
transform 1 0 41440 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1578_
timestamp 1698431365
transform 1 0 41552 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1579_
timestamp 1698431365
transform -1 0 46256 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1580_
timestamp 1698431365
transform -1 0 36624 0 1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1581_
timestamp 1698431365
transform 1 0 40096 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1582_
timestamp 1698431365
transform 1 0 41328 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1583_
timestamp 1698431365
transform 1 0 41104 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1584_
timestamp 1698431365
transform -1 0 43120 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1585_
timestamp 1698431365
transform -1 0 34944 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1586_
timestamp 1698431365
transform -1 0 40544 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1587_
timestamp 1698431365
transform 1 0 40544 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1588_
timestamp 1698431365
transform -1 0 42448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1589_
timestamp 1698431365
transform 1 0 42560 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1590_
timestamp 1698431365
transform 1 0 42784 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1591_
timestamp 1698431365
transform 1 0 41888 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1592_
timestamp 1698431365
transform 1 0 41440 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1593_
timestamp 1698431365
transform -1 0 43120 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1594_
timestamp 1698431365
transform 1 0 41664 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1595_
timestamp 1698431365
transform -1 0 47264 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1596_
timestamp 1698431365
transform -1 0 42000 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1597_
timestamp 1698431365
transform 1 0 36736 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1598_
timestamp 1698431365
transform 1 0 41216 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1599_
timestamp 1698431365
transform -1 0 43344 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1600_
timestamp 1698431365
transform 1 0 42000 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1601_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1602_
timestamp 1698431365
transform -1 0 44016 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1603_
timestamp 1698431365
transform -1 0 44128 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1604_
timestamp 1698431365
transform 1 0 42672 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1605_
timestamp 1698431365
transform 1 0 41888 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1606_
timestamp 1698431365
transform -1 0 43568 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1607_
timestamp 1698431365
transform -1 0 43008 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1608_
timestamp 1698431365
transform 1 0 37968 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1609_
timestamp 1698431365
transform -1 0 48048 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1610_
timestamp 1698431365
transform -1 0 43680 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1611_
timestamp 1698431365
transform 1 0 43680 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1612_
timestamp 1698431365
transform 1 0 31808 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1613_
timestamp 1698431365
transform -1 0 44016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1614_
timestamp 1698431365
transform -1 0 43568 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1615_
timestamp 1698431365
transform 1 0 43568 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1616_
timestamp 1698431365
transform 1 0 45024 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1617_
timestamp 1698431365
transform -1 0 46032 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1618_
timestamp 1698431365
transform -1 0 49728 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1619_
timestamp 1698431365
transform -1 0 46816 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1620_
timestamp 1698431365
transform -1 0 50624 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1621_
timestamp 1698431365
transform 1 0 45136 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1622_
timestamp 1698431365
transform 1 0 47712 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1698431365
transform 1 0 46144 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1624_
timestamp 1698431365
transform -1 0 46480 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1625_
timestamp 1698431365
transform 1 0 46368 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1626_
timestamp 1698431365
transform -1 0 47824 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1627_
timestamp 1698431365
transform -1 0 44688 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1628_
timestamp 1698431365
transform 1 0 44912 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1629_
timestamp 1698431365
transform -1 0 46592 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1630_
timestamp 1698431365
transform 1 0 45584 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1631_
timestamp 1698431365
transform -1 0 47712 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1632_
timestamp 1698431365
transform 1 0 51408 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1633_
timestamp 1698431365
transform 1 0 46256 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1634_
timestamp 1698431365
transform -1 0 47376 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1635_
timestamp 1698431365
transform 1 0 46480 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1636_
timestamp 1698431365
transform -1 0 49280 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1637_
timestamp 1698431365
transform 1 0 47264 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1638_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46928 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1639_
timestamp 1698431365
transform -1 0 48272 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1640_
timestamp 1698431365
transform 1 0 47264 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1641_
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1642_
timestamp 1698431365
transform -1 0 50176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1643_
timestamp 1698431365
transform 1 0 46592 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1644_
timestamp 1698431365
transform -1 0 47824 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1645_
timestamp 1698431365
transform 1 0 47824 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1646_
timestamp 1698431365
transform 1 0 48384 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1647_
timestamp 1698431365
transform 1 0 45584 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1648_
timestamp 1698431365
transform 1 0 46816 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1649_
timestamp 1698431365
transform 1 0 47376 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1650_
timestamp 1698431365
transform -1 0 48272 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1651_
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1652_
timestamp 1698431365
transform -1 0 49952 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1653_
timestamp 1698431365
transform 1 0 32256 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1654_
timestamp 1698431365
transform 1 0 47040 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1655_
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1656_
timestamp 1698431365
transform 1 0 48608 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1657_
timestamp 1698431365
transform -1 0 49616 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1658_
timestamp 1698431365
transform 1 0 48944 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1659_
timestamp 1698431365
transform -1 0 50848 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1660_
timestamp 1698431365
transform -1 0 49616 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1661_
timestamp 1698431365
transform 1 0 47264 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1662_
timestamp 1698431365
transform 1 0 50624 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1663_
timestamp 1698431365
transform -1 0 53200 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1664_
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1665_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48944 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1666_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44912 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1667_
timestamp 1698431365
transform 1 0 52864 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1668_
timestamp 1698431365
transform -1 0 50960 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1669_
timestamp 1698431365
transform 1 0 50960 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1670_
timestamp 1698431365
transform 1 0 33264 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1671_
timestamp 1698431365
transform 1 0 52080 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1672_
timestamp 1698431365
transform 1 0 54320 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1673_
timestamp 1698431365
transform 1 0 51968 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1674_
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1675_
timestamp 1698431365
transform -1 0 52640 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1676_
timestamp 1698431365
transform -1 0 53984 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1677_
timestamp 1698431365
transform 1 0 52752 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1678_
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1679_
timestamp 1698431365
transform 1 0 51632 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1680_
timestamp 1698431365
transform 1 0 52080 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1681_
timestamp 1698431365
transform -1 0 52416 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1682_
timestamp 1698431365
transform 1 0 50960 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1683_
timestamp 1698431365
transform 1 0 50848 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1684_
timestamp 1698431365
transform 1 0 51408 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1685_
timestamp 1698431365
transform -1 0 51184 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1686_
timestamp 1698431365
transform 1 0 51744 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1687_
timestamp 1698431365
transform -1 0 50176 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1688_
timestamp 1698431365
transform -1 0 52864 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1689_
timestamp 1698431365
transform 1 0 51072 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1690_
timestamp 1698431365
transform 1 0 51072 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1691_
timestamp 1698431365
transform 1 0 50176 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1692_
timestamp 1698431365
transform 1 0 51184 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1693_
timestamp 1698431365
transform 1 0 51408 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1694_
timestamp 1698431365
transform -1 0 53872 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1695_
timestamp 1698431365
transform -1 0 52752 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1696_
timestamp 1698431365
transform 1 0 51408 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1697_
timestamp 1698431365
transform 1 0 39872 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1698_
timestamp 1698431365
transform -1 0 51296 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1699_
timestamp 1698431365
transform 1 0 39424 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1700_
timestamp 1698431365
transform 1 0 39648 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1701_
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1702_
timestamp 1698431365
transform 1 0 39200 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1703_
timestamp 1698431365
transform -1 0 52304 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1704_
timestamp 1698431365
transform -1 0 40432 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1705_
timestamp 1698431365
transform 1 0 39200 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1706_
timestamp 1698431365
transform -1 0 41104 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1707_
timestamp 1698431365
transform -1 0 40208 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1708_
timestamp 1698431365
transform 1 0 38528 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1709_
timestamp 1698431365
transform 1 0 39984 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1710_
timestamp 1698431365
transform 1 0 38640 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1711_
timestamp 1698431365
transform 1 0 39200 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1712_
timestamp 1698431365
transform -1 0 39872 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1713_
timestamp 1698431365
transform -1 0 39200 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1714_
timestamp 1698431365
transform -1 0 40096 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1715_
timestamp 1698431365
transform -1 0 39200 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1716_
timestamp 1698431365
transform 1 0 25760 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1717_
timestamp 1698431365
transform -1 0 27104 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1718_
timestamp 1698431365
transform -1 0 26544 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1719_
timestamp 1698431365
transform 1 0 26544 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1720_
timestamp 1698431365
transform 1 0 29456 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1721_
timestamp 1698431365
transform -1 0 39872 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1722_
timestamp 1698431365
transform -1 0 29008 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1723_
timestamp 1698431365
transform -1 0 28448 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1724_
timestamp 1698431365
transform 1 0 26096 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1725_
timestamp 1698431365
transform -1 0 30128 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1726_
timestamp 1698431365
transform 1 0 30128 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1727_
timestamp 1698431365
transform 1 0 29120 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1728_
timestamp 1698431365
transform 1 0 26656 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1729_
timestamp 1698431365
transform 1 0 26768 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1730_
timestamp 1698431365
transform 1 0 28896 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1731_
timestamp 1698431365
transform -1 0 30576 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1732_
timestamp 1698431365
transform 1 0 25536 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1733_
timestamp 1698431365
transform -1 0 18032 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1734_
timestamp 1698431365
transform -1 0 25872 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1735_
timestamp 1698431365
transform 1 0 24192 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1736_
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1737_
timestamp 1698431365
transform 1 0 21952 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1738_
timestamp 1698431365
transform 1 0 23968 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1739_
timestamp 1698431365
transform -1 0 30128 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1740_
timestamp 1698431365
transform 1 0 25312 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1741_
timestamp 1698431365
transform -1 0 26432 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1742_
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1743_
timestamp 1698431365
transform 1 0 21728 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1744_
timestamp 1698431365
transform 1 0 23520 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1745_
timestamp 1698431365
transform 1 0 23184 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1746_
timestamp 1698431365
transform 1 0 26880 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1747_
timestamp 1698431365
transform 1 0 25424 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1748_
timestamp 1698431365
transform 1 0 28000 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1749_
timestamp 1698431365
transform 1 0 27888 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1750_
timestamp 1698431365
transform 1 0 17584 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1751_
timestamp 1698431365
transform 1 0 22848 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1752_
timestamp 1698431365
transform -1 0 20384 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1753_
timestamp 1698431365
transform 1 0 21168 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1754_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18592 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1755_
timestamp 1698431365
transform 1 0 19264 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1756_
timestamp 1698431365
transform 1 0 19376 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1757_
timestamp 1698431365
transform 1 0 18368 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1758_
timestamp 1698431365
transform 1 0 19376 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1759_
timestamp 1698431365
transform -1 0 19376 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1760_
timestamp 1698431365
transform 1 0 17920 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1761_
timestamp 1698431365
transform -1 0 17920 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1762_
timestamp 1698431365
transform 1 0 22624 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1763_
timestamp 1698431365
transform 1 0 31248 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1764_
timestamp 1698431365
transform 1 0 31808 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1698431365
transform 1 0 34048 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1766_
timestamp 1698431365
transform 1 0 33824 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1767_
timestamp 1698431365
transform 1 0 4928 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1768_
timestamp 1698431365
transform 1 0 4480 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1769_
timestamp 1698431365
transform 1 0 7952 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1770_
timestamp 1698431365
transform -1 0 9072 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1771_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7952 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1772_
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1773_
timestamp 1698431365
transform 1 0 5152 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1774_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4144 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1775_
timestamp 1698431365
transform 1 0 3696 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1776_
timestamp 1698431365
transform 1 0 3360 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1777_
timestamp 1698431365
transform 1 0 4480 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1778_
timestamp 1698431365
transform 1 0 6160 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1779_
timestamp 1698431365
transform 1 0 5936 0 1 40768
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1780_
timestamp 1698431365
transform -1 0 6720 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1781_
timestamp 1698431365
transform 1 0 5600 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1782_
timestamp 1698431365
transform 1 0 7168 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1783_
timestamp 1698431365
transform -1 0 6272 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1784_
timestamp 1698431365
transform -1 0 6272 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1785_
timestamp 1698431365
transform 1 0 5600 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1786_
timestamp 1698431365
transform 1 0 6832 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1787_
timestamp 1698431365
transform 1 0 11760 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1788_
timestamp 1698431365
transform -1 0 13104 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1789_
timestamp 1698431365
transform 1 0 11872 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1790_
timestamp 1698431365
transform -1 0 18144 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1791_
timestamp 1698431365
transform 1 0 17584 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1792_
timestamp 1698431365
transform 1 0 25312 0 -1 54880
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1793_
timestamp 1698431365
transform -1 0 17584 0 1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1794_
timestamp 1698431365
transform -1 0 15568 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1795_
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1796_
timestamp 1698431365
transform 1 0 14336 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1797_
timestamp 1698431365
transform 1 0 49616 0 -1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1798_
timestamp 1698431365
transform -1 0 40992 0 1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1799_
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1800_
timestamp 1698431365
transform 1 0 37856 0 1 51744
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1801_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41664 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1802_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1803_
timestamp 1698431365
transform -1 0 13888 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1804_
timestamp 1698431365
transform -1 0 11760 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1805_
timestamp 1698431365
transform 1 0 12432 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1806_
timestamp 1698431365
transform -1 0 13216 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1807_
timestamp 1698431365
transform 1 0 12208 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1808_
timestamp 1698431365
transform 1 0 13552 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1809_
timestamp 1698431365
transform 1 0 11760 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1810_
timestamp 1698431365
transform 1 0 12096 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1811_
timestamp 1698431365
transform -1 0 13664 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1812_
timestamp 1698431365
transform 1 0 20272 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1813_
timestamp 1698431365
transform -1 0 22176 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1814_
timestamp 1698431365
transform -1 0 20944 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1815_
timestamp 1698431365
transform 1 0 12432 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1816_
timestamp 1698431365
transform -1 0 14000 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1817_
timestamp 1698431365
transform 1 0 20272 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1818_
timestamp 1698431365
transform -1 0 25984 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1819_
timestamp 1698431365
transform -1 0 21616 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1820_
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1821_
timestamp 1698431365
transform -1 0 25872 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1822_
timestamp 1698431365
transform -1 0 22736 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1823_
timestamp 1698431365
transform 1 0 22176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1824_
timestamp 1698431365
transform -1 0 23296 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1825_
timestamp 1698431365
transform 1 0 21728 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1826_
timestamp 1698431365
transform -1 0 23856 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1827_
timestamp 1698431365
transform 1 0 20944 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1828_
timestamp 1698431365
transform -1 0 22624 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1829_
timestamp 1698431365
transform -1 0 21840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1830_
timestamp 1698431365
transform 1 0 22512 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1831_
timestamp 1698431365
transform -1 0 27776 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1832_
timestamp 1698431365
transform -1 0 24304 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1833_
timestamp 1698431365
transform -1 0 23744 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1834_
timestamp 1698431365
transform -1 0 29680 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1835_
timestamp 1698431365
transform -1 0 27440 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1836_
timestamp 1698431365
transform -1 0 26432 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1837_
timestamp 1698431365
transform -1 0 36400 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1838_
timestamp 1698431365
transform -1 0 28448 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1839_
timestamp 1698431365
transform -1 0 28784 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1840_
timestamp 1698431365
transform 1 0 13664 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1841_
timestamp 1698431365
transform 1 0 42784 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1842_
timestamp 1698431365
transform -1 0 43792 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1843_
timestamp 1698431365
transform -1 0 39200 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1844_
timestamp 1698431365
transform -1 0 35728 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1845_
timestamp 1698431365
transform -1 0 34944 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1846_
timestamp 1698431365
transform 1 0 14448 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1847_
timestamp 1698431365
transform 1 0 46032 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1848_
timestamp 1698431365
transform 1 0 40992 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1849_
timestamp 1698431365
transform 1 0 39424 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1850_
timestamp 1698431365
transform -1 0 38528 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1851_
timestamp 1698431365
transform -1 0 45360 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1852_
timestamp 1698431365
transform -1 0 41888 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1853_
timestamp 1698431365
transform -1 0 43232 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1854_
timestamp 1698431365
transform 1 0 43120 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1855_
timestamp 1698431365
transform -1 0 43792 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1856_
timestamp 1698431365
transform -1 0 50624 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1857_
timestamp 1698431365
transform 1 0 49280 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1858_
timestamp 1698431365
transform -1 0 47712 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1859_
timestamp 1698431365
transform 1 0 46816 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1860_
timestamp 1698431365
transform 1 0 52976 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1861_
timestamp 1698431365
transform 1 0 49280 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1862_
timestamp 1698431365
transform 1 0 50624 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1863_
timestamp 1698431365
transform 1 0 50400 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1864_
timestamp 1698431365
transform 1 0 51408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1865_
timestamp 1698431365
transform 1 0 50512 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1866_
timestamp 1698431365
transform 1 0 51520 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1867_
timestamp 1698431365
transform 1 0 54096 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1868_
timestamp 1698431365
transform -1 0 54096 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1869_
timestamp 1698431365
transform 1 0 53312 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1870_
timestamp 1698431365
transform 1 0 53312 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1871_
timestamp 1698431365
transform 1 0 54544 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1872_
timestamp 1698431365
transform 1 0 55552 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1873_
timestamp 1698431365
transform 1 0 54992 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1874_
timestamp 1698431365
transform -1 0 56896 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1875_
timestamp 1698431365
transform 1 0 54768 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1876_
timestamp 1698431365
transform -1 0 56224 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1877_
timestamp 1698431365
transform 1 0 53872 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1878_
timestamp 1698431365
transform -1 0 55888 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1879_
timestamp 1698431365
transform 1 0 54880 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1880_
timestamp 1698431365
transform -1 0 56896 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1881_
timestamp 1698431365
transform 1 0 53984 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1882_
timestamp 1698431365
transform -1 0 54656 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1883_
timestamp 1698431365
transform 1 0 54544 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1884_
timestamp 1698431365
transform 1 0 55664 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1885_
timestamp 1698431365
transform -1 0 55328 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1886_
timestamp 1698431365
transform 1 0 54208 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1887_
timestamp 1698431365
transform 1 0 55440 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1888_
timestamp 1698431365
transform 1 0 53648 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1889_
timestamp 1698431365
transform 1 0 54320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1890_
timestamp 1698431365
transform 1 0 16912 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1891_
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1892_
timestamp 1698431365
transform 1 0 40880 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1893_
timestamp 1698431365
transform 1 0 41888 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1894_
timestamp 1698431365
transform 1 0 16352 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1895_
timestamp 1698431365
transform 1 0 18592 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1896_
timestamp 1698431365
transform -1 0 32256 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1897_
timestamp 1698431365
transform -1 0 32704 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1898_
timestamp 1698431365
transform 1 0 29344 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1899_
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1900_
timestamp 1698431365
transform -1 0 21392 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1901_
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1902_
timestamp 1698431365
transform 1 0 24304 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1903_
timestamp 1698431365
transform -1 0 17808 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1904_
timestamp 1698431365
transform 1 0 18032 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1905_
timestamp 1698431365
transform 1 0 17584 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1906_
timestamp 1698431365
transform -1 0 16912 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1907_
timestamp 1698431365
transform 1 0 15792 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1908_
timestamp 1698431365
transform -1 0 16352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1909_
timestamp 1698431365
transform -1 0 14000 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1910_
timestamp 1698431365
transform 1 0 14784 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1911_
timestamp 1698431365
transform -1 0 14448 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1912_
timestamp 1698431365
transform 1 0 13328 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1913_
timestamp 1698431365
transform 1 0 15120 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1914_
timestamp 1698431365
transform -1 0 16464 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1915_
timestamp 1698431365
transform 1 0 16128 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1916_
timestamp 1698431365
transform 1 0 14000 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1917_
timestamp 1698431365
transform 1 0 49392 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1918_
timestamp 1698431365
transform -1 0 53984 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1919_
timestamp 1698431365
transform -1 0 50848 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1920_
timestamp 1698431365
transform -1 0 53424 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1921_
timestamp 1698431365
transform 1 0 51520 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1922_
timestamp 1698431365
transform -1 0 52976 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1923_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 50848 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1924_
timestamp 1698431365
transform 1 0 51520 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1925_
timestamp 1698431365
transform -1 0 52304 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1926_
timestamp 1698431365
transform 1 0 51520 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1927_
timestamp 1698431365
transform -1 0 53648 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1928_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 51856 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1929_
timestamp 1698431365
transform 1 0 50960 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1930_
timestamp 1698431365
transform -1 0 55216 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1931_
timestamp 1698431365
transform 1 0 53648 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1932_
timestamp 1698431365
transform 1 0 52640 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1933_
timestamp 1698431365
transform -1 0 54320 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1934_
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1935_
timestamp 1698431365
transform -1 0 56112 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1936_
timestamp 1698431365
transform -1 0 54432 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1937_
timestamp 1698431365
transform 1 0 54992 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1938_
timestamp 1698431365
transform 1 0 51856 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1939_
timestamp 1698431365
transform -1 0 52304 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1940_
timestamp 1698431365
transform -1 0 53424 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1941_
timestamp 1698431365
transform 1 0 53088 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1942_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 54208 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1943_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27664 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1944_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27776 0 -1 20384
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1945_
timestamp 1698431365
transform 1 0 27440 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1946_
timestamp 1698431365
transform 1 0 27888 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1947_
timestamp 1698431365
transform 1 0 22624 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1948_
timestamp 1698431365
transform 1 0 26320 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1949_
timestamp 1698431365
transform 1 0 27776 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1950_
timestamp 1698431365
transform 1 0 25648 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1951_
timestamp 1698431365
transform 1 0 25424 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1952_
timestamp 1698431365
transform 1 0 28224 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1953_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1954_
timestamp 1698431365
transform 1 0 29680 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1955_
timestamp 1698431365
transform 1 0 26656 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1956_
timestamp 1698431365
transform 1 0 29344 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1957_
timestamp 1698431365
transform 1 0 26320 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1958_
timestamp 1698431365
transform 1 0 23296 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1959_
timestamp 1698431365
transform 1 0 27552 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1960_
timestamp 1698431365
transform 1 0 28672 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1961_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30352 0 -1 18816
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1962_
timestamp 1698431365
transform -1 0 30240 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1963_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29344 0 -1 12544
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1964_
timestamp 1698431365
transform 1 0 25760 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1965_
timestamp 1698431365
transform -1 0 28000 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1966_
timestamp 1698431365
transform 1 0 25536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1967_
timestamp 1698431365
transform 1 0 26208 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1968_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27440 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1969_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1970_
timestamp 1698431365
transform -1 0 49952 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1971_
timestamp 1698431365
transform -1 0 48272 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1972_
timestamp 1698431365
transform -1 0 46928 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1973_
timestamp 1698431365
transform 1 0 42672 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1974_
timestamp 1698431365
transform 1 0 42224 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1975_
timestamp 1698431365
transform 1 0 43456 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1976_
timestamp 1698431365
transform -1 0 44464 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1977_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45920 0 -1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1978_
timestamp 1698431365
transform -1 0 42112 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1979_
timestamp 1698431365
transform 1 0 37408 0 -1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1980_
timestamp 1698431365
transform -1 0 36624 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1981_
timestamp 1698431365
transform 1 0 38976 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1982_
timestamp 1698431365
transform 1 0 40880 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1983_
timestamp 1698431365
transform -1 0 42672 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1984_
timestamp 1698431365
transform 1 0 39312 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1985_
timestamp 1698431365
transform 1 0 36848 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1986_
timestamp 1698431365
transform 1 0 35392 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1987_
timestamp 1698431365
transform 1 0 38080 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1988_
timestamp 1698431365
transform 1 0 42448 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1989_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42560 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1990_
timestamp 1698431365
transform 1 0 42560 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1991_
timestamp 1698431365
transform 1 0 43904 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1992_
timestamp 1698431365
transform -1 0 49840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1993_
timestamp 1698431365
transform -1 0 48944 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1994_
timestamp 1698431365
transform -1 0 49392 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1995_
timestamp 1698431365
transform 1 0 47488 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1996_
timestamp 1698431365
transform 1 0 45136 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1997_
timestamp 1698431365
transform 1 0 43120 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1998_
timestamp 1698431365
transform 1 0 45248 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1999_
timestamp 1698431365
transform 1 0 45248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2000_
timestamp 1698431365
transform -1 0 48272 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2001_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46368 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2002_
timestamp 1698431365
transform 1 0 46480 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2003_
timestamp 1698431365
transform -1 0 53424 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2004_
timestamp 1698431365
transform -1 0 52752 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2005_
timestamp 1698431365
transform -1 0 51408 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2006_
timestamp 1698431365
transform 1 0 50848 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2007_
timestamp 1698431365
transform 1 0 50848 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2008_
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2009_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 52192 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2010_
timestamp 1698431365
transform 1 0 49392 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2011_
timestamp 1698431365
transform 1 0 49728 0 -1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2012_
timestamp 1698431365
transform -1 0 48832 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2013_
timestamp 1698431365
transform 1 0 29568 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2014_
timestamp 1698431365
transform 1 0 29904 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2015_
timestamp 1698431365
transform 1 0 32256 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2016_
timestamp 1698431365
transform 1 0 30016 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2017_
timestamp 1698431365
transform -1 0 34048 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2018_
timestamp 1698431365
transform -1 0 38864 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2019_
timestamp 1698431365
transform -1 0 39312 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2020_
timestamp 1698431365
transform 1 0 36960 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2021_
timestamp 1698431365
transform -1 0 35392 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2022_
timestamp 1698431365
transform 1 0 34608 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2023_
timestamp 1698431365
transform -1 0 33376 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2024_
timestamp 1698431365
transform 1 0 29904 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2025_
timestamp 1698431365
transform -1 0 40320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2026_
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2027_
timestamp 1698431365
transform -1 0 39648 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2028_
timestamp 1698431365
transform 1 0 38640 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2029_
timestamp 1698431365
transform -1 0 39872 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2030_
timestamp 1698431365
transform 1 0 38304 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2031_
timestamp 1698431365
transform -1 0 32368 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2032_
timestamp 1698431365
transform -1 0 30016 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2033_
timestamp 1698431365
transform 1 0 19376 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2034_
timestamp 1698431365
transform 1 0 21392 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2035_
timestamp 1698431365
transform 1 0 22736 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2036_
timestamp 1698431365
transform -1 0 24640 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2037_
timestamp 1698431365
transform -1 0 19712 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2038_
timestamp 1698431365
transform 1 0 19712 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2039_
timestamp 1698431365
transform -1 0 20272 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2040_
timestamp 1698431365
transform 1 0 18480 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2041_
timestamp 1698431365
transform 1 0 13552 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2042_
timestamp 1698431365
transform 1 0 15792 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2043_
timestamp 1698431365
transform 1 0 15344 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2044_
timestamp 1698431365
transform 1 0 16128 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2045_
timestamp 1698431365
transform -1 0 17584 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2046_
timestamp 1698431365
transform 1 0 15568 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2047_
timestamp 1698431365
transform 1 0 14672 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2048_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2049_
timestamp 1698431365
transform 1 0 13664 0 -1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2050_
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2051_
timestamp 1698431365
transform 1 0 16800 0 1 10976
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2052_
timestamp 1698431365
transform -1 0 16128 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2053_
timestamp 1698431365
transform -1 0 6048 0 -1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2054_
timestamp 1698431365
transform 1 0 3920 0 -1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _2055_
timestamp 1698431365
transform 1 0 4816 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2056_
timestamp 1698431365
transform -1 0 7168 0 -1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2057_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6496 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2058_
timestamp 1698431365
transform 1 0 13776 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2059_
timestamp 1698431365
transform 1 0 14896 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2060_
timestamp 1698431365
transform 1 0 13216 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2061_
timestamp 1698431365
transform -1 0 14560 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2062_
timestamp 1698431365
transform 1 0 20944 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2063_
timestamp 1698431365
transform 1 0 22064 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2064_
timestamp 1698431365
transform -1 0 23408 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2065_
timestamp 1698431365
transform 1 0 18256 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2066_
timestamp 1698431365
transform -1 0 18480 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2067_
timestamp 1698431365
transform -1 0 21840 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2068_
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2069_
timestamp 1698431365
transform 1 0 17472 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2070_
timestamp 1698431365
transform -1 0 17584 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2071_
timestamp 1698431365
transform -1 0 16912 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2072_
timestamp 1698431365
transform 1 0 15456 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2073_
timestamp 1698431365
transform 1 0 19264 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2074_
timestamp 1698431365
transform 1 0 18368 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2075_
timestamp 1698431365
transform 1 0 18704 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2076_
timestamp 1698431365
transform 1 0 19376 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2077_
timestamp 1698431365
transform 1 0 20272 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2078_
timestamp 1698431365
transform 1 0 30464 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2079_
timestamp 1698431365
transform -1 0 30688 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2080_
timestamp 1698431365
transform 1 0 21840 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2081_
timestamp 1698431365
transform -1 0 22176 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2082_
timestamp 1698431365
transform 1 0 21728 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2083_
timestamp 1698431365
transform -1 0 20944 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2084_
timestamp 1698431365
transform 1 0 23072 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2085_
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2086_
timestamp 1698431365
transform 1 0 30352 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2087_
timestamp 1698431365
transform 1 0 23184 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2088_
timestamp 1698431365
transform 1 0 28784 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2089_
timestamp 1698431365
transform -1 0 28784 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2090_
timestamp 1698431365
transform 1 0 29344 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2091_
timestamp 1698431365
transform 1 0 30352 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2092_
timestamp 1698431365
transform -1 0 34944 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2093_
timestamp 1698431365
transform 1 0 31360 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2094_
timestamp 1698431365
transform -1 0 31808 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2095_
timestamp 1698431365
transform -1 0 33824 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2096_
timestamp 1698431365
transform 1 0 33824 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2097_
timestamp 1698431365
transform 1 0 16240 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2098_
timestamp 1698431365
transform -1 0 41664 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2099_
timestamp 1698431365
transform 1 0 39088 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2100_
timestamp 1698431365
transform -1 0 39312 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2101_
timestamp 1698431365
transform 1 0 39312 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2102_
timestamp 1698431365
transform 1 0 40992 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2103_
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2104_
timestamp 1698431365
transform -1 0 43232 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2105_
timestamp 1698431365
transform -1 0 42336 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2106_
timestamp 1698431365
transform 1 0 42896 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2107_
timestamp 1698431365
transform -1 0 42896 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2108_
timestamp 1698431365
transform 1 0 47264 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2109_
timestamp 1698431365
transform 1 0 45360 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2110_
timestamp 1698431365
transform 1 0 45696 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2111_
timestamp 1698431365
transform 1 0 46368 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2112_
timestamp 1698431365
transform 1 0 49280 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2113_
timestamp 1698431365
transform 1 0 44912 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2114_
timestamp 1698431365
transform 1 0 46480 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2115_
timestamp 1698431365
transform -1 0 46480 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2116_
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2117_
timestamp 1698431365
transform -1 0 48272 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2118_
timestamp 1698431365
transform 1 0 50400 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2119_
timestamp 1698431365
transform -1 0 53200 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2120_
timestamp 1698431365
transform 1 0 53760 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2121_
timestamp 1698431365
transform -1 0 54096 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2122_
timestamp 1698431365
transform 1 0 54432 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2123_
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2124_
timestamp 1698431365
transform 1 0 35056 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2125_
timestamp 1698431365
transform 1 0 51408 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2126_
timestamp 1698431365
transform 1 0 52192 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2127_
timestamp 1698431365
transform -1 0 51408 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2128_
timestamp 1698431365
transform 1 0 51520 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2129_
timestamp 1698431365
transform -1 0 35504 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2130_
timestamp 1698431365
transform 1 0 37632 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2131_
timestamp 1698431365
transform -1 0 36960 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2132_
timestamp 1698431365
transform 1 0 36736 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2133_
timestamp 1698431365
transform -1 0 36624 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2134_
timestamp 1698431365
transform 1 0 21280 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2135_
timestamp 1698431365
transform 1 0 26432 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2136_
timestamp 1698431365
transform -1 0 26880 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2137_
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2138_
timestamp 1698431365
transform 1 0 26656 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2139_
timestamp 1698431365
transform -1 0 15680 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2140_
timestamp 1698431365
transform 1 0 13776 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2141_
timestamp 1698431365
transform 1 0 14224 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2142_
timestamp 1698431365
transform -1 0 13104 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2143_
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2144_
timestamp 1698431365
transform 1 0 21728 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2145_
timestamp 1698431365
transform 1 0 13888 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2146_
timestamp 1698431365
transform -1 0 13776 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2147_
timestamp 1698431365
transform 1 0 14784 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2148_
timestamp 1698431365
transform 1 0 15680 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2149_
timestamp 1698431365
transform -1 0 15904 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2150_
timestamp 1698431365
transform -1 0 14896 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2151_
timestamp 1698431365
transform -1 0 17920 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2152_
timestamp 1698431365
transform -1 0 16464 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2153_
timestamp 1698431365
transform -1 0 13888 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2154_
timestamp 1698431365
transform -1 0 16688 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2155_
timestamp 1698431365
transform -1 0 14784 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2156_
timestamp 1698431365
transform 1 0 17920 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2157_
timestamp 1698431365
transform 1 0 16912 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2158_
timestamp 1698431365
transform -1 0 15792 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2159_
timestamp 1698431365
transform -1 0 18256 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2160_
timestamp 1698431365
transform -1 0 17024 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2161_
timestamp 1698431365
transform -1 0 23520 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2162_
timestamp 1698431365
transform -1 0 19600 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2163_
timestamp 1698431365
transform -1 0 19936 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2164_
timestamp 1698431365
transform -1 0 20608 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2165_
timestamp 1698431365
transform 1 0 18256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2166_
timestamp 1698431365
transform 1 0 22176 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2167_
timestamp 1698431365
transform -1 0 24864 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2168_
timestamp 1698431365
transform -1 0 24864 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2169_
timestamp 1698431365
transform -1 0 26096 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2170_
timestamp 1698431365
transform -1 0 24864 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2171_
timestamp 1698431365
transform 1 0 42112 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2172_
timestamp 1698431365
transform -1 0 42784 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2173_
timestamp 1698431365
transform -1 0 28560 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2174_
timestamp 1698431365
transform 1 0 27104 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2175_
timestamp 1698431365
transform -1 0 30016 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2176_
timestamp 1698431365
transform -1 0 28672 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2177_
timestamp 1698431365
transform 1 0 17584 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2178_
timestamp 1698431365
transform 1 0 37184 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2179_
timestamp 1698431365
transform -1 0 38864 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2180_
timestamp 1698431365
transform 1 0 35504 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2181_
timestamp 1698431365
transform -1 0 38416 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2182_
timestamp 1698431365
transform -1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2183_
timestamp 1698431365
transform -1 0 43456 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2184_
timestamp 1698431365
transform -1 0 40320 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2185_
timestamp 1698431365
transform -1 0 39312 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2186_
timestamp 1698431365
transform -1 0 41776 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2187_
timestamp 1698431365
transform 1 0 41776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2188_
timestamp 1698431365
transform -1 0 47488 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2189_
timestamp 1698431365
transform 1 0 43456 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2190_
timestamp 1698431365
transform -1 0 45136 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2191_
timestamp 1698431365
transform -1 0 46928 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2192_
timestamp 1698431365
transform -1 0 44128 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2193_
timestamp 1698431365
transform 1 0 45136 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2194_
timestamp 1698431365
transform 1 0 45808 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2195_
timestamp 1698431365
transform -1 0 48384 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2196_
timestamp 1698431365
transform -1 0 47936 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2197_
timestamp 1698431365
transform 1 0 47488 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2198_
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2199_
timestamp 1698431365
transform -1 0 50288 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2200_
timestamp 1698431365
transform 1 0 49168 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2201_
timestamp 1698431365
transform -1 0 51296 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2202_
timestamp 1698431365
transform 1 0 51296 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2203_
timestamp 1698431365
transform 1 0 43680 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2204_
timestamp 1698431365
transform 1 0 50624 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2205_
timestamp 1698431365
transform 1 0 51072 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2206_
timestamp 1698431365
transform 1 0 49616 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2207_
timestamp 1698431365
transform -1 0 52192 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2208_
timestamp 1698431365
transform 1 0 24976 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2209_
timestamp 1698431365
transform -1 0 36736 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2210_
timestamp 1698431365
transform -1 0 37184 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2211_
timestamp 1698431365
transform -1 0 35168 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2212_
timestamp 1698431365
transform 1 0 33712 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2213_
timestamp 1698431365
transform 1 0 15232 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2214_
timestamp 1698431365
transform -1 0 26992 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2215_
timestamp 1698431365
transform 1 0 25536 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2216_
timestamp 1698431365
transform -1 0 28000 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2217_
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2218_
timestamp 1698431365
transform -1 0 11760 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2219_
timestamp 1698431365
transform 1 0 9744 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2220_
timestamp 1698431365
transform -1 0 12656 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2221_
timestamp 1698431365
transform -1 0 11760 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2222_
timestamp 1698431365
transform -1 0 12320 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2223_
timestamp 1698431365
transform -1 0 11200 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2224_
timestamp 1698431365
transform -1 0 12432 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2225_
timestamp 1698431365
transform -1 0 10080 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2226_
timestamp 1698431365
transform -1 0 11424 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2227_
timestamp 1698431365
transform -1 0 9968 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2228_
timestamp 1698431365
transform 1 0 14000 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2229_
timestamp 1698431365
transform -1 0 11200 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2230_
timestamp 1698431365
transform -1 0 13104 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2231_
timestamp 1698431365
transform 1 0 16128 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2232_
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2233_
timestamp 1698431365
transform 1 0 14112 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2234_
timestamp 1698431365
transform -1 0 16128 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2235_
timestamp 1698431365
transform -1 0 15232 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2236_
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2237_
timestamp 1698431365
transform 1 0 14560 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2238_
timestamp 1698431365
transform 1 0 21840 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2239_
timestamp 1698431365
transform 1 0 24528 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2240_
timestamp 1698431365
transform 1 0 32032 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2241_
timestamp 1698431365
transform 1 0 22512 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2242_
timestamp 1698431365
transform 1 0 23184 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2243_
timestamp 1698431365
transform 1 0 30464 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2244_
timestamp 1698431365
transform -1 0 31920 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2245_
timestamp 1698431365
transform 1 0 25760 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2246_
timestamp 1698431365
transform 1 0 27104 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2247_
timestamp 1698431365
transform 1 0 25424 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2248_
timestamp 1698431365
transform 1 0 25536 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2249_
timestamp 1698431365
transform 1 0 25424 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2250_
timestamp 1698431365
transform 1 0 18368 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2251_
timestamp 1698431365
transform 1 0 19152 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2252_
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2253_
timestamp 1698431365
transform 1 0 11424 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2254_
timestamp 1698431365
transform 1 0 12432 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2255_
timestamp 1698431365
transform 1 0 19152 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2256_
timestamp 1698431365
transform 1 0 34608 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2257_
timestamp 1698431365
transform -1 0 35280 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2258_
timestamp 1698431365
transform -1 0 33040 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2259_
timestamp 1698431365
transform -1 0 34272 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2260_
timestamp 1698431365
transform 1 0 27888 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2261_
timestamp 1698431365
transform -1 0 17920 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2262_
timestamp 1698431365
transform 1 0 17920 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2263_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2264_
timestamp 1698431365
transform 1 0 29456 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2265_
timestamp 1698431365
transform -1 0 34720 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2266_
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2267_
timestamp 1698431365
transform -1 0 24192 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2268_
timestamp 1698431365
transform 1 0 30800 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2269_
timestamp 1698431365
transform 1 0 31248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2270_
timestamp 1698431365
transform 1 0 31360 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2271_
timestamp 1698431365
transform 1 0 19824 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2272_
timestamp 1698431365
transform 1 0 31360 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2273_
timestamp 1698431365
transform 1 0 35280 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2274_
timestamp 1698431365
transform 1 0 34160 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2275_
timestamp 1698431365
transform -1 0 34384 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2276_
timestamp 1698431365
transform 1 0 28560 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2277_
timestamp 1698431365
transform 1 0 30464 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2278_
timestamp 1698431365
transform 1 0 18032 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2279_
timestamp 1698431365
transform -1 0 30800 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2280_
timestamp 1698431365
transform 1 0 30464 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2281_
timestamp 1698431365
transform 1 0 31248 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2282_
timestamp 1698431365
transform 1 0 31808 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2283_
timestamp 1698431365
transform 1 0 31136 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2284_
timestamp 1698431365
transform 1 0 19264 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2285_
timestamp 1698431365
transform 1 0 35280 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2286_
timestamp 1698431365
transform 1 0 34272 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2287_
timestamp 1698431365
transform -1 0 34272 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2288_
timestamp 1698431365
transform 1 0 27888 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2289_
timestamp 1698431365
transform -1 0 30688 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2290_
timestamp 1698431365
transform 1 0 29344 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2291_
timestamp 1698431365
transform 1 0 29344 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2292_
timestamp 1698431365
transform -1 0 31696 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2293_
timestamp 1698431365
transform 1 0 32032 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2294_
timestamp 1698431365
transform 1 0 29680 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2295_
timestamp 1698431365
transform -1 0 24752 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2296_
timestamp 1698431365
transform -1 0 35728 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2297_
timestamp 1698431365
transform 1 0 35280 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2298_
timestamp 1698431365
transform 1 0 32816 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2299_
timestamp 1698431365
transform -1 0 33712 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2300_
timestamp 1698431365
transform 1 0 19600 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2301_
timestamp 1698431365
transform 1 0 35392 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2302_
timestamp 1698431365
transform -1 0 32928 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2303_
timestamp 1698431365
transform -1 0 32480 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2304_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2305_
timestamp 1698431365
transform 1 0 24528 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2306_
timestamp 1698431365
transform 1 0 25872 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2307_
timestamp 1698431365
transform -1 0 20272 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2308_
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2309_
timestamp 1698431365
transform -1 0 26544 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2310_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2311_
timestamp 1698431365
transform -1 0 19600 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2312_
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2313_
timestamp 1698431365
transform -1 0 32928 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2314_
timestamp 1698431365
transform -1 0 27776 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2315_
timestamp 1698431365
transform 1 0 26544 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2316_
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2317_
timestamp 1698431365
transform 1 0 29904 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2318_
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2319_
timestamp 1698431365
transform 1 0 28336 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2320_
timestamp 1698431365
transform -1 0 24192 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2321_
timestamp 1698431365
transform 1 0 32928 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2322_
timestamp 1698431365
transform -1 0 33376 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2323_
timestamp 1698431365
transform -1 0 31808 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2324_
timestamp 1698431365
transform -1 0 28224 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2325_
timestamp 1698431365
transform 1 0 28000 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2326_
timestamp 1698431365
transform 1 0 26544 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2327_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2328_
timestamp 1698431365
transform -1 0 26432 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2329_
timestamp 1698431365
transform 1 0 26432 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2330_
timestamp 1698431365
transform 1 0 26432 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2331_
timestamp 1698431365
transform 1 0 24864 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2332_
timestamp 1698431365
transform 1 0 23968 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2333_
timestamp 1698431365
transform 1 0 31136 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2334_
timestamp 1698431365
transform -1 0 34944 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2335_
timestamp 1698431365
transform -1 0 32704 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2336_
timestamp 1698431365
transform -1 0 31920 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2337_
timestamp 1698431365
transform 1 0 25760 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2338_
timestamp 1698431365
transform 1 0 30240 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2339_
timestamp 1698431365
transform 1 0 30128 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2340_
timestamp 1698431365
transform -1 0 31808 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2341_
timestamp 1698431365
transform 1 0 31808 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2342_
timestamp 1698431365
transform 1 0 31136 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2343_
timestamp 1698431365
transform 1 0 31696 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2344_
timestamp 1698431365
transform 1 0 33152 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2345_
timestamp 1698431365
transform -1 0 34048 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2346_
timestamp 1698431365
transform -1 0 39760 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2347_
timestamp 1698431365
transform -1 0 39088 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2348_
timestamp 1698431365
transform -1 0 34048 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2349_
timestamp 1698431365
transform 1 0 34496 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2350_
timestamp 1698431365
transform 1 0 33600 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2351_
timestamp 1698431365
transform 1 0 33040 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2352_
timestamp 1698431365
transform -1 0 33488 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2353_
timestamp 1698431365
transform 1 0 32032 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2354_
timestamp 1698431365
transform 1 0 34608 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2355_
timestamp 1698431365
transform 1 0 37408 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2356_
timestamp 1698431365
transform -1 0 34496 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2357_
timestamp 1698431365
transform 1 0 34272 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2358_
timestamp 1698431365
transform 1 0 34384 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2359_
timestamp 1698431365
transform 1 0 34048 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2360_
timestamp 1698431365
transform 1 0 34944 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2361_
timestamp 1698431365
transform 1 0 35728 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2362_
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2363_
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2364_
timestamp 1698431365
transform 1 0 35392 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2365_
timestamp 1698431365
transform -1 0 16128 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2366_
timestamp 1698431365
transform 1 0 10640 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2367_
timestamp 1698431365
transform 1 0 35952 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2368_
timestamp 1698431365
transform 1 0 33936 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2369_
timestamp 1698431365
transform 1 0 37408 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2370_
timestamp 1698431365
transform 1 0 36288 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2371_
timestamp 1698431365
transform -1 0 39312 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2372_
timestamp 1698431365
transform 1 0 37632 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2373_
timestamp 1698431365
transform 1 0 37296 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2374_
timestamp 1698431365
transform 1 0 37520 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2375_
timestamp 1698431365
transform 1 0 38864 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2376_
timestamp 1698431365
transform 1 0 38640 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2377_
timestamp 1698431365
transform -1 0 39088 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2378_
timestamp 1698431365
transform -1 0 38528 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2379_
timestamp 1698431365
transform -1 0 39536 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2380_
timestamp 1698431365
transform 1 0 38080 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2381_
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2382_
timestamp 1698431365
transform 1 0 35616 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2383_
timestamp 1698431365
transform -1 0 40096 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2384_
timestamp 1698431365
transform 1 0 40096 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2385_
timestamp 1698431365
transform -1 0 42448 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2386_
timestamp 1698431365
transform 1 0 42000 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2387_
timestamp 1698431365
transform 1 0 42000 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2388_
timestamp 1698431365
transform -1 0 35616 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2389_
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2390_
timestamp 1698431365
transform 1 0 34720 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2391_
timestamp 1698431365
transform 1 0 35056 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2392_
timestamp 1698431365
transform 1 0 42896 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2393_
timestamp 1698431365
transform -1 0 43904 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2394_
timestamp 1698431365
transform 1 0 41888 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2395_
timestamp 1698431365
transform 1 0 42448 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2396_
timestamp 1698431365
transform -1 0 43344 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2397_
timestamp 1698431365
transform -1 0 42672 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2398_
timestamp 1698431365
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2399_
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2400_
timestamp 1698431365
transform -1 0 39424 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2401_
timestamp 1698431365
transform -1 0 35504 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2402_
timestamp 1698431365
transform 1 0 35616 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2403_
timestamp 1698431365
transform 1 0 43568 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2404_
timestamp 1698431365
transform -1 0 43456 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2405_
timestamp 1698431365
transform -1 0 37744 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2406_
timestamp 1698431365
transform -1 0 38304 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2407_
timestamp 1698431365
transform 1 0 38080 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2408_
timestamp 1698431365
transform -1 0 40096 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2409_
timestamp 1698431365
transform 1 0 35504 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2410_
timestamp 1698431365
transform 1 0 39200 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2411_
timestamp 1698431365
transform 1 0 39088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2412_
timestamp 1698431365
transform 1 0 40768 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2413_
timestamp 1698431365
transform -1 0 45472 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2414_
timestamp 1698431365
transform 1 0 44352 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2415_
timestamp 1698431365
transform -1 0 45808 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2416_
timestamp 1698431365
transform 1 0 39760 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2417_
timestamp 1698431365
transform 1 0 42224 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2418_
timestamp 1698431365
transform 1 0 41664 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2419_
timestamp 1698431365
transform 1 0 45808 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2420_
timestamp 1698431365
transform 1 0 45472 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2421_
timestamp 1698431365
transform 1 0 46704 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2422_
timestamp 1698431365
transform -1 0 44464 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2423_
timestamp 1698431365
transform -1 0 39200 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2424_
timestamp 1698431365
transform 1 0 38416 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2425_
timestamp 1698431365
transform 1 0 43344 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2426_
timestamp 1698431365
transform 1 0 43568 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2427_
timestamp 1698431365
transform 1 0 45360 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2428_
timestamp 1698431365
transform 1 0 44912 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2429_
timestamp 1698431365
transform -1 0 39088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2430_
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2431_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2432_
timestamp 1698431365
transform -1 0 39984 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2433_
timestamp 1698431365
transform 1 0 38416 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2434_
timestamp 1698431365
transform 1 0 31360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2435_
timestamp 1698431365
transform 1 0 38528 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2436_
timestamp 1698431365
transform 1 0 42336 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2437_
timestamp 1698431365
transform 1 0 47376 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2438_
timestamp 1698431365
transform -1 0 49952 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2439_
timestamp 1698431365
transform 1 0 42448 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2440_
timestamp 1698431365
transform -1 0 44128 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2441_
timestamp 1698431365
transform 1 0 44688 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2442_
timestamp 1698431365
transform 1 0 45360 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2443_
timestamp 1698431365
transform -1 0 38416 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2444_
timestamp 1698431365
transform 1 0 38640 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2445_
timestamp 1698431365
transform 1 0 47488 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2446_
timestamp 1698431365
transform 1 0 49952 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2447_
timestamp 1698431365
transform 1 0 49952 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2448_
timestamp 1698431365
transform -1 0 51408 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2449_
timestamp 1698431365
transform -1 0 40544 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2450_
timestamp 1698431365
transform -1 0 41664 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2451_
timestamp 1698431365
transform 1 0 45248 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2452_
timestamp 1698431365
transform 1 0 46928 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2453_
timestamp 1698431365
transform 1 0 42000 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2454_
timestamp 1698431365
transform -1 0 53984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2455_
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2456_
timestamp 1698431365
transform -1 0 51520 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2457_
timestamp 1698431365
transform -1 0 53536 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2458_
timestamp 1698431365
transform -1 0 42112 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2459_
timestamp 1698431365
transform 1 0 40656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2460_
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2461_
timestamp 1698431365
transform 1 0 41216 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2462_
timestamp 1698431365
transform 1 0 42896 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2463_
timestamp 1698431365
transform -1 0 44464 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2464_
timestamp 1698431365
transform -1 0 47040 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2465_
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2466_
timestamp 1698431365
transform 1 0 49840 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2467_
timestamp 1698431365
transform -1 0 52192 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2468_
timestamp 1698431365
transform 1 0 22176 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2469_
timestamp 1698431365
transform 1 0 42784 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2470_
timestamp 1698431365
transform 1 0 41328 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2471_
timestamp 1698431365
transform 1 0 42672 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2472_
timestamp 1698431365
transform -1 0 44688 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2473_
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2474_
timestamp 1698431365
transform 1 0 45024 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2475_
timestamp 1698431365
transform -1 0 54992 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2476_
timestamp 1698431365
transform -1 0 50848 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2477_
timestamp 1698431365
transform 1 0 50736 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2478_
timestamp 1698431365
transform -1 0 51072 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2479_
timestamp 1698431365
transform -1 0 41216 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2480_
timestamp 1698431365
transform 1 0 38080 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2481_
timestamp 1698431365
transform 1 0 40096 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2482_
timestamp 1698431365
transform 1 0 38752 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2483_
timestamp 1698431365
transform 1 0 42336 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2484_
timestamp 1698431365
transform -1 0 44464 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2485_
timestamp 1698431365
transform -1 0 48272 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2486_
timestamp 1698431365
transform -1 0 38752 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2487_
timestamp 1698431365
transform 1 0 38752 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2488_
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2489_
timestamp 1698431365
transform -1 0 46480 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2490_
timestamp 1698431365
transform 1 0 45136 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2491_
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2492_
timestamp 1698431365
transform 1 0 43008 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2493_
timestamp 1698431365
transform 1 0 44576 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2494_
timestamp 1698431365
transform 1 0 43792 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2495_
timestamp 1698431365
transform 1 0 51072 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2496_
timestamp 1698431365
transform -1 0 50288 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2497_
timestamp 1698431365
transform -1 0 44016 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2498_
timestamp 1698431365
transform 1 0 38976 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2499_
timestamp 1698431365
transform 1 0 39984 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2500_
timestamp 1698431365
transform -1 0 19712 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2501_
timestamp 1698431365
transform 1 0 40880 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2502_
timestamp 1698431365
transform 1 0 40432 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2503_
timestamp 1698431365
transform 1 0 42672 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2504_
timestamp 1698431365
transform -1 0 48272 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2505_
timestamp 1698431365
transform 1 0 50736 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2506_
timestamp 1698431365
transform 1 0 50736 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2507_
timestamp 1698431365
transform -1 0 49392 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2508_
timestamp 1698431365
transform 1 0 42000 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2509_
timestamp 1698431365
transform 1 0 41328 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2510_
timestamp 1698431365
transform -1 0 45584 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2511_
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2512_
timestamp 1698431365
transform 1 0 44128 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2513_
timestamp 1698431365
transform -1 0 42000 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2514_
timestamp 1698431365
transform -1 0 36736 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2515_
timestamp 1698431365
transform -1 0 37072 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2516_
timestamp 1698431365
transform -1 0 36624 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2517_
timestamp 1698431365
transform -1 0 36848 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2518_
timestamp 1698431365
transform -1 0 36064 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2519_
timestamp 1698431365
transform -1 0 18256 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2520_
timestamp 1698431365
transform 1 0 36064 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2521_
timestamp 1698431365
transform -1 0 37744 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2522_
timestamp 1698431365
transform -1 0 37184 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2523_
timestamp 1698431365
transform 1 0 38304 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2524_
timestamp 1698431365
transform -1 0 38752 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2525_
timestamp 1698431365
transform -1 0 38864 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2526_
timestamp 1698431365
transform -1 0 39648 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2527_
timestamp 1698431365
transform -1 0 38976 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2528_
timestamp 1698431365
transform -1 0 36624 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2529_
timestamp 1698431365
transform 1 0 37072 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2530_
timestamp 1698431365
transform 1 0 38416 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2531_
timestamp 1698431365
transform -1 0 40544 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2532_
timestamp 1698431365
transform 1 0 40544 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2533_
timestamp 1698431365
transform -1 0 37968 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2534_
timestamp 1698431365
transform -1 0 34944 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2535_
timestamp 1698431365
transform -1 0 34496 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2536_
timestamp 1698431365
transform 1 0 34944 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2537_
timestamp 1698431365
transform -1 0 33600 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2538_
timestamp 1698431365
transform -1 0 34608 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2539_
timestamp 1698431365
transform 1 0 34048 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2540_
timestamp 1698431365
transform -1 0 34048 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2541_
timestamp 1698431365
transform 1 0 21952 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2542_
timestamp 1698431365
transform 1 0 26544 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2543_
timestamp 1698431365
transform -1 0 26992 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2544_
timestamp 1698431365
transform 1 0 31360 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2545_
timestamp 1698431365
transform 1 0 31248 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2546_
timestamp 1698431365
transform -1 0 34384 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2547_
timestamp 1698431365
transform -1 0 32816 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2548_
timestamp 1698431365
transform 1 0 31136 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2549_
timestamp 1698431365
transform 1 0 32816 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2550_
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2551_
timestamp 1698431365
transform 1 0 26992 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2552_
timestamp 1698431365
transform 1 0 26880 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2553_
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2554_
timestamp 1698431365
transform -1 0 24864 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2555_
timestamp 1698431365
transform 1 0 23744 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2556_
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2557_
timestamp 1698431365
transform -1 0 24976 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2558_
timestamp 1698431365
transform -1 0 22736 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2559_
timestamp 1698431365
transform 1 0 23408 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2560_
timestamp 1698431365
transform 1 0 22624 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2561_
timestamp 1698431365
transform -1 0 21840 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2562_
timestamp 1698431365
transform 1 0 22400 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2563_
timestamp 1698431365
transform 1 0 22848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2564_
timestamp 1698431365
transform -1 0 23744 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2565_
timestamp 1698431365
transform -1 0 24528 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2566_
timestamp 1698431365
transform -1 0 23296 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2567_
timestamp 1698431365
transform 1 0 20384 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2568_
timestamp 1698431365
transform 1 0 21840 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2569_
timestamp 1698431365
transform 1 0 22176 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2570_
timestamp 1698431365
transform -1 0 21840 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2571_
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2572_
timestamp 1698431365
transform -1 0 20384 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2573_
timestamp 1698431365
transform 1 0 18592 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2574_
timestamp 1698431365
transform -1 0 19152 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2575_
timestamp 1698431365
transform -1 0 18256 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2576_
timestamp 1698431365
transform 1 0 17920 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2577_
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2578_
timestamp 1698431365
transform -1 0 14000 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2579_
timestamp 1698431365
transform 1 0 16016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2580_
timestamp 1698431365
transform -1 0 17360 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2581_
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2582_
timestamp 1698431365
transform -1 0 19600 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2583_
timestamp 1698431365
transform 1 0 19488 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2584_
timestamp 1698431365
transform -1 0 19376 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2585_
timestamp 1698431365
transform 1 0 17920 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2586_
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2587_
timestamp 1698431365
transform -1 0 16912 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2588_
timestamp 1698431365
transform -1 0 15456 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _2589_
timestamp 1698431365
transform 1 0 8512 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2590_
timestamp 1698431365
transform 1 0 7280 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2591_
timestamp 1698431365
transform 1 0 8288 0 1 26656
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2592_
timestamp 1698431365
transform 1 0 8736 0 1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2593_
timestamp 1698431365
transform -1 0 8288 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2594_
timestamp 1698431365
transform 1 0 8624 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2595_
timestamp 1698431365
transform 1 0 7952 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2596_
timestamp 1698431365
transform 1 0 7392 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2597_
timestamp 1698431365
transform -1 0 10528 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2598_
timestamp 1698431365
transform 1 0 12208 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2599_
timestamp 1698431365
transform 1 0 14672 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2600_
timestamp 1698431365
transform -1 0 14784 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2601_
timestamp 1698431365
transform 1 0 14560 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2602_
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2603_
timestamp 1698431365
transform -1 0 18256 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2604_
timestamp 1698431365
transform -1 0 15904 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2605_
timestamp 1698431365
transform -1 0 15008 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2606_
timestamp 1698431365
transform 1 0 12320 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2607_
timestamp 1698431365
transform -1 0 14448 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2608_
timestamp 1698431365
transform -1 0 14112 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2609_
timestamp 1698431365
transform -1 0 12992 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2610_
timestamp 1698431365
transform -1 0 13552 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2611_
timestamp 1698431365
transform -1 0 14224 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2612_
timestamp 1698431365
transform 1 0 15120 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2613_
timestamp 1698431365
transform 1 0 15008 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2614_
timestamp 1698431365
transform -1 0 7168 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2615_
timestamp 1698431365
transform -1 0 16800 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2616_
timestamp 1698431365
transform 1 0 14448 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2617_
timestamp 1698431365
transform -1 0 15232 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2618_
timestamp 1698431365
transform 1 0 15456 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2619_
timestamp 1698431365
transform -1 0 13104 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2620_
timestamp 1698431365
transform 1 0 7840 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2621_
timestamp 1698431365
transform 1 0 11200 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2622_
timestamp 1698431365
transform -1 0 12992 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2623_
timestamp 1698431365
transform 1 0 10080 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2624_
timestamp 1698431365
transform 1 0 11424 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2625_
timestamp 1698431365
transform 1 0 10976 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2626_
timestamp 1698431365
transform -1 0 12208 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2627_
timestamp 1698431365
transform -1 0 12432 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2628_
timestamp 1698431365
transform -1 0 10528 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2629_
timestamp 1698431365
transform -1 0 9632 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2630_
timestamp 1698431365
transform -1 0 9184 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2631_
timestamp 1698431365
transform -1 0 9296 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2632_
timestamp 1698431365
transform -1 0 7952 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2633_
timestamp 1698431365
transform -1 0 10304 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2634_
timestamp 1698431365
transform -1 0 8848 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2635_
timestamp 1698431365
transform -1 0 8736 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2636_
timestamp 1698431365
transform 1 0 11536 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2637_
timestamp 1698431365
transform -1 0 10304 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2638_
timestamp 1698431365
transform -1 0 10752 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2639_
timestamp 1698431365
transform -1 0 9968 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2640_
timestamp 1698431365
transform 1 0 5824 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2641_
timestamp 1698431365
transform -1 0 7392 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2642_
timestamp 1698431365
transform 1 0 5936 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2643_
timestamp 1698431365
transform -1 0 12992 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2644_
timestamp 1698431365
transform -1 0 3808 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2645_
timestamp 1698431365
transform 1 0 10080 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2646_
timestamp 1698431365
transform 1 0 7840 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2647_
timestamp 1698431365
transform 1 0 9968 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2648_
timestamp 1698431365
transform 1 0 4368 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2649_
timestamp 1698431365
transform -1 0 6048 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2650_
timestamp 1698431365
transform 1 0 3472 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2651_
timestamp 1698431365
transform -1 0 7280 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2652_
timestamp 1698431365
transform -1 0 8288 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2653_
timestamp 1698431365
transform -1 0 7728 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2654_
timestamp 1698431365
transform -1 0 6384 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2655_
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2656_
timestamp 1698431365
transform 1 0 4032 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2657_
timestamp 1698431365
transform -1 0 5264 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2658_
timestamp 1698431365
transform 1 0 2576 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2659_
timestamp 1698431365
transform -1 0 17024 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2660_
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2661_
timestamp 1698431365
transform 1 0 7840 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2662_
timestamp 1698431365
transform -1 0 7840 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2663_
timestamp 1698431365
transform -1 0 6496 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2664_
timestamp 1698431365
transform 1 0 4368 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2665_
timestamp 1698431365
transform -1 0 4816 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2666_
timestamp 1698431365
transform 1 0 3360 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2667_
timestamp 1698431365
transform 1 0 8288 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2668_
timestamp 1698431365
transform 1 0 7728 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2669_
timestamp 1698431365
transform -1 0 9184 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2670_
timestamp 1698431365
transform -1 0 6944 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2671_
timestamp 1698431365
transform 1 0 4368 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2672_
timestamp 1698431365
transform -1 0 5824 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2673_
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2674_
timestamp 1698431365
transform 1 0 2912 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2675_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2676_
timestamp 1698431365
transform -1 0 10752 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2677_
timestamp 1698431365
transform -1 0 7504 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2678_
timestamp 1698431365
transform 1 0 5936 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2679_
timestamp 1698431365
transform 1 0 3808 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2680_
timestamp 1698431365
transform 1 0 3584 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2681_
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2682_
timestamp 1698431365
transform 1 0 9744 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2683_
timestamp 1698431365
transform 1 0 13104 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2684_
timestamp 1698431365
transform -1 0 13776 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2685_
timestamp 1698431365
transform -1 0 11536 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2686_
timestamp 1698431365
transform 1 0 10304 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2687_
timestamp 1698431365
transform 1 0 11200 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2688_
timestamp 1698431365
transform -1 0 12880 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2689_
timestamp 1698431365
transform -1 0 13552 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2690_
timestamp 1698431365
transform 1 0 11760 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2691_
timestamp 1698431365
transform 1 0 11200 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2692_
timestamp 1698431365
transform -1 0 6944 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2693_
timestamp 1698431365
transform 1 0 9856 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2694_
timestamp 1698431365
transform -1 0 10864 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2695_
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2696_
timestamp 1698431365
transform 1 0 7280 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2697_
timestamp 1698431365
transform -1 0 9072 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2698_
timestamp 1698431365
transform -1 0 6832 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2699_
timestamp 1698431365
transform -1 0 4032 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2700_
timestamp 1698431365
transform 1 0 4256 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2701_
timestamp 1698431365
transform 1 0 6048 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2702_
timestamp 1698431365
transform 1 0 5152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2703_
timestamp 1698431365
transform 1 0 9072 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2704_
timestamp 1698431365
transform 1 0 7840 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2705_
timestamp 1698431365
transform -1 0 9184 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2706_
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2707_
timestamp 1698431365
transform 1 0 6048 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2708_
timestamp 1698431365
transform -1 0 3136 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2709_
timestamp 1698431365
transform 1 0 3136 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2710_
timestamp 1698431365
transform 1 0 7840 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2711_
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2712_
timestamp 1698431365
transform -1 0 10864 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2713_
timestamp 1698431365
transform -1 0 6384 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2714_
timestamp 1698431365
transform 1 0 4144 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2715_
timestamp 1698431365
transform -1 0 5040 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2716_
timestamp 1698431365
transform 1 0 3584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2717_
timestamp 1698431365
transform -1 0 9184 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2718_
timestamp 1698431365
transform -1 0 7616 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2719_
timestamp 1698431365
transform -1 0 6832 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2720_
timestamp 1698431365
transform -1 0 6272 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2721_
timestamp 1698431365
transform 1 0 3808 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2722_
timestamp 1698431365
transform -1 0 5376 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2723_
timestamp 1698431365
transform 1 0 3248 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2724_
timestamp 1698431365
transform 1 0 2352 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2725_
timestamp 1698431365
transform -1 0 10416 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2726_
timestamp 1698431365
transform 1 0 7728 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2727_
timestamp 1698431365
transform -1 0 7728 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2728_
timestamp 1698431365
transform -1 0 5600 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2729_
timestamp 1698431365
transform 1 0 3808 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2730_
timestamp 1698431365
transform -1 0 5264 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2731_
timestamp 1698431365
transform 1 0 3024 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2732_
timestamp 1698431365
transform -1 0 10976 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2733_
timestamp 1698431365
transform -1 0 7952 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2734_
timestamp 1698431365
transform -1 0 10416 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2735_
timestamp 1698431365
transform -1 0 7168 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2736_
timestamp 1698431365
transform -1 0 7728 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2737_
timestamp 1698431365
transform -1 0 6384 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2738_
timestamp 1698431365
transform 1 0 3808 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2739_
timestamp 1698431365
transform -1 0 5376 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2740_
timestamp 1698431365
transform -1 0 5264 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2741_
timestamp 1698431365
transform 1 0 2912 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2742_
timestamp 1698431365
transform 1 0 4368 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2743_
timestamp 1698431365
transform 1 0 7728 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2744_
timestamp 1698431365
transform -1 0 7840 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2745_
timestamp 1698431365
transform -1 0 6496 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2746_
timestamp 1698431365
transform 1 0 4816 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2747_
timestamp 1698431365
transform -1 0 4368 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2748_
timestamp 1698431365
transform 1 0 3136 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2749_
timestamp 1698431365
transform -1 0 9184 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2750_
timestamp 1698431365
transform -1 0 8400 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2751_
timestamp 1698431365
transform -1 0 7504 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2752_
timestamp 1698431365
transform -1 0 6608 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2753_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2754_
timestamp 1698431365
transform -1 0 4592 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2755_
timestamp 1698431365
transform 1 0 3024 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2756_
timestamp 1698431365
transform 1 0 5376 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2757_
timestamp 1698431365
transform 1 0 6496 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2758_
timestamp 1698431365
transform 1 0 5936 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2759_
timestamp 1698431365
transform -1 0 7280 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2760_
timestamp 1698431365
transform 1 0 6048 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2761_
timestamp 1698431365
transform 1 0 4144 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2762_
timestamp 1698431365
transform -1 0 6384 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2763_
timestamp 1698431365
transform 1 0 7504 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2764_
timestamp 1698431365
transform 1 0 7280 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2765_
timestamp 1698431365
transform 1 0 8960 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2766_
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2767_
timestamp 1698431365
transform 1 0 6496 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2768_
timestamp 1698431365
transform -1 0 6496 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2769_
timestamp 1698431365
transform -1 0 11200 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2770_
timestamp 1698431365
transform -1 0 10304 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2771_
timestamp 1698431365
transform -1 0 10752 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2772_
timestamp 1698431365
transform 1 0 9856 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2773_
timestamp 1698431365
transform 1 0 8288 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2774_
timestamp 1698431365
transform 1 0 10304 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2775_
timestamp 1698431365
transform -1 0 10976 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2776_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2777_
timestamp 1698431365
transform 1 0 11648 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2778_
timestamp 1698431365
transform 1 0 10640 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2779_
timestamp 1698431365
transform -1 0 12320 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2780_
timestamp 1698431365
transform 1 0 10864 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2781_
timestamp 1698431365
transform 1 0 11648 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2782_
timestamp 1698431365
transform 1 0 11424 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2783_
timestamp 1698431365
transform 1 0 16128 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2784_
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2785_
timestamp 1698431365
transform -1 0 12208 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2786_
timestamp 1698431365
transform 1 0 11424 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2787_
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2788_
timestamp 1698431365
transform 1 0 12208 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2789_
timestamp 1698431365
transform -1 0 12880 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2790_
timestamp 1698431365
transform 1 0 11872 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2791_
timestamp 1698431365
transform -1 0 14672 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2792_
timestamp 1698431365
transform 1 0 12768 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2793_
timestamp 1698431365
transform -1 0 14672 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2794_
timestamp 1698431365
transform -1 0 13328 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2795_
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2796_
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2797_
timestamp 1698431365
transform -1 0 14560 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2798_
timestamp 1698431365
transform 1 0 13328 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2799_
timestamp 1698431365
transform 1 0 14336 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2800_
timestamp 1698431365
transform 1 0 13440 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2801_
timestamp 1698431365
transform -1 0 14784 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2802_
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2803_
timestamp 1698431365
transform -1 0 14784 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2804_
timestamp 1698431365
transform 1 0 12880 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2805_
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2806_
timestamp 1698431365
transform 1 0 14784 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2807_
timestamp 1698431365
transform -1 0 13440 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2808_
timestamp 1698431365
transform -1 0 14336 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2809_
timestamp 1698431365
transform 1 0 18928 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2810_
timestamp 1698431365
transform -1 0 15232 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2811_
timestamp 1698431365
transform 1 0 14784 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2812_
timestamp 1698431365
transform -1 0 16016 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2813_
timestamp 1698431365
transform -1 0 17024 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2814_
timestamp 1698431365
transform 1 0 15792 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2815_
timestamp 1698431365
transform -1 0 17920 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2816_
timestamp 1698431365
transform 1 0 16576 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2817_
timestamp 1698431365
transform 1 0 16016 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2818_
timestamp 1698431365
transform 1 0 15904 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2819_
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2820_
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2821_
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2822_
timestamp 1698431365
transform -1 0 18816 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2823_
timestamp 1698431365
transform 1 0 17808 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2824_
timestamp 1698431365
transform 1 0 16576 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2825_
timestamp 1698431365
transform 1 0 17248 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2826_
timestamp 1698431365
transform 1 0 19264 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2827_
timestamp 1698431365
transform 1 0 18704 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2828_
timestamp 1698431365
transform 1 0 20496 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2829_
timestamp 1698431365
transform 1 0 19600 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2830_
timestamp 1698431365
transform -1 0 17024 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2831_
timestamp 1698431365
transform 1 0 17360 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2832_
timestamp 1698431365
transform 1 0 18592 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2833_
timestamp 1698431365
transform -1 0 19824 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2834_
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2835_
timestamp 1698431365
transform -1 0 20496 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2836_
timestamp 1698431365
transform 1 0 15904 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2837_
timestamp 1698431365
transform 1 0 15344 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2838_
timestamp 1698431365
transform 1 0 17136 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2839_
timestamp 1698431365
transform -1 0 18704 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2840_
timestamp 1698431365
transform 1 0 18592 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2841_
timestamp 1698431365
transform 1 0 18816 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2842_
timestamp 1698431365
transform 1 0 14224 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2843_
timestamp 1698431365
transform 1 0 13776 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2844_
timestamp 1698431365
transform -1 0 18704 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2845_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2846_
timestamp 1698431365
transform 1 0 15344 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2847_
timestamp 1698431365
transform 1 0 15792 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2848_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7840 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2849_
timestamp 1698431365
transform 1 0 4928 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2850_
timestamp 1698431365
transform 1 0 7504 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2851_
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2852_
timestamp 1698431365
transform 1 0 30464 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2853_
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2854_
timestamp 1698431365
transform 1 0 27328 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2855_
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2856_
timestamp 1698431365
transform 1 0 21616 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2857_
timestamp 1698431365
transform -1 0 30352 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2858_
timestamp 1698431365
transform 1 0 37296 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2859_
timestamp 1698431365
transform 1 0 34608 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2860_
timestamp 1698431365
transform 1 0 34272 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2861_
timestamp 1698431365
transform 1 0 34944 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2862_
timestamp 1698431365
transform 1 0 33040 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2863_
timestamp 1698431365
transform 1 0 42448 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2864_
timestamp 1698431365
transform 1 0 41216 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2865_
timestamp 1698431365
transform 1 0 42224 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2866_
timestamp 1698431365
transform 1 0 45024 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2867_
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2868_
timestamp 1698431365
transform 1 0 48160 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2869_
timestamp 1698431365
transform 1 0 48608 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2870_
timestamp 1698431365
transform 1 0 49168 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2871_
timestamp 1698431365
transform 1 0 53536 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2872_
timestamp 1698431365
transform -1 0 56336 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2873_
timestamp 1698431365
transform 1 0 52864 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2874_
timestamp 1698431365
transform 1 0 52528 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2875_
timestamp 1698431365
transform 1 0 41104 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2876_
timestamp 1698431365
transform 1 0 38640 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2877_
timestamp 1698431365
transform 1 0 25536 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2878_
timestamp 1698431365
transform 1 0 29456 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2879_
timestamp 1698431365
transform -1 0 27888 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2880_
timestamp 1698431365
transform 1 0 26208 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2881_
timestamp 1698431365
transform -1 0 21168 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2882_
timestamp 1698431365
transform 1 0 33600 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2883_
timestamp 1698431365
transform -1 0 8848 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2884_
timestamp 1698431365
transform 1 0 19152 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2885_
timestamp 1698431365
transform 1 0 18928 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2886_
timestamp 1698431365
transform 1 0 21616 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2887_
timestamp 1698431365
transform 1 0 21392 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2888_
timestamp 1698431365
transform 1 0 20272 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2889_
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2890_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2891_
timestamp 1698431365
transform 1 0 27216 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2892_
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2893_
timestamp 1698431365
transform 1 0 36624 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2894_
timestamp 1698431365
transform -1 0 42784 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2895_
timestamp 1698431365
transform 1 0 42560 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2896_
timestamp 1698431365
transform -1 0 48944 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2897_
timestamp 1698431365
transform -1 0 51968 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2898_
timestamp 1698431365
transform -1 0 53536 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2899_
timestamp 1698431365
transform -1 0 53200 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2900_
timestamp 1698431365
transform -1 0 55440 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2901_
timestamp 1698431365
transform -1 0 57120 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2902_
timestamp 1698431365
transform 1 0 55104 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2903_
timestamp 1698431365
transform 1 0 54880 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2904_
timestamp 1698431365
transform 1 0 55104 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2905_
timestamp 1698431365
transform 1 0 55104 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2906_
timestamp 1698431365
transform 1 0 55104 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2907_
timestamp 1698431365
transform -1 0 56224 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2908_
timestamp 1698431365
transform 1 0 41552 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2909_
timestamp 1698431365
transform 1 0 31360 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2910_
timestamp 1698431365
transform -1 0 32256 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2911_
timestamp 1698431365
transform 1 0 24752 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2912_
timestamp 1698431365
transform 1 0 17248 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2913_
timestamp 1698431365
transform 1 0 14896 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2914_
timestamp 1698431365
transform 1 0 12432 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2915_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2916_
timestamp 1698431365
transform 1 0 16912 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2917_
timestamp 1698431365
transform 1 0 13776 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2918_
timestamp 1698431365
transform 1 0 17472 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2919_
timestamp 1698431365
transform 1 0 19376 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2920_
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2921_
timestamp 1698431365
transform 1 0 20496 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2922_
timestamp 1698431365
transform 1 0 29792 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2923_
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2924_
timestamp 1698431365
transform 1 0 29456 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2925_
timestamp 1698431365
transform 1 0 30464 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2926_
timestamp 1698431365
transform 1 0 30688 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2927_
timestamp 1698431365
transform 1 0 38864 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2928_
timestamp 1698431365
transform 1 0 37296 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2929_
timestamp 1698431365
transform 1 0 41216 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2930_
timestamp 1698431365
transform 1 0 41440 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2931_
timestamp 1698431365
transform 1 0 44912 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2932_
timestamp 1698431365
transform -1 0 49952 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2933_
timestamp 1698431365
transform 1 0 45136 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2934_
timestamp 1698431365
transform 1 0 47152 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2935_
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2936_
timestamp 1698431365
transform -1 0 55776 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2937_
timestamp 1698431365
transform -1 0 54320 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2938_
timestamp 1698431365
transform -1 0 53648 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2939_
timestamp 1698431365
transform 1 0 36960 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2940_
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2941_
timestamp 1698431365
transform 1 0 22960 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2942_
timestamp 1698431365
transform 1 0 23968 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2943_
timestamp 1698431365
transform 1 0 13776 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2944_
timestamp 1698431365
transform 1 0 10416 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2945_
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2946_
timestamp 1698431365
transform 1 0 13776 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2947_
timestamp 1698431365
transform 1 0 12992 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2948_
timestamp 1698431365
transform 1 0 11984 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2949_
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2950_
timestamp 1698431365
transform 1 0 13664 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2951_
timestamp 1698431365
transform -1 0 17696 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2952_
timestamp 1698431365
transform 1 0 18704 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2953_
timestamp 1698431365
transform 1 0 17696 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2954_
timestamp 1698431365
transform 1 0 23296 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2955_
timestamp 1698431365
transform 1 0 23520 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2956_
timestamp 1698431365
transform 1 0 26656 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2957_
timestamp 1698431365
transform 1 0 27440 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2958_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35840 0 -1 56448
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2959_
timestamp 1698431365
transform 1 0 34608 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2960_
timestamp 1698431365
transform 1 0 37520 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2961_
timestamp 1698431365
transform -1 0 43120 0 -1 56448
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2962_
timestamp 1698431365
transform -1 0 45136 0 -1 53312
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2963_
timestamp 1698431365
transform 1 0 42448 0 -1 54880
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2964_
timestamp 1698431365
transform -1 0 48608 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2965_
timestamp 1698431365
transform -1 0 48720 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2966_
timestamp 1698431365
transform 1 0 48608 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2967_
timestamp 1698431365
transform -1 0 53312 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2968_
timestamp 1698431365
transform 1 0 51520 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2969_
timestamp 1698431365
transform -1 0 52304 0 -1 51744
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2970_
timestamp 1698431365
transform 1 0 35168 0 -1 51744
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2971_
timestamp 1698431365
transform 1 0 33152 0 1 51744
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2972_
timestamp 1698431365
transform 1 0 25424 0 -1 51744
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2973_
timestamp 1698431365
transform 1 0 24416 0 1 50176
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2974_
timestamp 1698431365
transform 1 0 9856 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2975_
timestamp 1698431365
transform 1 0 9408 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2976_
timestamp 1698431365
transform 1 0 8176 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2977_
timestamp 1698431365
transform 1 0 7952 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2978_
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2979_
timestamp 1698431365
transform 1 0 11312 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2980_
timestamp 1698431365
transform 1 0 24528 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2981_
timestamp 1698431365
transform 1 0 22624 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2982_
timestamp 1698431365
transform -1 0 34160 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2983_
timestamp 1698431365
transform 1 0 23632 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2984_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2985_
timestamp 1698431365
transform 1 0 22288 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2986_
timestamp 1698431365
transform 1 0 21616 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2987_
timestamp 1698431365
transform -1 0 32816 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2988_
timestamp 1698431365
transform 1 0 31248 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2989_
timestamp 1698431365
transform 1 0 34272 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2990_
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2991_
timestamp 1698431365
transform 1 0 42672 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2992_
timestamp 1698431365
transform 1 0 38864 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2993_
timestamp 1698431365
transform 1 0 39424 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2994_
timestamp 1698431365
transform 1 0 41776 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2995_
timestamp 1698431365
transform 1 0 45136 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2996_
timestamp 1698431365
transform 1 0 45136 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2997_
timestamp 1698431365
transform 1 0 46928 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2998_
timestamp 1698431365
transform 1 0 45136 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2999_
timestamp 1698431365
transform 1 0 44912 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3000_
timestamp 1698431365
transform 1 0 47936 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3001_
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3002_
timestamp 1698431365
transform 1 0 47264 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3003_
timestamp 1698431365
transform 1 0 44800 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3004_
timestamp 1698431365
transform 1 0 37296 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3005_
timestamp 1698431365
transform -1 0 44016 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3006_
timestamp 1698431365
transform 1 0 25536 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3007_
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3008_
timestamp 1698431365
transform 1 0 19264 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3009_
timestamp 1698431365
transform -1 0 22176 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3010_
timestamp 1698431365
transform 1 0 12096 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3011_
timestamp 1698431365
transform 1 0 15120 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3012_
timestamp 1698431365
transform -1 0 10192 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3013_
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3014_
timestamp 1698431365
transform 1 0 15680 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3015_
timestamp 1698431365
transform 1 0 4368 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3016_
timestamp 1698431365
transform 1 0 14672 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3017_
timestamp 1698431365
transform 1 0 10304 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3018_
timestamp 1698431365
transform 1 0 7392 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3019_
timestamp 1698431365
transform 1 0 4480 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3020_
timestamp 1698431365
transform 1 0 1680 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3021_
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3022_
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3023_
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3024_
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3025_
timestamp 1698431365
transform -1 0 12656 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3026_
timestamp 1698431365
transform 1 0 6160 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3027_
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3028_
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3029_
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3030_
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3031_
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3032_
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3033_
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3034_
timestamp 1698431365
transform 1 0 1792 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3035_
timestamp 1698431365
transform 1 0 4816 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3036_
timestamp 1698431365
transform 1 0 7168 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3037_
timestamp 1698431365
transform -1 0 11648 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3038_
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3039_
timestamp 1698431365
transform -1 0 16128 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3040_
timestamp 1698431365
transform 1 0 11648 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3041_
timestamp 1698431365
transform 1 0 11536 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3042_
timestamp 1698431365
transform -1 0 18704 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3043_
timestamp 1698431365
transform -1 0 20496 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3044_
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3045_
timestamp 1698431365
transform -1 0 22512 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3046_
timestamp 1698431365
transform -1 0 20496 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3047_
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3048_
timestamp 1698431365
transform -1 0 8624 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1425__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31472 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1428__A3
timestamp 1698431365
transform -1 0 9072 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1435__I
timestamp 1698431365
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__I0
timestamp 1698431365
transform -1 0 21952 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__S
timestamp 1698431365
transform -1 0 22400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1439__I
timestamp 1698431365
transform 1 0 38416 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1440__I
timestamp 1698431365
transform -1 0 31360 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1445__A1
timestamp 1698431365
transform 1 0 30576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1447__I
timestamp 1698431365
transform 1 0 33600 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1449__I
timestamp 1698431365
transform 1 0 33600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__A2
timestamp 1698431365
transform 1 0 31584 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__I
timestamp 1698431365
transform -1 0 35728 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A2
timestamp 1698431365
transform 1 0 20048 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__B
timestamp 1698431365
transform -1 0 20496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1465__I
timestamp 1698431365
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__B
timestamp 1698431365
transform 1 0 30688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A1
timestamp 1698431365
transform -1 0 29792 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__B
timestamp 1698431365
transform 1 0 31584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1470__A1
timestamp 1698431365
transform 1 0 31808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1473__B
timestamp 1698431365
transform -1 0 19712 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__B
timestamp 1698431365
transform 1 0 30128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1479__B
timestamp 1698431365
transform -1 0 30352 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1481__B
timestamp 1698431365
transform 1 0 29232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1485__A1
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__I
timestamp 1698431365
transform 1 0 24528 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A1
timestamp 1698431365
transform 1 0 24976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1493__A2
timestamp 1698431365
transform 1 0 27664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__A1
timestamp 1698431365
transform 1 0 26432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1495__I
timestamp 1698431365
transform 1 0 21616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__A1
timestamp 1698431365
transform 1 0 24192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A1
timestamp 1698431365
transform 1 0 25872 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A2
timestamp 1698431365
transform 1 0 27216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__A1
timestamp 1698431365
transform 1 0 28112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__I
timestamp 1698431365
transform 1 0 38864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1509__B
timestamp 1698431365
transform 1 0 24976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__A1
timestamp 1698431365
transform 1 0 27552 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__A1
timestamp 1698431365
transform -1 0 27888 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__B
timestamp 1698431365
transform -1 0 27888 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1515__A1
timestamp 1698431365
transform -1 0 28672 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__I
timestamp 1698431365
transform 1 0 33152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A2
timestamp 1698431365
transform 1 0 37968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A4
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A1
timestamp 1698431365
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A2
timestamp 1698431365
transform 1 0 36512 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__B
timestamp 1698431365
transform 1 0 36064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A1
timestamp 1698431365
transform -1 0 35168 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A3
timestamp 1698431365
transform -1 0 36736 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__A1
timestamp 1698431365
transform -1 0 37520 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__I
timestamp 1698431365
transform -1 0 25200 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__A1
timestamp 1698431365
transform 1 0 34160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__A2
timestamp 1698431365
transform 1 0 33712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1534__A1
timestamp 1698431365
transform -1 0 35392 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1534__A2
timestamp 1698431365
transform 1 0 32704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1538__A1
timestamp 1698431365
transform -1 0 35840 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1541__A2
timestamp 1698431365
transform 1 0 31808 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1542__A1
timestamp 1698431365
transform 1 0 35056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__B
timestamp 1698431365
transform -1 0 31808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1549__I
timestamp 1698431365
transform 1 0 37408 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A1
timestamp 1698431365
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__A1
timestamp 1698431365
transform -1 0 37744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A1
timestamp 1698431365
transform -1 0 37296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A2
timestamp 1698431365
transform 1 0 34720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A1
timestamp 1698431365
transform 1 0 33824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__A1
timestamp 1698431365
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__A1
timestamp 1698431365
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1567__A1
timestamp 1698431365
transform 1 0 36736 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__A1
timestamp 1698431365
transform 1 0 37184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__I
timestamp 1698431365
transform 1 0 46256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1572__I
timestamp 1698431365
transform 1 0 41440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1573__A1
timestamp 1698431365
transform -1 0 38864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__A2
timestamp 1698431365
transform 1 0 37968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__A1
timestamp 1698431365
transform -1 0 44128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__A2
timestamp 1698431365
transform 1 0 40880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__A1
timestamp 1698431365
transform -1 0 43568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1581__A2
timestamp 1698431365
transform -1 0 40096 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__B
timestamp 1698431365
transform -1 0 39648 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__I
timestamp 1698431365
transform -1 0 42784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1591__A1
timestamp 1698431365
transform 1 0 44912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1592__A1
timestamp 1698431365
transform 1 0 43680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1594__A1
timestamp 1698431365
transform -1 0 41664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1596__A2
timestamp 1698431365
transform 1 0 43568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A1
timestamp 1698431365
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A2
timestamp 1698431365
transform 1 0 37520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A3
timestamp 1698431365
transform 1 0 38304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__A1
timestamp 1698431365
transform 1 0 42000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__A2
timestamp 1698431365
transform 1 0 40992 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__A1
timestamp 1698431365
transform -1 0 43568 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__A2
timestamp 1698431365
transform 1 0 42112 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__B
timestamp 1698431365
transform 1 0 43792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__I
timestamp 1698431365
transform 1 0 38416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A1
timestamp 1698431365
transform 1 0 44128 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A2
timestamp 1698431365
transform 1 0 42560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__B
timestamp 1698431365
transform -1 0 43904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__A1
timestamp 1698431365
transform -1 0 46032 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A1
timestamp 1698431365
transform -1 0 45136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__A1
timestamp 1698431365
transform 1 0 45360 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__A2
timestamp 1698431365
transform 1 0 46368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__A3
timestamp 1698431365
transform 1 0 44912 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__B
timestamp 1698431365
transform 1 0 49504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1635__A1
timestamp 1698431365
transform 1 0 48832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__A1
timestamp 1698431365
transform 1 0 47488 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__A1
timestamp 1698431365
transform 1 0 48048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A2
timestamp 1698431365
transform -1 0 47040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__B
timestamp 1698431365
transform 1 0 45360 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__B
timestamp 1698431365
transform -1 0 49952 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__A1
timestamp 1698431365
transform 1 0 48832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__A1
timestamp 1698431365
transform 1 0 49056 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__A3
timestamp 1698431365
transform 1 0 47040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A2
timestamp 1698431365
transform 1 0 49952 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__B2
timestamp 1698431365
transform -1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__B
timestamp 1698431365
transform 1 0 55440 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A1
timestamp 1698431365
transform 1 0 56672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A1
timestamp 1698431365
transform 1 0 56560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A2
timestamp 1698431365
transform 1 0 50400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__B2
timestamp 1698431365
transform 1 0 50848 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__B
timestamp 1698431365
transform 1 0 50848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A1
timestamp 1698431365
transform 1 0 50736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__A1
timestamp 1698431365
transform 1 0 50288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__A1
timestamp 1698431365
transform 1 0 40208 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__A1
timestamp 1698431365
transform 1 0 40992 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__B2
timestamp 1698431365
transform -1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__B
timestamp 1698431365
transform 1 0 41104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__A1
timestamp 1698431365
transform 1 0 38416 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__A1
timestamp 1698431365
transform 1 0 27328 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__B
timestamp 1698431365
transform -1 0 31248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__A1
timestamp 1698431365
transform 1 0 28672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__A1
timestamp 1698431365
transform 1 0 30800 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1744__B
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__A1
timestamp 1698431365
transform 1 0 29232 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__A1
timestamp 1698431365
transform 1 0 29232 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__B
timestamp 1698431365
transform 1 0 23296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__B
timestamp 1698431365
transform 1 0 22288 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A1
timestamp 1698431365
transform 1 0 20160 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__B2
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__B
timestamp 1698431365
transform -1 0 18480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__A1
timestamp 1698431365
transform 1 0 31584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__A1
timestamp 1698431365
transform -1 0 34048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A1
timestamp 1698431365
transform -1 0 33824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__A4
timestamp 1698431365
transform -1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__A1
timestamp 1698431365
transform 1 0 15792 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__A4
timestamp 1698431365
transform 1 0 41888 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__A3
timestamp 1698431365
transform -1 0 15904 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__I
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__A2
timestamp 1698431365
transform 1 0 14784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__I
timestamp 1698431365
transform 1 0 19376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__A2
timestamp 1698431365
transform 1 0 19040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__I
timestamp 1698431365
transform 1 0 12208 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__I
timestamp 1698431365
transform -1 0 13552 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__I
timestamp 1698431365
transform 1 0 20048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__I
timestamp 1698431365
transform -1 0 20944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__I
timestamp 1698431365
transform -1 0 22512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__I
timestamp 1698431365
transform 1 0 43008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__I
timestamp 1698431365
transform 1 0 44912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__I
timestamp 1698431365
transform -1 0 46032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__I
timestamp 1698431365
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__I
timestamp 1698431365
transform 1 0 52752 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__I
timestamp 1698431365
transform 1 0 53872 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__I
timestamp 1698431365
transform 1 0 53312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__I
timestamp 1698431365
transform 1 0 53648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__I
timestamp 1698431365
transform 1 0 53760 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__A2
timestamp 1698431365
transform 1 0 56336 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1886__A2
timestamp 1698431365
transform 1 0 56672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__A2
timestamp 1698431365
transform -1 0 55776 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__I
timestamp 1698431365
transform 1 0 16016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__I
timestamp 1698431365
transform -1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__A2
timestamp 1698431365
transform -1 0 42784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__B1
timestamp 1698431365
transform 1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__I
timestamp 1698431365
transform 1 0 16128 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__I
timestamp 1698431365
transform -1 0 18592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__B1
timestamp 1698431365
transform 1 0 31024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__B1
timestamp 1698431365
transform 1 0 29120 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__B1
timestamp 1698431365
transform 1 0 27216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1903__I
timestamp 1698431365
transform 1 0 18032 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__I
timestamp 1698431365
transform 1 0 17808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__A2
timestamp 1698431365
transform 1 0 16576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A2
timestamp 1698431365
transform -1 0 16576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A2
timestamp 1698431365
transform 1 0 14896 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A2
timestamp 1698431365
transform -1 0 14000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A2
timestamp 1698431365
transform 1 0 52864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1963__B
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__A2
timestamp 1698431365
transform 1 0 28896 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A2
timestamp 1698431365
transform -1 0 42112 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A2
timestamp 1698431365
transform 1 0 42336 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1979__A2
timestamp 1698431365
transform 1 0 37184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__A2
timestamp 1698431365
transform -1 0 33824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__A2
timestamp 1698431365
transform -1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A2
timestamp 1698431365
transform -1 0 37296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__B1
timestamp 1698431365
transform -1 0 34272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A2
timestamp 1698431365
transform 1 0 42224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__A2
timestamp 1698431365
transform 1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__A2
timestamp 1698431365
transform -1 0 45136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__A2
timestamp 1698431365
transform 1 0 44016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__A2
timestamp 1698431365
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A1
timestamp 1698431365
transform 1 0 46928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__A1
timestamp 1698431365
transform -1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A2
timestamp 1698431365
transform 1 0 14896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A2
timestamp 1698431365
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__I
timestamp 1698431365
transform -1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2065__A2
timestamp 1698431365
transform 1 0 19376 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__I
timestamp 1698431365
transform 1 0 19040 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__I
timestamp 1698431365
transform -1 0 30464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__A2
timestamp 1698431365
transform -1 0 29456 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__I
timestamp 1698431365
transform 1 0 22960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2098__I
timestamp 1698431365
transform 1 0 40320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2108__I
timestamp 1698431365
transform 1 0 48160 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2118__I
timestamp 1698431365
transform 1 0 51296 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__I
timestamp 1698431365
transform 1 0 34832 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__A1
timestamp 1698431365
transform -1 0 50512 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__I
timestamp 1698431365
transform 1 0 35728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2134__I
timestamp 1698431365
transform 1 0 21392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A1
timestamp 1698431365
transform 1 0 24640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2144__I
timestamp 1698431365
transform -1 0 20944 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2145__A2
timestamp 1698431365
transform -1 0 15008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__A2
timestamp 1698431365
transform 1 0 16576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2151__I
timestamp 1698431365
transform 1 0 18144 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2152__A2
timestamp 1698431365
transform -1 0 15456 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__A2
timestamp 1698431365
transform 1 0 16800 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__I
timestamp 1698431365
transform 1 0 18592 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2161__I
timestamp 1698431365
transform -1 0 22176 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__I
timestamp 1698431365
transform -1 0 21728 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2171__I
timestamp 1698431365
transform 1 0 43008 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2177__I
timestamp 1698431365
transform 1 0 18368 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2178__I
timestamp 1698431365
transform 1 0 40208 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__I
timestamp 1698431365
transform 1 0 46592 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2198__I
timestamp 1698431365
transform 1 0 48160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2204__B1
timestamp 1698431365
transform 1 0 50400 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2206__B1
timestamp 1698431365
transform 1 0 49504 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2206__B2
timestamp 1698431365
transform -1 0 49392 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__I
timestamp 1698431365
transform 1 0 24192 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2209__A1
timestamp 1698431365
transform 1 0 37520 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2209__B1
timestamp 1698431365
transform -1 0 37296 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2211__B1
timestamp 1698431365
transform -1 0 37296 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2213__I
timestamp 1698431365
transform -1 0 15008 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__B1
timestamp 1698431365
transform 1 0 24640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2216__B1
timestamp 1698431365
transform -1 0 27664 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2216__B2
timestamp 1698431365
transform 1 0 28224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__I
timestamp 1698431365
transform 1 0 11760 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2219__I
timestamp 1698431365
transform 1 0 10416 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2220__A1
timestamp 1698431365
transform 1 0 12880 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2220__B1
timestamp 1698431365
transform 1 0 13328 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2222__B1
timestamp 1698431365
transform 1 0 12880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2224__B1
timestamp 1698431365
transform -1 0 12768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2226__B1
timestamp 1698431365
transform 1 0 11424 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2228__A2
timestamp 1698431365
transform 1 0 15120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2228__B
timestamp 1698431365
transform 1 0 15568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2230__I
timestamp 1698431365
transform -1 0 11424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2232__I
timestamp 1698431365
transform 1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__I
timestamp 1698431365
transform 1 0 15456 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__A1
timestamp 1698431365
transform 1 0 14224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__I
timestamp 1698431365
transform -1 0 20720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2240__I
timestamp 1698431365
transform -1 0 32032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2242__I
timestamp 1698431365
transform 1 0 22960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2244__I
timestamp 1698431365
transform -1 0 31024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__A1
timestamp 1698431365
transform 1 0 27776 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2247__A2
timestamp 1698431365
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__A1
timestamp 1698431365
transform 1 0 26432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__A2
timestamp 1698431365
transform 1 0 25312 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__A1
timestamp 1698431365
transform -1 0 26768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2250__I
timestamp 1698431365
transform 1 0 17920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2255__A1
timestamp 1698431365
transform 1 0 20272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2259__A1
timestamp 1698431365
transform -1 0 34048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__I
timestamp 1698431365
transform 1 0 17024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2263__A1
timestamp 1698431365
transform 1 0 28336 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2264__A1
timestamp 1698431365
transform -1 0 30016 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__I
timestamp 1698431365
transform -1 0 33824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__I
timestamp 1698431365
transform -1 0 30464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2270__I
timestamp 1698431365
transform -1 0 31360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2272__I
timestamp 1698431365
transform -1 0 31360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2274__A2
timestamp 1698431365
transform 1 0 33936 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2275__A1
timestamp 1698431365
transform -1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2280__A1
timestamp 1698431365
transform 1 0 28000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2281__A1
timestamp 1698431365
transform 1 0 32592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2283__A1
timestamp 1698431365
transform 1 0 29120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2286__A2
timestamp 1698431365
transform 1 0 35728 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2286__A3
timestamp 1698431365
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2287__A1
timestamp 1698431365
transform 1 0 36176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2288__A2
timestamp 1698431365
transform -1 0 27888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__B
timestamp 1698431365
transform 1 0 31024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__A1
timestamp 1698431365
transform 1 0 30576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2298__A1
timestamp 1698431365
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2298__A2
timestamp 1698431365
transform 1 0 34384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2298__A3
timestamp 1698431365
transform 1 0 34832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2298__A4
timestamp 1698431365
transform 1 0 35280 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2303__A1
timestamp 1698431365
transform 1 0 30912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2309__A1
timestamp 1698431365
transform 1 0 27216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2309__A2
timestamp 1698431365
transform -1 0 26992 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2310__A1
timestamp 1698431365
transform 1 0 24192 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2314__A2
timestamp 1698431365
transform 1 0 27440 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2316__B
timestamp 1698431365
transform -1 0 28336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2318__A1
timestamp 1698431365
transform 1 0 28000 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2319__I0
timestamp 1698431365
transform 1 0 30240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__B
timestamp 1698431365
transform 1 0 29344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2330__A1
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2331__A2
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2332__A1
timestamp 1698431365
transform -1 0 23968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2333__I
timestamp 1698431365
transform -1 0 31136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__B
timestamp 1698431365
transform -1 0 32704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2337__A2
timestamp 1698431365
transform -1 0 26880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2338__B
timestamp 1698431365
transform -1 0 31360 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2349__B
timestamp 1698431365
transform 1 0 34272 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__A1
timestamp 1698431365
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2355__I
timestamp 1698431365
transform -1 0 36512 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2356__B
timestamp 1698431365
transform 1 0 34720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2358__A2
timestamp 1698431365
transform -1 0 34720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2361__A1
timestamp 1698431365
transform 1 0 35168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2364__A1
timestamp 1698431365
transform 1 0 38192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2365__I
timestamp 1698431365
transform 1 0 15232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2377__A1
timestamp 1698431365
transform 1 0 39984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__A1
timestamp 1698431365
transform -1 0 37408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__S
timestamp 1698431365
transform -1 0 40768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2386__A2
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2387__A1
timestamp 1698431365
transform 1 0 41776 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__A1
timestamp 1698431365
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2396__A1
timestamp 1698431365
transform 1 0 43568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2400__A1
timestamp 1698431365
transform 1 0 39424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2401__A1
timestamp 1698431365
transform -1 0 35952 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2402__A1
timestamp 1698431365
transform 1 0 37184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2405__A1
timestamp 1698431365
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2406__A1
timestamp 1698431365
transform 1 0 38528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2408__A1
timestamp 1698431365
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2409__A1
timestamp 1698431365
transform -1 0 36848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2409__A2
timestamp 1698431365
transform -1 0 37296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2410__A1
timestamp 1698431365
transform 1 0 40432 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2411__B
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2412__A1
timestamp 1698431365
transform 1 0 41440 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__B2
timestamp 1698431365
transform 1 0 39536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2417__A1
timestamp 1698431365
transform -1 0 45136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2417__A2
timestamp 1698431365
transform 1 0 44016 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2418__A1
timestamp 1698431365
transform 1 0 41440 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2422__A1
timestamp 1698431365
transform 1 0 44688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__A1
timestamp 1698431365
transform 1 0 39088 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2424__A1
timestamp 1698431365
transform 1 0 39984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2425__B2
timestamp 1698431365
transform -1 0 43120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2426__I
timestamp 1698431365
transform -1 0 43568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2427__I0
timestamp 1698431365
transform 1 0 48832 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2429__A1
timestamp 1698431365
transform -1 0 38192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2429__A2
timestamp 1698431365
transform -1 0 37744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2430__A1
timestamp 1698431365
transform 1 0 38080 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2430__A2
timestamp 1698431365
transform 1 0 37632 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2432__I
timestamp 1698431365
transform 1 0 40208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2434__I
timestamp 1698431365
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2436__A1
timestamp 1698431365
transform 1 0 43904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__A1
timestamp 1698431365
transform 1 0 46592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__I
timestamp 1698431365
transform 1 0 40208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2440__B2
timestamp 1698431365
transform 1 0 44912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__A1
timestamp 1698431365
transform 1 0 40208 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A1
timestamp 1698431365
transform 1 0 47264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2449__A1
timestamp 1698431365
transform 1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2450__A1
timestamp 1698431365
transform 1 0 40992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2451__I0
timestamp 1698431365
transform 1 0 47824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2453__I
timestamp 1698431365
transform 1 0 40992 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2458__A2
timestamp 1698431365
transform 1 0 41216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__A1
timestamp 1698431365
transform 1 0 44576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__A1
timestamp 1698431365
transform 1 0 42896 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__C
timestamp 1698431365
transform -1 0 43568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2464__A2
timestamp 1698431365
transform 1 0 45920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2469__B
timestamp 1698431365
transform 1 0 43792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__A1
timestamp 1698431365
transform 1 0 43456 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2471__A1
timestamp 1698431365
transform 1 0 44352 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2472__A1
timestamp 1698431365
transform 1 0 44240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A1
timestamp 1698431365
transform 1 0 41440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A2
timestamp 1698431365
transform 1 0 41888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A4
timestamp 1698431365
transform 1 0 42336 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2482__A1
timestamp 1698431365
transform -1 0 41216 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__A1
timestamp 1698431365
transform 1 0 44128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__A1
timestamp 1698431365
transform 1 0 44688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__C
timestamp 1698431365
transform 1 0 43680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__A2
timestamp 1698431365
transform 1 0 48496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__A1
timestamp 1698431365
transform -1 0 37856 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2487__A1
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2489__B
timestamp 1698431365
transform 1 0 45472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2491__A1
timestamp 1698431365
transform 1 0 45024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2492__I
timestamp 1698431365
transform 1 0 44128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2497__A1
timestamp 1698431365
transform 1 0 43232 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A1
timestamp 1698431365
transform -1 0 39872 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A2
timestamp 1698431365
transform -1 0 41216 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2501__A1
timestamp 1698431365
transform -1 0 42000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2501__B
timestamp 1698431365
transform 1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2502__A1
timestamp 1698431365
transform -1 0 41552 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2503__A1
timestamp 1698431365
transform 1 0 42448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__A2
timestamp 1698431365
transform 1 0 47152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A1
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__B
timestamp 1698431365
transform 1 0 42000 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__S
timestamp 1698431365
transform 1 0 43680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2513__A1
timestamp 1698431365
transform 1 0 43120 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2515__A1
timestamp 1698431365
transform -1 0 37296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A1
timestamp 1698431365
transform -1 0 37296 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2521__A1
timestamp 1698431365
transform 1 0 37968 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__A1
timestamp 1698431365
transform 1 0 37520 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2527__A1
timestamp 1698431365
transform -1 0 39424 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2528__A1
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2528__B
timestamp 1698431365
transform 1 0 35056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2529__A1
timestamp 1698431365
transform -1 0 39088 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2530__B2
timestamp 1698431365
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__A1
timestamp 1698431365
transform -1 0 38192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__A2
timestamp 1698431365
transform 1 0 38416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__A1
timestamp 1698431365
transform 1 0 35168 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__A1
timestamp 1698431365
transform -1 0 34048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2540__A1
timestamp 1698431365
transform 1 0 33824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2546__A1
timestamp 1698431365
transform -1 0 35392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2547__B
timestamp 1698431365
transform 1 0 30912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__A1
timestamp 1698431365
transform -1 0 31136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__A1
timestamp 1698431365
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2550__A1
timestamp 1698431365
transform 1 0 34720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__A1
timestamp 1698431365
transform 1 0 24976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__B
timestamp 1698431365
transform 1 0 26208 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2554__A1
timestamp 1698431365
transform 1 0 23968 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2558__A1
timestamp 1698431365
transform 1 0 21504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2559__A1
timestamp 1698431365
transform -1 0 24976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__A1
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__A2
timestamp 1698431365
transform -1 0 22512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2566__A1
timestamp 1698431365
transform 1 0 23520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2567__A1
timestamp 1698431365
transform -1 0 20384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2568__S
timestamp 1698431365
transform -1 0 23744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__A1
timestamp 1698431365
transform -1 0 21168 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__B
timestamp 1698431365
transform -1 0 21840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__A1
timestamp 1698431365
transform -1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__B
timestamp 1698431365
transform -1 0 19600 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__A1
timestamp 1698431365
transform 1 0 19264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__I
timestamp 1698431365
transform 1 0 18704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__A1
timestamp 1698431365
transform -1 0 20048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__A2
timestamp 1698431365
transform -1 0 19152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__A2
timestamp 1698431365
transform 1 0 18368 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__A1
timestamp 1698431365
transform -1 0 17920 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__I0
timestamp 1698431365
transform 1 0 17472 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__A2
timestamp 1698431365
transform 1 0 16016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__A2
timestamp 1698431365
transform -1 0 14448 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2619__I
timestamp 1698431365
transform 1 0 14224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__A2
timestamp 1698431365
transform -1 0 11200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2622__A2
timestamp 1698431365
transform 1 0 13216 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2623__I
timestamp 1698431365
transform 1 0 10976 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__A1
timestamp 1698431365
transform 1 0 12096 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__I
timestamp 1698431365
transform -1 0 12656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__A1
timestamp 1698431365
transform -1 0 7280 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__A1
timestamp 1698431365
transform 1 0 7616 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__A1
timestamp 1698431365
transform -1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2642__A1
timestamp 1698431365
transform -1 0 5936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__I
timestamp 1698431365
transform 1 0 3808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__A1
timestamp 1698431365
transform 1 0 10640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__I
timestamp 1698431365
transform -1 0 7728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2656__I
timestamp 1698431365
transform 1 0 3808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__I
timestamp 1698431365
transform -1 0 7056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2674__I
timestamp 1698431365
transform 1 0 2688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2688__I
timestamp 1698431365
transform 1 0 13104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__I
timestamp 1698431365
transform 1 0 6944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__I
timestamp 1698431365
transform -1 0 3584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__A2
timestamp 1698431365
transform -1 0 8512 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__A1
timestamp 1698431365
transform 1 0 10528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__S
timestamp 1698431365
transform 1 0 7504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2709__I
timestamp 1698431365
transform 1 0 3584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__I
timestamp 1698431365
transform -1 0 4032 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2742__I
timestamp 1698431365
transform -1 0 5936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2756__I
timestamp 1698431365
transform -1 0 7392 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2765__A2
timestamp 1698431365
transform -1 0 10080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2766__A1
timestamp 1698431365
transform -1 0 9856 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2767__S
timestamp 1698431365
transform -1 0 8512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2783__I
timestamp 1698431365
transform 1 0 16800 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2806__A1
timestamp 1698431365
transform -1 0 16576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2808__A2
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2809__I
timestamp 1698431365
transform 1 0 19824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2841__A1
timestamp 1698431365
transform 1 0 18928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2844__A2
timestamp 1698431365
transform 1 0 18704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2845__A1
timestamp 1698431365
transform -1 0 19376 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2846__S
timestamp 1698431365
transform 1 0 17472 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2848__CLK
timestamp 1698431365
transform 1 0 11088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2849__CLK
timestamp 1698431365
transform 1 0 8400 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2850__CLK
timestamp 1698431365
transform 1 0 10976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2851__CLK
timestamp 1698431365
transform -1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2852__CLK
timestamp 1698431365
transform 1 0 33712 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2853__CLK
timestamp 1698431365
transform 1 0 32480 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2854__CLK
timestamp 1698431365
transform -1 0 31024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2855__CLK
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2856__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2857__CLK
timestamp 1698431365
transform 1 0 31360 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2858__CLK
timestamp 1698431365
transform 1 0 37968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2859__CLK
timestamp 1698431365
transform 1 0 38080 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2860__CLK
timestamp 1698431365
transform 1 0 38192 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2861__CLK
timestamp 1698431365
transform 1 0 34720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2862__CLK
timestamp 1698431365
transform 1 0 36288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2863__CLK
timestamp 1698431365
transform 1 0 45920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2864__CLK
timestamp 1698431365
transform 1 0 44912 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2865__CLK
timestamp 1698431365
transform 1 0 46480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2866__CLK
timestamp 1698431365
transform 1 0 48832 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2867__CLK
timestamp 1698431365
transform 1 0 51184 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2868__CLK
timestamp 1698431365
transform 1 0 51632 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2869__CLK
timestamp 1698431365
transform 1 0 52752 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2870__CLK
timestamp 1698431365
transform 1 0 48944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2871__CLK
timestamp 1698431365
transform 1 0 54096 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2872__CLK
timestamp 1698431365
transform 1 0 52080 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2873__CLK
timestamp 1698431365
transform 1 0 50400 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2874__CLK
timestamp 1698431365
transform 1 0 56000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2875__CLK
timestamp 1698431365
transform -1 0 45136 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2876__CLK
timestamp 1698431365
transform 1 0 38864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2877__CLK
timestamp 1698431365
transform 1 0 28784 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2878__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2879__CLK
timestamp 1698431365
transform 1 0 27888 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2880__CLK
timestamp 1698431365
transform 1 0 29456 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2881__CLK
timestamp 1698431365
transform 1 0 21392 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2882__CLK
timestamp 1698431365
transform 1 0 36400 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2884__CLK
timestamp 1698431365
transform 1 0 23296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2885__CLK
timestamp 1698431365
transform 1 0 22400 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2886__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2887__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2888__CLK
timestamp 1698431365
transform 1 0 24416 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2889__CLK
timestamp 1698431365
transform 1 0 21840 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2890__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2891__CLK
timestamp 1698431365
transform 1 0 26992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2892__CLK
timestamp 1698431365
transform 1 0 36400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2893__CLK
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2894__CLK
timestamp 1698431365
transform 1 0 42784 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2895__CLK
timestamp 1698431365
transform 1 0 46032 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2896__CLK
timestamp 1698431365
transform -1 0 49392 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2897__CLK
timestamp 1698431365
transform 1 0 48496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2898__CLK
timestamp 1698431365
transform 1 0 50064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2899__CLK
timestamp 1698431365
transform 1 0 49728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2900__CLK
timestamp 1698431365
transform 1 0 51968 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2901__CLK
timestamp 1698431365
transform 1 0 53648 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2902__CLK
timestamp 1698431365
transform 1 0 54880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2903__CLK
timestamp 1698431365
transform -1 0 54880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2904__CLK
timestamp 1698431365
transform 1 0 54880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2905__CLK
timestamp 1698431365
transform 1 0 54880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2906__CLK
timestamp 1698431365
transform 1 0 54880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2907__CLK
timestamp 1698431365
transform 1 0 53200 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2908__CLK
timestamp 1698431365
transform 1 0 45024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2909__CLK
timestamp 1698431365
transform -1 0 34832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2910__CLK
timestamp 1698431365
transform 1 0 32928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2911__CLK
timestamp 1698431365
transform 1 0 24080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2912__CLK
timestamp 1698431365
transform 1 0 17024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2913__CLK
timestamp 1698431365
transform 1 0 14672 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2914__CLK
timestamp 1698431365
transform 1 0 12208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2915__CLK
timestamp 1698431365
transform 1 0 20720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2922__CLK
timestamp 1698431365
transform -1 0 33824 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2923__CLK
timestamp 1698431365
transform 1 0 31808 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2924__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2925__CLK
timestamp 1698431365
transform 1 0 34608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2926__CLK
timestamp 1698431365
transform -1 0 35392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2927__CLK
timestamp 1698431365
transform 1 0 41440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2928__CLK
timestamp 1698431365
transform 1 0 38752 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2929__CLK
timestamp 1698431365
transform 1 0 44912 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2930__CLK
timestamp 1698431365
transform 1 0 44912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2931__CLK
timestamp 1698431365
transform 1 0 49168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2932__CLK
timestamp 1698431365
transform 1 0 50176 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2933__CLK
timestamp 1698431365
transform -1 0 47152 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2934__CLK
timestamp 1698431365
transform 1 0 51744 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2935__CLK
timestamp 1698431365
transform 1 0 52752 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2936__CLK
timestamp 1698431365
transform 1 0 53088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2937__CLK
timestamp 1698431365
transform 1 0 50848 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2938__CLK
timestamp 1698431365
transform 1 0 53872 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2939__CLK
timestamp 1698431365
transform -1 0 36288 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2940__CLK
timestamp 1698431365
transform 1 0 36512 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2941__CLK
timestamp 1698431365
transform 1 0 27104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2945__CLK
timestamp 1698431365
transform 1 0 12880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2946__CLK
timestamp 1698431365
transform 1 0 14112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2956__CLK
timestamp 1698431365
transform 1 0 30128 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2957__CLK
timestamp 1698431365
transform 1 0 30912 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2958__CLK
timestamp 1698431365
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2959__CLK
timestamp 1698431365
transform 1 0 35056 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2960__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2961__CLK
timestamp 1698431365
transform 1 0 44912 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2962__CLK
timestamp 1698431365
transform 1 0 45136 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2963__CLK
timestamp 1698431365
transform 1 0 48832 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2964__CLK
timestamp 1698431365
transform 1 0 49840 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2965__CLK
timestamp 1698431365
transform 1 0 48944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2966__CLK
timestamp 1698431365
transform 1 0 52080 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2967__CLK
timestamp 1698431365
transform 1 0 53536 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2968__CLK
timestamp 1698431365
transform 1 0 50848 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2969__CLK
timestamp 1698431365
transform 1 0 53200 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2970__CLK
timestamp 1698431365
transform 1 0 35168 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2971__CLK
timestamp 1698431365
transform 1 0 38640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2972__CLK
timestamp 1698431365
transform 1 0 29120 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2978__CLK
timestamp 1698431365
transform 1 0 12880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2979__CLK
timestamp 1698431365
transform 1 0 11088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2980__CLK
timestamp 1698431365
transform 1 0 24080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2981__CLK
timestamp 1698431365
transform 1 0 22400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2982__CLK
timestamp 1698431365
transform 1 0 34384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2983__CLK
timestamp 1698431365
transform 1 0 23408 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2984__CLK
timestamp 1698431365
transform -1 0 23968 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2985__CLK
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2986__CLK
timestamp 1698431365
transform 1 0 24864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2987__CLK
timestamp 1698431365
transform 1 0 33040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2988__CLK
timestamp 1698431365
transform -1 0 35392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2989__CLK
timestamp 1698431365
transform 1 0 37744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2990__CLK
timestamp 1698431365
transform 1 0 41216 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2991__CLK
timestamp 1698431365
transform 1 0 46144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2992__CLK
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2993__CLK
timestamp 1698431365
transform 1 0 44016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2994__CLK
timestamp 1698431365
transform 1 0 46704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2995__CLK
timestamp 1698431365
transform 1 0 48832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2996__CLK
timestamp 1698431365
transform 1 0 48832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2997__CLK
timestamp 1698431365
transform 1 0 50400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2998__CLK
timestamp 1698431365
transform 1 0 48832 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2999__CLK
timestamp 1698431365
transform -1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3000__CLK
timestamp 1698431365
transform 1 0 51856 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3001__CLK
timestamp 1698431365
transform 1 0 47936 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3002__CLK
timestamp 1698431365
transform 1 0 50512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3003__CLK
timestamp 1698431365
transform 1 0 48832 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3004__CLK
timestamp 1698431365
transform -1 0 37744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3005__CLK
timestamp 1698431365
transform 1 0 44016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3006__CLK
timestamp 1698431365
transform -1 0 25536 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3007__CLK
timestamp 1698431365
transform -1 0 26432 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3008__CLK
timestamp 1698431365
transform 1 0 22960 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3009__CLK
timestamp 1698431365
transform 1 0 22176 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3010__CLK
timestamp 1698431365
transform 1 0 11872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3011__CLK
timestamp 1698431365
transform 1 0 17920 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3012__CLK
timestamp 1698431365
transform 1 0 10192 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3013__CLK
timestamp 1698431365
transform 1 0 11536 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3014__CLK
timestamp 1698431365
transform 1 0 14784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3015__CLK
timestamp 1698431365
transform 1 0 7616 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3016__CLK
timestamp 1698431365
transform 1 0 17920 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3017__CLK
timestamp 1698431365
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3018__CLK
timestamp 1698431365
transform 1 0 10864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3019__CLK
timestamp 1698431365
transform 1 0 7952 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3020__CLK
timestamp 1698431365
transform 1 0 4256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3021__CLK
timestamp 1698431365
transform -1 0 5712 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3022__CLK
timestamp 1698431365
transform 1 0 5040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3023__CLK
timestamp 1698431365
transform 1 0 5488 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3024__CLK
timestamp 1698431365
transform 1 0 4816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3025__CLK
timestamp 1698431365
transform 1 0 10080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3026__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3027__CLK
timestamp 1698431365
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3028__CLK
timestamp 1698431365
transform 1 0 5712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3029__CLK
timestamp 1698431365
transform 1 0 6048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3030__CLK
timestamp 1698431365
transform -1 0 5936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3031__CLK
timestamp 1698431365
transform 1 0 5488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3032__CLK
timestamp 1698431365
transform 1 0 4816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3033__CLK
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3034__CLK
timestamp 1698431365
transform 1 0 4592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3035__CLK
timestamp 1698431365
transform 1 0 8064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3036__CLK
timestamp 1698431365
transform 1 0 11200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3037__CLK
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3038__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3039__CLK
timestamp 1698431365
transform 1 0 16352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3040__CLK
timestamp 1698431365
transform 1 0 11424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3041__CLK
timestamp 1698431365
transform 1 0 11312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3042__CLK
timestamp 1698431365
transform 1 0 18928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3043__CLK
timestamp 1698431365
transform 1 0 20720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3044__CLK
timestamp 1698431365
transform 1 0 22512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3045__CLK
timestamp 1698431365
transform 1 0 22736 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3046__CLK
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3047__CLK
timestamp 1698431365
transform 1 0 18368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform -1 0 29568 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_clk_I
timestamp 1698431365
transform -1 0 9744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_clk_I
timestamp 1698431365
transform 1 0 11088 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_clk_I
timestamp 1698431365
transform -1 0 25200 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_clk_I
timestamp 1698431365
transform 1 0 24080 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_clk_I
timestamp 1698431365
transform 1 0 14224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_clk_I
timestamp 1698431365
transform 1 0 13552 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_clk_I
timestamp 1698431365
transform 1 0 25312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_clk_I
timestamp 1698431365
transform 1 0 24416 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_clk_I
timestamp 1698431365
transform 1 0 43120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_clk_I
timestamp 1698431365
transform 1 0 46144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_clk_I
timestamp 1698431365
transform 1 0 49392 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_clk_I
timestamp 1698431365
transform 1 0 45920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_clk_I
timestamp 1698431365
transform 1 0 35840 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_clk_I
timestamp 1698431365
transform 1 0 35504 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_clk_I
timestamp 1698431365
transform 1 0 50176 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_clk_I
timestamp 1698431365
transform -1 0 48832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 2464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 2464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 2912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 2464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 2464 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 2464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 2464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 2464 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 2464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 2464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 2912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 2464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 3136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 2464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 3136 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 2912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 2464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 29232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 38416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 37184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 37856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 39312 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 39760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 40432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 57232 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 57904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 54768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 58352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 33376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 57680 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 57232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 57680 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 57680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 57232 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 5040 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform 1 0 3360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 34944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform 1 0 7952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform 1 0 7280 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 34272 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform -1 0 32032 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform -1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform -1 0 29680 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform -1 0 31024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform -1 0 35840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform -1 0 36512 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform 1 0 6384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform 1 0 6160 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698431365
transform 1 0 6160 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698431365
transform 1 0 3136 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698431365
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698431365
transform 1 0 4592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698431365
transform 1 0 3808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1698431365
transform 1 0 5264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1698431365
transform 1 0 2464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1698431365
transform 1 0 5712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1698431365
transform 1 0 1792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1698431365
transform 1 0 5936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1698431365
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1698431365
transform 1 0 4144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1698431365
transform -1 0 2240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1698431365
transform 1 0 3136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1698431365
transform 1 0 3584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1698431365
transform -1 0 17696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1698431365
transform -1 0 18256 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1698431365
transform 1 0 5600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1698431365
transform 1 0 3136 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1698431365
transform 1 0 5264 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1698431365
transform 1 0 5712 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1698431365
transform 1 0 5936 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1698431365
transform 1 0 3136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1698431365
transform 1 0 5040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1698431365
transform 1 0 7728 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1698431365
transform 1 0 5712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1698431365
transform 1 0 2688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1698431365
transform 1 0 3136 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output85_I
timestamp 1698431365
transform 1 0 50400 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output101_I
timestamp 1698431365
transform 1 0 55216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output102_I
timestamp 1698431365
transform 1 0 34160 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output108_I
timestamp 1698431365
transform 1 0 46592 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output114_I
timestamp 1698431365
transform -1 0 55440 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30016 0 1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1698431365
transform 1 0 6832 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1698431365
transform 1 0 20944 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1698431365
transform 1 0 20496 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1698431365
transform 1 0 10192 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1698431365
transform 1 0 11424 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1698431365
transform 1 0 21952 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1698431365
transform -1 0 24192 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1698431365
transform 1 0 42448 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1698431365
transform 1 0 46368 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1698431365
transform 1 0 49616 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1698431365
transform 1 0 46816 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1698431365
transform 1 0 32704 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1698431365
transform 1 0 32368 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1698431365
transform 1 0 48832 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_104 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_120 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14784 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_128 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15680 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_132 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_157
timestamp 1698431365
transform 1 0 18928 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165
timestamp 1698431365
transform 1 0 19824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_188
timestamp 1698431365
transform 1 0 22400 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_196
timestamp 1698431365
transform 1 0 23296 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_200
timestamp 1698431365
transform 1 0 23744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_214
timestamp 1698431365
transform 1 0 25312 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_230
timestamp 1698431365
transform 1 0 27104 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_244
timestamp 1698431365
transform 1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_246
timestamp 1698431365
transform 1 0 28896 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_249
timestamp 1698431365
transform 1 0 29232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698431365
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_338
timestamp 1698431365
transform 1 0 39200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_354
timestamp 1698431365
transform 1 0 40992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_370
timestamp 1698431365
transform 1 0 42784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494
timestamp 1698431365
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502
timestamp 1698431365
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_146
timestamp 1698431365
transform 1 0 17696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_148
timestamp 1698431365
transform 1 0 17920 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_151
timestamp 1698431365
transform 1 0 18256 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183
timestamp 1698431365
transform 1 0 21840 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698431365
transform 1 0 23632 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698431365
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_244
timestamp 1698431365
transform 1 0 28672 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_260
timestamp 1698431365
transform 1 0 30464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_262
timestamp 1698431365
transform 1 0 30688 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_265
timestamp 1698431365
transform 1 0 31024 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_269
timestamp 1698431365
transform 1 0 31472 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_271
timestamp 1698431365
transform 1 0 31696 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_274
timestamp 1698431365
transform 1 0 32032 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_286
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_290
timestamp 1698431365
transform 1 0 33824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_294
timestamp 1698431365
transform 1 0 34272 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_300
timestamp 1698431365
transform 1 0 34944 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_304
timestamp 1698431365
transform 1 0 35392 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_308
timestamp 1698431365
transform 1 0 35840 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_314
timestamp 1698431365
transform 1 0 36512 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_320
timestamp 1698431365
transform 1 0 37184 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_326
timestamp 1698431365
transform 1 0 37856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_328
timestamp 1698431365
transform 1 0 38080 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_337
timestamp 1698431365
transform 1 0 39088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_341
timestamp 1698431365
transform 1 0 39536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_345
timestamp 1698431365
transform 1 0 39984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698431365
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_508
timestamp 1698431365
transform 1 0 58240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698431365
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698431365
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_88
timestamp 1698431365
transform 1 0 11200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_121
timestamp 1698431365
transform 1 0 14896 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_137
timestamp 1698431365
transform 1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_279
timestamp 1698431365
transform 1 0 32592 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_295
timestamp 1698431365
transform 1 0 34384 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_300
timestamp 1698431365
transform 1 0 34944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_304
timestamp 1698431365
transform 1 0 35392 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_312
timestamp 1698431365
transform 1 0 36288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_314
timestamp 1698431365
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_489
timestamp 1698431365
transform 1 0 56112 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698431365
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_34
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_50
timestamp 1698431365
transform 1 0 6944 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_58
timestamp 1698431365
transform 1 0 7840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_62
timestamp 1698431365
transform 1 0 8288 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_132
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_228
timestamp 1698431365
transform 1 0 26880 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_260
timestamp 1698431365
transform 1 0 30464 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_311
timestamp 1698431365
transform 1 0 36176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_344
timestamp 1698431365
transform 1 0 39872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_348
timestamp 1698431365
transform 1 0 40320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_362
timestamp 1698431365
transform 1 0 41888 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_372
timestamp 1698431365
transform 1 0 43008 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_404
timestamp 1698431365
transform 1 0 46592 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_39
timestamp 1698431365
transform 1 0 5712 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_46
timestamp 1698431365
transform 1 0 6496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_50
timestamp 1698431365
transform 1 0 6944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_86
timestamp 1698431365
transform 1 0 10976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_90
timestamp 1698431365
transform 1 0 11424 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_102
timestamp 1698431365
transform 1 0 12768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_120
timestamp 1698431365
transform 1 0 14784 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_124
timestamp 1698431365
transform 1 0 15232 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_155
timestamp 1698431365
transform 1 0 18704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_159
timestamp 1698431365
transform 1 0 19152 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_209
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_217
timestamp 1698431365
transform 1 0 25648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_219
timestamp 1698431365
transform 1 0 25872 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_224
timestamp 1698431365
transform 1 0 26432 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_240
timestamp 1698431365
transform 1 0 28224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_263
timestamp 1698431365
transform 1 0 30800 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_296
timestamp 1698431365
transform 1 0 34496 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_327
timestamp 1698431365
transform 1 0 37968 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_338
timestamp 1698431365
transform 1 0 39200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_340
timestamp 1698431365
transform 1 0 39424 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_374
timestamp 1698431365
transform 1 0 43232 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_379
timestamp 1698431365
transform 1 0 43792 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_383
timestamp 1698431365
transform 1 0 44240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_489
timestamp 1698431365
transform 1 0 56112 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_505
timestamp 1698431365
transform 1 0 57904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_8
timestamp 1698431365
transform 1 0 2240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_12
timestamp 1698431365
transform 1 0 2688 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_20
timestamp 1698431365
transform 1 0 3584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_24
timestamp 1698431365
transform 1 0 4032 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_28
timestamp 1698431365
transform 1 0 4480 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_60
timestamp 1698431365
transform 1 0 8064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_64
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_68
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_86
timestamp 1698431365
transform 1 0 10976 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_94
timestamp 1698431365
transform 1 0 11872 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_103
timestamp 1698431365
transform 1 0 12880 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_119
timestamp 1698431365
transform 1 0 14672 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_127
timestamp 1698431365
transform 1 0 15568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_134
timestamp 1698431365
transform 1 0 16352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_138
timestamp 1698431365
transform 1 0 16800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_171
timestamp 1698431365
transform 1 0 20496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_175
timestamp 1698431365
transform 1 0 20944 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_183
timestamp 1698431365
transform 1 0 21840 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_195
timestamp 1698431365
transform 1 0 23184 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_205
timestamp 1698431365
transform 1 0 24304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_207
timestamp 1698431365
transform 1 0 24528 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_245
timestamp 1698431365
transform 1 0 28784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_266
timestamp 1698431365
transform 1 0 31136 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_274
timestamp 1698431365
transform 1 0 32032 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_278
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_286
timestamp 1698431365
transform 1 0 33376 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_313
timestamp 1698431365
transform 1 0 36400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_317
timestamp 1698431365
transform 1 0 36848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_319
timestamp 1698431365
transform 1 0 37072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_349
timestamp 1698431365
transform 1 0 40432 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_364
timestamp 1698431365
transform 1 0 42112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_397
timestamp 1698431365
transform 1 0 45808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_401
timestamp 1698431365
transform 1 0 46256 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_417
timestamp 1698431365
transform 1 0 48048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_419
timestamp 1698431365
transform 1 0 48272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_33
timestamp 1698431365
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_61
timestamp 1698431365
transform 1 0 8176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_96
timestamp 1698431365
transform 1 0 12096 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_119
timestamp 1698431365
transform 1 0 14672 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_127
timestamp 1698431365
transform 1 0 15568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_131
timestamp 1698431365
transform 1 0 16016 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_148
timestamp 1698431365
transform 1 0 17920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_150
timestamp 1698431365
transform 1 0 18144 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_156
timestamp 1698431365
transform 1 0 18816 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_163
timestamp 1698431365
transform 1 0 19600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_167
timestamp 1698431365
transform 1 0 20048 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_181
timestamp 1698431365
transform 1 0 21616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_214
timestamp 1698431365
transform 1 0 25312 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_222
timestamp 1698431365
transform 1 0 26208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_242
timestamp 1698431365
transform 1 0 28448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_251
timestamp 1698431365
transform 1 0 29456 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_281
timestamp 1698431365
transform 1 0 32816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_285
timestamp 1698431365
transform 1 0 33264 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_289
timestamp 1698431365
transform 1 0 33712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_291
timestamp 1698431365
transform 1 0 33936 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_294
timestamp 1698431365
transform 1 0 34272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_310
timestamp 1698431365
transform 1 0 36064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_312
timestamp 1698431365
transform 1 0 36288 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_326
timestamp 1698431365
transform 1 0 37856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_330
timestamp 1698431365
transform 1 0 38304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_332
timestamp 1698431365
transform 1 0 38528 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_335
timestamp 1698431365
transform 1 0 38864 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_382
timestamp 1698431365
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_393
timestamp 1698431365
transform 1 0 45360 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_425
timestamp 1698431365
transform 1 0 48944 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_441
timestamp 1698431365
transform 1 0 50736 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_449
timestamp 1698431365
transform 1 0 51632 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_453
timestamp 1698431365
transform 1 0 52080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_489
timestamp 1698431365
transform 1 0 56112 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_505
timestamp 1698431365
transform 1 0 57904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_20
timestamp 1698431365
transform 1 0 3584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_24
timestamp 1698431365
transform 1 0 4032 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_50
timestamp 1698431365
transform 1 0 6944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_54
timestamp 1698431365
transform 1 0 7392 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_109
timestamp 1698431365
transform 1 0 13552 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_128
timestamp 1698431365
transform 1 0 15680 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_155
timestamp 1698431365
transform 1 0 18704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_157
timestamp 1698431365
transform 1 0 18928 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_187
timestamp 1698431365
transform 1 0 22288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_191
timestamp 1698431365
transform 1 0 22736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_195
timestamp 1698431365
transform 1 0 23184 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_200
timestamp 1698431365
transform 1 0 23744 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_208
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_224
timestamp 1698431365
transform 1 0 26432 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_228
timestamp 1698431365
transform 1 0 26880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_236
timestamp 1698431365
transform 1 0 27776 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_252
timestamp 1698431365
transform 1 0 29568 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_260
timestamp 1698431365
transform 1 0 30464 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_264
timestamp 1698431365
transform 1 0 30912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_268
timestamp 1698431365
transform 1 0 31360 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_286
timestamp 1698431365
transform 1 0 33376 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_292
timestamp 1698431365
transform 1 0 34048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_294
timestamp 1698431365
transform 1 0 34272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_301
timestamp 1698431365
transform 1 0 35056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_303
timestamp 1698431365
transform 1 0 35280 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_314
timestamp 1698431365
transform 1 0 36512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_316
timestamp 1698431365
transform 1 0 36736 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_322
timestamp 1698431365
transform 1 0 37408 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_334
timestamp 1698431365
transform 1 0 38752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_345
timestamp 1698431365
transform 1 0 39984 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_360
timestamp 1698431365
transform 1 0 41664 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_364
timestamp 1698431365
transform 1 0 42112 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_379
timestamp 1698431365
transform 1 0 43792 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_398
timestamp 1698431365
transform 1 0 45920 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_414
timestamp 1698431365
transform 1 0 47712 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_418
timestamp 1698431365
transform 1 0 48160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_31
timestamp 1698431365
transform 1 0 4816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_61
timestamp 1698431365
transform 1 0 8176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_65
timestamp 1698431365
transform 1 0 8624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_67
timestamp 1698431365
transform 1 0 8848 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_74
timestamp 1698431365
transform 1 0 9632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_78
timestamp 1698431365
transform 1 0 10080 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_86
timestamp 1698431365
transform 1 0 10976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_132
timestamp 1698431365
transform 1 0 16128 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_136
timestamp 1698431365
transform 1 0 16576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_209
timestamp 1698431365
transform 1 0 24752 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_239
timestamp 1698431365
transform 1 0 28112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_253
timestamp 1698431365
transform 1 0 29680 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_290
timestamp 1698431365
transform 1 0 33824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_312
timestamp 1698431365
transform 1 0 36288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_314
timestamp 1698431365
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_380
timestamp 1698431365
transform 1 0 43904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_391
timestamp 1698431365
transform 1 0 45136 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_395
timestamp 1698431365
transform 1 0 45584 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_425
timestamp 1698431365
transform 1 0 48944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_429
timestamp 1698431365
transform 1 0 49392 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_445
timestamp 1698431365
transform 1 0 51184 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_453
timestamp 1698431365
transform 1 0 52080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_489
timestamp 1698431365
transform 1 0 56112 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_505
timestamp 1698431365
transform 1 0 57904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_8
timestamp 1698431365
transform 1 0 2240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_23
timestamp 1698431365
transform 1 0 3920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_33
timestamp 1698431365
transform 1 0 5040 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_37
timestamp 1698431365
transform 1 0 5488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_53
timestamp 1698431365
transform 1 0 7280 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_61
timestamp 1698431365
transform 1 0 8176 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_82
timestamp 1698431365
transform 1 0 10528 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_90
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_122
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_124
timestamp 1698431365
transform 1 0 15232 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_131
timestamp 1698431365
transform 1 0 16016 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_156
timestamp 1698431365
transform 1 0 18816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_176
timestamp 1698431365
transform 1 0 21056 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_180
timestamp 1698431365
transform 1 0 21504 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_224
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_255
timestamp 1698431365
transform 1 0 29904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_265
timestamp 1698431365
transform 1 0 31024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_267
timestamp 1698431365
transform 1 0 31248 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_287
timestamp 1698431365
transform 1 0 33488 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_304
timestamp 1698431365
transform 1 0 35392 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_308
timestamp 1698431365
transform 1 0 35840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_322
timestamp 1698431365
transform 1 0 37408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_341
timestamp 1698431365
transform 1 0 39536 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_345
timestamp 1698431365
transform 1 0 39984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_347
timestamp 1698431365
transform 1 0 40208 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_356
timestamp 1698431365
transform 1 0 41216 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_360
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_362
timestamp 1698431365
transform 1 0 41888 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_398
timestamp 1698431365
transform 1 0 45920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_402
timestamp 1698431365
transform 1 0 46368 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_418
timestamp 1698431365
transform 1 0 48160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_14
timestamp 1698431365
transform 1 0 2912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_29
timestamp 1698431365
transform 1 0 4592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_33
timestamp 1698431365
transform 1 0 5040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_65
timestamp 1698431365
transform 1 0 8624 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_81
timestamp 1698431365
transform 1 0 10416 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_88
timestamp 1698431365
transform 1 0 11200 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_113
timestamp 1698431365
transform 1 0 14000 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_129
timestamp 1698431365
transform 1 0 15792 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_137
timestamp 1698431365
transform 1 0 16688 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_140
timestamp 1698431365
transform 1 0 17024 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_148
timestamp 1698431365
transform 1 0 17920 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_152
timestamp 1698431365
transform 1 0 18368 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_154
timestamp 1698431365
transform 1 0 18592 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_193
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_197
timestamp 1698431365
transform 1 0 23408 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_199
timestamp 1698431365
transform 1 0 23632 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_216
timestamp 1698431365
transform 1 0 25536 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_257
timestamp 1698431365
transform 1 0 30128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_261
timestamp 1698431365
transform 1 0 30576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_263
timestamp 1698431365
transform 1 0 30800 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_277
timestamp 1698431365
transform 1 0 32368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_281
timestamp 1698431365
transform 1 0 32816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_291
timestamp 1698431365
transform 1 0 33936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_293
timestamp 1698431365
transform 1 0 34160 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_296
timestamp 1698431365
transform 1 0 34496 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_312
timestamp 1698431365
transform 1 0 36288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_321
timestamp 1698431365
transform 1 0 37296 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_324
timestamp 1698431365
transform 1 0 37632 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_328
timestamp 1698431365
transform 1 0 38080 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_330
timestamp 1698431365
transform 1 0 38304 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_337
timestamp 1698431365
transform 1 0 39088 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_345
timestamp 1698431365
transform 1 0 39984 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_349
timestamp 1698431365
transform 1 0 40432 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_352
timestamp 1698431365
transform 1 0 40768 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_358
timestamp 1698431365
transform 1 0 41440 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_360
timestamp 1698431365
transform 1 0 41664 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_376
timestamp 1698431365
transform 1 0 43456 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_378
timestamp 1698431365
transform 1 0 43680 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_403
timestamp 1698431365
transform 1 0 46480 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_405
timestamp 1698431365
transform 1 0 46704 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_410
timestamp 1698431365
transform 1 0 47264 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_442
timestamp 1698431365
transform 1 0 50848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_450
timestamp 1698431365
transform 1 0 51744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_454
timestamp 1698431365
transform 1 0 52192 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_489
timestamp 1698431365
transform 1 0 56112 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_505
timestamp 1698431365
transform 1 0 57904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_39
timestamp 1698431365
transform 1 0 5712 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_84
timestamp 1698431365
transform 1 0 10752 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_100
timestamp 1698431365
transform 1 0 12544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_119
timestamp 1698431365
transform 1 0 14672 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_135
timestamp 1698431365
transform 1 0 16464 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_156
timestamp 1698431365
transform 1 0 18816 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_189
timestamp 1698431365
transform 1 0 22512 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_193
timestamp 1698431365
transform 1 0 22960 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_201
timestamp 1698431365
transform 1 0 23856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_205
timestamp 1698431365
transform 1 0 24304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_207
timestamp 1698431365
transform 1 0 24528 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_244
timestamp 1698431365
transform 1 0 28672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_248
timestamp 1698431365
transform 1 0 29120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_252
timestamp 1698431365
transform 1 0 29568 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_260
timestamp 1698431365
transform 1 0 30464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_262
timestamp 1698431365
transform 1 0 30688 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_273
timestamp 1698431365
transform 1 0 31920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698431365
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_289
timestamp 1698431365
transform 1 0 33712 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_301
timestamp 1698431365
transform 1 0 35056 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_305
timestamp 1698431365
transform 1 0 35504 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_318
timestamp 1698431365
transform 1 0 36960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_337
timestamp 1698431365
transform 1 0 39088 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_343
timestamp 1698431365
transform 1 0 39760 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_347
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_390
timestamp 1698431365
transform 1 0 45024 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_394
timestamp 1698431365
transform 1 0 45472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_396
timestamp 1698431365
transform 1 0 45696 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_414
timestamp 1698431365
transform 1 0 47712 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_418
timestamp 1698431365
transform 1 0 48160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_444
timestamp 1698431365
transform 1 0 51072 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_476
timestamp 1698431365
transform 1 0 54656 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_484
timestamp 1698431365
transform 1 0 55552 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_488
timestamp 1698431365
transform 1 0 56000 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_14
timestamp 1698431365
transform 1 0 2912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_27
timestamp 1698431365
transform 1 0 4368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_31
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_39
timestamp 1698431365
transform 1 0 5712 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_64
timestamp 1698431365
transform 1 0 8512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_82
timestamp 1698431365
transform 1 0 10528 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_84
timestamp 1698431365
transform 1 0 10752 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_102
timestamp 1698431365
transform 1 0 12768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_125
timestamp 1698431365
transform 1 0 15344 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_129
timestamp 1698431365
transform 1 0 15792 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_166
timestamp 1698431365
transform 1 0 19936 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_183
timestamp 1698431365
transform 1 0 21840 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_216
timestamp 1698431365
transform 1 0 25536 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_231
timestamp 1698431365
transform 1 0 27216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_233
timestamp 1698431365
transform 1 0 27440 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_240
timestamp 1698431365
transform 1 0 28224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_259
timestamp 1698431365
transform 1 0 30352 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_273
timestamp 1698431365
transform 1 0 31920 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_277
timestamp 1698431365
transform 1 0 32368 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_292
timestamp 1698431365
transform 1 0 34048 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_397
timestamp 1698431365
transform 1 0 45808 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_401
timestamp 1698431365
transform 1 0 46256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_411
timestamp 1698431365
transform 1 0 47376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_419
timestamp 1698431365
transform 1 0 48272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_452
timestamp 1698431365
transform 1 0 51968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_454
timestamp 1698431365
transform 1 0 52192 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_489
timestamp 1698431365
transform 1 0 56112 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_505
timestamp 1698431365
transform 1 0 57904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_35
timestamp 1698431365
transform 1 0 5264 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_39
timestamp 1698431365
transform 1 0 5712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_43
timestamp 1698431365
transform 1 0 6160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_45
timestamp 1698431365
transform 1 0 6384 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_63
timestamp 1698431365
transform 1 0 8400 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_98
timestamp 1698431365
transform 1 0 12320 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_128
timestamp 1698431365
transform 1 0 15680 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_155
timestamp 1698431365
transform 1 0 18704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_165
timestamp 1698431365
transform 1 0 19824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_204
timestamp 1698431365
transform 1 0 24192 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_220
timestamp 1698431365
transform 1 0 25984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_222
timestamp 1698431365
transform 1 0 26208 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_250
timestamp 1698431365
transform 1 0 29344 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_258
timestamp 1698431365
transform 1 0 30240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_306
timestamp 1698431365
transform 1 0 35616 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_324
timestamp 1698431365
transform 1 0 37632 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_341
timestamp 1698431365
transform 1 0 39536 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_358
timestamp 1698431365
transform 1 0 41440 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_400
timestamp 1698431365
transform 1 0 46144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_419
timestamp 1698431365
transform 1 0 48272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_426
timestamp 1698431365
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_466
timestamp 1698431365
transform 1 0 53536 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_482
timestamp 1698431365
transform 1 0 55328 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1698431365
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_31
timestamp 1698431365
transform 1 0 4816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_71
timestamp 1698431365
transform 1 0 9296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_75
timestamp 1698431365
transform 1 0 9744 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_132
timestamp 1698431365
transform 1 0 16128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_151
timestamp 1698431365
transform 1 0 18256 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_167
timestamp 1698431365
transform 1 0 20048 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_209
timestamp 1698431365
transform 1 0 24752 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_213
timestamp 1698431365
transform 1 0 25200 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_215
timestamp 1698431365
transform 1 0 25424 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_239
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_263
timestamp 1698431365
transform 1 0 30800 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_286
timestamp 1698431365
transform 1 0 33376 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_296
timestamp 1698431365
transform 1 0 34496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_300
timestamp 1698431365
transform 1 0 34944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_327
timestamp 1698431365
transform 1 0 37968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_331
timestamp 1698431365
transform 1 0 38416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_364
timestamp 1698431365
transform 1 0 42112 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_383
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_389
timestamp 1698431365
transform 1 0 44912 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_397
timestamp 1698431365
transform 1 0 45808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_433
timestamp 1698431365
transform 1 0 49840 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_437
timestamp 1698431365
transform 1 0 50288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_467
timestamp 1698431365
transform 1 0 53648 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_499
timestamp 1698431365
transform 1 0 57232 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_507
timestamp 1698431365
transform 1 0 58128 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_14
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_41
timestamp 1698431365
transform 1 0 5936 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_43
timestamp 1698431365
transform 1 0 6160 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_74
timestamp 1698431365
transform 1 0 9632 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_81
timestamp 1698431365
transform 1 0 10416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_85
timestamp 1698431365
transform 1 0 10864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_87
timestamp 1698431365
transform 1 0 11088 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_94
timestamp 1698431365
transform 1 0 11872 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_102
timestamp 1698431365
transform 1 0 12768 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_108
timestamp 1698431365
transform 1 0 13440 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_124
timestamp 1698431365
transform 1 0 15232 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_128
timestamp 1698431365
transform 1 0 15680 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_130
timestamp 1698431365
transform 1 0 15904 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_150
timestamp 1698431365
transform 1 0 18144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_159
timestamp 1698431365
transform 1 0 19152 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_201
timestamp 1698431365
transform 1 0 23856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_203
timestamp 1698431365
transform 1 0 24080 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_220
timestamp 1698431365
transform 1 0 25984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_224
timestamp 1698431365
transform 1 0 26432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_233
timestamp 1698431365
transform 1 0 27440 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_237
timestamp 1698431365
transform 1 0 27888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_256
timestamp 1698431365
transform 1 0 30016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_260
timestamp 1698431365
transform 1 0 30464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_266
timestamp 1698431365
transform 1 0 31136 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_274
timestamp 1698431365
transform 1 0 32032 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698431365
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_290
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_323
timestamp 1698431365
transform 1 0 37520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_327
timestamp 1698431365
transform 1 0 37968 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_335
timestamp 1698431365
transform 1 0 38864 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_339
timestamp 1698431365
transform 1 0 39312 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_342
timestamp 1698431365
transform 1 0 39648 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_379
timestamp 1698431365
transform 1 0 43792 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_383
timestamp 1698431365
transform 1 0 44240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_402
timestamp 1698431365
transform 1 0 46368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_404
timestamp 1698431365
transform 1 0 46592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_417
timestamp 1698431365
transform 1 0 48048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_463
timestamp 1698431365
transform 1 0 53200 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_479
timestamp 1698431365
transform 1 0 54992 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_487
timestamp 1698431365
transform 1 0 55888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_489
timestamp 1698431365
transform 1 0 56112 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_508
timestamp 1698431365
transform 1 0 58240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_31
timestamp 1698431365
transform 1 0 4816 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_41
timestamp 1698431365
transform 1 0 5936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_45
timestamp 1698431365
transform 1 0 6384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_81
timestamp 1698431365
transform 1 0 10416 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_91
timestamp 1698431365
transform 1 0 11536 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_99
timestamp 1698431365
transform 1 0 12432 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_103
timestamp 1698431365
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_120
timestamp 1698431365
transform 1 0 14784 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_132
timestamp 1698431365
transform 1 0 16128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_206
timestamp 1698431365
transform 1 0 24416 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_236
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_269
timestamp 1698431365
transform 1 0 31472 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_292
timestamp 1698431365
transform 1 0 34048 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_296
timestamp 1698431365
transform 1 0 34496 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_303
timestamp 1698431365
transform 1 0 35280 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_319
timestamp 1698431365
transform 1 0 37072 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_330
timestamp 1698431365
transform 1 0 38304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_375
timestamp 1698431365
transform 1 0 43344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_379
timestamp 1698431365
transform 1 0 43792 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_383
timestamp 1698431365
transform 1 0 44240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_389
timestamp 1698431365
transform 1 0 44912 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_428
timestamp 1698431365
transform 1 0 49280 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_434
timestamp 1698431365
transform 1 0 49952 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_438
timestamp 1698431365
transform 1 0 50400 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_452
timestamp 1698431365
transform 1 0 51968 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_454
timestamp 1698431365
transform 1 0 52192 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_461
timestamp 1698431365
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_463
timestamp 1698431365
transform 1 0 53200 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_468
timestamp 1698431365
transform 1 0 53760 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_500
timestamp 1698431365
transform 1 0 57344 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_508
timestamp 1698431365
transform 1 0 58240 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_8
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_14
timestamp 1698431365
transform 1 0 2912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_18
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_30
timestamp 1698431365
transform 1 0 4704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_44
timestamp 1698431365
transform 1 0 6272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_82
timestamp 1698431365
transform 1 0 10528 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_86
timestamp 1698431365
transform 1 0 10976 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_88
timestamp 1698431365
transform 1 0 11200 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698431365
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_164
timestamp 1698431365
transform 1 0 19712 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_172
timestamp 1698431365
transform 1 0 20608 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_181
timestamp 1698431365
transform 1 0 21616 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_191
timestamp 1698431365
transform 1 0 22736 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_199
timestamp 1698431365
transform 1 0 23632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_202
timestamp 1698431365
transform 1 0 23968 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_206
timestamp 1698431365
transform 1 0 24416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_231
timestamp 1698431365
transform 1 0 27216 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_235
timestamp 1698431365
transform 1 0 27664 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_237
timestamp 1698431365
transform 1 0 27888 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_259
timestamp 1698431365
transform 1 0 30352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_263
timestamp 1698431365
transform 1 0 30800 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698431365
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_290
timestamp 1698431365
transform 1 0 33824 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_306
timestamp 1698431365
transform 1 0 35616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_310
timestamp 1698431365
transform 1 0 36064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_333
timestamp 1698431365
transform 1 0 38640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_337
timestamp 1698431365
transform 1 0 39088 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_360
timestamp 1698431365
transform 1 0 41664 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_369
timestamp 1698431365
transform 1 0 42672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_373
timestamp 1698431365
transform 1 0 43120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_377
timestamp 1698431365
transform 1 0 43568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_379
timestamp 1698431365
transform 1 0 43792 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_385
timestamp 1698431365
transform 1 0 44464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_389
timestamp 1698431365
transform 1 0 44912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_426
timestamp 1698431365
transform 1 0 49056 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_442
timestamp 1698431365
transform 1 0 50848 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_450
timestamp 1698431365
transform 1 0 51744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_483
timestamp 1698431365
transform 1 0 55440 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_487
timestamp 1698431365
transform 1 0 55888 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_489
timestamp 1698431365
transform 1 0 56112 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_14
timestamp 1698431365
transform 1 0 2912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_85
timestamp 1698431365
transform 1 0 10864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_89
timestamp 1698431365
transform 1 0 11312 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_97
timestamp 1698431365
transform 1 0 12208 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_120
timestamp 1698431365
transform 1 0 14784 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_135
timestamp 1698431365
transform 1 0 16464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_139
timestamp 1698431365
transform 1 0 16912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_155
timestamp 1698431365
transform 1 0 18704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_159
timestamp 1698431365
transform 1 0 19152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_208
timestamp 1698431365
transform 1 0 24640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_210
timestamp 1698431365
transform 1 0 24864 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_225
timestamp 1698431365
transform 1 0 26544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_229
timestamp 1698431365
transform 1 0 26992 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_233
timestamp 1698431365
transform 1 0 27440 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_261
timestamp 1698431365
transform 1 0 30576 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_265
timestamp 1698431365
transform 1 0 31024 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_289
timestamp 1698431365
transform 1 0 33712 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_297
timestamp 1698431365
transform 1 0 34608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_313
timestamp 1698431365
transform 1 0 36400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_321
timestamp 1698431365
transform 1 0 37296 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_330
timestamp 1698431365
transform 1 0 38304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_334
timestamp 1698431365
transform 1 0 38752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_336
timestamp 1698431365
transform 1 0 38976 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_339
timestamp 1698431365
transform 1 0 39312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_343
timestamp 1698431365
transform 1 0 39760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_347
timestamp 1698431365
transform 1 0 40208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_351
timestamp 1698431365
transform 1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_353
timestamp 1698431365
transform 1 0 40880 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_356
timestamp 1698431365
transform 1 0 41216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_360
timestamp 1698431365
transform 1 0 41664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_362
timestamp 1698431365
transform 1 0 41888 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_371
timestamp 1698431365
transform 1 0 42896 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_395
timestamp 1698431365
transform 1 0 45584 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_399
timestamp 1698431365
transform 1 0 46032 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_402
timestamp 1698431365
transform 1 0 46368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_406
timestamp 1698431365
transform 1 0 46816 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_436
timestamp 1698431365
transform 1 0 50176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_440
timestamp 1698431365
transform 1 0 50624 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_448
timestamp 1698431365
transform 1 0 51520 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_452
timestamp 1698431365
transform 1 0 51968 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_454
timestamp 1698431365
transform 1 0 52192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_461
timestamp 1698431365
transform 1 0 52976 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_477
timestamp 1698431365
transform 1 0 54768 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_36
timestamp 1698431365
transform 1 0 5376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_40
timestamp 1698431365
transform 1 0 5824 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_50
timestamp 1698431365
transform 1 0 6944 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_62
timestamp 1698431365
transform 1 0 8288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_64
timestamp 1698431365
transform 1 0 8512 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_97
timestamp 1698431365
transform 1 0 12208 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_104
timestamp 1698431365
transform 1 0 12992 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_111
timestamp 1698431365
transform 1 0 13776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_121
timestamp 1698431365
transform 1 0 14896 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698431365
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_146
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_154
timestamp 1698431365
transform 1 0 18592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_201
timestamp 1698431365
transform 1 0 23856 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_205
timestamp 1698431365
transform 1 0 24304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_228
timestamp 1698431365
transform 1 0 26880 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_303
timestamp 1698431365
transform 1 0 35280 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_305
timestamp 1698431365
transform 1 0 35504 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_318
timestamp 1698431365
transform 1 0 36960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_322
timestamp 1698431365
transform 1 0 37408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_326
timestamp 1698431365
transform 1 0 37856 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_345
timestamp 1698431365
transform 1 0 39984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_356
timestamp 1698431365
transform 1 0 41216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_360
timestamp 1698431365
transform 1 0 41664 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_362
timestamp 1698431365
transform 1 0 41888 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_408
timestamp 1698431365
transform 1 0 47040 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_417
timestamp 1698431365
transform 1 0 48048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_419
timestamp 1698431365
transform 1 0 48272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_426
timestamp 1698431365
transform 1 0 49056 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_434
timestamp 1698431365
transform 1 0 49952 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_459
timestamp 1698431365
transform 1 0 52752 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_467
timestamp 1698431365
transform 1 0 53648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_471
timestamp 1698431365
transform 1 0 54096 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_487
timestamp 1698431365
transform 1 0 55888 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_489
timestamp 1698431365
transform 1 0 56112 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_508
timestamp 1698431365
transform 1 0 58240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_16
timestamp 1698431365
transform 1 0 3136 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_33
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_45
timestamp 1698431365
transform 1 0 6384 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_49
timestamp 1698431365
transform 1 0 6832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_52
timestamp 1698431365
transform 1 0 7168 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_103
timestamp 1698431365
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_158
timestamp 1698431365
transform 1 0 19040 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698431365
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_181
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_191
timestamp 1698431365
transform 1 0 22736 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_195
timestamp 1698431365
transform 1 0 23184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_232
timestamp 1698431365
transform 1 0 27328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_234
timestamp 1698431365
transform 1 0 27552 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_261
timestamp 1698431365
transform 1 0 30576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_263
timestamp 1698431365
transform 1 0 30800 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_293
timestamp 1698431365
transform 1 0 34160 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_329
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_358
timestamp 1698431365
transform 1 0 41440 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_376
timestamp 1698431365
transform 1 0 43456 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_391
timestamp 1698431365
transform 1 0 45136 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_413
timestamp 1698431365
transform 1 0 47600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_417
timestamp 1698431365
transform 1 0 48048 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_433
timestamp 1698431365
transform 1 0 49840 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_465
timestamp 1698431365
transform 1 0 53424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_498
timestamp 1698431365
transform 1 0 57120 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_502
timestamp 1698431365
transform 1 0 57568 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_505
timestamp 1698431365
transform 1 0 57904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_16
timestamp 1698431365
transform 1 0 3136 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_33
timestamp 1698431365
transform 1 0 5040 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_37
timestamp 1698431365
transform 1 0 5488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_41
timestamp 1698431365
transform 1 0 5936 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_49
timestamp 1698431365
transform 1 0 6832 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_57
timestamp 1698431365
transform 1 0 7728 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_92
timestamp 1698431365
transform 1 0 11648 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_96
timestamp 1698431365
transform 1 0 12096 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_155
timestamp 1698431365
transform 1 0 18704 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_164
timestamp 1698431365
transform 1 0 19712 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_216
timestamp 1698431365
transform 1 0 25536 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_230
timestamp 1698431365
transform 1 0 27104 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_245
timestamp 1698431365
transform 1 0 28784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_247
timestamp 1698431365
transform 1 0 29008 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_258
timestamp 1698431365
transform 1 0 30240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_265
timestamp 1698431365
transform 1 0 31024 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_286
timestamp 1698431365
transform 1 0 33376 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_290
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_293
timestamp 1698431365
transform 1 0 34160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_297
timestamp 1698431365
transform 1 0 34608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_301
timestamp 1698431365
transform 1 0 35056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_305
timestamp 1698431365
transform 1 0 35504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_309
timestamp 1698431365
transform 1 0 35952 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_313
timestamp 1698431365
transform 1 0 36400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_317
timestamp 1698431365
transform 1 0 36848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_321
timestamp 1698431365
transform 1 0 37296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_325
timestamp 1698431365
transform 1 0 37744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_360
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_390
timestamp 1698431365
transform 1 0 45024 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_432
timestamp 1698431365
transform 1 0 49728 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_458
timestamp 1698431365
transform 1 0 52640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_462
timestamp 1698431365
transform 1 0 53088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_466
timestamp 1698431365
transform 1 0 53536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_470
timestamp 1698431365
transform 1 0 53984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_474
timestamp 1698431365
transform 1 0 54432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_488
timestamp 1698431365
transform 1 0 56000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_496
timestamp 1698431365
transform 1 0 56896 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_499
timestamp 1698431365
transform 1 0 57232 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_31
timestamp 1698431365
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_41
timestamp 1698431365
transform 1 0 5936 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_45
timestamp 1698431365
transform 1 0 6384 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_53
timestamp 1698431365
transform 1 0 7280 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_77
timestamp 1698431365
transform 1 0 9968 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_85
timestamp 1698431365
transform 1 0 10864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_87
timestamp 1698431365
transform 1 0 11088 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_113
timestamp 1698431365
transform 1 0 14000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_126
timestamp 1698431365
transform 1 0 15456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_128
timestamp 1698431365
transform 1 0 15680 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_135
timestamp 1698431365
transform 1 0 16464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_139
timestamp 1698431365
transform 1 0 16912 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_142
timestamp 1698431365
transform 1 0 17248 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_146
timestamp 1698431365
transform 1 0 17696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_150
timestamp 1698431365
transform 1 0 18144 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_154
timestamp 1698431365
transform 1 0 18592 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_157
timestamp 1698431365
transform 1 0 18928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_161
timestamp 1698431365
transform 1 0 19376 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_169
timestamp 1698431365
transform 1 0 20272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_185
timestamp 1698431365
transform 1 0 22064 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_190
timestamp 1698431365
transform 1 0 22624 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_206
timestamp 1698431365
transform 1 0 24416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_210
timestamp 1698431365
transform 1 0 24864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_220
timestamp 1698431365
transform 1 0 25984 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_228
timestamp 1698431365
transform 1 0 26880 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_232
timestamp 1698431365
transform 1 0 27328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_234
timestamp 1698431365
transform 1 0 27552 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_266
timestamp 1698431365
transform 1 0 31136 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_277
timestamp 1698431365
transform 1 0 32368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_301
timestamp 1698431365
transform 1 0 35056 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_303
timestamp 1698431365
transform 1 0 35280 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_310
timestamp 1698431365
transform 1 0 36064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698431365
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_325
timestamp 1698431365
transform 1 0 37744 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_345
timestamp 1698431365
transform 1 0 39984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_349
timestamp 1698431365
transform 1 0 40432 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_353
timestamp 1698431365
transform 1 0 40880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_355
timestamp 1698431365
transform 1 0 41104 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_363
timestamp 1698431365
transform 1 0 42000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_375
timestamp 1698431365
transform 1 0 43344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_379
timestamp 1698431365
transform 1 0 43792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_383
timestamp 1698431365
transform 1 0 44240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_391
timestamp 1698431365
transform 1 0 45136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_399
timestamp 1698431365
transform 1 0 46032 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_403
timestamp 1698431365
transform 1 0 46480 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_407
timestamp 1698431365
transform 1 0 46928 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_423
timestamp 1698431365
transform 1 0 48720 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_431
timestamp 1698431365
transform 1 0 49616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_433
timestamp 1698431365
transform 1 0 49840 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_440
timestamp 1698431365
transform 1 0 50624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_454
timestamp 1698431365
transform 1 0 52192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_463
timestamp 1698431365
transform 1 0 53200 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_476
timestamp 1698431365
transform 1 0 54656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_57
timestamp 1698431365
transform 1 0 7728 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_61
timestamp 1698431365
transform 1 0 8176 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_80
timestamp 1698431365
transform 1 0 10304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_84
timestamp 1698431365
transform 1 0 10752 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_103
timestamp 1698431365
transform 1 0 12880 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_107
timestamp 1698431365
transform 1 0 13328 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_123
timestamp 1698431365
transform 1 0 15120 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_131
timestamp 1698431365
transform 1 0 16016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_133
timestamp 1698431365
transform 1 0 16240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_148
timestamp 1698431365
transform 1 0 17920 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_186
timestamp 1698431365
transform 1 0 22176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_190
timestamp 1698431365
transform 1 0 22624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_192
timestamp 1698431365
transform 1 0 22848 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698431365
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_228
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_232
timestamp 1698431365
transform 1 0 27328 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_237
timestamp 1698431365
transform 1 0 27888 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_248
timestamp 1698431365
transform 1 0 29120 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_271
timestamp 1698431365
transform 1 0 31696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_273
timestamp 1698431365
transform 1 0 31920 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_305
timestamp 1698431365
transform 1 0 35504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_309
timestamp 1698431365
transform 1 0 35952 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_313
timestamp 1698431365
transform 1 0 36400 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_315
timestamp 1698431365
transform 1 0 36624 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_330
timestamp 1698431365
transform 1 0 38304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_332
timestamp 1698431365
transform 1 0 38528 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_345
timestamp 1698431365
transform 1 0 39984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_356
timestamp 1698431365
transform 1 0 41216 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_360
timestamp 1698431365
transform 1 0 41664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_364
timestamp 1698431365
transform 1 0 42112 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_368
timestamp 1698431365
transform 1 0 42560 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_374
timestamp 1698431365
transform 1 0 43232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_378
timestamp 1698431365
transform 1 0 43680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_382
timestamp 1698431365
transform 1 0 44128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_386
timestamp 1698431365
transform 1 0 44576 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_402
timestamp 1698431365
transform 1 0 46368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_406
timestamp 1698431365
transform 1 0 46816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_410
timestamp 1698431365
transform 1 0 47264 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_419
timestamp 1698431365
transform 1 0 48272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_434
timestamp 1698431365
transform 1 0 49952 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_438
timestamp 1698431365
transform 1 0 50400 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_462
timestamp 1698431365
transform 1 0 53088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_478
timestamp 1698431365
transform 1 0 54880 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_488
timestamp 1698431365
transform 1 0 56000 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_496
timestamp 1698431365
transform 1 0 56896 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_113
timestamp 1698431365
transform 1 0 14000 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_117
timestamp 1698431365
transform 1 0 14448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_156
timestamp 1698431365
transform 1 0 18816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_168
timestamp 1698431365
transform 1 0 20160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_170
timestamp 1698431365
transform 1 0 20384 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_186
timestamp 1698431365
transform 1 0 22176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_252
timestamp 1698431365
transform 1 0 29568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_256
timestamp 1698431365
transform 1 0 30016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_260
timestamp 1698431365
transform 1 0 30464 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_263
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_267
timestamp 1698431365
transform 1 0 31248 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_271
timestamp 1698431365
transform 1 0 31696 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_274
timestamp 1698431365
transform 1 0 32032 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_295
timestamp 1698431365
transform 1 0 34384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_309
timestamp 1698431365
transform 1 0 35952 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_313
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_339
timestamp 1698431365
transform 1 0 39312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_341
timestamp 1698431365
transform 1 0 39536 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_364
timestamp 1698431365
transform 1 0 42112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_371
timestamp 1698431365
transform 1 0 42896 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_382
timestamp 1698431365
transform 1 0 44128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_424
timestamp 1698431365
transform 1 0 48832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_428
timestamp 1698431365
transform 1 0 49280 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_436
timestamp 1698431365
transform 1 0 50176 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_470
timestamp 1698431365
transform 1 0 53984 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_474
timestamp 1698431365
transform 1 0 54432 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_507
timestamp 1698431365
transform 1 0 58128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_14
timestamp 1698431365
transform 1 0 2912 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_20
timestamp 1698431365
transform 1 0 3584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_24
timestamp 1698431365
transform 1 0 4032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_32
timestamp 1698431365
transform 1 0 4928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_47
timestamp 1698431365
transform 1 0 6608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_51
timestamp 1698431365
transform 1 0 7056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_55
timestamp 1698431365
transform 1 0 7504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_59
timestamp 1698431365
transform 1 0 7952 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_67
timestamp 1698431365
transform 1 0 8848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_76
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698431365
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698431365
transform 1 0 10752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_86
timestamp 1698431365
transform 1 0 10976 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_124
timestamp 1698431365
transform 1 0 15232 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_131
timestamp 1698431365
transform 1 0 16016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698431365
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_151
timestamp 1698431365
transform 1 0 18256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_157
timestamp 1698431365
transform 1 0 18928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_188
timestamp 1698431365
transform 1 0 22400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_194
timestamp 1698431365
transform 1 0 23072 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_204
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_214
timestamp 1698431365
transform 1 0 25312 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_261
timestamp 1698431365
transform 1 0 30576 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698431365
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_294
timestamp 1698431365
transform 1 0 34272 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_296
timestamp 1698431365
transform 1 0 34496 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_315
timestamp 1698431365
transform 1 0 36624 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_323
timestamp 1698431365
transform 1 0 37520 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_327
timestamp 1698431365
transform 1 0 37968 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_348
timestamp 1698431365
transform 1 0 40320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_378
timestamp 1698431365
transform 1 0 43680 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_387
timestamp 1698431365
transform 1 0 44688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_418
timestamp 1698431365
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_426
timestamp 1698431365
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_428
timestamp 1698431365
transform 1 0 49280 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_470
timestamp 1698431365
transform 1 0 53984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_474
timestamp 1698431365
transform 1 0 54432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_494
timestamp 1698431365
transform 1 0 56672 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_10
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_30
timestamp 1698431365
transform 1 0 4704 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_33
timestamp 1698431365
transform 1 0 5040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_46
timestamp 1698431365
transform 1 0 6496 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_53
timestamp 1698431365
transform 1 0 7280 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_57
timestamp 1698431365
transform 1 0 7728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_61
timestamp 1698431365
transform 1 0 8176 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_69
timestamp 1698431365
transform 1 0 9072 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_73
timestamp 1698431365
transform 1 0 9520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_75
timestamp 1698431365
transform 1 0 9744 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_82
timestamp 1698431365
transform 1 0 10528 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_98
timestamp 1698431365
transform 1 0 12320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_102
timestamp 1698431365
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_117
timestamp 1698431365
transform 1 0 14448 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_124
timestamp 1698431365
transform 1 0 15232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_128
timestamp 1698431365
transform 1 0 15680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_130
timestamp 1698431365
transform 1 0 15904 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_133
timestamp 1698431365
transform 1 0 16240 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_141
timestamp 1698431365
transform 1 0 17136 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_145
timestamp 1698431365
transform 1 0 17584 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_147
timestamp 1698431365
transform 1 0 17808 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_150
timestamp 1698431365
transform 1 0 18144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_154
timestamp 1698431365
transform 1 0 18592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_156
timestamp 1698431365
transform 1 0 18816 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_167
timestamp 1698431365
transform 1 0 20048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_192
timestamp 1698431365
transform 1 0 22848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_200
timestamp 1698431365
transform 1 0 23744 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_209
timestamp 1698431365
transform 1 0 24752 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_213
timestamp 1698431365
transform 1 0 25200 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_217
timestamp 1698431365
transform 1 0 25648 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_236
timestamp 1698431365
transform 1 0 27776 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_264
timestamp 1698431365
transform 1 0 30912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_276
timestamp 1698431365
transform 1 0 32256 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_284
timestamp 1698431365
transform 1 0 33152 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_288
timestamp 1698431365
transform 1 0 33600 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_300
timestamp 1698431365
transform 1 0 34944 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_307
timestamp 1698431365
transform 1 0 35728 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698431365
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_323
timestamp 1698431365
transform 1 0 37520 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_355
timestamp 1698431365
transform 1 0 41104 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_368
timestamp 1698431365
transform 1 0 42560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_370
timestamp 1698431365
transform 1 0 42784 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_373
timestamp 1698431365
transform 1 0 43120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_377
timestamp 1698431365
transform 1 0 43568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_381
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_389
timestamp 1698431365
transform 1 0 44912 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_396
timestamp 1698431365
transform 1 0 45696 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_412
timestamp 1698431365
transform 1 0 47488 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_431
timestamp 1698431365
transform 1 0 49616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_467
timestamp 1698431365
transform 1 0 53648 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_475
timestamp 1698431365
transform 1 0 54544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_477
timestamp 1698431365
transform 1 0 54768 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_55
timestamp 1698431365
transform 1 0 7504 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_57
timestamp 1698431365
transform 1 0 7728 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_84
timestamp 1698431365
transform 1 0 10752 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_88
timestamp 1698431365
transform 1 0 11200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_90
timestamp 1698431365
transform 1 0 11424 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_99
timestamp 1698431365
transform 1 0 12432 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_103
timestamp 1698431365
transform 1 0 12880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_110
timestamp 1698431365
transform 1 0 13664 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_114
timestamp 1698431365
transform 1 0 14112 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_132
timestamp 1698431365
transform 1 0 16128 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_163
timestamp 1698431365
transform 1 0 19600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_167
timestamp 1698431365
transform 1 0 20048 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_173
timestamp 1698431365
transform 1 0 20720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_177
timestamp 1698431365
transform 1 0 21168 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_196
timestamp 1698431365
transform 1 0 23296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_200
timestamp 1698431365
transform 1 0 23744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_202
timestamp 1698431365
transform 1 0 23968 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_205
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_220
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_224
timestamp 1698431365
transform 1 0 26432 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_232
timestamp 1698431365
transform 1 0 27328 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_255
timestamp 1698431365
transform 1 0 29904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_259
timestamp 1698431365
transform 1 0 30352 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_272
timestamp 1698431365
transform 1 0 31808 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_286
timestamp 1698431365
transform 1 0 33376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_298
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_300
timestamp 1698431365
transform 1 0 34944 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_309
timestamp 1698431365
transform 1 0 35952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_316
timestamp 1698431365
transform 1 0 36736 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_318
timestamp 1698431365
transform 1 0 36960 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_321
timestamp 1698431365
transform 1 0 37296 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_325
timestamp 1698431365
transform 1 0 37744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_329
timestamp 1698431365
transform 1 0 38192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_333
timestamp 1698431365
transform 1 0 38640 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_356
timestamp 1698431365
transform 1 0 41216 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_363
timestamp 1698431365
transform 1 0 42000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_365
timestamp 1698431365
transform 1 0 42224 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_376
timestamp 1698431365
transform 1 0 43456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_380
timestamp 1698431365
transform 1 0 43904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_384
timestamp 1698431365
transform 1 0 44352 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_388
timestamp 1698431365
transform 1 0 44800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_392
timestamp 1698431365
transform 1 0 45248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_396
timestamp 1698431365
transform 1 0 45696 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_404
timestamp 1698431365
transform 1 0 46592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_408
timestamp 1698431365
transform 1 0 47040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_418
timestamp 1698431365
transform 1 0 48160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_428
timestamp 1698431365
transform 1 0 49280 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_442
timestamp 1698431365
transform 1 0 50848 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_453
timestamp 1698431365
transform 1 0 52080 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_457
timestamp 1698431365
transform 1 0 52528 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_463
timestamp 1698431365
transform 1 0 53200 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_475
timestamp 1698431365
transform 1 0 54544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_477
timestamp 1698431365
transform 1 0 54768 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_487
timestamp 1698431365
transform 1 0 55888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_489
timestamp 1698431365
transform 1 0 56112 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_496
timestamp 1698431365
transform 1 0 56896 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_14
timestamp 1698431365
transform 1 0 2912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_41
timestamp 1698431365
transform 1 0 5936 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_43
timestamp 1698431365
transform 1 0 6160 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_50
timestamp 1698431365
transform 1 0 6944 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_54
timestamp 1698431365
transform 1 0 7392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_56
timestamp 1698431365
transform 1 0 7616 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_122
timestamp 1698431365
transform 1 0 15008 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_152
timestamp 1698431365
transform 1 0 18368 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_161
timestamp 1698431365
transform 1 0 19376 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_185
timestamp 1698431365
transform 1 0 22064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_236
timestamp 1698431365
transform 1 0 27776 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_262
timestamp 1698431365
transform 1 0 30688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_286
timestamp 1698431365
transform 1 0 33376 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_300
timestamp 1698431365
transform 1 0 34944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_304
timestamp 1698431365
transform 1 0 35392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_306
timestamp 1698431365
transform 1 0 35616 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_327
timestamp 1698431365
transform 1 0 37968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_336
timestamp 1698431365
transform 1 0 38976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_340
timestamp 1698431365
transform 1 0 39424 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_344
timestamp 1698431365
transform 1 0 39872 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_346
timestamp 1698431365
transform 1 0 40096 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_349
timestamp 1698431365
transform 1 0 40432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_361
timestamp 1698431365
transform 1 0 41776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_365
timestamp 1698431365
transform 1 0 42224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_403
timestamp 1698431365
transform 1 0 46480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_424
timestamp 1698431365
transform 1 0 48832 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_440
timestamp 1698431365
transform 1 0 50624 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_475
timestamp 1698431365
transform 1 0 54544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_477
timestamp 1698431365
transform 1 0 54768 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_14
timestamp 1698431365
transform 1 0 2912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_26
timestamp 1698431365
transform 1 0 4256 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_40
timestamp 1698431365
transform 1 0 5824 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_48
timestamp 1698431365
transform 1 0 6720 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_52
timestamp 1698431365
transform 1 0 7168 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_61
timestamp 1698431365
transform 1 0 8176 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_80
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_88
timestamp 1698431365
transform 1 0 11200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_120
timestamp 1698431365
transform 1 0 14784 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_156
timestamp 1698431365
transform 1 0 18816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_214
timestamp 1698431365
transform 1 0 25312 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_223
timestamp 1698431365
transform 1 0 26320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_227
timestamp 1698431365
transform 1 0 26768 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_235
timestamp 1698431365
transform 1 0 27664 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_255
timestamp 1698431365
transform 1 0 29904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_259
timestamp 1698431365
transform 1 0 30352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_263
timestamp 1698431365
transform 1 0 30800 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_266
timestamp 1698431365
transform 1 0 31136 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_296
timestamp 1698431365
transform 1 0 34496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_300
timestamp 1698431365
transform 1 0 34944 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_304
timestamp 1698431365
transform 1 0 35392 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_306
timestamp 1698431365
transform 1 0 35616 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_341
timestamp 1698431365
transform 1 0 39536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_371
timestamp 1698431365
transform 1 0 42896 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_385
timestamp 1698431365
transform 1 0 44464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_389
timestamp 1698431365
transform 1 0 44912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_426
timestamp 1698431365
transform 1 0 49056 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_430
timestamp 1698431365
transform 1 0 49504 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_487
timestamp 1698431365
transform 1 0 55888 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_489
timestamp 1698431365
transform 1 0 56112 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_496
timestamp 1698431365
transform 1 0 56896 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_499
timestamp 1698431365
transform 1 0 57232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_31
timestamp 1698431365
transform 1 0 4816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_39
timestamp 1698431365
transform 1 0 5712 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_66
timestamp 1698431365
transform 1 0 8736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_74
timestamp 1698431365
transform 1 0 9632 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_90
timestamp 1698431365
transform 1 0 11424 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_98
timestamp 1698431365
transform 1 0 12320 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_115
timestamp 1698431365
transform 1 0 14224 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_131
timestamp 1698431365
transform 1 0 16016 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_139
timestamp 1698431365
transform 1 0 16912 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_143
timestamp 1698431365
transform 1 0 17360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_145
timestamp 1698431365
transform 1 0 17584 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_158
timestamp 1698431365
transform 1 0 19040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_162
timestamp 1698431365
transform 1 0 19488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_166
timestamp 1698431365
transform 1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_170
timestamp 1698431365
transform 1 0 20384 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_188
timestamp 1698431365
transform 1 0 22400 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_196
timestamp 1698431365
transform 1 0 23296 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_200
timestamp 1698431365
transform 1 0 23744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_204
timestamp 1698431365
transform 1 0 24192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_206
timestamp 1698431365
transform 1 0 24416 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_215
timestamp 1698431365
transform 1 0 25424 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_222
timestamp 1698431365
transform 1 0 26208 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_226
timestamp 1698431365
transform 1 0 26656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_228
timestamp 1698431365
transform 1 0 26880 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_265
timestamp 1698431365
transform 1 0 31024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_267
timestamp 1698431365
transform 1 0 31248 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_280
timestamp 1698431365
transform 1 0 32704 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_288
timestamp 1698431365
transform 1 0 33600 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_292
timestamp 1698431365
transform 1 0 34048 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_296
timestamp 1698431365
transform 1 0 34496 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_321
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_329
timestamp 1698431365
transform 1 0 38192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_333
timestamp 1698431365
transform 1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_337
timestamp 1698431365
transform 1 0 39088 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_345
timestamp 1698431365
transform 1 0 39984 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_370
timestamp 1698431365
transform 1 0 42784 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_381
timestamp 1698431365
transform 1 0 44016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_399
timestamp 1698431365
transform 1 0 46032 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_408
timestamp 1698431365
transform 1 0 47040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_410
timestamp 1698431365
transform 1 0 47264 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_419
timestamp 1698431365
transform 1 0 48272 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_423
timestamp 1698431365
transform 1 0 48720 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_431
timestamp 1698431365
transform 1 0 49616 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_452
timestamp 1698431365
transform 1 0 51968 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_454
timestamp 1698431365
transform 1 0 52192 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_473
timestamp 1698431365
transform 1 0 54320 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_484
timestamp 1698431365
transform 1 0 55552 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_489
timestamp 1698431365
transform 1 0 56112 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_493
timestamp 1698431365
transform 1 0 56560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_499
timestamp 1698431365
transform 1 0 57232 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_14
timestamp 1698431365
transform 1 0 2912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_31
timestamp 1698431365
transform 1 0 4816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_35
timestamp 1698431365
transform 1 0 5264 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_62
timestamp 1698431365
transform 1 0 8288 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_64
timestamp 1698431365
transform 1 0 8512 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_80
timestamp 1698431365
transform 1 0 10304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_82
timestamp 1698431365
transform 1 0 10528 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_85
timestamp 1698431365
transform 1 0 10864 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_93
timestamp 1698431365
transform 1 0 11760 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_125
timestamp 1698431365
transform 1 0 15344 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_133
timestamp 1698431365
transform 1 0 16240 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_137
timestamp 1698431365
transform 1 0 16688 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_201
timestamp 1698431365
transform 1 0 23856 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_216
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_253
timestamp 1698431365
transform 1 0 29680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_297
timestamp 1698431365
transform 1 0 34608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_299
timestamp 1698431365
transform 1 0 34832 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_308
timestamp 1698431365
transform 1 0 35840 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_325
timestamp 1698431365
transform 1 0 37744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_342
timestamp 1698431365
transform 1 0 39648 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_356
timestamp 1698431365
transform 1 0 41216 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_359
timestamp 1698431365
transform 1 0 41552 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_376
timestamp 1698431365
transform 1 0 43456 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_395
timestamp 1698431365
transform 1 0 45584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_397
timestamp 1698431365
transform 1 0 45808 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_400
timestamp 1698431365
transform 1 0 46144 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_408
timestamp 1698431365
transform 1 0 47040 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698431365
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_424
timestamp 1698431365
transform 1 0 48832 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_437
timestamp 1698431365
transform 1 0 50288 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_449
timestamp 1698431365
transform 1 0 51632 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_465
timestamp 1698431365
transform 1 0 53424 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_489
timestamp 1698431365
transform 1 0 56112 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_494
timestamp 1698431365
transform 1 0 56672 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_31
timestamp 1698431365
transform 1 0 4816 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_45
timestamp 1698431365
transform 1 0 6384 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_53
timestamp 1698431365
transform 1 0 7280 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_57
timestamp 1698431365
transform 1 0 7728 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_89
timestamp 1698431365
transform 1 0 11312 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_97
timestamp 1698431365
transform 1 0 12208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_113
timestamp 1698431365
transform 1 0 14000 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_129
timestamp 1698431365
transform 1 0 15792 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_159
timestamp 1698431365
transform 1 0 19152 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_163
timestamp 1698431365
transform 1 0 19600 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_183
timestamp 1698431365
transform 1 0 21840 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_185
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_207
timestamp 1698431365
transform 1 0 24528 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_211
timestamp 1698431365
transform 1 0 24976 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_227
timestamp 1698431365
transform 1 0 26768 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_234
timestamp 1698431365
transform 1 0 27552 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_242
timestamp 1698431365
transform 1 0 28448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_265
timestamp 1698431365
transform 1 0 31024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_267
timestamp 1698431365
transform 1 0 31248 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_324
timestamp 1698431365
transform 1 0 37632 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_348
timestamp 1698431365
transform 1 0 40320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_356
timestamp 1698431365
transform 1 0 41216 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_372
timestamp 1698431365
transform 1 0 43008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_380
timestamp 1698431365
transform 1 0 43904 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_383
timestamp 1698431365
transform 1 0 44240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_402
timestamp 1698431365
transform 1 0 46368 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_410
timestamp 1698431365
transform 1 0 47264 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_414
timestamp 1698431365
transform 1 0 47712 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_416
timestamp 1698431365
transform 1 0 47936 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_441
timestamp 1698431365
transform 1 0 50736 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_454
timestamp 1698431365
transform 1 0 52192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_467
timestamp 1698431365
transform 1 0 53648 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_469
timestamp 1698431365
transform 1 0 53872 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_476
timestamp 1698431365
transform 1 0 54656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_20
timestamp 1698431365
transform 1 0 3584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_35
timestamp 1698431365
transform 1 0 5264 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_39
timestamp 1698431365
transform 1 0 5712 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_43
timestamp 1698431365
transform 1 0 6160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_47
timestamp 1698431365
transform 1 0 6608 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_55
timestamp 1698431365
transform 1 0 7504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_57
timestamp 1698431365
transform 1 0 7728 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_84
timestamp 1698431365
transform 1 0 10752 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_104
timestamp 1698431365
transform 1 0 12992 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_108
timestamp 1698431365
transform 1 0 13440 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_116
timestamp 1698431365
transform 1 0 14336 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_120
timestamp 1698431365
transform 1 0 14784 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_123
timestamp 1698431365
transform 1 0 15120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_137
timestamp 1698431365
transform 1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_159
timestamp 1698431365
transform 1 0 19152 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_172
timestamp 1698431365
transform 1 0 20608 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_208
timestamp 1698431365
transform 1 0 24640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_218
timestamp 1698431365
transform 1 0 25760 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_222
timestamp 1698431365
transform 1 0 26208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_224
timestamp 1698431365
transform 1 0 26432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_240
timestamp 1698431365
transform 1 0 28224 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_248
timestamp 1698431365
transform 1 0 29120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_250
timestamp 1698431365
transform 1 0 29344 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_277
timestamp 1698431365
transform 1 0 32368 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_279
timestamp 1698431365
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_297
timestamp 1698431365
transform 1 0 34608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_299
timestamp 1698431365
transform 1 0 34832 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_310
timestamp 1698431365
transform 1 0 36064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_312
timestamp 1698431365
transform 1 0 36288 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_317
timestamp 1698431365
transform 1 0 36848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_321
timestamp 1698431365
transform 1 0 37296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_381
timestamp 1698431365
transform 1 0 44016 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_417
timestamp 1698431365
transform 1 0 48048 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_419
timestamp 1698431365
transform 1 0 48272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_426
timestamp 1698431365
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_428
timestamp 1698431365
transform 1 0 49280 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_481
timestamp 1698431365
transform 1 0 55216 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_487
timestamp 1698431365
transform 1 0 55888 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_489
timestamp 1698431365
transform 1 0 56112 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_496
timestamp 1698431365
transform 1 0 56896 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_504
timestamp 1698431365
transform 1 0 57792 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_508
timestamp 1698431365
transform 1 0 58240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_8
timestamp 1698431365
transform 1 0 2240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_10
timestamp 1698431365
transform 1 0 2464 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_39
timestamp 1698431365
transform 1 0 5712 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_48
timestamp 1698431365
transform 1 0 6720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_50
timestamp 1698431365
transform 1 0 6944 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_83
timestamp 1698431365
transform 1 0 10640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_85
timestamp 1698431365
transform 1 0 10864 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_94
timestamp 1698431365
transform 1 0 11872 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_98
timestamp 1698431365
transform 1 0 12320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_102
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_151
timestamp 1698431365
transform 1 0 18256 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_173
timestamp 1698431365
transform 1 0 20720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_185
timestamp 1698431365
transform 1 0 22064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_187
timestamp 1698431365
transform 1 0 22288 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_211
timestamp 1698431365
transform 1 0 24976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_213
timestamp 1698431365
transform 1 0 25200 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_249
timestamp 1698431365
transform 1 0 29232 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_306
timestamp 1698431365
transform 1 0 35616 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_312
timestamp 1698431365
transform 1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_325
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_339
timestamp 1698431365
transform 1 0 39312 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_347
timestamp 1698431365
transform 1 0 40208 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_366
timestamp 1698431365
transform 1 0 42336 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_370
timestamp 1698431365
transform 1 0 42784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_380
timestamp 1698431365
transform 1 0 43904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698431365
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_403
timestamp 1698431365
transform 1 0 46480 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_407
timestamp 1698431365
transform 1 0 46928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_409
timestamp 1698431365
transform 1 0 47152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_439
timestamp 1698431365
transform 1 0 50512 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_445
timestamp 1698431365
transform 1 0 51184 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_465
timestamp 1698431365
transform 1 0 53424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_482
timestamp 1698431365
transform 1 0 55328 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_486
timestamp 1698431365
transform 1 0 55776 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_502
timestamp 1698431365
transform 1 0 57568 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_506
timestamp 1698431365
transform 1 0 58016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_508
timestamp 1698431365
transform 1 0 58240 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_31
timestamp 1698431365
transform 1 0 4816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_33
timestamp 1698431365
transform 1 0 5040 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_52
timestamp 1698431365
transform 1 0 7168 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_109
timestamp 1698431365
transform 1 0 13552 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_132
timestamp 1698431365
transform 1 0 16128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_158
timestamp 1698431365
transform 1 0 19040 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_162
timestamp 1698431365
transform 1 0 19488 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_169
timestamp 1698431365
transform 1 0 20272 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_179
timestamp 1698431365
transform 1 0 21392 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_195
timestamp 1698431365
transform 1 0 23184 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_203
timestamp 1698431365
transform 1 0 24080 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_207
timestamp 1698431365
transform 1 0 24528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698431365
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_221
timestamp 1698431365
transform 1 0 26096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_229
timestamp 1698431365
transform 1 0 26992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_233
timestamp 1698431365
transform 1 0 27440 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_241
timestamp 1698431365
transform 1 0 28336 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_245
timestamp 1698431365
transform 1 0 28784 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_247
timestamp 1698431365
transform 1 0 29008 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_259
timestamp 1698431365
transform 1 0 30352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_263
timestamp 1698431365
transform 1 0 30800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_292
timestamp 1698431365
transform 1 0 34048 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_296
timestamp 1698431365
transform 1 0 34496 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_300
timestamp 1698431365
transform 1 0 34944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_314
timestamp 1698431365
transform 1 0 36512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_318
timestamp 1698431365
transform 1 0 36960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_322
timestamp 1698431365
transform 1 0 37408 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_330
timestamp 1698431365
transform 1 0 38304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_332
timestamp 1698431365
transform 1 0 38528 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_342
timestamp 1698431365
transform 1 0 39648 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_356
timestamp 1698431365
transform 1 0 41216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_358
timestamp 1698431365
transform 1 0 41440 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_388
timestamp 1698431365
transform 1 0 44800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_392
timestamp 1698431365
transform 1 0 45248 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_408
timestamp 1698431365
transform 1 0 47040 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_418
timestamp 1698431365
transform 1 0 48160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_438
timestamp 1698431365
transform 1 0 50400 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_441
timestamp 1698431365
transform 1 0 50736 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_459
timestamp 1698431365
transform 1 0 52752 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_508
timestamp 1698431365
transform 1 0 58240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_83
timestamp 1698431365
transform 1 0 10640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_87
timestamp 1698431365
transform 1 0 11088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_89
timestamp 1698431365
transform 1 0 11312 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_95
timestamp 1698431365
transform 1 0 11984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_113
timestamp 1698431365
transform 1 0 14000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_117
timestamp 1698431365
transform 1 0 14448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_119
timestamp 1698431365
transform 1 0 14672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_133
timestamp 1698431365
transform 1 0 16240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_135
timestamp 1698431365
transform 1 0 16464 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_138
timestamp 1698431365
transform 1 0 16800 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_191
timestamp 1698431365
transform 1 0 22736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_195
timestamp 1698431365
transform 1 0 23184 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_238
timestamp 1698431365
transform 1 0 28000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_240
timestamp 1698431365
transform 1 0 28224 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_280
timestamp 1698431365
transform 1 0 32704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_284
timestamp 1698431365
transform 1 0 33152 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_288
timestamp 1698431365
transform 1 0 33600 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_321
timestamp 1698431365
transform 1 0 37296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_329
timestamp 1698431365
transform 1 0 38192 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_345
timestamp 1698431365
transform 1 0 39984 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_361
timestamp 1698431365
transform 1 0 41776 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_365
timestamp 1698431365
transform 1 0 42224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_367
timestamp 1698431365
transform 1 0 42448 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_370
timestamp 1698431365
transform 1 0 42784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_374
timestamp 1698431365
transform 1 0 43232 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_378
timestamp 1698431365
transform 1 0 43680 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_449
timestamp 1698431365
transform 1 0 51632 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_453
timestamp 1698431365
transform 1 0 52080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_461
timestamp 1698431365
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_465
timestamp 1698431365
transform 1 0 53424 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_477
timestamp 1698431365
transform 1 0 54768 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_6
timestamp 1698431365
transform 1 0 2016 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_22
timestamp 1698431365
transform 1 0 3808 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_57
timestamp 1698431365
transform 1 0 7728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_61
timestamp 1698431365
transform 1 0 8176 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_67
timestamp 1698431365
transform 1 0 8848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698431365
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_76
timestamp 1698431365
transform 1 0 9856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_84
timestamp 1698431365
transform 1 0 10752 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_88
timestamp 1698431365
transform 1 0 11200 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_96
timestamp 1698431365
transform 1 0 12096 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_128
timestamp 1698431365
transform 1 0 15680 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_138
timestamp 1698431365
transform 1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_144
timestamp 1698431365
transform 1 0 17472 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_158
timestamp 1698431365
transform 1 0 19040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_189
timestamp 1698431365
transform 1 0 22512 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_205
timestamp 1698431365
transform 1 0 24304 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_207
timestamp 1698431365
transform 1 0 24528 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_218
timestamp 1698431365
transform 1 0 25760 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_222
timestamp 1698431365
transform 1 0 26208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_226
timestamp 1698431365
transform 1 0 26656 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_242
timestamp 1698431365
transform 1 0 28448 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_250
timestamp 1698431365
transform 1 0 29344 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_257
timestamp 1698431365
transform 1 0 30128 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_267
timestamp 1698431365
transform 1 0 31248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_269
timestamp 1698431365
transform 1 0 31472 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_272
timestamp 1698431365
transform 1 0 31808 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_286
timestamp 1698431365
transform 1 0 33376 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_288
timestamp 1698431365
transform 1 0 33600 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_291
timestamp 1698431365
transform 1 0 33936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_295
timestamp 1698431365
transform 1 0 34384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_356
timestamp 1698431365
transform 1 0 41216 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_376
timestamp 1698431365
transform 1 0 43456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_380
timestamp 1698431365
transform 1 0 43904 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_384
timestamp 1698431365
transform 1 0 44352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_401
timestamp 1698431365
transform 1 0 46256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_405
timestamp 1698431365
transform 1 0 46704 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_430
timestamp 1698431365
transform 1 0 49504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_434
timestamp 1698431365
transform 1 0 49952 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_456
timestamp 1698431365
transform 1 0 52416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_470
timestamp 1698431365
transform 1 0 53984 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698431365
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_508
timestamp 1698431365
transform 1 0 58240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_42
timestamp 1698431365
transform 1 0 6048 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_74
timestamp 1698431365
transform 1 0 9632 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_82
timestamp 1698431365
transform 1 0 10528 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_88
timestamp 1698431365
transform 1 0 11200 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_111
timestamp 1698431365
transform 1 0 13776 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_117
timestamp 1698431365
transform 1 0 14448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_150
timestamp 1698431365
transform 1 0 18144 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_166
timestamp 1698431365
transform 1 0 19936 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_174
timestamp 1698431365
transform 1 0 20832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_183
timestamp 1698431365
transform 1 0 21840 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_208
timestamp 1698431365
transform 1 0 24640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_210
timestamp 1698431365
transform 1 0 24864 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_213
timestamp 1698431365
transform 1 0 25200 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_217
timestamp 1698431365
transform 1 0 25648 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_229
timestamp 1698431365
transform 1 0 26992 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_233
timestamp 1698431365
transform 1 0 27440 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_237
timestamp 1698431365
transform 1 0 27888 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_265
timestamp 1698431365
transform 1 0 31024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_284
timestamp 1698431365
transform 1 0 33152 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_290
timestamp 1698431365
transform 1 0 33824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_321
timestamp 1698431365
transform 1 0 37296 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_325
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_327
timestamp 1698431365
transform 1 0 37968 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_350
timestamp 1698431365
transform 1 0 40544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_352
timestamp 1698431365
transform 1 0 40768 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_378
timestamp 1698431365
transform 1 0 43680 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_382
timestamp 1698431365
transform 1 0 44128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_391
timestamp 1698431365
transform 1 0 45136 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_395
timestamp 1698431365
transform 1 0 45584 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_397
timestamp 1698431365
transform 1 0 45808 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_436
timestamp 1698431365
transform 1 0 50176 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_469
timestamp 1698431365
transform 1 0 53872 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_473
timestamp 1698431365
transform 1 0 54320 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_481
timestamp 1698431365
transform 1 0 55216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_28
timestamp 1698431365
transform 1 0 4480 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_61
timestamp 1698431365
transform 1 0 8176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_65
timestamp 1698431365
transform 1 0 8624 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_101
timestamp 1698431365
transform 1 0 12656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_105
timestamp 1698431365
transform 1 0 13104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_109
timestamp 1698431365
transform 1 0 13552 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_121
timestamp 1698431365
transform 1 0 14896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_125
timestamp 1698431365
transform 1 0 15344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_129
timestamp 1698431365
transform 1 0 15792 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_134
timestamp 1698431365
transform 1 0 16352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_138
timestamp 1698431365
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_150
timestamp 1698431365
transform 1 0 18144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_160
timestamp 1698431365
transform 1 0 19264 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_192
timestamp 1698431365
transform 1 0 22848 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_229
timestamp 1698431365
transform 1 0 26992 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_247
timestamp 1698431365
transform 1 0 29008 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_268
timestamp 1698431365
transform 1 0 31360 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_272
timestamp 1698431365
transform 1 0 31808 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_288
timestamp 1698431365
transform 1 0 33600 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_326
timestamp 1698431365
transform 1 0 37856 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_330
timestamp 1698431365
transform 1 0 38304 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_338
timestamp 1698431365
transform 1 0 39200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_345
timestamp 1698431365
transform 1 0 39984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_396
timestamp 1698431365
transform 1 0 45696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_400
timestamp 1698431365
transform 1 0 46144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1698431365
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_440
timestamp 1698431365
transform 1 0 50624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_442
timestamp 1698431365
transform 1 0 50848 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_463
timestamp 1698431365
transform 1 0 53200 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_508
timestamp 1698431365
transform 1 0 58240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_14
timestamp 1698431365
transform 1 0 2912 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_18
timestamp 1698431365
transform 1 0 3360 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_84
timestamp 1698431365
transform 1 0 10752 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_88
timestamp 1698431365
transform 1 0 11200 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_92
timestamp 1698431365
transform 1 0 11648 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_95
timestamp 1698431365
transform 1 0 11984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_113
timestamp 1698431365
transform 1 0 14000 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_129
timestamp 1698431365
transform 1 0 15792 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_145
timestamp 1698431365
transform 1 0 17584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_149
timestamp 1698431365
transform 1 0 18032 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_157
timestamp 1698431365
transform 1 0 18928 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_170
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_181
timestamp 1698431365
transform 1 0 21616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_183
timestamp 1698431365
transform 1 0 21840 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_211
timestamp 1698431365
transform 1 0 24976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_213
timestamp 1698431365
transform 1 0 25200 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_219
timestamp 1698431365
transform 1 0 25872 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_233
timestamp 1698431365
transform 1 0 27440 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_251
timestamp 1698431365
transform 1 0 29456 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_270
timestamp 1698431365
transform 1 0 31584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_274
timestamp 1698431365
transform 1 0 32032 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_278
timestamp 1698431365
transform 1 0 32480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_288
timestamp 1698431365
transform 1 0 33600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_312
timestamp 1698431365
transform 1 0 36288 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1698431365
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_321
timestamp 1698431365
transform 1 0 37296 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_329
timestamp 1698431365
transform 1 0 38192 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_353
timestamp 1698431365
transform 1 0 40880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_357
timestamp 1698431365
transform 1 0 41328 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_373
timestamp 1698431365
transform 1 0 43120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_377
timestamp 1698431365
transform 1 0 43568 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_401
timestamp 1698431365
transform 1 0 46256 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_428
timestamp 1698431365
transform 1 0 49280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_432
timestamp 1698431365
transform 1 0 49728 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_436
timestamp 1698431365
transform 1 0 50176 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_465
timestamp 1698431365
transform 1 0 53424 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_495
timestamp 1698431365
transform 1 0 56784 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_503
timestamp 1698431365
transform 1 0 57680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_507
timestamp 1698431365
transform 1 0 58128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_8
timestamp 1698431365
transform 1 0 2240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_12
timestamp 1698431365
transform 1 0 2688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_16
timestamp 1698431365
transform 1 0 3136 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_32
timestamp 1698431365
transform 1 0 4928 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_36
timestamp 1698431365
transform 1 0 5376 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_48
timestamp 1698431365
transform 1 0 6720 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_55
timestamp 1698431365
transform 1 0 7504 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_63
timestamp 1698431365
transform 1 0 8400 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_67
timestamp 1698431365
transform 1 0 8848 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_69
timestamp 1698431365
transform 1 0 9072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_80
timestamp 1698431365
transform 1 0 10304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_84
timestamp 1698431365
transform 1 0 10752 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_86
timestamp 1698431365
transform 1 0 10976 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_93
timestamp 1698431365
transform 1 0 11760 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_95
timestamp 1698431365
transform 1 0 11984 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_118
timestamp 1698431365
transform 1 0 14560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_122
timestamp 1698431365
transform 1 0 15008 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_138
timestamp 1698431365
transform 1 0 16800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_146
timestamp 1698431365
transform 1 0 17696 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_185
timestamp 1698431365
transform 1 0 22064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_189
timestamp 1698431365
transform 1 0 22512 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_193
timestamp 1698431365
transform 1 0 22960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698431365
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698431365
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_224
timestamp 1698431365
transform 1 0 26432 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_231
timestamp 1698431365
transform 1 0 27216 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_233
timestamp 1698431365
transform 1 0 27440 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_252
timestamp 1698431365
transform 1 0 29568 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_256
timestamp 1698431365
transform 1 0 30016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_260
timestamp 1698431365
transform 1 0 30464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_264
timestamp 1698431365
transform 1 0 30912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_266
timestamp 1698431365
transform 1 0 31136 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698431365
transform 1 0 32144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_284
timestamp 1698431365
transform 1 0 33152 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_293
timestamp 1698431365
transform 1 0 34160 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_300
timestamp 1698431365
transform 1 0 34944 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_304
timestamp 1698431365
transform 1 0 35392 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_308
timestamp 1698431365
transform 1 0 35840 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_312
timestamp 1698431365
transform 1 0 36288 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_332
timestamp 1698431365
transform 1 0 38528 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_336
timestamp 1698431365
transform 1 0 38976 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_347
timestamp 1698431365
transform 1 0 40208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_366
timestamp 1698431365
transform 1 0 42336 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_382
timestamp 1698431365
transform 1 0 44128 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_390
timestamp 1698431365
transform 1 0 45024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_392
timestamp 1698431365
transform 1 0 45248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_415
timestamp 1698431365
transform 1 0 47824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_419
timestamp 1698431365
transform 1 0 48272 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_426
timestamp 1698431365
transform 1 0 49056 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_434
timestamp 1698431365
transform 1 0 49952 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_440
timestamp 1698431365
transform 1 0 50624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_462
timestamp 1698431365
transform 1 0 53088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_508
timestamp 1698431365
transform 1 0 58240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_8
timestamp 1698431365
transform 1 0 2240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_12
timestamp 1698431365
transform 1 0 2688 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_28
timestamp 1698431365
transform 1 0 4480 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_32
timestamp 1698431365
transform 1 0 4928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_48
timestamp 1698431365
transform 1 0 6720 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_87
timestamp 1698431365
transform 1 0 11088 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_102
timestamp 1698431365
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698431365
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_109
timestamp 1698431365
transform 1 0 13552 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_118
timestamp 1698431365
transform 1 0 14560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_157
timestamp 1698431365
transform 1 0 18928 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_161
timestamp 1698431365
transform 1 0 19376 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_170
timestamp 1698431365
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_172
timestamp 1698431365
transform 1 0 20608 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_191
timestamp 1698431365
transform 1 0 22736 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_193
timestamp 1698431365
transform 1 0 22960 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_202
timestamp 1698431365
transform 1 0 23968 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_234
timestamp 1698431365
transform 1 0 27552 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_237
timestamp 1698431365
transform 1 0 27888 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_261
timestamp 1698431365
transform 1 0 30576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_265
timestamp 1698431365
transform 1 0 31024 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_269
timestamp 1698431365
transform 1 0 31472 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_271
timestamp 1698431365
transform 1 0 31696 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_280
timestamp 1698431365
transform 1 0 32704 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_286
timestamp 1698431365
transform 1 0 33376 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_319
timestamp 1698431365
transform 1 0 37072 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_330
timestamp 1698431365
transform 1 0 38304 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_338
timestamp 1698431365
transform 1 0 39200 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_342
timestamp 1698431365
transform 1 0 39648 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_391
timestamp 1698431365
transform 1 0 45136 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_399
timestamp 1698431365
transform 1 0 46032 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_414
timestamp 1698431365
transform 1 0 47712 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_451
timestamp 1698431365
transform 1 0 51856 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_459
timestamp 1698431365
transform 1 0 52752 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_489
timestamp 1698431365
transform 1 0 56112 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_505
timestamp 1698431365
transform 1 0 57904 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_8
timestamp 1698431365
transform 1 0 2240 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_12
timestamp 1698431365
transform 1 0 2688 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_52
timestamp 1698431365
transform 1 0 7168 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_58
timestamp 1698431365
transform 1 0 7840 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_76
timestamp 1698431365
transform 1 0 9856 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_78
timestamp 1698431365
transform 1 0 10080 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_81
timestamp 1698431365
transform 1 0 10416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_85
timestamp 1698431365
transform 1 0 10864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_89
timestamp 1698431365
transform 1 0 11312 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_97
timestamp 1698431365
transform 1 0 12208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_99
timestamp 1698431365
transform 1 0 12432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_112
timestamp 1698431365
transform 1 0 13888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_116
timestamp 1698431365
transform 1 0 14336 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_124
timestamp 1698431365
transform 1 0 15232 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_132
timestamp 1698431365
transform 1 0 16128 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_158
timestamp 1698431365
transform 1 0 19040 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_166
timestamp 1698431365
transform 1 0 19936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_170
timestamp 1698431365
transform 1 0 20384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_172
timestamp 1698431365
transform 1 0 20608 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_181
timestamp 1698431365
transform 1 0 21616 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_190
timestamp 1698431365
transform 1 0 22624 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_208
timestamp 1698431365
transform 1 0 24640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_286
timestamp 1698431365
transform 1 0 33376 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_297
timestamp 1698431365
transform 1 0 34608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_299
timestamp 1698431365
transform 1 0 34832 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_312
timestamp 1698431365
transform 1 0 36288 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_356
timestamp 1698431365
transform 1 0 41216 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_373
timestamp 1698431365
transform 1 0 43120 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_377
timestamp 1698431365
transform 1 0 43568 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_380
timestamp 1698431365
transform 1 0 43904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_384
timestamp 1698431365
transform 1 0 44352 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_392
timestamp 1698431365
transform 1 0 45248 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_399
timestamp 1698431365
transform 1 0 46032 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_401
timestamp 1698431365
transform 1 0 46256 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_406
timestamp 1698431365
transform 1 0 46816 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_414
timestamp 1698431365
transform 1 0 47712 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_418
timestamp 1698431365
transform 1 0 48160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_451
timestamp 1698431365
transform 1 0 51856 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_453
timestamp 1698431365
transform 1 0 52080 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_496
timestamp 1698431365
transform 1 0 56896 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_504
timestamp 1698431365
transform 1 0 57792 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_508
timestamp 1698431365
transform 1 0 58240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_28
timestamp 1698431365
transform 1 0 4480 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_32
timestamp 1698431365
transform 1 0 4928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_48
timestamp 1698431365
transform 1 0 6720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_87
timestamp 1698431365
transform 1 0 11088 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_136
timestamp 1698431365
transform 1 0 16576 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_144
timestamp 1698431365
transform 1 0 17472 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_160
timestamp 1698431365
transform 1 0 19264 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_168
timestamp 1698431365
transform 1 0 20160 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_172
timestamp 1698431365
transform 1 0 20608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698431365
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_206
timestamp 1698431365
transform 1 0 24416 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_251
timestamp 1698431365
transform 1 0 29456 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_259
timestamp 1698431365
transform 1 0 30352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_263
timestamp 1698431365
transform 1 0 30800 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_280
timestamp 1698431365
transform 1 0 32704 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_304
timestamp 1698431365
transform 1 0 35392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_306
timestamp 1698431365
transform 1 0 35616 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_313
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_325
timestamp 1698431365
transform 1 0 37744 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_329
timestamp 1698431365
transform 1 0 38192 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_333
timestamp 1698431365
transform 1 0 38640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_337
timestamp 1698431365
transform 1 0 39088 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_353
timestamp 1698431365
transform 1 0 40880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_355
timestamp 1698431365
transform 1 0 41104 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_399
timestamp 1698431365
transform 1 0 46032 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_415
timestamp 1698431365
transform 1 0 47824 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_423
timestamp 1698431365
transform 1 0 48720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_427
timestamp 1698431365
transform 1 0 49168 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_435
timestamp 1698431365
transform 1 0 50064 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_439
timestamp 1698431365
transform 1 0 50512 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_443
timestamp 1698431365
transform 1 0 50960 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_461
timestamp 1698431365
transform 1 0 52976 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_491
timestamp 1698431365
transform 1 0 56336 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_495
timestamp 1698431365
transform 1 0 56784 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_503
timestamp 1698431365
transform 1 0 57680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_507
timestamp 1698431365
transform 1 0 58128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_8
timestamp 1698431365
transform 1 0 2240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_12
timestamp 1698431365
transform 1 0 2688 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_20
timestamp 1698431365
transform 1 0 3584 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_24
timestamp 1698431365
transform 1 0 4032 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_26
timestamp 1698431365
transform 1 0 4256 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_67
timestamp 1698431365
transform 1 0 8848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_69
timestamp 1698431365
transform 1 0 9072 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_150
timestamp 1698431365
transform 1 0 18144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_164
timestamp 1698431365
transform 1 0 19712 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_172
timestamp 1698431365
transform 1 0 20608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_174
timestamp 1698431365
transform 1 0 20832 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_231
timestamp 1698431365
transform 1 0 27216 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_235
timestamp 1698431365
transform 1 0 27664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_239
timestamp 1698431365
transform 1 0 28112 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_243
timestamp 1698431365
transform 1 0 28560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_247
timestamp 1698431365
transform 1 0 29008 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_251
timestamp 1698431365
transform 1 0 29456 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_268
timestamp 1698431365
transform 1 0 31360 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_286
timestamp 1698431365
transform 1 0 33376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_317
timestamp 1698431365
transform 1 0 36848 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_323
timestamp 1698431365
transform 1 0 37520 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_330
timestamp 1698431365
transform 1 0 38304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_361
timestamp 1698431365
transform 1 0 41776 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_365
timestamp 1698431365
transform 1 0 42224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_367
timestamp 1698431365
transform 1 0 42448 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_419
timestamp 1698431365
transform 1 0 48272 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_426
timestamp 1698431365
transform 1 0 49056 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_456
timestamp 1698431365
transform 1 0 52416 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_486
timestamp 1698431365
transform 1 0 55776 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_500
timestamp 1698431365
transform 1 0 57344 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_14
timestamp 1698431365
transform 1 0 2912 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_18
timestamp 1698431365
transform 1 0 3360 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_78
timestamp 1698431365
transform 1 0 10080 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_134
timestamp 1698431365
transform 1 0 16352 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_138
timestamp 1698431365
transform 1 0 16800 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_146
timestamp 1698431365
transform 1 0 17696 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_150
timestamp 1698431365
transform 1 0 18144 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_166
timestamp 1698431365
transform 1 0 19936 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_170
timestamp 1698431365
transform 1 0 20384 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_183
timestamp 1698431365
transform 1 0 21840 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_209
timestamp 1698431365
transform 1 0 24752 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_213
timestamp 1698431365
transform 1 0 25200 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_215
timestamp 1698431365
transform 1 0 25424 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_249
timestamp 1698431365
transform 1 0 29232 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_258
timestamp 1698431365
transform 1 0 30240 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_289
timestamp 1698431365
transform 1 0 33712 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_291
timestamp 1698431365
transform 1 0 33936 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_300
timestamp 1698431365
transform 1 0 34944 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_304
timestamp 1698431365
transform 1 0 35392 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_307
timestamp 1698431365
transform 1 0 35728 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_362
timestamp 1698431365
transform 1 0 41888 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_383
timestamp 1698431365
transform 1 0 44240 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_389
timestamp 1698431365
transform 1 0 44912 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_395
timestamp 1698431365
transform 1 0 45584 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_399
timestamp 1698431365
transform 1 0 46032 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_407
timestamp 1698431365
transform 1 0 46928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_409
timestamp 1698431365
transform 1 0 47152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_447
timestamp 1698431365
transform 1 0 51408 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_451
timestamp 1698431365
transform 1 0 51856 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_8
timestamp 1698431365
transform 1 0 2240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_12
timestamp 1698431365
transform 1 0 2688 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_16
timestamp 1698431365
transform 1 0 3136 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_20
timestamp 1698431365
transform 1 0 3584 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_56
timestamp 1698431365
transform 1 0 7616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_58
timestamp 1698431365
transform 1 0 7840 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_68
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_76
timestamp 1698431365
transform 1 0 9856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_78
timestamp 1698431365
transform 1 0 10080 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_85
timestamp 1698431365
transform 1 0 10864 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_92
timestamp 1698431365
transform 1 0 11648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_104
timestamp 1698431365
transform 1 0 12992 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_106
timestamp 1698431365
transform 1 0 13216 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_113
timestamp 1698431365
transform 1 0 14000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_117
timestamp 1698431365
transform 1 0 14448 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_119
timestamp 1698431365
transform 1 0 14672 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_122
timestamp 1698431365
transform 1 0 15008 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_186
timestamp 1698431365
transform 1 0 22176 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_188
timestamp 1698431365
transform 1 0 22400 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_202
timestamp 1698431365
transform 1 0 23968 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_216
timestamp 1698431365
transform 1 0 25536 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_230
timestamp 1698431365
transform 1 0 27104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_234
timestamp 1698431365
transform 1 0 27552 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_242
timestamp 1698431365
transform 1 0 28448 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_252
timestamp 1698431365
transform 1 0 29568 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_256
timestamp 1698431365
transform 1 0 30016 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_275
timestamp 1698431365
transform 1 0 32144 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_286
timestamp 1698431365
transform 1 0 33376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_288
timestamp 1698431365
transform 1 0 33600 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_291
timestamp 1698431365
transform 1 0 33936 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_295
timestamp 1698431365
transform 1 0 34384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_297
timestamp 1698431365
transform 1 0 34608 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_329
timestamp 1698431365
transform 1 0 38192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_333
timestamp 1698431365
transform 1 0 38640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_337
timestamp 1698431365
transform 1 0 39088 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_346
timestamp 1698431365
transform 1 0 40096 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_354
timestamp 1698431365
transform 1 0 40992 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_361
timestamp 1698431365
transform 1 0 41776 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_394
timestamp 1698431365
transform 1 0 45472 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_401
timestamp 1698431365
transform 1 0 46256 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_405
timestamp 1698431365
transform 1 0 46704 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_409
timestamp 1698431365
transform 1 0 47152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_411
timestamp 1698431365
transform 1 0 47376 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698431365
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_424
timestamp 1698431365
transform 1 0 48832 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_433
timestamp 1698431365
transform 1 0 49840 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_441
timestamp 1698431365
transform 1 0 50736 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_8
timestamp 1698431365
transform 1 0 2240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_12
timestamp 1698431365
transform 1 0 2688 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_16
timestamp 1698431365
transform 1 0 3136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_25
timestamp 1698431365
transform 1 0 4144 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_33
timestamp 1698431365
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_45
timestamp 1698431365
transform 1 0 6384 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_69
timestamp 1698431365
transform 1 0 9072 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_77
timestamp 1698431365
transform 1 0 9968 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_83
timestamp 1698431365
transform 1 0 10640 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_97
timestamp 1698431365
transform 1 0 12208 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_113
timestamp 1698431365
transform 1 0 14000 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_121
timestamp 1698431365
transform 1 0 14896 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_128
timestamp 1698431365
transform 1 0 15680 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_144
timestamp 1698431365
transform 1 0 17472 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_164
timestamp 1698431365
transform 1 0 19712 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_166
timestamp 1698431365
transform 1 0 19936 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_181
timestamp 1698431365
transform 1 0 21616 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_184
timestamp 1698431365
transform 1 0 21952 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_195
timestamp 1698431365
transform 1 0 23184 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_219
timestamp 1698431365
transform 1 0 25872 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_221
timestamp 1698431365
transform 1 0 26096 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_230
timestamp 1698431365
transform 1 0 27104 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_243
timestamp 1698431365
transform 1 0 28560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_251
timestamp 1698431365
transform 1 0 29456 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_255
timestamp 1698431365
transform 1 0 29904 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_257
timestamp 1698431365
transform 1 0 30128 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_264
timestamp 1698431365
transform 1 0 30912 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_268
timestamp 1698431365
transform 1 0 31360 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_282
timestamp 1698431365
transform 1 0 32928 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_286
timestamp 1698431365
transform 1 0 33376 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_300
timestamp 1698431365
transform 1 0 34944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_310
timestamp 1698431365
transform 1 0 36064 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_314
timestamp 1698431365
transform 1 0 36512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_325
timestamp 1698431365
transform 1 0 37744 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_329
timestamp 1698431365
transform 1 0 38192 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_350
timestamp 1698431365
transform 1 0 40544 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_358
timestamp 1698431365
transform 1 0 41440 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_362
timestamp 1698431365
transform 1 0 41888 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_372
timestamp 1698431365
transform 1 0 43008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_374
timestamp 1698431365
transform 1 0 43232 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_377
timestamp 1698431365
transform 1 0 43568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_391
timestamp 1698431365
transform 1 0 45136 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_404
timestamp 1698431365
transform 1 0 46592 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_408
timestamp 1698431365
transform 1 0 47040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_418
timestamp 1698431365
transform 1 0 48160 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_422
timestamp 1698431365
transform 1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_431
timestamp 1698431365
transform 1 0 49616 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_435
timestamp 1698431365
transform 1 0 50064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_437
timestamp 1698431365
transform 1 0 50288 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_8
timestamp 1698431365
transform 1 0 2240 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_12
timestamp 1698431365
transform 1 0 2688 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_67
timestamp 1698431365
transform 1 0 8848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_74
timestamp 1698431365
transform 1 0 9632 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_110
timestamp 1698431365
transform 1 0 13664 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_149
timestamp 1698431365
transform 1 0 18032 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_157
timestamp 1698431365
transform 1 0 18928 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_181
timestamp 1698431365
transform 1 0 21616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_185
timestamp 1698431365
transform 1 0 22064 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_207
timestamp 1698431365
transform 1 0 24528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_214
timestamp 1698431365
transform 1 0 25312 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_236
timestamp 1698431365
transform 1 0 27776 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_259
timestamp 1698431365
transform 1 0 30352 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_275
timestamp 1698431365
transform 1 0 32144 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_290
timestamp 1698431365
transform 1 0 33824 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_327
timestamp 1698431365
transform 1 0 37968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_349
timestamp 1698431365
transform 1 0 40432 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_356
timestamp 1698431365
transform 1 0 41216 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_360
timestamp 1698431365
transform 1 0 41664 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_377
timestamp 1698431365
transform 1 0 43568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_381
timestamp 1698431365
transform 1 0 44016 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_389
timestamp 1698431365
transform 1 0 44912 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_393
timestamp 1698431365
transform 1 0 45360 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_427
timestamp 1698431365
transform 1 0 49168 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1698431365
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_28
timestamp 1698431365
transform 1 0 4480 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_32
timestamp 1698431365
transform 1 0 4928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_53
timestamp 1698431365
transform 1 0 7280 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_57
timestamp 1698431365
transform 1 0 7728 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_88
timestamp 1698431365
transform 1 0 11200 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_92
timestamp 1698431365
transform 1 0 11648 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_96
timestamp 1698431365
transform 1 0 12096 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_119
timestamp 1698431365
transform 1 0 14672 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_135
timestamp 1698431365
transform 1 0 16464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_139
timestamp 1698431365
transform 1 0 16912 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_147
timestamp 1698431365
transform 1 0 17808 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_159
timestamp 1698431365
transform 1 0 19152 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_163
timestamp 1698431365
transform 1 0 19600 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_167
timestamp 1698431365
transform 1 0 20048 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_205
timestamp 1698431365
transform 1 0 24304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_209
timestamp 1698431365
transform 1 0 24752 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_213
timestamp 1698431365
transform 1 0 25200 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_215
timestamp 1698431365
transform 1 0 25424 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_226
timestamp 1698431365
transform 1 0 26656 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_240
timestamp 1698431365
transform 1 0 28224 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_244
timestamp 1698431365
transform 1 0 28672 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_276
timestamp 1698431365
transform 1 0 32256 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_308
timestamp 1698431365
transform 1 0 35840 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_312
timestamp 1698431365
transform 1 0 36288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_325
timestamp 1698431365
transform 1 0 37744 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_327
timestamp 1698431365
transform 1 0 37968 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_346
timestamp 1698431365
transform 1 0 40096 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_354
timestamp 1698431365
transform 1 0 40992 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_356
timestamp 1698431365
transform 1 0 41216 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_362
timestamp 1698431365
transform 1 0 41888 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_366
timestamp 1698431365
transform 1 0 42336 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_368
timestamp 1698431365
transform 1 0 42560 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_381
timestamp 1698431365
transform 1 0 44016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_391
timestamp 1698431365
transform 1 0 45136 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_418
timestamp 1698431365
transform 1 0 48160 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_435
timestamp 1698431365
transform 1 0 50064 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_8
timestamp 1698431365
transform 1 0 2240 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_12
timestamp 1698431365
transform 1 0 2688 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_44
timestamp 1698431365
transform 1 0 6272 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_60
timestamp 1698431365
transform 1 0 8064 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_68
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_77
timestamp 1698431365
transform 1 0 9968 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_127
timestamp 1698431365
transform 1 0 15568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_131
timestamp 1698431365
transform 1 0 16016 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_138
timestamp 1698431365
transform 1 0 16800 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_177
timestamp 1698431365
transform 1 0 21168 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_216
timestamp 1698431365
transform 1 0 25536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_224
timestamp 1698431365
transform 1 0 26432 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_234
timestamp 1698431365
transform 1 0 27552 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_242
timestamp 1698431365
transform 1 0 28448 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_246
timestamp 1698431365
transform 1 0 28896 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_248
timestamp 1698431365
transform 1 0 29120 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_263
timestamp 1698431365
transform 1 0 30800 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_276
timestamp 1698431365
transform 1 0 32256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_299
timestamp 1698431365
transform 1 0 34832 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_303
timestamp 1698431365
transform 1 0 35280 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_305
timestamp 1698431365
transform 1 0 35504 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_314
timestamp 1698431365
transform 1 0 36512 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_316
timestamp 1698431365
transform 1 0 36736 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_337
timestamp 1698431365
transform 1 0 39088 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_345
timestamp 1698431365
transform 1 0 39984 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_349
timestamp 1698431365
transform 1 0 40432 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_354
timestamp 1698431365
transform 1 0 40992 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_367
timestamp 1698431365
transform 1 0 42448 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_394
timestamp 1698431365
transform 1 0 45472 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_402
timestamp 1698431365
transform 1 0 46368 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_406
timestamp 1698431365
transform 1 0 46816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_438
timestamp 1698431365
transform 1 0 50400 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_481
timestamp 1698431365
transform 1 0 55216 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_485
timestamp 1698431365
transform 1 0 55664 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_489
timestamp 1698431365
transform 1 0 56112 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698431365
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_14
timestamp 1698431365
transform 1 0 2912 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_18
timestamp 1698431365
transform 1 0 3360 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_53
timestamp 1698431365
transform 1 0 7280 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_99
timestamp 1698431365
transform 1 0 12432 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_130
timestamp 1698431365
transform 1 0 15904 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_146
timestamp 1698431365
transform 1 0 17696 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_153
timestamp 1698431365
transform 1 0 18480 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_161
timestamp 1698431365
transform 1 0 19376 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_228
timestamp 1698431365
transform 1 0 26880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_232
timestamp 1698431365
transform 1 0 27328 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_236
timestamp 1698431365
transform 1 0 27776 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_251
timestamp 1698431365
transform 1 0 29456 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_267
timestamp 1698431365
transform 1 0 31248 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_269
timestamp 1698431365
transform 1 0 31472 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_306
timestamp 1698431365
transform 1 0 35616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_310
timestamp 1698431365
transform 1 0 36064 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_314
timestamp 1698431365
transform 1 0 36512 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_325
timestamp 1698431365
transform 1 0 37744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_329
timestamp 1698431365
transform 1 0 38192 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_337
timestamp 1698431365
transform 1 0 39088 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_339
timestamp 1698431365
transform 1 0 39312 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_362
timestamp 1698431365
transform 1 0 41888 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_366
timestamp 1698431365
transform 1 0 42336 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_374
timestamp 1698431365
transform 1 0 43232 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_381
timestamp 1698431365
transform 1 0 44016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_399
timestamp 1698431365
transform 1 0 46032 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_407
timestamp 1698431365
transform 1 0 46928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_425
timestamp 1698431365
transform 1 0 48944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_429
timestamp 1698431365
transform 1 0 49392 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_439
timestamp 1698431365
transform 1 0 50512 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_447
timestamp 1698431365
transform 1 0 51408 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_449
timestamp 1698431365
transform 1 0 51632 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_8
timestamp 1698431365
transform 1 0 2240 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_12
timestamp 1698431365
transform 1 0 2688 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_16
timestamp 1698431365
transform 1 0 3136 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_48
timestamp 1698431365
transform 1 0 6720 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_64
timestamp 1698431365
transform 1 0 8512 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_68
timestamp 1698431365
transform 1 0 8960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_78
timestamp 1698431365
transform 1 0 10080 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_82
timestamp 1698431365
transform 1 0 10528 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_88
timestamp 1698431365
transform 1 0 11200 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_98
timestamp 1698431365
transform 1 0 12320 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_102
timestamp 1698431365
transform 1 0 12768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_139
timestamp 1698431365
transform 1 0 16912 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_150
timestamp 1698431365
transform 1 0 18144 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_158
timestamp 1698431365
transform 1 0 19040 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_162
timestamp 1698431365
transform 1 0 19488 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_204
timestamp 1698431365
transform 1 0 24192 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_208
timestamp 1698431365
transform 1 0 24640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_261
timestamp 1698431365
transform 1 0 30576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_265
timestamp 1698431365
transform 1 0 31024 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_269
timestamp 1698431365
transform 1 0 31472 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_271
timestamp 1698431365
transform 1 0 31696 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_279
timestamp 1698431365
transform 1 0 32592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_286
timestamp 1698431365
transform 1 0 33376 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_294
timestamp 1698431365
transform 1 0 34272 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_298
timestamp 1698431365
transform 1 0 34720 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_307
timestamp 1698431365
transform 1 0 35728 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_309
timestamp 1698431365
transform 1 0 35952 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_347
timestamp 1698431365
transform 1 0 40208 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_349
timestamp 1698431365
transform 1 0 40432 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_369
timestamp 1698431365
transform 1 0 42672 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_377
timestamp 1698431365
transform 1 0 43568 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_387
timestamp 1698431365
transform 1 0 44688 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_418
timestamp 1698431365
transform 1 0 48160 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_434
timestamp 1698431365
transform 1 0 49952 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_467
timestamp 1698431365
transform 1 0 53648 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_471
timestamp 1698431365
transform 1 0 54096 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_487
timestamp 1698431365
transform 1 0 55888 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_489
timestamp 1698431365
transform 1 0 56112 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_508
timestamp 1698431365
transform 1 0 58240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_8
timestamp 1698431365
transform 1 0 2240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_12
timestamp 1698431365
transform 1 0 2688 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_28
timestamp 1698431365
transform 1 0 4480 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_32
timestamp 1698431365
transform 1 0 4928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_69
timestamp 1698431365
transform 1 0 9072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_71
timestamp 1698431365
transform 1 0 9296 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_101
timestamp 1698431365
transform 1 0 12656 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_123
timestamp 1698431365
transform 1 0 15120 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_131
timestamp 1698431365
transform 1 0 16016 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_174
timestamp 1698431365
transform 1 0 20832 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_183
timestamp 1698431365
transform 1 0 21840 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_187
timestamp 1698431365
transform 1 0 22288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_232
timestamp 1698431365
transform 1 0 27328 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_242
timestamp 1698431365
transform 1 0 28448 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_244
timestamp 1698431365
transform 1 0 28672 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_252
timestamp 1698431365
transform 1 0 29568 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_288
timestamp 1698431365
transform 1 0 33600 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_290
timestamp 1698431365
transform 1 0 33824 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_305
timestamp 1698431365
transform 1 0 35504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_353
timestamp 1698431365
transform 1 0 40880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_355
timestamp 1698431365
transform 1 0 41104 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_391
timestamp 1698431365
transform 1 0 45136 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_395
timestamp 1698431365
transform 1 0 45584 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_402
timestamp 1698431365
transform 1 0 46368 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_404
timestamp 1698431365
transform 1 0 46592 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_434
timestamp 1698431365
transform 1 0 49952 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_438
timestamp 1698431365
transform 1 0 50400 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_457
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_473
timestamp 1698431365
transform 1 0 54320 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_8
timestamp 1698431365
transform 1 0 2240 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_12
timestamp 1698431365
transform 1 0 2688 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_44
timestamp 1698431365
transform 1 0 6272 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_60
timestamp 1698431365
transform 1 0 8064 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_68
timestamp 1698431365
transform 1 0 8960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_88
timestamp 1698431365
transform 1 0 11200 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_101
timestamp 1698431365
transform 1 0 12656 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_105
timestamp 1698431365
transform 1 0 13104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_109
timestamp 1698431365
transform 1 0 13552 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_150
timestamp 1698431365
transform 1 0 18144 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_158
timestamp 1698431365
transform 1 0 19040 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_160
timestamp 1698431365
transform 1 0 19264 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_190
timestamp 1698431365
transform 1 0 22624 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_206
timestamp 1698431365
transform 1 0 24416 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_220
timestamp 1698431365
transform 1 0 25984 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_228
timestamp 1698431365
transform 1 0 26880 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_267
timestamp 1698431365
transform 1 0 31248 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_312
timestamp 1698431365
transform 1 0 36288 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_332
timestamp 1698431365
transform 1 0 38528 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_336
timestamp 1698431365
transform 1 0 38976 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_346
timestamp 1698431365
transform 1 0 40096 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_374
timestamp 1698431365
transform 1 0 43232 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_382
timestamp 1698431365
transform 1 0 44128 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_390
timestamp 1698431365
transform 1 0 45024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_392
timestamp 1698431365
transform 1 0 45248 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_401
timestamp 1698431365
transform 1 0 46256 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_416
timestamp 1698431365
transform 1 0 47936 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_460
timestamp 1698431365
transform 1 0 52864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_464
timestamp 1698431365
transform 1 0 53312 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_480
timestamp 1698431365
transform 1 0 55104 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_488
timestamp 1698431365
transform 1 0 56000 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698431365
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_8
timestamp 1698431365
transform 1 0 2240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_12
timestamp 1698431365
transform 1 0 2688 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_28
timestamp 1698431365
transform 1 0 4480 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_32
timestamp 1698431365
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_69
timestamp 1698431365
transform 1 0 9072 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_73
timestamp 1698431365
transform 1 0 9520 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_75
timestamp 1698431365
transform 1 0 9744 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_111
timestamp 1698431365
transform 1 0 13776 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_126
timestamp 1698431365
transform 1 0 15456 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_130
timestamp 1698431365
transform 1 0 15904 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_134
timestamp 1698431365
transform 1 0 16352 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_136
timestamp 1698431365
transform 1 0 16576 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_145
timestamp 1698431365
transform 1 0 17584 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_161
timestamp 1698431365
transform 1 0 19376 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_169
timestamp 1698431365
transform 1 0 20272 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_173
timestamp 1698431365
transform 1 0 20720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_185
timestamp 1698431365
transform 1 0 22064 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_187
timestamp 1698431365
transform 1 0 22288 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_194
timestamp 1698431365
transform 1 0 23072 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_231
timestamp 1698431365
transform 1 0 27216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_235
timestamp 1698431365
transform 1 0 27664 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_243
timestamp 1698431365
transform 1 0 28560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_251
timestamp 1698431365
transform 1 0 29456 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_255
timestamp 1698431365
transform 1 0 29904 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_257
timestamp 1698431365
transform 1 0 30128 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_266
timestamp 1698431365
transform 1 0 31136 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_270
timestamp 1698431365
transform 1 0 31584 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_274
timestamp 1698431365
transform 1 0 32032 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_276
timestamp 1698431365
transform 1 0 32256 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_303
timestamp 1698431365
transform 1 0 35280 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_307
timestamp 1698431365
transform 1 0 35728 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_311
timestamp 1698431365
transform 1 0 36176 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_314
timestamp 1698431365
transform 1 0 36512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_321
timestamp 1698431365
transform 1 0 37296 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_325
timestamp 1698431365
transform 1 0 37744 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_327
timestamp 1698431365
transform 1 0 37968 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_360
timestamp 1698431365
transform 1 0 41664 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_364
timestamp 1698431365
transform 1 0 42112 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_379
timestamp 1698431365
transform 1 0 43792 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_383
timestamp 1698431365
transform 1 0 44240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_393
timestamp 1698431365
transform 1 0 45360 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_401
timestamp 1698431365
transform 1 0 46256 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_405
timestamp 1698431365
transform 1 0 46704 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_444
timestamp 1698431365
transform 1 0 51072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_448
timestamp 1698431365
transform 1 0 51520 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_452
timestamp 1698431365
transform 1 0 51968 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_454
timestamp 1698431365
transform 1 0 52192 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_486
timestamp 1698431365
transform 1 0 55776 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_502
timestamp 1698431365
transform 1 0 57568 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_506
timestamp 1698431365
transform 1 0 58016 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_508
timestamp 1698431365
transform 1 0 58240 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_8
timestamp 1698431365
transform 1 0 2240 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_12
timestamp 1698431365
transform 1 0 2688 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_44
timestamp 1698431365
transform 1 0 6272 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_60
timestamp 1698431365
transform 1 0 8064 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_68
timestamp 1698431365
transform 1 0 8960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_88
timestamp 1698431365
transform 1 0 11200 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_93
timestamp 1698431365
transform 1 0 11760 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_130
timestamp 1698431365
transform 1 0 15904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_150
timestamp 1698431365
transform 1 0 18144 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_154
timestamp 1698431365
transform 1 0 18592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_160
timestamp 1698431365
transform 1 0 19264 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_175
timestamp 1698431365
transform 1 0 20944 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_179
timestamp 1698431365
transform 1 0 21392 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_186
timestamp 1698431365
transform 1 0 22176 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_200
timestamp 1698431365
transform 1 0 23744 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_238
timestamp 1698431365
transform 1 0 28000 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_242
timestamp 1698431365
transform 1 0 28448 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_244
timestamp 1698431365
transform 1 0 28672 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_253
timestamp 1698431365
transform 1 0 29680 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_255
timestamp 1698431365
transform 1 0 29904 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_262
timestamp 1698431365
transform 1 0 30688 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_270
timestamp 1698431365
transform 1 0 31584 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_300
timestamp 1698431365
transform 1 0 34944 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_304
timestamp 1698431365
transform 1 0 35392 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_306
timestamp 1698431365
transform 1 0 35616 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_320
timestamp 1698431365
transform 1 0 37184 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_356
timestamp 1698431365
transform 1 0 41216 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_387
timestamp 1698431365
transform 1 0 44688 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_430
timestamp 1698431365
transform 1 0 49504 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_480
timestamp 1698431365
transform 1 0 55104 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_488
timestamp 1698431365
transform 1 0 56000 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_508
timestamp 1698431365
transform 1 0 58240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_28
timestamp 1698431365
transform 1 0 4480 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_32
timestamp 1698431365
transform 1 0 4928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_112
timestamp 1698431365
transform 1 0 13888 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_122
timestamp 1698431365
transform 1 0 15008 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_135
timestamp 1698431365
transform 1 0 16464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_137
timestamp 1698431365
transform 1 0 16688 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_151
timestamp 1698431365
transform 1 0 18256 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_166
timestamp 1698431365
transform 1 0 19936 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_174
timestamp 1698431365
transform 1 0 20832 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_237
timestamp 1698431365
transform 1 0 27888 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_276
timestamp 1698431365
transform 1 0 32256 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_360
timestamp 1698431365
transform 1 0 41664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_370
timestamp 1698431365
transform 1 0 42784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_374
timestamp 1698431365
transform 1 0 43232 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_382
timestamp 1698431365
transform 1 0 44128 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1698431365
transform 1 0 44352 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_454
timestamp 1698431365
transform 1 0 52192 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_486
timestamp 1698431365
transform 1 0 55776 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_502
timestamp 1698431365
transform 1 0 57568 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_506
timestamp 1698431365
transform 1 0 58016 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_508
timestamp 1698431365
transform 1 0 58240 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_66
timestamp 1698431365
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_104
timestamp 1698431365
transform 1 0 12992 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_112
timestamp 1698431365
transform 1 0 13888 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_120
timestamp 1698431365
transform 1 0 14784 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_137
timestamp 1698431365
transform 1 0 16688 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_139
timestamp 1698431365
transform 1 0 16912 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_173
timestamp 1698431365
transform 1 0 20720 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_181
timestamp 1698431365
transform 1 0 21616 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_191
timestamp 1698431365
transform 1 0 22736 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_201
timestamp 1698431365
transform 1 0 23856 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_209
timestamp 1698431365
transform 1 0 24752 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_214
timestamp 1698431365
transform 1 0 25312 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_246
timestamp 1698431365
transform 1 0 28896 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_250
timestamp 1698431365
transform 1 0 29344 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_288
timestamp 1698431365
transform 1 0 33600 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_347
timestamp 1698431365
transform 1 0 40208 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_349
timestamp 1698431365
transform 1 0 40432 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_384
timestamp 1698431365
transform 1 0 44352 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_388
timestamp 1698431365
transform 1 0 44800 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_395
timestamp 1698431365
transform 1 0 45584 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_411
timestamp 1698431365
transform 1 0 47376 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_419
timestamp 1698431365
transform 1 0 48272 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_422
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_471
timestamp 1698431365
transform 1 0 54096 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_487
timestamp 1698431365
transform 1 0 55888 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_489
timestamp 1698431365
transform 1 0 56112 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1698431365
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698431365
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_136
timestamp 1698431365
transform 1 0 16576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_140
timestamp 1698431365
transform 1 0 17024 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_144
timestamp 1698431365
transform 1 0 17472 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_161
timestamp 1698431365
transform 1 0 19376 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_181
timestamp 1698431365
transform 1 0 21616 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_190
timestamp 1698431365
transform 1 0 22624 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_198
timestamp 1698431365
transform 1 0 23520 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_202
timestamp 1698431365
transform 1 0 23968 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_210
timestamp 1698431365
transform 1 0 24864 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_243
timestamp 1698431365
transform 1 0 28560 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_249
timestamp 1698431365
transform 1 0 29232 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_319
timestamp 1698431365
transform 1 0 37072 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_363
timestamp 1698431365
transform 1 0 42000 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_379
timestamp 1698431365
transform 1 0 43792 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_383
timestamp 1698431365
transform 1 0 44240 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_393
timestamp 1698431365
transform 1 0 45360 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_401
timestamp 1698431365
transform 1 0 46256 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_403
timestamp 1698431365
transform 1 0 46480 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_406
timestamp 1698431365
transform 1 0 46816 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_424
timestamp 1698431365
transform 1 0 48832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_426
timestamp 1698431365
transform 1 0 49056 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_429
timestamp 1698431365
transform 1 0 49392 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_449
timestamp 1698431365
transform 1 0 51632 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_453
timestamp 1698431365
transform 1 0 52080 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_461
timestamp 1698431365
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_465
timestamp 1698431365
transform 1 0 53424 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_497
timestamp 1698431365
transform 1 0 57008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_505
timestamp 1698431365
transform 1 0 57904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1698431365
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_104
timestamp 1698431365
transform 1 0 12992 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_120
timestamp 1698431365
transform 1 0 14784 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_124
timestamp 1698431365
transform 1 0 15232 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_129
timestamp 1698431365
transform 1 0 15792 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_137
timestamp 1698431365
transform 1 0 16688 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_139
timestamp 1698431365
transform 1 0 16912 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_148
timestamp 1698431365
transform 1 0 17920 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_152
timestamp 1698431365
transform 1 0 18368 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_156
timestamp 1698431365
transform 1 0 18816 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_160
timestamp 1698431365
transform 1 0 19264 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_166
timestamp 1698431365
transform 1 0 19936 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_170
timestamp 1698431365
transform 1 0 20384 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_200
timestamp 1698431365
transform 1 0 23744 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_221
timestamp 1698431365
transform 1 0 26096 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_225
timestamp 1698431365
transform 1 0 26544 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_255
timestamp 1698431365
transform 1 0 29904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_265
timestamp 1698431365
transform 1 0 31024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_267
timestamp 1698431365
transform 1 0 31248 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_276
timestamp 1698431365
transform 1 0 32256 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_334
timestamp 1698431365
transform 1 0 38752 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_336
timestamp 1698431365
transform 1 0 38976 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_345
timestamp 1698431365
transform 1 0 39984 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_349
timestamp 1698431365
transform 1 0 40432 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_356
timestamp 1698431365
transform 1 0 41216 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_416
timestamp 1698431365
transform 1 0 47936 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_428
timestamp 1698431365
transform 1 0 49280 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_432
timestamp 1698431365
transform 1 0 49728 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_436
timestamp 1698431365
transform 1 0 50176 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_440
timestamp 1698431365
transform 1 0 50624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_477
timestamp 1698431365
transform 1 0 54768 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_485
timestamp 1698431365
transform 1 0 55664 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_489
timestamp 1698431365
transform 1 0 56112 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_508
timestamp 1698431365
transform 1 0 58240 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698431365
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_109
timestamp 1698431365
transform 1 0 13552 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_172
timestamp 1698431365
transform 1 0 20608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_174
timestamp 1698431365
transform 1 0 20832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_179
timestamp 1698431365
transform 1 0 21392 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_182
timestamp 1698431365
transform 1 0 21728 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_227
timestamp 1698431365
transform 1 0 26768 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_229
timestamp 1698431365
transform 1 0 26992 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_243
timestamp 1698431365
transform 1 0 28560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_256
timestamp 1698431365
transform 1 0 30016 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_321
timestamp 1698431365
transform 1 0 37296 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_331
timestamp 1698431365
transform 1 0 38416 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_391
timestamp 1698431365
transform 1 0 45136 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_393
timestamp 1698431365
transform 1 0 45360 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_423
timestamp 1698431365
transform 1 0 48720 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_427
timestamp 1698431365
transform 1 0 49168 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_450
timestamp 1698431365
transform 1 0 51744 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_454
timestamp 1698431365
transform 1 0 52192 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_489
timestamp 1698431365
transform 1 0 56112 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_505
timestamp 1698431365
transform 1 0 57904 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_232
timestamp 1698431365
transform 1 0 27328 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_262
timestamp 1698431365
transform 1 0 30688 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_272
timestamp 1698431365
transform 1 0 31808 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_296
timestamp 1698431365
transform 1 0 34496 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_348
timestamp 1698431365
transform 1 0 40320 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_365
timestamp 1698431365
transform 1 0 42224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_426
timestamp 1698431365
transform 1 0 49056 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_431
timestamp 1698431365
transform 1 0 49616 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_464
timestamp 1698431365
transform 1 0 53312 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_468
timestamp 1698431365
transform 1 0 53760 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_484
timestamp 1698431365
transform 1 0 55552 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_488
timestamp 1698431365
transform 1 0 56000 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698431365
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_115
timestamp 1698431365
transform 1 0 14224 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_193
timestamp 1698431365
transform 1 0 22960 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_195
timestamp 1698431365
transform 1 0 23184 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_225
timestamp 1698431365
transform 1 0 26544 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_233
timestamp 1698431365
transform 1 0 27440 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_237
timestamp 1698431365
transform 1 0 27888 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_239
timestamp 1698431365
transform 1 0 28112 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_244
timestamp 1698431365
transform 1 0 28672 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_255
timestamp 1698431365
transform 1 0 29904 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_259
timestamp 1698431365
transform 1 0 30352 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_261
timestamp 1698431365
transform 1 0 30576 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_291
timestamp 1698431365
transform 1 0 33936 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_295
timestamp 1698431365
transform 1 0 34384 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_299
timestamp 1698431365
transform 1 0 34832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_303
timestamp 1698431365
transform 1 0 35280 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_309
timestamp 1698431365
transform 1 0 35952 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_314
timestamp 1698431365
transform 1 0 36512 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_321
timestamp 1698431365
transform 1 0 37296 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_382
timestamp 1698431365
transform 1 0 44128 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_384
timestamp 1698431365
transform 1 0 44352 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_391
timestamp 1698431365
transform 1 0 45136 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_451
timestamp 1698431365
transform 1 0 51856 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_489
timestamp 1698431365
transform 1 0 56112 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_505
timestamp 1698431365
transform 1 0 57904 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_36
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_104
timestamp 1698431365
transform 1 0 12992 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_138
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_142
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_172
timestamp 1698431365
transform 1 0 20608 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_176
timestamp 1698431365
transform 1 0 21056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_210
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_240
timestamp 1698431365
transform 1 0 28224 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_244
timestamp 1698431365
transform 1 0 28672 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_300
timestamp 1698431365
transform 1 0 34944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_304
timestamp 1698431365
transform 1 0 35392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_339
timestamp 1698431365
transform 1 0 39312 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_373
timestamp 1698431365
transform 1 0 43120 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_402
timestamp 1698431365
transform 1 0 46368 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_406
timestamp 1698431365
transform 1 0 46816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_436
timestamp 1698431365
transform 1 0 50176 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_440
timestamp 1698431365
transform 1 0 50624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_444
timestamp 1698431365
transform 1 0 51072 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_478
timestamp 1698431365
transform 1 0 54880 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_494
timestamp 1698431365
transform 1 0 56672 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_502
timestamp 1698431365
transform 1 0 57568 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_506
timestamp 1698431365
transform 1 0 58016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_508
timestamp 1698431365
transform 1 0 58240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 2240 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 2240 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 29680 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input20
timestamp 1698431365
transform -1 0 39088 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 37856 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input22
timestamp 1698431365
transform -1 0 38528 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input23
timestamp 1698431365
transform -1 0 39200 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input24
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 40992 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 57680 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input27
timestamp 1698431365
transform -1 0 58352 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input28
timestamp 1698431365
transform -1 0 57680 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform -1 0 58352 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input30
timestamp 1698431365
transform 1 0 33376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input31
timestamp 1698431365
transform -1 0 58352 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 57680 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input33
timestamp 1698431365
transform -1 0 58352 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 57680 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input35
timestamp 1698431365
transform -1 0 58352 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform -1 0 58352 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform -1 0 58352 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input38
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 2240 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input40
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input41
timestamp 1698431365
transform 1 0 34944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 2240 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698431365
transform 1 0 2240 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input44
timestamp 1698431365
transform 1 0 34272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input45
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform 1 0 32704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input47
timestamp 1698431365
transform 1 0 30352 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform 1 0 31024 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input49
timestamp 1698431365
transform -1 0 36512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform -1 0 37184 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1698431365
transform 1 0 2912 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input52
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input53
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1698431365
transform 1 0 2240 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input58
timestamp 1698431365
transform 1 0 2912 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1698431365
transform 1 0 2240 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input62
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input63
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1698431365
transform 1 0 2240 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input65
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input66
timestamp 1698431365
transform 1 0 2240 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input67
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input68
timestamp 1698431365
transform 1 0 2240 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input69
timestamp 1698431365
transform 1 0 16912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input70
timestamp 1698431365
transform 1 0 17584 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input71
timestamp 1698431365
transform -1 0 18928 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input72
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input73
timestamp 1698431365
transform 1 0 2240 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1698431365
transform 1 0 2240 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input76
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input77
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input78
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input79
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input80
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input81
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input82
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input83
timestamp 1698431365
transform 1 0 2240 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output84 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20384 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output85
timestamp 1698431365
transform -1 0 50176 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output86
timestamp 1698431365
transform 1 0 40768 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output87
timestamp 1698431365
transform 1 0 55440 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output88
timestamp 1698431365
transform 1 0 53312 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output89
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output90
timestamp 1698431365
transform 1 0 53312 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output91
timestamp 1698431365
transform 1 0 55440 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output92
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output93
timestamp 1698431365
transform 1 0 53312 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output94
timestamp 1698431365
transform 1 0 55440 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output95
timestamp 1698431365
transform 1 0 35840 0 -1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output96
timestamp 1698431365
transform -1 0 56224 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output97
timestamp 1698431365
transform -1 0 55440 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output98
timestamp 1698431365
transform 1 0 55440 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output99
timestamp 1698431365
transform 1 0 55440 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output100
timestamp 1698431365
transform 1 0 53312 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output101
timestamp 1698431365
transform 1 0 55440 0 1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output102
timestamp 1698431365
transform 1 0 33712 0 1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output103
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output104
timestamp 1698431365
transform -1 0 24192 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output105
timestamp 1698431365
transform 1 0 30240 0 1 51744
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output106
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output107
timestamp 1698431365
transform -1 0 4480 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output108
timestamp 1698431365
transform -1 0 46368 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output109
timestamp 1698431365
transform 1 0 28896 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output110
timestamp 1698431365
transform -1 0 24864 0 -1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output111
timestamp 1698431365
transform 1 0 25648 0 1 51744
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output112
timestamp 1698431365
transform -1 0 28000 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output113
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output114
timestamp 1698431365
transform 1 0 55440 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output115
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output116
timestamp 1698431365
transform -1 0 4480 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output117
timestamp 1698431365
transform -1 0 4480 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output118
timestamp 1698431365
transform -1 0 4480 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_152
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_153
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_154
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_155
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_156
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_157
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_158
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_159
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_160
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_161
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_162
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_163
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_164
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_165
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_166
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_167
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_168
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_169
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_170
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_171
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_172
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_173
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_174
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_175
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_176
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_177
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_178
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_179
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_180
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_181
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_182
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_183
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_184
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_185
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_186
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_187
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_188
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_189
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_190
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_191
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_192
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_193
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_194
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_195
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_196
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_197
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_198
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_199
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_200
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_201
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_202
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_203
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_204
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_205
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_206
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_207
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_208
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_209
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_210
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_211
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_212
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_213
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_214
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_215
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_216
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_217
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_218
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_219
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_220
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_221
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_222
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_223
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_224
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_225
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_226
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_227
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_228
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_229
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_230
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_231
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_232
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_233
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_234
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_235
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_236
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_237
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_238
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_239
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_240
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_241
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_242
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_243
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_244
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_245
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_246
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_247
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_248
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_249
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_250
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_251
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_252
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_253
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_254
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_258
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_259
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_260
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_261
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_267
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_268
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_276
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_283
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_284
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_285
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_290
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_291
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_292
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_293
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_294
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_295
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_297
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_298
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_299
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_300
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_301
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_302
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_303
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_304
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_305
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_306
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_307
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_308
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_309
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_310
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_311
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_312
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_313
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_314
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_315
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_316
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_317
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_318
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_319
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_320
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_321
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_322
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_323
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_324
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_325
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_326
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_327
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_328
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_329
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_330
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_331
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_332
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_333
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_334
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_335
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_336
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_337
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_338
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_339
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_340
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_341
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_342
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_343
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_344
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_345
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_346
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_347
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_348
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_349
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_350
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_351
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_352
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_353
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_354
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_355
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_356
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_357
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_358
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_360
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_361
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_362
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_363
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_364
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_365
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_367
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_368
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_369
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_370
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_371
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_372
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_374
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_375
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_376
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_377
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_378
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_379
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_381
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_382
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_383
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_384
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_385
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_386
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_387
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_388
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_389
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_390
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_391
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_392
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_393
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_394
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_395
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_396
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_397
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_398
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_399
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_400
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_402
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_403
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_404
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_405
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_406
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_407
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_409
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_410
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_411
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_412
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_416
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_417
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_422
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_427
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_428
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_429
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_431
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_432
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_433
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_434
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_437
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_442
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_445
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_446
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_447
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_448
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_449
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_450
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_451
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_452
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_453
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_454
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_455
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_456
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_457
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_458
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_459
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_460
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_461
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_462
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_463
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_464
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_465
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_466
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_467
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_468
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_469
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_470
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_471
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_472
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_473
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_474
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_475
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_476
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_477
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_478
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_479
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_480
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_481
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_482
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_483
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_484
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_485
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_486
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_487
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_488
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_489
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_490
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_491
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_492
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_493
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_494
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_495
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_496
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_497
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_498
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_499
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_500
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_501
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_502
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_503
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_504
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_505
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_506
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_507
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_508
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_509
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_510
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_511
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_512
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_513
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_514
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_515
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_516
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_517
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_518
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_519
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_520
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_521
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_522
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_523
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_524
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_525
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_526
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_527
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_528
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_529
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_530
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_531
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_532
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_533
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_534
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_535
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_536
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_537
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_538
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_539
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_540
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_541
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_542
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_543
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_544
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_545
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_546
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_547
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_548
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_549
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_550
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_551
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_552
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_553
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_554
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_555
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_556
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_557
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_558
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_559
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_560
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_561
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_562
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_563
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_564
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_565
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_566
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_567
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_568
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_569
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_570
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_571
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_572
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_573
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_574
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_575
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_576
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_577
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_578
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_579
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_580
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_581
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_582
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_583
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_584
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_585
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_586
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_587
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_588
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_589
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_590
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_591
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_592
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_593
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_594
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_595
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_596
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_597
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_598
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_599
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_600
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_601
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_602
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_603
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_604
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_605
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_606
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_607
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_608
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_609
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_610
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_611
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_612
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_613
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_614
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_615
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_616
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_617
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_618
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_619
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_620
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_621
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_622
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_623
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_624
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_625
timestamp 1698431365
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 55104 800 55216 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 20160 59200 20272 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[0]
port 1 nsew signal tristate
flabel metal2 s 38304 59200 38416 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[10]
port 2 nsew signal tristate
flabel metal2 s 36288 59200 36400 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[11]
port 3 nsew signal tristate
flabel metal3 s 59200 34272 60000 34384 0 FreeSans 448 0 0 0 pcpi_div_rd[12]
port 4 nsew signal tristate
flabel metal3 s 59200 39648 60000 39760 0 FreeSans 448 0 0 0 pcpi_div_rd[13]
port 5 nsew signal tristate
flabel metal3 s 59200 44352 60000 44464 0 FreeSans 448 0 0 0 pcpi_div_rd[14]
port 6 nsew signal tristate
flabel metal3 s 59200 41664 60000 41776 0 FreeSans 448 0 0 0 pcpi_div_rd[15]
port 7 nsew signal tristate
flabel metal3 s 59200 38304 60000 38416 0 FreeSans 448 0 0 0 pcpi_div_rd[16]
port 8 nsew signal tristate
flabel metal3 s 59200 43008 60000 43120 0 FreeSans 448 0 0 0 pcpi_div_rd[17]
port 9 nsew signal tristate
flabel metal3 s 59200 34944 60000 35056 0 FreeSans 448 0 0 0 pcpi_div_rd[18]
port 10 nsew signal tristate
flabel metal3 s 59200 42336 60000 42448 0 FreeSans 448 0 0 0 pcpi_div_rd[19]
port 11 nsew signal tristate
flabel metal2 s 33600 59200 33712 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[1]
port 12 nsew signal tristate
flabel metal3 s 59200 35616 60000 35728 0 FreeSans 448 0 0 0 pcpi_div_rd[20]
port 13 nsew signal tristate
flabel metal3 s 59200 40992 60000 41104 0 FreeSans 448 0 0 0 pcpi_div_rd[21]
port 14 nsew signal tristate
flabel metal3 s 59200 37632 60000 37744 0 FreeSans 448 0 0 0 pcpi_div_rd[22]
port 15 nsew signal tristate
flabel metal3 s 59200 40320 60000 40432 0 FreeSans 448 0 0 0 pcpi_div_rd[23]
port 16 nsew signal tristate
flabel metal3 s 59200 36960 60000 37072 0 FreeSans 448 0 0 0 pcpi_div_rd[24]
port 17 nsew signal tristate
flabel metal3 s 59200 43680 60000 43792 0 FreeSans 448 0 0 0 pcpi_div_rd[25]
port 18 nsew signal tristate
flabel metal2 s 28896 59200 29008 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[26]
port 19 nsew signal tristate
flabel metal2 s 32256 59200 32368 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[27]
port 20 nsew signal tristate
flabel metal2 s 27552 59200 27664 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[28]
port 21 nsew signal tristate
flabel metal2 s 30240 59200 30352 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[29]
port 22 nsew signal tristate
flabel metal2 s 31584 59200 31696 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[2]
port 23 nsew signal tristate
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 pcpi_div_rd[30]
port 24 nsew signal tristate
flabel metal2 s 36960 59200 37072 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[31]
port 25 nsew signal tristate
flabel metal2 s 30912 59200 31024 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[3]
port 26 nsew signal tristate
flabel metal2 s 23520 59200 23632 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[4]
port 27 nsew signal tristate
flabel metal2 s 25536 59200 25648 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[5]
port 28 nsew signal tristate
flabel metal2 s 29568 59200 29680 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[6]
port 29 nsew signal tristate
flabel metal3 s 59200 38976 60000 39088 0 FreeSans 448 0 0 0 pcpi_div_rd[7]
port 30 nsew signal tristate
flabel metal3 s 59200 36288 60000 36400 0 FreeSans 448 0 0 0 pcpi_div_rd[8]
port 31 nsew signal tristate
flabel metal2 s 37632 59200 37744 60000 0 FreeSans 448 90 0 0 pcpi_div_rd[9]
port 32 nsew signal tristate
flabel metal3 s 0 49728 800 49840 0 FreeSans 448 0 0 0 pcpi_div_ready
port 33 nsew signal tristate
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 pcpi_div_valid
port 34 nsew signal input
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 pcpi_div_wait
port 35 nsew signal tristate
flabel metal3 s 0 43680 800 43792 0 FreeSans 448 0 0 0 pcpi_div_wr
port 36 nsew signal tristate
flabel metal3 s 0 43008 800 43120 0 FreeSans 448 0 0 0 pcpi_insn[0]
port 37 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 pcpi_insn[10]
port 38 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 pcpi_insn[11]
port 39 nsew signal input
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 pcpi_insn[12]
port 40 nsew signal input
flabel metal3 s 0 37632 800 37744 0 FreeSans 448 0 0 0 pcpi_insn[13]
port 41 nsew signal input
flabel metal3 s 0 38304 800 38416 0 FreeSans 448 0 0 0 pcpi_insn[14]
port 42 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 pcpi_insn[15]
port 43 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 pcpi_insn[16]
port 44 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 pcpi_insn[17]
port 45 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 pcpi_insn[18]
port 46 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 pcpi_insn[19]
port 47 nsew signal input
flabel metal3 s 0 44352 800 44464 0 FreeSans 448 0 0 0 pcpi_insn[1]
port 48 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 pcpi_insn[20]
port 49 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 pcpi_insn[21]
port 50 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 pcpi_insn[22]
port 51 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 pcpi_insn[23]
port 52 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 pcpi_insn[24]
port 53 nsew signal input
flabel metal3 s 0 45024 800 45136 0 FreeSans 448 0 0 0 pcpi_insn[25]
port 54 nsew signal input
flabel metal3 s 0 47712 800 47824 0 FreeSans 448 0 0 0 pcpi_insn[26]
port 55 nsew signal input
flabel metal3 s 0 49056 800 49168 0 FreeSans 448 0 0 0 pcpi_insn[27]
port 56 nsew signal input
flabel metal3 s 0 48384 800 48496 0 FreeSans 448 0 0 0 pcpi_insn[28]
port 57 nsew signal input
flabel metal3 s 0 41664 800 41776 0 FreeSans 448 0 0 0 pcpi_insn[29]
port 58 nsew signal input
flabel metal3 s 0 47040 800 47152 0 FreeSans 448 0 0 0 pcpi_insn[2]
port 59 nsew signal input
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 pcpi_insn[30]
port 60 nsew signal input
flabel metal3 s 0 35616 800 35728 0 FreeSans 448 0 0 0 pcpi_insn[31]
port 61 nsew signal input
flabel metal3 s 0 38976 800 39088 0 FreeSans 448 0 0 0 pcpi_insn[3]
port 62 nsew signal input
flabel metal3 s 0 45696 800 45808 0 FreeSans 448 0 0 0 pcpi_insn[4]
port 63 nsew signal input
flabel metal3 s 0 46368 800 46480 0 FreeSans 448 0 0 0 pcpi_insn[5]
port 64 nsew signal input
flabel metal3 s 0 42336 800 42448 0 FreeSans 448 0 0 0 pcpi_insn[6]
port 65 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 pcpi_insn[7]
port 66 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 pcpi_insn[8]
port 67 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 pcpi_insn[9]
port 68 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 pcpi_rs1[0]
port 69 nsew signal input
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 pcpi_rs1[10]
port 70 nsew signal input
flabel metal2 s 36288 0 36400 800 0 FreeSans 448 90 0 0 pcpi_rs1[11]
port 71 nsew signal input
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 pcpi_rs1[12]
port 72 nsew signal input
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 pcpi_rs1[13]
port 73 nsew signal input
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 pcpi_rs1[14]
port 74 nsew signal input
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 pcpi_rs1[15]
port 75 nsew signal input
flabel metal3 s 59200 23520 60000 23632 0 FreeSans 448 0 0 0 pcpi_rs1[16]
port 76 nsew signal input
flabel metal3 s 59200 22848 60000 22960 0 FreeSans 448 0 0 0 pcpi_rs1[17]
port 77 nsew signal input
flabel metal3 s 59200 24864 60000 24976 0 FreeSans 448 0 0 0 pcpi_rs1[18]
port 78 nsew signal input
flabel metal3 s 59200 24192 60000 24304 0 FreeSans 448 0 0 0 pcpi_rs1[19]
port 79 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 pcpi_rs1[1]
port 80 nsew signal input
flabel metal3 s 59200 25536 60000 25648 0 FreeSans 448 0 0 0 pcpi_rs1[20]
port 81 nsew signal input
flabel metal3 s 59200 26208 60000 26320 0 FreeSans 448 0 0 0 pcpi_rs1[21]
port 82 nsew signal input
flabel metal3 s 59200 29568 60000 29680 0 FreeSans 448 0 0 0 pcpi_rs1[22]
port 83 nsew signal input
flabel metal3 s 59200 28896 60000 29008 0 FreeSans 448 0 0 0 pcpi_rs1[23]
port 84 nsew signal input
flabel metal3 s 59200 27552 60000 27664 0 FreeSans 448 0 0 0 pcpi_rs1[24]
port 85 nsew signal input
flabel metal3 s 59200 26880 60000 26992 0 FreeSans 448 0 0 0 pcpi_rs1[25]
port 86 nsew signal input
flabel metal3 s 59200 28224 60000 28336 0 FreeSans 448 0 0 0 pcpi_rs1[26]
port 87 nsew signal input
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 pcpi_rs1[27]
port 88 nsew signal input
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 pcpi_rs1[28]
port 89 nsew signal input
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 pcpi_rs1[29]
port 90 nsew signal input
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 pcpi_rs1[2]
port 91 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 pcpi_rs1[30]
port 92 nsew signal input
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 pcpi_rs1[31]
port 93 nsew signal input
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 pcpi_rs1[3]
port 94 nsew signal input
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 pcpi_rs1[4]
port 95 nsew signal input
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 pcpi_rs1[5]
port 96 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 pcpi_rs1[6]
port 97 nsew signal input
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 pcpi_rs1[7]
port 98 nsew signal input
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 pcpi_rs1[8]
port 99 nsew signal input
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 pcpi_rs1[9]
port 100 nsew signal input
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 pcpi_rs2[0]
port 101 nsew signal input
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 pcpi_rs2[10]
port 102 nsew signal input
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 pcpi_rs2[11]
port 103 nsew signal input
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 pcpi_rs2[12]
port 104 nsew signal input
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 pcpi_rs2[13]
port 105 nsew signal input
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 pcpi_rs2[14]
port 106 nsew signal input
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 pcpi_rs2[15]
port 107 nsew signal input
flabel metal3 s 0 10080 800 10192 0 FreeSans 448 0 0 0 pcpi_rs2[16]
port 108 nsew signal input
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 pcpi_rs2[17]
port 109 nsew signal input
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 pcpi_rs2[18]
port 110 nsew signal input
flabel metal3 s 0 12768 800 12880 0 FreeSans 448 0 0 0 pcpi_rs2[19]
port 111 nsew signal input
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 pcpi_rs2[1]
port 112 nsew signal input
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 pcpi_rs2[20]
port 113 nsew signal input
flabel metal3 s 0 14112 800 14224 0 FreeSans 448 0 0 0 pcpi_rs2[21]
port 114 nsew signal input
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 pcpi_rs2[22]
port 115 nsew signal input
flabel metal3 s 0 10752 800 10864 0 FreeSans 448 0 0 0 pcpi_rs2[23]
port 116 nsew signal input
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 pcpi_rs2[24]
port 117 nsew signal input
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 pcpi_rs2[25]
port 118 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 pcpi_rs2[26]
port 119 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 pcpi_rs2[27]
port 120 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 pcpi_rs2[28]
port 121 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 pcpi_rs2[29]
port 122 nsew signal input
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 pcpi_rs2[2]
port 123 nsew signal input
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 pcpi_rs2[30]
port 124 nsew signal input
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 pcpi_rs2[31]
port 125 nsew signal input
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 pcpi_rs2[3]
port 126 nsew signal input
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 pcpi_rs2[4]
port 127 nsew signal input
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 pcpi_rs2[5]
port 128 nsew signal input
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 pcpi_rs2[6]
port 129 nsew signal input
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 pcpi_rs2[7]
port 130 nsew signal input
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 pcpi_rs2[8]
port 131 nsew signal input
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 pcpi_rs2[9]
port 132 nsew signal input
flabel metal3 s 0 40992 800 41104 0 FreeSans 448 0 0 0 resetn
port 133 nsew signal input
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 134 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 134 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 135 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 135 nsew ground bidirectional
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 18200 42224 18200 42224 0 _0000_
rlabel metal2 35840 42056 35840 42056 0 _0001_
rlabel metal2 34104 47208 34104 47208 0 _0002_
rlabel metal2 43400 36232 43400 36232 0 _0003_
rlabel metal2 42000 39032 42000 39032 0 _0004_
rlabel metal2 43176 42112 43176 42112 0 _0005_
rlabel metal2 45752 39984 45752 39984 0 _0006_
rlabel metal3 48384 38696 48384 38696 0 _0007_
rlabel metal3 48328 41048 48328 41048 0 _0008_
rlabel metal2 47880 37240 47880 37240 0 _0009_
rlabel metal2 50120 40936 50120 40936 0 _0010_
rlabel metal2 31416 41328 31416 41328 0 _0011_
rlabel metal3 53536 36568 53536 36568 0 _0012_
rlabel metal2 55384 39984 55384 39984 0 _0013_
rlabel metal3 52696 37240 52696 37240 0 _0014_
rlabel metal2 51688 40040 51688 40040 0 _0015_
rlabel metal3 41328 37912 41328 37912 0 _0016_
rlabel metal2 39592 41328 39592 41328 0 _0017_
rlabel metal2 26824 40824 26824 40824 0 _0018_
rlabel metal2 30408 38668 30408 38668 0 _0019_
rlabel metal2 26936 39144 26936 39144 0 _0020_
rlabel metal2 27160 38976 27160 38976 0 _0021_
rlabel metal2 29736 43960 29736 43960 0 _0022_
rlabel metal2 20104 36848 20104 36848 0 _0023_
rlabel metal2 34104 39984 34104 39984 0 _0024_
rlabel metal2 28168 45920 28168 45920 0 _0025_
rlabel metal2 22120 39928 22120 39928 0 _0026_
rlabel metal3 23016 40488 23016 40488 0 _0027_
rlabel metal2 27832 47824 27832 47824 0 _0028_
rlabel metal2 38248 38668 38248 38668 0 _0029_
rlabel metal2 35504 35784 35504 35784 0 _0030_
rlabel metal2 35224 43848 35224 43848 0 _0031_
rlabel metal2 9240 40712 9240 40712 0 _0032_
rlabel metal2 10360 41272 10360 41272 0 _0033_
rlabel metal3 8232 37912 8232 37912 0 _0034_
rlabel metal2 5544 37184 5544 37184 0 _0035_
rlabel metal3 7896 36568 7896 36568 0 _0036_
rlabel metal2 7896 43176 7896 43176 0 _0037_
rlabel metal2 20664 24360 20664 24360 0 _0038_
rlabel metal2 20664 22792 20664 22792 0 _0039_
rlabel metal2 22512 21672 22512 21672 0 _0040_
rlabel metal2 22344 19544 22344 19544 0 _0041_
rlabel metal2 21224 15148 21224 15148 0 _0042_
rlabel metal2 23016 10136 23016 10136 0 _0043_
rlabel metal2 26096 8456 26096 8456 0 _0044_
rlabel metal2 28224 7560 28224 7560 0 _0045_
rlabel metal2 34664 7112 34664 7112 0 _0046_
rlabel metal2 37576 7784 37576 7784 0 _0047_
rlabel metal3 42392 8120 42392 8120 0 _0048_
rlabel metal2 43512 8680 43512 8680 0 _0049_
rlabel metal2 47656 11368 47656 11368 0 _0050_
rlabel metal2 50960 13944 50960 13944 0 _0051_
rlabel metal2 52584 15624 52584 15624 0 _0052_
rlabel metal2 52248 17192 52248 17192 0 _0053_
rlabel metal2 53592 18088 53592 18088 0 _0054_
rlabel metal2 56168 21112 56168 21112 0 _0055_
rlabel metal2 56056 22680 56056 22680 0 _0056_
rlabel metal2 55832 24248 55832 24248 0 _0057_
rlabel metal2 56056 25816 56056 25816 0 _0058_
rlabel metal2 56056 27776 56056 27776 0 _0059_
rlabel metal2 56056 30520 56056 30520 0 _0060_
rlabel metal2 55272 32872 55272 32872 0 _0061_
rlabel metal2 42224 31976 42224 31976 0 _0062_
rlabel metal2 32312 31640 32312 31640 0 _0063_
rlabel metal3 29960 33208 29960 33208 0 _0064_
rlabel metal3 25144 33208 25144 33208 0 _0065_
rlabel metal2 18200 33656 18200 33656 0 _0066_
rlabel metal2 15848 35224 15848 35224 0 _0067_
rlabel metal2 13384 34440 13384 34440 0 _0068_
rlabel metal2 18200 45416 18200 45416 0 _0069_
rlabel metal2 17864 47824 17864 47824 0 _0070_
rlabel metal2 16408 47880 16408 47880 0 _0071_
rlabel metal2 18424 51688 18424 51688 0 _0072_
rlabel metal2 20440 48328 20440 48328 0 _0073_
rlabel metal3 21952 50456 21952 50456 0 _0074_
rlabel metal3 21056 52248 21056 52248 0 _0075_
rlabel metal2 30744 47992 30744 47992 0 _0076_
rlabel metal3 29232 50456 29232 50456 0 _0077_
rlabel metal2 30520 51464 30520 51464 0 _0078_
rlabel metal2 31416 54096 31416 54096 0 _0079_
rlabel metal3 34216 54432 34216 54432 0 _0080_
rlabel metal2 39032 51632 39032 51632 0 _0081_
rlabel metal2 38248 50176 38248 50176 0 _0082_
rlabel metal2 42112 47544 42112 47544 0 _0083_
rlabel metal2 42392 49448 42392 49448 0 _0084_
rlabel metal2 45920 46760 45920 46760 0 _0085_
rlabel metal2 49560 47152 49560 47152 0 _0086_
rlabel metal2 46088 50568 46088 50568 0 _0087_
rlabel metal2 48048 49112 48048 49112 0 _0088_
rlabel metal2 53592 50456 53592 50456 0 _0089_
rlabel metal2 54824 49392 54824 49392 0 _0090_
rlabel metal2 53368 45808 53368 45808 0 _0091_
rlabel metal3 52360 46760 52360 46760 0 _0092_
rlabel metal3 37296 46648 37296 46648 0 _0093_
rlabel metal3 37072 47320 37072 47320 0 _0094_
rlabel metal3 25200 45976 25200 45976 0 _0095_
rlabel metal2 24920 48440 24920 48440 0 _0096_
rlabel metal2 14728 43176 14728 43176 0 _0097_
rlabel metal2 13608 43120 13608 43120 0 _0098_
rlabel metal2 14280 39984 14280 39984 0 _0099_
rlabel metal2 14728 40712 14728 40712 0 _0100_
rlabel metal2 14616 46312 14616 46312 0 _0101_
rlabel metal2 12936 50176 12936 50176 0 _0102_
rlabel metal2 14504 51800 14504 51800 0 _0103_
rlabel metal2 15512 53368 15512 53368 0 _0104_
rlabel metal2 16744 54936 16744 54936 0 _0105_
rlabel metal2 19656 53760 19656 53760 0 _0106_
rlabel metal2 18536 54936 18536 54936 0 _0107_
rlabel metal2 24416 55832 24416 55832 0 _0108_
rlabel metal2 24584 52976 24584 52976 0 _0109_
rlabel metal2 27608 53256 27608 53256 0 _0110_
rlabel metal2 28392 54824 28392 54824 0 _0111_
rlabel metal3 36288 55496 36288 55496 0 _0112_
rlabel metal2 35560 54656 35560 54656 0 _0113_
rlabel metal2 39032 54936 39032 54936 0 _0114_
rlabel metal2 42112 55944 42112 55944 0 _0115_
rlabel metal2 44240 53032 44240 53032 0 _0116_
rlabel metal2 43400 54824 43400 54824 0 _0117_
rlabel metal2 48104 54936 48104 54936 0 _0118_
rlabel metal2 47768 53368 47768 53368 0 _0119_
rlabel metal2 49448 54936 49448 54936 0 _0120_
rlabel metal2 51576 54040 51576 54040 0 _0121_
rlabel metal3 51912 52920 51912 52920 0 _0122_
rlabel metal2 51912 51016 51912 51016 0 _0123_
rlabel metal2 36512 51240 36512 51240 0 _0124_
rlabel metal2 34048 51352 34048 51352 0 _0125_
rlabel metal2 26320 51240 26320 51240 0 _0126_
rlabel metal2 25368 50232 25368 50232 0 _0127_
rlabel metal2 10808 49336 10808 49336 0 _0128_
rlabel metal2 10920 47096 10920 47096 0 _0129_
rlabel metal2 9128 46200 9128 46200 0 _0130_
rlabel metal2 8904 44632 8904 44632 0 _0131_
rlabel metal2 10808 35112 10808 35112 0 _0132_
rlabel metal3 13552 24584 13552 24584 0 _0133_
rlabel metal2 25480 27216 25480 27216 0 _0134_
rlabel metal2 23632 24024 23632 24024 0 _0135_
rlabel metal3 32312 20888 32312 20888 0 _0136_
rlabel metal3 27272 20664 27272 20664 0 _0137_
rlabel metal2 22120 17808 22120 17808 0 _0138_
rlabel metal2 23464 15400 23464 15400 0 _0139_
rlabel metal2 22568 12488 22568 12488 0 _0140_
rlabel metal3 31640 9688 31640 9688 0 _0141_
rlabel metal2 32256 8344 32256 8344 0 _0142_
rlabel metal2 35672 16520 35672 16520 0 _0143_
rlabel metal2 38696 15120 38696 15120 0 _0144_
rlabel metal2 43624 12488 43624 12488 0 _0145_
rlabel metal2 39816 16408 39816 16408 0 _0146_
rlabel metal2 40376 17864 40376 17864 0 _0147_
rlabel metal2 41944 21168 41944 21168 0 _0148_
rlabel metal2 46088 18760 46088 18760 0 _0149_
rlabel metal2 46088 21896 46088 21896 0 _0150_
rlabel metal2 47824 19320 47824 19320 0 _0151_
rlabel metal2 46088 28056 46088 28056 0 _0152_
rlabel metal2 45864 25032 45864 25032 0 _0153_
rlabel metal2 47992 29008 47992 29008 0 _0154_
rlabel metal3 44968 33208 44968 33208 0 _0155_
rlabel metal2 47992 30632 47992 30632 0 _0156_
rlabel metal3 45192 31080 45192 31080 0 _0157_
rlabel metal2 38248 34440 38248 34440 0 _0158_
rlabel metal2 41048 30464 41048 30464 0 _0159_
rlabel metal2 26488 32256 26488 32256 0 _0160_
rlabel metal2 27384 29736 27384 29736 0 _0161_
rlabel metal2 20216 34440 20216 34440 0 _0162_
rlabel metal2 21224 29736 21224 29736 0 _0163_
rlabel metal2 13048 29736 13048 29736 0 _0164_
rlabel metal2 16408 26684 16408 26684 0 _0165_
rlabel metal3 16072 37912 16072 37912 0 _0166_
rlabel metal2 6440 39032 6440 39032 0 _0167_
rlabel metal2 15680 24024 15680 24024 0 _0168_
rlabel metal2 11256 32144 11256 32144 0 _0169_
rlabel metal2 8400 32760 8400 32760 0 _0170_
rlabel metal2 6216 33488 6216 33488 0 _0171_
rlabel metal2 2856 33208 2856 33208 0 _0172_
rlabel metal2 2856 31892 2856 31892 0 _0173_
rlabel metal2 3640 29848 3640 29848 0 _0174_
rlabel metal2 3640 28280 3640 28280 0 _0175_
rlabel metal2 3864 25872 3864 25872 0 _0176_
rlabel metal2 11704 23520 11704 23520 0 _0177_
rlabel metal2 7112 24304 7112 24304 0 _0178_
rlabel metal2 2576 23352 2576 23352 0 _0179_
rlabel metal2 2520 22008 2520 22008 0 _0180_
rlabel metal2 2520 20328 2520 20328 0 _0181_
rlabel metal2 3304 16800 3304 16800 0 _0182_
rlabel metal2 3192 15736 3192 15736 0 _0183_
rlabel metal2 2520 13328 2520 13328 0 _0184_
rlabel metal2 2576 11480 2576 11480 0 _0185_
rlabel metal3 4424 9688 4424 9688 0 _0186_
rlabel metal2 5992 8512 5992 8512 0 _0187_
rlabel metal2 8120 8624 8120 8624 0 _0188_
rlabel metal2 10696 10528 10696 10528 0 _0189_
rlabel metal2 10584 7784 10584 7784 0 _0190_
rlabel metal2 15176 8624 15176 8624 0 _0191_
rlabel metal2 12600 7000 12600 7000 0 _0192_
rlabel metal2 12488 18480 12488 18480 0 _0193_
rlabel metal2 17696 8344 17696 8344 0 _0194_
rlabel metal3 18816 9128 18816 9128 0 _0195_
rlabel metal2 19824 10696 19824 10696 0 _0196_
rlabel metal2 20216 13328 20216 13328 0 _0197_
rlabel metal2 19544 17864 19544 17864 0 _0198_
rlabel metal2 16072 21504 16072 21504 0 _0199_
rlabel metal3 45752 15288 45752 15288 0 _0200_
rlabel metal3 43288 15288 43288 15288 0 _0201_
rlabel metal2 43400 15904 43400 15904 0 _0202_
rlabel metal2 44464 15512 44464 15512 0 _0203_
rlabel metal3 42672 12824 42672 12824 0 _0204_
rlabel metal2 42840 10080 42840 10080 0 _0205_
rlabel metal2 40936 9464 40936 9464 0 _0206_
rlabel metal2 39144 9464 39144 9464 0 _0207_
rlabel metal2 39256 9968 39256 9968 0 _0208_
rlabel metal2 41048 12488 41048 12488 0 _0209_
rlabel metal2 41160 13384 41160 13384 0 _0210_
rlabel metal2 47320 24640 47320 24640 0 _0211_
rlabel metal2 39592 11536 39592 11536 0 _0212_
rlabel metal2 37352 11480 37352 11480 0 _0213_
rlabel metal2 37464 9660 37464 9660 0 _0214_
rlabel metal2 43176 12544 43176 12544 0 _0215_
rlabel metal2 42952 10808 42952 10808 0 _0216_
rlabel metal3 42504 11256 42504 11256 0 _0217_
rlabel metal2 43064 13328 43064 13328 0 _0218_
rlabel metal2 46648 14168 46648 14168 0 _0219_
rlabel metal3 49056 15848 49056 15848 0 _0220_
rlabel metal2 47600 15288 47600 15288 0 _0221_
rlabel metal2 49112 16352 49112 16352 0 _0222_
rlabel metal2 47096 17248 47096 17248 0 _0223_
rlabel metal2 45640 15120 45640 15120 0 _0224_
rlabel metal2 43960 16296 43960 16296 0 _0225_
rlabel metal2 45808 15512 45808 15512 0 _0226_
rlabel metal2 46536 15232 46536 15232 0 _0227_
rlabel metal3 47376 15400 47376 15400 0 _0228_
rlabel metal3 47096 15288 47096 15288 0 _0229_
rlabel metal2 47768 22848 47768 22848 0 _0230_
rlabel metal2 53088 29176 53088 29176 0 _0231_
rlabel metal2 50904 21448 50904 21448 0 _0232_
rlabel metal2 50120 22792 50120 22792 0 _0233_
rlabel metal2 51352 23632 51352 23632 0 _0234_
rlabel metal3 51408 26264 51408 26264 0 _0235_
rlabel metal3 52528 30072 52528 30072 0 _0236_
rlabel metal2 49784 29680 49784 29680 0 _0237_
rlabel metal2 48776 30128 48776 30128 0 _0238_
rlabel metal2 48664 27496 48664 27496 0 _0239_
rlabel metal2 47544 25984 47544 25984 0 _0240_
rlabel metal2 30296 30800 30296 30800 0 _0241_
rlabel metal2 31864 29064 31864 29064 0 _0242_
rlabel metal2 32536 29288 32536 29288 0 _0243_
rlabel metal3 32536 30856 32536 30856 0 _0244_
rlabel metal2 33544 30296 33544 30296 0 _0245_
rlabel metal2 39032 29736 39032 29736 0 _0246_
rlabel metal2 36680 31136 36680 31136 0 _0247_
rlabel metal2 35112 29904 35112 29904 0 _0248_
rlabel metal2 34888 28616 34888 28616 0 _0249_
rlabel metal2 24248 30576 24248 30576 0 _0250_
rlabel metal2 30856 30128 30856 30128 0 _0251_
rlabel metal2 29736 30688 29736 30688 0 _0252_
rlabel metal3 39760 29960 39760 29960 0 _0253_
rlabel metal3 38472 30184 38472 30184 0 _0254_
rlabel metal3 39144 32760 39144 32760 0 _0255_
rlabel metal2 39256 29680 39256 29680 0 _0256_
rlabel metal2 39368 30240 39368 30240 0 _0257_
rlabel metal2 35672 29624 35672 29624 0 _0258_
rlabel metal3 30856 30968 30856 30968 0 _0259_
rlabel metal3 24248 31640 24248 31640 0 _0260_
rlabel metal2 22960 30968 22960 30968 0 _0261_
rlabel metal2 24808 31584 24808 31584 0 _0262_
rlabel metal2 23128 30632 23128 30632 0 _0263_
rlabel metal2 19040 31192 19040 31192 0 _0264_
rlabel metal2 19432 31248 19432 31248 0 _0265_
rlabel metal2 20104 31192 20104 31192 0 _0266_
rlabel metal2 19208 31920 19208 31920 0 _0267_
rlabel metal3 18088 31640 18088 31640 0 _0268_
rlabel metal2 16408 31248 16408 31248 0 _0269_
rlabel metal2 15848 32928 15848 32928 0 _0270_
rlabel metal2 16520 31416 16520 31416 0 _0271_
rlabel metal2 16744 31640 16744 31640 0 _0272_
rlabel metal2 17192 31584 17192 31584 0 _0273_
rlabel metal2 15904 32312 15904 32312 0 _0274_
rlabel metal2 14952 32144 14952 32144 0 _0275_
rlabel metal2 15736 11088 15736 11088 0 _0276_
rlabel metal2 15064 10920 15064 10920 0 _0277_
rlabel metal3 16520 16632 16520 16632 0 _0278_
rlabel metal2 14728 11256 14728 11256 0 _0279_
rlabel metal2 14448 17080 14448 17080 0 _0280_
rlabel metal2 5656 24808 5656 24808 0 _0281_
rlabel metal2 1624 21560 1624 21560 0 _0282_
rlabel metal2 6104 25760 6104 25760 0 _0283_
rlabel metal2 6328 26180 6328 26180 0 _0284_
rlabel metal3 10080 25704 10080 25704 0 _0285_
rlabel metal2 14280 25984 14280 25984 0 _0286_
rlabel metal2 15176 32424 15176 32424 0 _0287_
rlabel metal2 13832 38584 13832 38584 0 _0288_
rlabel metal2 21224 38724 21224 38724 0 _0289_
rlabel metal2 21896 38724 21896 38724 0 _0290_
rlabel metal2 23128 44240 23128 44240 0 _0291_
rlabel metal2 22568 22680 22568 22680 0 _0292_
rlabel metal2 18536 45080 18536 45080 0 _0293_
rlabel metal3 20440 49784 20440 49784 0 _0294_
rlabel metal2 17696 46872 17696 46872 0 _0295_
rlabel metal2 16744 48216 16744 48216 0 _0296_
rlabel metal2 23464 51296 23464 51296 0 _0297_
rlabel metal2 19712 50456 19712 50456 0 _0298_
rlabel metal2 18648 51352 18648 51352 0 _0299_
rlabel metal3 20048 49672 20048 49672 0 _0300_
rlabel metal2 44912 51352 44912 51352 0 _0301_
rlabel metal2 21896 51688 21896 51688 0 _0302_
rlabel metal2 22064 50680 22064 50680 0 _0303_
rlabel metal3 21392 52136 21392 52136 0 _0304_
rlabel metal2 26376 23156 26376 23156 0 _0305_
rlabel metal2 29288 47936 29288 47936 0 _0306_
rlabel metal3 32816 54712 32816 54712 0 _0307_
rlabel metal2 29064 49616 29064 49616 0 _0308_
rlabel metal2 29624 52192 29624 52192 0 _0309_
rlabel metal2 39256 52472 39256 52472 0 _0310_
rlabel metal2 31640 53704 31640 53704 0 _0311_
rlabel metal3 33768 54376 33768 54376 0 _0312_
rlabel metal2 40432 48104 40432 48104 0 _0313_
rlabel metal2 41384 50904 41384 50904 0 _0314_
rlabel metal2 39256 51464 39256 51464 0 _0315_
rlabel metal2 41160 51016 41160 51016 0 _0316_
rlabel metal2 43064 48608 43064 48608 0 _0317_
rlabel metal2 42168 48384 42168 48384 0 _0318_
rlabel metal2 42952 49112 42952 49112 0 _0319_
rlabel metal3 46984 51464 46984 51464 0 _0320_
rlabel metal2 45808 47656 45808 47656 0 _0321_
rlabel metal3 48048 46760 48048 46760 0 _0322_
rlabel metal3 53536 51352 53536 51352 0 _0323_
rlabel metal2 46536 51128 46536 51128 0 _0324_
rlabel metal3 48496 50008 48496 50008 0 _0325_
rlabel metal3 54488 50008 54488 50008 0 _0326_
rlabel metal3 53424 49896 53424 49896 0 _0327_
rlabel metal2 53816 50820 53816 50820 0 _0328_
rlabel metal2 22008 26096 22008 26096 0 _0329_
rlabel metal2 36904 47936 36904 47936 0 _0330_
rlabel metal2 51800 47376 51800 47376 0 _0331_
rlabel metal2 51128 47768 51128 47768 0 _0332_
rlabel metal2 26376 46200 26376 46200 0 _0333_
rlabel metal2 36792 46984 36792 46984 0 _0334_
rlabel metal2 36456 47880 36456 47880 0 _0335_
rlabel metal2 13944 44520 13944 44520 0 _0336_
rlabel metal2 26712 46312 26712 46312 0 _0337_
rlabel metal2 26824 48048 26824 48048 0 _0338_
rlabel metal2 13552 42504 13552 42504 0 _0339_
rlabel metal3 14224 42952 14224 42952 0 _0340_
rlabel metal3 13160 42952 13160 42952 0 _0341_
rlabel metal2 14952 40824 14952 40824 0 _0342_
rlabel metal2 13608 40600 13608 40600 0 _0343_
rlabel metal3 15456 41160 15456 41160 0 _0344_
rlabel metal3 14952 45976 14952 45976 0 _0345_
rlabel metal2 17416 52584 17416 52584 0 _0346_
rlabel metal3 14784 50680 14784 50680 0 _0347_
rlabel metal3 15400 51240 15400 51240 0 _0348_
rlabel metal2 17584 53704 17584 53704 0 _0349_
rlabel metal2 15624 53424 15624 53424 0 _0350_
rlabel metal2 16856 54656 16856 54656 0 _0351_
rlabel metal3 25088 53032 25088 53032 0 _0352_
rlabel metal2 19656 52920 19656 52920 0 _0353_
rlabel metal2 19880 54096 19880 54096 0 _0354_
rlabel metal2 25368 53368 25368 53368 0 _0355_
rlabel metal2 24360 54292 24360 54292 0 _0356_
rlabel metal3 25032 52248 25032 52248 0 _0357_
rlabel metal2 45416 53200 45416 53200 0 _0358_
rlabel metal2 42280 53872 42280 53872 0 _0359_
rlabel metal2 27832 53872 27832 53872 0 _0360_
rlabel metal2 29288 54488 29288 54488 0 _0361_
rlabel metal2 25256 52696 25256 52696 0 _0362_
rlabel metal2 39592 54432 39592 54432 0 _0363_
rlabel metal2 38360 54936 38360 54936 0 _0364_
rlabel metal3 37016 53816 37016 53816 0 _0365_
rlabel metal2 46536 54264 46536 54264 0 _0366_
rlabel metal2 39144 54656 39144 54656 0 _0367_
rlabel metal2 41944 54656 41944 54656 0 _0368_
rlabel metal2 46088 54040 46088 54040 0 _0369_
rlabel metal2 44576 53816 44576 53816 0 _0370_
rlabel metal2 46424 54936 46424 54936 0 _0371_
rlabel metal2 49952 53480 49952 53480 0 _0372_
rlabel metal2 46312 53648 46312 53648 0 _0373_
rlabel metal2 47544 53032 47544 53032 0 _0374_
rlabel metal3 50848 52136 50848 52136 0 _0375_
rlabel metal2 49560 54096 49560 54096 0 _0376_
rlabel metal2 51128 53816 51128 53816 0 _0377_
rlabel metal2 44184 51688 44184 51688 0 _0378_
rlabel metal2 51240 52528 51240 52528 0 _0379_
rlabel metal3 51072 50680 51072 50680 0 _0380_
rlabel metal3 25816 49784 25816 49784 0 _0381_
rlabel metal3 36624 49672 36624 49672 0 _0382_
rlabel metal2 33880 51520 33880 51520 0 _0383_
rlabel metal2 13384 49112 13384 49112 0 _0384_
rlabel metal2 25704 49616 25704 49616 0 _0385_
rlabel metal3 26376 49672 26376 49672 0 _0386_
rlabel metal3 10248 42840 10248 42840 0 _0387_
rlabel metal2 11592 47432 11592 47432 0 _0388_
rlabel metal2 11928 48440 11928 48440 0 _0389_
rlabel metal3 11424 46760 11424 46760 0 _0390_
rlabel metal2 11816 46256 11816 46256 0 _0391_
rlabel metal3 10360 44968 10360 44968 0 _0392_
rlabel metal2 11032 35168 11032 35168 0 _0393_
rlabel metal2 16296 10080 16296 10080 0 _0394_
rlabel metal3 16632 9912 16632 9912 0 _0395_
rlabel metal2 13832 20664 13832 20664 0 _0396_
rlabel metal2 22792 27216 22792 27216 0 _0397_
rlabel metal2 44184 29456 44184 29456 0 _0398_
rlabel metal2 11536 22120 11536 22120 0 _0399_
rlabel metal2 13832 24248 13832 24248 0 _0400_
rlabel metal2 18088 26432 18088 26432 0 _0401_
rlabel metal2 26712 30016 26712 30016 0 _0402_
rlabel metal2 25928 24472 25928 24472 0 _0403_
rlabel metal2 23464 23072 23464 23072 0 _0404_
rlabel metal3 24360 23016 24360 23016 0 _0405_
rlabel metal2 30576 20552 30576 20552 0 _0406_
rlabel metal2 42616 26208 42616 26208 0 _0407_
rlabel metal3 27104 25368 27104 25368 0 _0408_
rlabel metal2 26152 25032 26152 25032 0 _0409_
rlabel metal2 25704 25900 25704 25900 0 _0410_
rlabel metal2 26040 27944 26040 27944 0 _0411_
rlabel metal2 19432 21168 19432 21168 0 _0412_
rlabel metal2 19544 24640 19544 24640 0 _0413_
rlabel metal2 21784 25648 21784 25648 0 _0414_
rlabel metal2 12096 27608 12096 27608 0 _0415_
rlabel metal2 19600 25704 19600 25704 0 _0416_
rlabel via2 22456 25256 22456 25256 0 _0417_
rlabel metal2 35112 25088 35112 25088 0 _0418_
rlabel metal2 33656 17584 33656 17584 0 _0419_
rlabel metal2 32760 24192 32760 24192 0 _0420_
rlabel metal3 31696 24696 31696 24696 0 _0421_
rlabel metal2 28672 25368 28672 25368 0 _0422_
rlabel metal2 18088 24304 18088 24304 0 _0423_
rlabel metal2 18536 21952 18536 21952 0 _0424_
rlabel metal2 29512 24192 29512 24192 0 _0425_
rlabel metal2 30072 24920 30072 24920 0 _0426_
rlabel metal2 30408 25816 30408 25816 0 _0427_
rlabel metal3 29512 24920 29512 24920 0 _0428_
rlabel metal2 31248 17416 31248 17416 0 _0429_
rlabel metal2 43736 20328 43736 20328 0 _0430_
rlabel metal2 31864 18928 31864 18928 0 _0431_
rlabel metal2 20552 20552 20552 20552 0 _0432_
rlabel metal2 43064 18928 43064 18928 0 _0433_
rlabel metal2 40376 24976 40376 24976 0 _0434_
rlabel metal2 34384 22456 34384 22456 0 _0435_
rlabel metal2 33096 23800 33096 23800 0 _0436_
rlabel metal3 29792 23240 29792 23240 0 _0437_
rlabel metal2 30968 22400 30968 22400 0 _0438_
rlabel metal2 18872 22288 18872 22288 0 _0439_
rlabel metal2 30576 21672 30576 21672 0 _0440_
rlabel metal2 30968 21952 30968 21952 0 _0441_
rlabel metal2 31976 21112 31976 21112 0 _0442_
rlabel metal2 32088 19824 32088 19824 0 _0443_
rlabel metal2 24920 29624 24920 29624 0 _0444_
rlabel metal2 35728 23688 35728 23688 0 _0445_
rlabel metal3 34272 23016 34272 23016 0 _0446_
rlabel metal3 32312 23128 32312 23128 0 _0447_
rlabel metal2 29904 21560 29904 21560 0 _0448_
rlabel metal2 45528 26684 45528 26684 0 _0449_
rlabel metal2 29960 22568 29960 22568 0 _0450_
rlabel metal2 29624 21952 29624 21952 0 _0451_
rlabel metal2 32200 21756 32200 21756 0 _0452_
rlabel metal2 30520 21056 30520 21056 0 _0453_
rlabel metal2 24136 18424 24136 18424 0 _0454_
rlabel metal2 40152 28056 40152 28056 0 _0455_
rlabel metal2 38920 24808 38920 24808 0 _0456_
rlabel metal2 33544 20664 33544 20664 0 _0457_
rlabel metal2 26824 18816 26824 18816 0 _0458_
rlabel metal2 20328 18984 20328 18984 0 _0459_
rlabel metal2 39592 21952 39592 21952 0 _0460_
rlabel metal2 32312 18592 32312 18592 0 _0461_
rlabel metal2 27048 18368 27048 18368 0 _0462_
rlabel metal2 26600 17696 26600 17696 0 _0463_
rlabel metal2 25928 17640 25928 17640 0 _0464_
rlabel metal2 26824 17976 26824 17976 0 _0465_
rlabel metal2 26376 18312 26376 18312 0 _0466_
rlabel metal3 25984 18424 25984 18424 0 _0467_
rlabel metal2 25816 18928 25816 18928 0 _0468_
rlabel metal2 19096 19880 19096 19880 0 _0469_
rlabel metal2 32648 18032 32648 18032 0 _0470_
rlabel metal3 30464 17528 30464 17528 0 _0471_
rlabel metal2 27272 17192 27272 17192 0 _0472_
rlabel metal3 27776 17528 27776 17528 0 _0473_
rlabel metal3 29512 17416 29512 17416 0 _0474_
rlabel metal2 30016 17640 30016 17640 0 _0475_
rlabel metal2 29120 16856 29120 16856 0 _0476_
rlabel metal2 24024 16016 24024 16016 0 _0477_
rlabel metal2 33208 16744 33208 16744 0 _0478_
rlabel metal2 31192 15736 31192 15736 0 _0479_
rlabel metal2 27272 14000 27272 14000 0 _0480_
rlabel metal2 27384 13720 27384 13720 0 _0481_
rlabel metal2 26264 13272 26264 13272 0 _0482_
rlabel metal2 26824 12544 26824 12544 0 _0483_
rlabel metal2 26376 12264 26376 12264 0 _0484_
rlabel metal2 26152 13328 26152 13328 0 _0485_
rlabel metal2 26712 13272 26712 13272 0 _0486_
rlabel metal3 24136 12880 24136 12880 0 _0487_
rlabel metal3 24920 12824 24920 12824 0 _0488_
rlabel metal2 31640 18368 31640 18368 0 _0489_
rlabel metal2 26264 25984 26264 25984 0 _0490_
rlabel metal3 32032 15176 32032 15176 0 _0491_
rlabel metal3 31192 12936 31192 12936 0 _0492_
rlabel metal2 30296 11760 30296 11760 0 _0493_
rlabel metal2 30632 11704 30632 11704 0 _0494_
rlabel metal2 30408 12544 30408 12544 0 _0495_
rlabel metal2 31976 12712 31976 12712 0 _0496_
rlabel metal2 31864 11592 31864 11592 0 _0497_
rlabel metal3 33544 15848 33544 15848 0 _0498_
rlabel metal2 33320 13496 33320 13496 0 _0499_
rlabel metal2 33040 12824 33040 12824 0 _0500_
rlabel metal2 39480 13608 39480 13608 0 _0501_
rlabel metal2 37800 12488 37800 12488 0 _0502_
rlabel metal2 34104 11088 34104 11088 0 _0503_
rlabel metal2 34608 12376 34608 12376 0 _0504_
rlabel metal2 33880 12656 33880 12656 0 _0505_
rlabel metal2 33320 12488 33320 12488 0 _0506_
rlabel metal2 32928 11368 32928 11368 0 _0507_
rlabel metal2 39088 17640 39088 17640 0 _0508_
rlabel metal2 39256 16128 39256 16128 0 _0509_
rlabel metal2 34216 15568 34216 15568 0 _0510_
rlabel metal3 35616 15176 35616 15176 0 _0511_
rlabel metal2 34664 11088 34664 11088 0 _0512_
rlabel metal3 34776 11480 34776 11480 0 _0513_
rlabel metal3 36120 14784 36120 14784 0 _0514_
rlabel metal2 36232 14840 36232 14840 0 _0515_
rlabel metal3 36344 15960 36344 15960 0 _0516_
rlabel metal3 36680 15848 36680 15848 0 _0517_
rlabel metal3 16184 17416 16184 17416 0 _0518_
rlabel metal2 23128 14952 23128 14952 0 _0519_
rlabel metal2 37688 15680 37688 15680 0 _0520_
rlabel metal3 36008 14280 36008 14280 0 _0521_
rlabel metal2 37352 15400 37352 15400 0 _0522_
rlabel metal2 37576 13944 37576 13944 0 _0523_
rlabel metal2 38920 11760 38920 11760 0 _0524_
rlabel metal2 37912 11312 37912 11312 0 _0525_
rlabel metal2 37576 10192 37576 10192 0 _0526_
rlabel metal3 38696 11424 38696 11424 0 _0527_
rlabel metal2 38136 12824 38136 12824 0 _0528_
rlabel metal2 39368 12544 39368 12544 0 _0529_
rlabel metal2 38472 13720 38472 13720 0 _0530_
rlabel metal2 39368 14616 39368 14616 0 _0531_
rlabel metal2 39032 15344 39032 15344 0 _0532_
rlabel metal2 36680 13832 36680 13832 0 _0533_
rlabel metal3 36792 13776 36792 13776 0 _0534_
rlabel metal3 40096 11368 40096 11368 0 _0535_
rlabel metal2 41272 11648 41272 11648 0 _0536_
rlabel metal2 42168 13216 42168 13216 0 _0537_
rlabel metal2 42504 12152 42504 12152 0 _0538_
rlabel metal2 34048 14728 34048 14728 0 _0539_
rlabel metal2 35336 20384 35336 20384 0 _0540_
rlabel metal2 35336 19376 35336 19376 0 _0541_
rlabel metal2 36680 18704 36680 18704 0 _0542_
rlabel metal2 43456 12936 43456 12936 0 _0543_
rlabel metal3 42280 16632 42280 16632 0 _0544_
rlabel metal3 42504 17080 42504 17080 0 _0545_
rlabel metal2 43008 16744 43008 16744 0 _0546_
rlabel metal2 42840 17920 42840 17920 0 _0547_
rlabel metal3 38136 18144 38136 18144 0 _0548_
rlabel metal3 37352 17640 37352 17640 0 _0549_
rlabel metal2 38416 17640 38416 17640 0 _0550_
rlabel metal3 35560 20552 35560 20552 0 _0551_
rlabel metal3 37464 19208 37464 19208 0 _0552_
rlabel metal2 43176 15568 43176 15568 0 _0553_
rlabel metal2 42280 15960 42280 15960 0 _0554_
rlabel metal2 37464 18536 37464 18536 0 _0555_
rlabel metal2 38136 18536 38136 18536 0 _0556_
rlabel metal3 38920 18424 38920 18424 0 _0557_
rlabel metal2 39088 20216 39088 20216 0 _0558_
rlabel metal2 39984 20104 39984 20104 0 _0559_
rlabel metal3 40152 20664 40152 20664 0 _0560_
rlabel metal2 40600 20664 40600 20664 0 _0561_
rlabel metal2 45192 17136 45192 17136 0 _0562_
rlabel metal2 44968 16016 44968 16016 0 _0563_
rlabel metal2 44632 17808 44632 17808 0 _0564_
rlabel metal3 41160 20776 41160 20776 0 _0565_
rlabel metal2 42448 20776 42448 20776 0 _0566_
rlabel metal2 45976 16632 45976 16632 0 _0567_
rlabel metal3 44800 17416 44800 17416 0 _0568_
rlabel metal2 44296 18088 44296 18088 0 _0569_
rlabel metal2 44016 18648 44016 18648 0 _0570_
rlabel metal2 38864 20216 38864 20216 0 _0571_
rlabel metal2 43736 19600 43736 19600 0 _0572_
rlabel metal2 44072 19376 44072 19376 0 _0573_
rlabel metal2 46312 20440 46312 20440 0 _0574_
rlabel metal2 45192 19488 45192 19488 0 _0575_
rlabel metal3 38024 21000 38024 21000 0 _0576_
rlabel metal2 39592 24136 39592 24136 0 _0577_
rlabel metal2 38584 23072 38584 23072 0 _0578_
rlabel metal3 40320 23912 40320 23912 0 _0579_
rlabel metal3 41160 23688 41160 23688 0 _0580_
rlabel metal2 42952 22568 42952 22568 0 _0581_
rlabel metal2 39256 22736 39256 22736 0 _0582_
rlabel metal2 43064 23688 43064 23688 0 _0583_
rlabel metal2 48104 23072 48104 23072 0 _0584_
rlabel metal3 46256 23240 46256 23240 0 _0585_
rlabel metal2 44016 23912 44016 23912 0 _0586_
rlabel metal3 44352 23128 44352 23128 0 _0587_
rlabel metal2 45528 22624 45528 22624 0 _0588_
rlabel metal3 38780 23128 38780 23128 0 _0589_
rlabel metal3 40712 21672 40712 21672 0 _0590_
rlabel metal2 50344 26208 50344 26208 0 _0591_
rlabel metal2 50232 21896 50232 21896 0 _0592_
rlabel metal2 50344 21280 50344 21280 0 _0593_
rlabel metal3 45304 20888 45304 20888 0 _0594_
rlabel metal3 40544 21784 40544 21784 0 _0595_
rlabel metal3 43624 21000 43624 21000 0 _0596_
rlabel metal3 46312 20664 46312 20664 0 _0597_
rlabel metal2 16576 17752 16576 17752 0 _0598_
rlabel metal3 53256 24696 53256 24696 0 _0599_
rlabel metal2 52808 22568 52808 22568 0 _0600_
rlabel metal2 52472 24248 52472 24248 0 _0601_
rlabel metal2 44352 26824 44352 26824 0 _0602_
rlabel metal2 40824 24752 40824 24752 0 _0603_
rlabel metal3 41944 24696 41944 24696 0 _0604_
rlabel metal2 41272 25200 41272 25200 0 _0605_
rlabel metal2 42392 25704 42392 25704 0 _0606_
rlabel metal3 43680 26488 43680 26488 0 _0607_
rlabel metal2 46200 28728 46200 28728 0 _0608_
rlabel metal3 51688 25368 51688 25368 0 _0609_
rlabel metal2 50232 25144 50232 25144 0 _0610_
rlabel metal3 47768 24696 47768 24696 0 _0611_
rlabel metal2 23576 26096 23576 26096 0 _0612_
rlabel metal2 42952 24920 42952 24920 0 _0613_
rlabel metal2 42784 23240 42784 23240 0 _0614_
rlabel metal2 43176 23408 43176 23408 0 _0615_
rlabel metal3 44856 24136 44856 24136 0 _0616_
rlabel metal2 44968 24584 44968 24584 0 _0617_
rlabel metal2 52920 28840 52920 28840 0 _0618_
rlabel metal2 50736 26488 50736 26488 0 _0619_
rlabel metal2 51240 28336 51240 28336 0 _0620_
rlabel metal2 44352 28056 44352 28056 0 _0621_
rlabel metal2 39928 24304 39928 24304 0 _0622_
rlabel metal2 38808 25144 38808 25144 0 _0623_
rlabel metal3 40208 25480 40208 25480 0 _0624_
rlabel metal2 39984 25592 39984 25592 0 _0625_
rlabel metal3 43344 27832 43344 27832 0 _0626_
rlabel metal3 45808 28616 45808 28616 0 _0627_
rlabel metal2 38528 25592 38528 25592 0 _0628_
rlabel metal3 42392 27160 42392 27160 0 _0629_
rlabel metal2 46424 27328 46424 27328 0 _0630_
rlabel metal2 46200 27384 46200 27384 0 _0631_
rlabel metal2 45528 27608 45528 27608 0 _0632_
rlabel metal2 45080 27160 45080 27160 0 _0633_
rlabel metal3 44520 31864 44520 31864 0 _0634_
rlabel metal2 44072 33600 44072 33600 0 _0635_
rlabel metal2 50904 29064 50904 29064 0 _0636_
rlabel metal2 43848 28896 43848 28896 0 _0637_
rlabel metal2 43512 28784 43512 28784 0 _0638_
rlabel metal2 40208 24920 40208 24920 0 _0639_
rlabel metal2 40488 27608 40488 27608 0 _0640_
rlabel metal2 40712 25704 40712 25704 0 _0641_
rlabel metal2 41160 27888 41160 27888 0 _0642_
rlabel metal2 40712 29064 40712 29064 0 _0643_
rlabel metal3 45416 29400 45416 29400 0 _0644_
rlabel metal2 51352 30464 51352 30464 0 _0645_
rlabel metal2 49112 30240 49112 30240 0 _0646_
rlabel metal2 44408 29792 44408 29792 0 _0647_
rlabel metal2 42280 28392 42280 28392 0 _0648_
rlabel metal2 42616 28896 42616 28896 0 _0649_
rlabel metal2 45304 29904 45304 29904 0 _0650_
rlabel metal2 44968 30464 44968 30464 0 _0651_
rlabel metal2 37296 27048 37296 27048 0 _0652_
rlabel metal2 36176 26488 36176 26488 0 _0653_
rlabel metal2 35896 28168 35896 28168 0 _0654_
rlabel metal2 35448 29680 35448 29680 0 _0655_
rlabel metal3 36400 28504 36400 28504 0 _0656_
rlabel metal2 35728 28728 35728 28728 0 _0657_
rlabel metal2 17472 24696 17472 24696 0 _0658_
rlabel metal2 37576 29008 37576 29008 0 _0659_
rlabel metal2 37128 29400 37128 29400 0 _0660_
rlabel metal2 38696 32704 38696 32704 0 _0661_
rlabel metal2 38584 34160 38584 34160 0 _0662_
rlabel metal2 39088 28056 39088 28056 0 _0663_
rlabel metal2 38864 27048 38864 27048 0 _0664_
rlabel metal2 38696 27552 38696 27552 0 _0665_
rlabel metal2 36344 27216 36344 27216 0 _0666_
rlabel metal3 38528 27720 38528 27720 0 _0667_
rlabel metal2 39144 27664 39144 27664 0 _0668_
rlabel metal3 40488 30184 40488 30184 0 _0669_
rlabel metal3 35840 26936 35840 26936 0 _0670_
rlabel metal2 34440 27384 34440 27384 0 _0671_
rlabel metal2 33320 28056 33320 28056 0 _0672_
rlabel metal3 34832 29400 34832 29400 0 _0673_
rlabel metal2 33320 28840 33320 28840 0 _0674_
rlabel metal2 34104 29848 34104 29848 0 _0675_
rlabel metal2 33936 29400 33936 29400 0 _0676_
rlabel metal3 30296 29512 30296 29512 0 _0677_
rlabel metal2 23464 29512 23464 29512 0 _0678_
rlabel metal2 26824 31864 26824 31864 0 _0679_
rlabel metal2 31640 29008 31640 29008 0 _0680_
rlabel metal2 31920 28056 31920 28056 0 _0681_
rlabel metal3 24584 27048 24584 27048 0 _0682_
rlabel metal2 32480 27160 32480 27160 0 _0683_
rlabel metal3 32424 26936 32424 26936 0 _0684_
rlabel metal2 33096 27440 33096 27440 0 _0685_
rlabel metal3 29792 27832 29792 27832 0 _0686_
rlabel metal2 27216 28840 27216 28840 0 _0687_
rlabel metal3 24976 26488 24976 26488 0 _0688_
rlabel metal2 23744 27944 23744 27944 0 _0689_
rlabel metal2 24696 31360 24696 31360 0 _0690_
rlabel metal2 23744 30296 23744 30296 0 _0691_
rlabel metal2 22568 30408 22568 30408 0 _0692_
rlabel metal2 22456 30352 22456 30352 0 _0693_
rlabel metal2 24136 30800 24136 30800 0 _0694_
rlabel metal2 22904 34552 22904 34552 0 _0695_
rlabel metal2 23240 31808 23240 31808 0 _0696_
rlabel metal2 23240 31192 23240 31192 0 _0697_
rlabel metal2 22624 30856 22624 30856 0 _0698_
rlabel metal3 20888 27048 20888 27048 0 _0699_
rlabel metal3 22008 26488 22008 26488 0 _0700_
rlabel metal3 22064 27832 22064 27832 0 _0701_
rlabel metal2 22232 28056 22232 28056 0 _0702_
rlabel metal3 22064 29624 22064 29624 0 _0703_
rlabel metal2 21448 27440 21448 27440 0 _0704_
rlabel metal2 19208 28224 19208 28224 0 _0705_
rlabel metal2 18984 30520 18984 30520 0 _0706_
rlabel metal2 18312 29064 18312 29064 0 _0707_
rlabel metal2 18032 28840 18032 28840 0 _0708_
rlabel metal2 18648 28952 18648 28952 0 _0709_
rlabel metal2 17640 29624 17640 29624 0 _0710_
rlabel metal2 16464 30072 16464 30072 0 _0711_
rlabel metal2 17080 30576 17080 30576 0 _0712_
rlabel metal2 18088 28280 18088 28280 0 _0713_
rlabel metal2 18928 26488 18928 26488 0 _0714_
rlabel metal2 19320 27160 19320 27160 0 _0715_
rlabel metal2 18648 27552 18648 27552 0 _0716_
rlabel metal2 17752 26264 17752 26264 0 _0717_
rlabel metal3 17136 26264 17136 26264 0 _0718_
rlabel metal2 14728 21952 14728 21952 0 _0719_
rlabel metal2 8008 29792 8008 29792 0 _0720_
rlabel metal2 8624 27608 8624 27608 0 _0721_
rlabel metal4 9912 21336 9912 21336 0 _0722_
rlabel metal2 9016 18648 9016 18648 0 _0723_
rlabel metal3 7952 17528 7952 17528 0 _0724_
rlabel metal2 9128 16968 9128 16968 0 _0725_
rlabel metal2 9408 17416 9408 17416 0 _0726_
rlabel metal3 9296 15176 9296 15176 0 _0727_
rlabel metal2 11032 15736 11032 15736 0 _0728_
rlabel metal2 12824 15736 12824 15736 0 _0729_
rlabel metal2 14728 15624 14728 15624 0 _0730_
rlabel metal2 15176 15848 15176 15848 0 _0731_
rlabel metal2 16352 16968 16352 16968 0 _0732_
rlabel metal2 16856 16016 16856 16016 0 _0733_
rlabel metal2 16184 18480 16184 18480 0 _0734_
rlabel metal2 15400 19712 15400 19712 0 _0735_
rlabel metal2 14560 26936 14560 26936 0 _0736_
rlabel metal2 14000 26712 14000 26712 0 _0737_
rlabel metal2 14168 27664 14168 27664 0 _0738_
rlabel metal2 13608 28280 13608 28280 0 _0739_
rlabel metal2 12544 28616 12544 28616 0 _0740_
rlabel metal2 13048 28336 13048 28336 0 _0741_
rlabel metal2 16968 34272 16968 34272 0 _0742_
rlabel metal2 15400 37744 15400 37744 0 _0743_
rlabel metal2 16016 24808 16016 24808 0 _0744_
rlabel metal2 14952 26600 14952 26600 0 _0745_
rlabel metal2 15624 24976 15624 24976 0 _0746_
rlabel metal2 12936 20384 12936 20384 0 _0747_
rlabel metal2 10808 30688 10808 30688 0 _0748_
rlabel metal2 12096 30968 12096 30968 0 _0749_
rlabel metal2 12600 31360 12600 31360 0 _0750_
rlabel metal2 7224 33600 7224 33600 0 _0751_
rlabel metal2 11704 32032 11704 32032 0 _0752_
rlabel metal2 10248 32200 10248 32200 0 _0753_
rlabel metal2 10360 25760 10360 25760 0 _0754_
rlabel metal2 9968 25368 9968 25368 0 _0755_
rlabel metal2 7560 20104 7560 20104 0 _0756_
rlabel metal2 8736 29624 8736 29624 0 _0757_
rlabel metal2 7952 31640 7952 31640 0 _0758_
rlabel metal2 7672 31920 7672 31920 0 _0759_
rlabel metal3 9296 32536 9296 32536 0 _0760_
rlabel metal2 8120 33432 8120 33432 0 _0761_
rlabel metal2 10248 27608 10248 27608 0 _0762_
rlabel metal2 9968 29624 9968 29624 0 _0763_
rlabel metal2 9688 31080 9688 31080 0 _0764_
rlabel metal2 9464 31808 9464 31808 0 _0765_
rlabel metal2 6048 31864 6048 31864 0 _0766_
rlabel metal2 6776 33320 6776 33320 0 _0767_
rlabel metal2 2520 11928 2520 11928 0 _0768_
rlabel metal2 3304 27440 3304 27440 0 _0769_
rlabel metal3 9408 30184 9408 30184 0 _0770_
rlabel metal2 9016 31360 9016 31360 0 _0771_
rlabel metal2 5096 31584 5096 31584 0 _0772_
rlabel metal2 3640 31696 3640 31696 0 _0773_
rlabel metal2 4088 31752 4088 31752 0 _0774_
rlabel metal2 7112 26544 7112 26544 0 _0775_
rlabel metal2 7616 29400 7616 29400 0 _0776_
rlabel metal2 6384 29288 6384 29288 0 _0777_
rlabel metal2 6104 29904 6104 29904 0 _0778_
rlabel metal2 2856 30856 2856 30856 0 _0779_
rlabel metal2 5656 28224 5656 28224 0 _0780_
rlabel metal2 4760 31360 4760 31360 0 _0781_
rlabel metal2 16520 21896 16520 21896 0 _0782_
rlabel metal3 4984 23688 4984 23688 0 _0783_
rlabel metal2 7672 28728 7672 28728 0 _0784_
rlabel metal2 6496 28616 6496 28616 0 _0785_
rlabel metal3 5544 27944 5544 27944 0 _0786_
rlabel metal2 4648 28168 4648 28168 0 _0787_
rlabel metal2 4312 29456 4312 29456 0 _0788_
rlabel metal2 9016 27272 9016 27272 0 _0789_
rlabel metal2 8232 26544 8232 26544 0 _0790_
rlabel metal2 8008 26432 8008 26432 0 _0791_
rlabel metal2 6440 27104 6440 27104 0 _0792_
rlabel metal2 4648 27104 4648 27104 0 _0793_
rlabel metal3 4760 27832 4760 27832 0 _0794_
rlabel metal2 3976 21896 3976 21896 0 _0795_
rlabel metal2 9688 26992 9688 26992 0 _0796_
rlabel metal3 8456 26152 8456 26152 0 _0797_
rlabel metal2 6664 26208 6664 26208 0 _0798_
rlabel metal2 3752 25760 3752 25760 0 _0799_
rlabel metal2 4312 26152 4312 26152 0 _0800_
rlabel metal2 11816 23072 11816 23072 0 _0801_
rlabel metal2 9128 19992 9128 19992 0 _0802_
rlabel metal2 13608 23184 13608 23184 0 _0803_
rlabel metal2 11424 19768 11424 19768 0 _0804_
rlabel metal2 11256 20888 11256 20888 0 _0805_
rlabel metal2 11424 21672 11424 21672 0 _0806_
rlabel metal2 11480 22848 11480 22848 0 _0807_
rlabel metal2 13384 10416 13384 10416 0 _0808_
rlabel metal2 12768 10696 12768 10696 0 _0809_
rlabel metal3 11704 22456 11704 22456 0 _0810_
rlabel metal2 5880 18592 5880 18592 0 _0811_
rlabel metal2 13048 17528 13048 17528 0 _0812_
rlabel metal2 10584 19768 10584 19768 0 _0813_
rlabel metal2 8680 21112 8680 21112 0 _0814_
rlabel metal2 7784 21112 7784 21112 0 _0815_
rlabel metal2 6664 21952 6664 21952 0 _0816_
rlabel metal2 3304 22232 3304 22232 0 _0817_
rlabel metal2 3752 23576 3752 23576 0 _0818_
rlabel metal3 5488 24808 5488 24808 0 _0819_
rlabel metal2 5768 24640 5768 24640 0 _0820_
rlabel metal2 8904 21728 8904 21728 0 _0821_
rlabel metal2 9016 21728 9016 21728 0 _0822_
rlabel metal3 9464 23128 9464 23128 0 _0823_
rlabel metal3 8568 23240 8568 23240 0 _0824_
rlabel metal3 4648 23128 4648 23128 0 _0825_
rlabel metal2 3864 16856 3864 16856 0 _0826_
rlabel metal2 8568 21280 8568 21280 0 _0827_
rlabel metal2 9800 20888 9800 20888 0 _0828_
rlabel metal2 6272 20664 6272 20664 0 _0829_
rlabel metal2 5992 20832 5992 20832 0 _0830_
rlabel metal2 4368 20888 4368 20888 0 _0831_
rlabel metal2 4536 21616 4536 21616 0 _0832_
rlabel metal2 7896 19040 7896 19040 0 _0833_
rlabel metal2 6552 19376 6552 19376 0 _0834_
rlabel metal2 6104 18704 6104 18704 0 _0835_
rlabel metal2 5768 18368 5768 18368 0 _0836_
rlabel metal2 4088 19600 4088 19600 0 _0837_
rlabel metal2 4872 20272 4872 20272 0 _0838_
rlabel metal2 3304 15120 3304 15120 0 _0839_
rlabel metal2 8344 15120 8344 15120 0 _0840_
rlabel metal2 8008 18256 8008 18256 0 _0841_
rlabel metal2 6552 18088 6552 18088 0 _0842_
rlabel metal2 4424 18368 4424 18368 0 _0843_
rlabel metal2 4088 17696 4088 17696 0 _0844_
rlabel metal2 3640 17752 3640 17752 0 _0845_
rlabel metal2 5992 15680 5992 15680 0 _0846_
rlabel metal2 7784 17752 7784 17752 0 _0847_
rlabel metal2 16184 16688 16184 16688 0 _0848_
rlabel metal2 6832 17864 6832 17864 0 _0849_
rlabel metal2 6384 15960 6384 15960 0 _0850_
rlabel metal3 5320 15288 5320 15288 0 _0851_
rlabel metal3 3584 15288 3584 15288 0 _0852_
rlabel metal2 5096 15204 5096 15204 0 _0853_
rlabel metal2 4760 15624 4760 15624 0 _0854_
rlabel metal2 6216 10528 6216 10528 0 _0855_
rlabel metal2 8008 15568 8008 15568 0 _0856_
rlabel metal2 6664 15148 6664 15148 0 _0857_
rlabel metal2 5544 14224 5544 14224 0 _0858_
rlabel metal2 3304 13216 3304 13216 0 _0859_
rlabel metal2 3864 13608 3864 13608 0 _0860_
rlabel metal3 7728 15288 7728 15288 0 _0861_
rlabel metal2 8120 14560 8120 14560 0 _0862_
rlabel metal2 6384 12264 6384 12264 0 _0863_
rlabel metal2 6104 11648 6104 11648 0 _0864_
rlabel metal2 3192 11816 3192 11816 0 _0865_
rlabel metal2 3864 12432 3864 12432 0 _0866_
rlabel metal2 5936 9800 5936 9800 0 _0867_
rlabel metal2 6720 14280 6720 14280 0 _0868_
rlabel metal2 7112 12544 7112 12544 0 _0869_
rlabel metal2 6776 11312 6776 11312 0 _0870_
rlabel metal2 6272 9800 6272 9800 0 _0871_
rlabel metal2 5544 9856 5544 9856 0 _0872_
rlabel metal2 8008 13328 8008 13328 0 _0873_
rlabel metal2 8456 12544 8456 12544 0 _0874_
rlabel metal2 9240 11816 9240 11816 0 _0875_
rlabel metal2 7784 10248 7784 10248 0 _0876_
rlabel metal2 6328 8904 6328 8904 0 _0877_
rlabel metal2 15512 12264 15512 12264 0 _0878_
rlabel metal2 10080 14392 10080 14392 0 _0879_
rlabel metal2 9968 12264 9968 12264 0 _0880_
rlabel metal2 9016 11200 9016 11200 0 _0881_
rlabel metal2 9576 9520 9576 9520 0 _0882_
rlabel metal2 15960 8736 15960 8736 0 _0883_
rlabel metal2 10416 8232 10416 8232 0 _0884_
rlabel metal2 11984 10024 11984 10024 0 _0885_
rlabel metal2 11424 15960 11424 15960 0 _0886_
rlabel metal2 11144 15148 11144 15148 0 _0887_
rlabel metal2 11704 11144 11704 11144 0 _0888_
rlabel metal2 11704 11592 11704 11592 0 _0889_
rlabel metal2 16632 12040 16632 12040 0 _0890_
rlabel metal2 14392 16072 14392 16072 0 _0891_
rlabel metal2 11816 15232 11816 15232 0 _0892_
rlabel metal3 13048 13160 13048 13160 0 _0893_
rlabel metal2 12992 9800 12992 9800 0 _0894_
rlabel metal2 12040 8512 12040 8512 0 _0895_
rlabel metal2 12600 8512 12600 8512 0 _0896_
rlabel metal2 14392 10472 14392 10472 0 _0897_
rlabel metal3 13440 15288 13440 15288 0 _0898_
rlabel metal2 13160 14112 13160 14112 0 _0899_
rlabel metal2 13776 11368 13776 11368 0 _0900_
rlabel metal2 13608 10640 13608 10640 0 _0901_
rlabel metal2 14280 14448 14280 14448 0 _0902_
rlabel metal2 14504 12936 14504 12936 0 _0903_
rlabel metal2 14504 12040 14504 12040 0 _0904_
rlabel metal2 13496 9912 13496 9912 0 _0905_
rlabel metal2 14168 8232 14168 8232 0 _0906_
rlabel metal3 14112 19096 14112 19096 0 _0907_
rlabel metal2 13384 17416 13384 17416 0 _0908_
rlabel metal2 14952 18032 14952 18032 0 _0909_
rlabel metal3 14504 18200 14504 18200 0 _0910_
rlabel metal2 14224 15736 14224 15736 0 _0911_
rlabel metal2 20104 12376 20104 12376 0 _0912_
rlabel metal2 15008 16184 15008 16184 0 _0913_
rlabel metal2 15904 12264 15904 12264 0 _0914_
rlabel metal2 15960 10584 15960 10584 0 _0915_
rlabel metal3 17248 9800 17248 9800 0 _0916_
rlabel metal3 16688 9240 16688 9240 0 _0917_
rlabel metal2 17080 18088 17080 18088 0 _0918_
rlabel metal2 16296 15624 16296 15624 0 _0919_
rlabel metal2 18312 13944 18312 13944 0 _0920_
rlabel metal2 18032 12264 18032 12264 0 _0921_
rlabel metal2 17920 10808 17920 10808 0 _0922_
rlabel metal2 18648 13552 18648 13552 0 _0923_
rlabel metal2 18536 10304 18536 10304 0 _0924_
rlabel metal2 17080 15484 17080 15484 0 _0925_
rlabel metal3 18928 14392 18928 14392 0 _0926_
rlabel metal2 19488 12936 19488 12936 0 _0927_
rlabel metal3 19432 12376 19432 12376 0 _0928_
rlabel metal2 20440 12040 20440 12040 0 _0929_
rlabel metal3 17192 15176 17192 15176 0 _0930_
rlabel metal3 18648 14504 18648 14504 0 _0931_
rlabel metal2 19096 15008 19096 15008 0 _0932_
rlabel metal2 20328 13720 20328 13720 0 _0933_
rlabel metal2 19544 12432 19544 12432 0 _0934_
rlabel metal2 16408 18704 16408 18704 0 _0935_
rlabel metal2 16520 18760 16520 18760 0 _0936_
rlabel metal2 17640 19264 17640 19264 0 _0937_
rlabel metal2 18984 18704 18984 18704 0 _0938_
rlabel metal2 19096 17304 19096 17304 0 _0939_
rlabel metal2 14504 20552 14504 20552 0 _0940_
rlabel metal2 14952 21224 14952 21224 0 _0941_
rlabel metal2 18200 21616 18200 21616 0 _0942_
rlabel metal3 17136 21672 17136 21672 0 _0943_
rlabel metal2 15624 22008 15624 22008 0 _0944_
rlabel metal2 31528 39480 31528 39480 0 _0945_
rlabel metal2 32536 43120 32536 43120 0 _0946_
rlabel metal2 8568 40096 8568 40096 0 _0947_
rlabel metal2 8344 41272 8344 41272 0 _0948_
rlabel metal2 8624 40600 8624 40600 0 _0949_
rlabel metal2 10416 39816 10416 39816 0 _0950_
rlabel metal2 28952 26488 28952 26488 0 _0951_
rlabel metal2 21672 41944 21672 41944 0 _0952_
rlabel metal3 20440 43624 20440 43624 0 _0953_
rlabel metal2 41832 37128 41832 37128 0 _0954_
rlabel metal2 38248 40824 38248 40824 0 _0955_
rlabel metal3 19936 41944 19936 41944 0 _0956_
rlabel metal2 41272 41328 41272 41328 0 _0957_
rlabel metal2 30408 43848 30408 43848 0 _0958_
rlabel metal2 29512 40824 29512 40824 0 _0959_
rlabel metal3 24584 42616 24584 42616 0 _0960_
rlabel metal3 30352 26264 30352 26264 0 _0961_
rlabel metal2 31304 27384 31304 27384 0 _0962_
rlabel metal2 29960 41328 29960 41328 0 _0963_
rlabel metal2 11480 37632 11480 37632 0 _0964_
rlabel metal3 43624 37464 43624 37464 0 _0965_
rlabel metal3 33656 39368 33656 39368 0 _0966_
rlabel metal3 34944 34664 34944 34664 0 _0967_
rlabel metal2 34104 36456 34104 36456 0 _0968_
rlabel metal2 32312 39872 32312 39872 0 _0969_
rlabel metal2 32424 40880 32424 40880 0 _0970_
rlabel metal2 20216 46368 20216 46368 0 _0971_
rlabel metal2 36232 38864 36232 38864 0 _0972_
rlabel metal2 24584 44464 24584 44464 0 _0973_
rlabel metal2 20552 43176 20552 43176 0 _0974_
rlabel metal2 21448 42728 21448 42728 0 _0975_
rlabel metal3 40516 42616 40516 42616 0 _0976_
rlabel metal2 20216 41384 20216 41384 0 _0977_
rlabel metal2 19992 43680 19992 43680 0 _0978_
rlabel metal3 25256 43624 25256 43624 0 _0979_
rlabel metal2 29624 20552 29624 20552 0 _0980_
rlabel metal2 28056 22568 28056 22568 0 _0981_
rlabel metal2 47880 43120 47880 43120 0 _0982_
rlabel metal2 24360 36288 24360 36288 0 _0983_
rlabel metal2 30632 36456 30632 36456 0 _0984_
rlabel metal2 42056 42168 42056 42168 0 _0985_
rlabel metal2 30856 35952 30856 35952 0 _0986_
rlabel metal2 30968 37408 30968 37408 0 _0987_
rlabel metal2 28280 45528 28280 45528 0 _0988_
rlabel metal3 21168 45864 21168 45864 0 _0989_
rlabel metal3 22792 45696 22792 45696 0 _0990_
rlabel metal2 27944 20384 27944 20384 0 _0991_
rlabel metal2 30128 20776 30128 20776 0 _0992_
rlabel metal2 29960 26376 29960 26376 0 _0993_
rlabel metal2 29064 27776 29064 27776 0 _0994_
rlabel metal3 28840 28056 28840 28056 0 _0995_
rlabel metal2 28728 30632 28728 30632 0 _0996_
rlabel metal2 23016 41888 23016 41888 0 _0997_
rlabel metal2 25368 47096 25368 47096 0 _0998_
rlabel metal3 21336 48888 21336 48888 0 _0999_
rlabel metal2 22680 41160 22680 41160 0 _1000_
rlabel metal3 25368 42504 25368 42504 0 _1001_
rlabel metal3 23744 41160 23744 41160 0 _1002_
rlabel metal2 24640 41048 24640 41048 0 _1003_
rlabel metal2 25592 16464 25592 16464 0 _1004_
rlabel metal2 26152 21560 26152 21560 0 _1005_
rlabel metal2 26656 35896 26656 35896 0 _1006_
rlabel metal2 26824 16520 26824 16520 0 _1007_
rlabel metal2 26320 35672 26320 35672 0 _1008_
rlabel metal2 25536 38920 25536 38920 0 _1009_
rlabel metal3 26264 40320 26264 40320 0 _1010_
rlabel metal2 23240 43848 23240 43848 0 _1011_
rlabel metal2 22568 50876 22568 50876 0 _1012_
rlabel metal2 23576 41328 23576 41328 0 _1013_
rlabel metal2 23576 42728 23576 42728 0 _1014_
rlabel metal2 23352 41440 23352 41440 0 _1015_
rlabel metal3 28616 16968 28616 16968 0 _1016_
rlabel metal2 26824 35280 26824 35280 0 _1017_
rlabel metal2 26488 36848 26488 36848 0 _1018_
rlabel metal3 25032 39928 25032 39928 0 _1019_
rlabel metal2 38696 40656 38696 40656 0 _1020_
rlabel metal2 24248 44352 24248 44352 0 _1021_
rlabel metal2 23744 44408 23744 44408 0 _1022_
rlabel metal2 26264 46984 26264 46984 0 _1023_
rlabel metal2 25592 11508 25592 11508 0 _1024_
rlabel metal2 20272 24360 20272 24360 0 _1025_
rlabel metal3 28448 37240 28448 37240 0 _1026_
rlabel metal2 28504 36792 28504 36792 0 _1027_
rlabel metal2 28952 37968 28952 37968 0 _1028_
rlabel metal2 42840 38472 42840 38472 0 _1029_
rlabel metal2 38920 44800 38920 44800 0 _1030_
rlabel metal2 26376 47096 26376 47096 0 _1031_
rlabel metal2 37912 45136 37912 45136 0 _1032_
rlabel metal2 38136 40376 38136 40376 0 _1033_
rlabel metal2 37576 22512 37576 22512 0 _1034_
rlabel metal2 37128 22008 37128 22008 0 _1035_
rlabel metal2 37352 37744 37352 37744 0 _1036_
rlabel metal2 37408 40264 37408 40264 0 _1037_
rlabel metal2 36736 38360 36736 38360 0 _1038_
rlabel metal2 37016 38416 37016 38416 0 _1039_
rlabel metal2 35896 10472 35896 10472 0 _1040_
rlabel metal2 34496 10696 34496 10696 0 _1041_
rlabel metal2 24808 36680 24808 36680 0 _1042_
rlabel metal2 36120 32312 36120 32312 0 _1043_
rlabel metal2 36512 33992 36512 33992 0 _1044_
rlabel metal2 34608 35896 34608 35896 0 _1045_
rlabel metal2 21224 16632 21224 16632 0 _1046_
rlabel metal3 34944 36344 34944 36344 0 _1047_
rlabel metal2 25928 40488 25928 40488 0 _1048_
rlabel metal3 35392 36232 35392 36232 0 _1049_
rlabel metal3 31024 49896 31024 49896 0 _1050_
rlabel metal2 40936 46704 40936 46704 0 _1051_
rlabel metal2 32312 46480 32312 46480 0 _1052_
rlabel metal2 33880 45024 33880 45024 0 _1053_
rlabel metal2 34496 41048 34496 41048 0 _1054_
rlabel metal3 42280 36456 42280 36456 0 _1055_
rlabel metal2 31696 45080 31696 45080 0 _1056_
rlabel metal2 32984 44688 32984 44688 0 _1057_
rlabel metal2 35000 44184 35000 44184 0 _1058_
rlabel metal2 37240 11592 37240 11592 0 _1059_
rlabel metal2 37016 10752 37016 10752 0 _1060_
rlabel metal2 34944 34888 34944 34888 0 _1061_
rlabel metal2 36176 35000 36176 35000 0 _1062_
rlabel metal2 35784 40208 35784 40208 0 _1063_
rlabel metal2 34440 33264 34440 33264 0 _1064_
rlabel metal2 34328 33488 34328 33488 0 _1065_
rlabel metal3 35840 36344 35840 36344 0 _1066_
rlabel metal2 33432 43680 33432 43680 0 _1067_
rlabel metal2 33656 44352 33656 44352 0 _1068_
rlabel metal3 33880 43624 33880 43624 0 _1069_
rlabel metal3 35112 42728 35112 42728 0 _1070_
rlabel metal2 33208 47712 33208 47712 0 _1071_
rlabel metal2 33320 48664 33320 48664 0 _1072_
rlabel metal2 34104 48552 34104 48552 0 _1073_
rlabel metal2 38808 10360 38808 10360 0 _1074_
rlabel metal2 36120 33712 36120 33712 0 _1075_
rlabel metal2 35336 32592 35336 32592 0 _1076_
rlabel metal3 35336 47208 35336 47208 0 _1077_
rlabel metal2 41832 22792 41832 22792 0 _1078_
rlabel metal3 40488 11144 40488 11144 0 _1079_
rlabel metal2 38360 22176 38360 22176 0 _1080_
rlabel metal2 41160 34608 41160 34608 0 _1081_
rlabel metal2 41832 35672 41832 35672 0 _1082_
rlabel metal2 41496 35728 41496 35728 0 _1083_
rlabel metal3 45528 36344 45528 36344 0 _1084_
rlabel metal2 42000 35896 42000 35896 0 _1085_
rlabel metal2 45752 42560 45752 42560 0 _1086_
rlabel metal2 40152 47712 40152 47712 0 _1087_
rlabel metal2 40376 46592 40376 46592 0 _1088_
rlabel metal2 41832 44632 41832 44632 0 _1089_
rlabel metal2 42504 41608 42504 41608 0 _1090_
rlabel metal2 42112 38808 42112 38808 0 _1091_
rlabel metal3 40544 45976 40544 45976 0 _1092_
rlabel metal2 41832 40656 41832 40656 0 _1093_
rlabel metal2 42504 20552 42504 20552 0 _1094_
rlabel metal2 43288 21728 43288 21728 0 _1095_
rlabel metal2 50344 35560 50344 35560 0 _1096_
rlabel metal2 42168 34328 42168 34328 0 _1097_
rlabel metal2 42952 38724 42952 38724 0 _1098_
rlabel metal2 42616 38864 42616 38864 0 _1099_
rlabel metal2 45080 22176 45080 22176 0 _1100_
rlabel metal3 41720 22624 41720 22624 0 _1101_
rlabel metal3 45920 23016 45920 23016 0 _1102_
rlabel metal3 42000 40600 42000 40600 0 _1103_
rlabel metal2 42168 42000 42168 42000 0 _1104_
rlabel metal2 42000 46648 42000 46648 0 _1105_
rlabel metal2 43736 46144 43736 46144 0 _1106_
rlabel metal2 43512 45136 43512 45136 0 _1107_
rlabel metal2 43624 48160 43624 48160 0 _1108_
rlabel metal2 42672 42728 42672 42728 0 _1109_
rlabel metal2 42952 43680 42952 43680 0 _1110_
rlabel metal2 42896 42728 42896 42728 0 _1111_
rlabel metal2 39704 41832 39704 41832 0 _1112_
rlabel metal3 46984 23912 46984 23912 0 _1113_
rlabel metal3 43680 40264 43680 40264 0 _1114_
rlabel metal3 45360 39592 45360 39592 0 _1115_
rlabel metal2 45080 41776 45080 41776 0 _1116_
rlabel metal2 43736 44800 43736 44800 0 _1117_
rlabel metal3 43568 44968 43568 44968 0 _1118_
rlabel metal2 45192 42000 45192 42000 0 _1119_
rlabel metal2 45304 39872 45304 39872 0 _1120_
rlabel metal2 48776 26208 48776 26208 0 _1121_
rlabel metal4 46088 28896 46088 28896 0 _1122_
rlabel metal2 48048 35784 48048 35784 0 _1123_
rlabel metal3 46704 36232 46704 36232 0 _1124_
rlabel metal3 46424 37352 46424 37352 0 _1125_
rlabel metal3 46872 38024 46872 38024 0 _1126_
rlabel metal2 46536 38668 46536 38668 0 _1127_
rlabel metal3 46816 38584 46816 38584 0 _1128_
rlabel metal2 47320 45808 47320 45808 0 _1129_
rlabel metal2 45304 46088 45304 46088 0 _1130_
rlabel metal2 46536 44688 46536 44688 0 _1131_
rlabel metal2 46312 43176 46312 43176 0 _1132_
rlabel metal2 46816 43400 46816 43400 0 _1133_
rlabel metal3 47152 20552 47152 20552 0 _1134_
rlabel metal2 46760 41440 46760 41440 0 _1135_
rlabel metal2 47040 36568 47040 36568 0 _1136_
rlabel metal2 47432 39788 47432 39788 0 _1137_
rlabel metal3 47936 46872 47936 46872 0 _1138_
rlabel metal2 47544 43120 47544 43120 0 _1139_
rlabel metal2 48104 42672 48104 42672 0 _1140_
rlabel metal2 47992 41440 47992 41440 0 _1141_
rlabel metal2 49112 26320 49112 26320 0 _1142_
rlabel metal2 47152 34216 47152 34216 0 _1143_
rlabel metal2 47656 34832 47656 34832 0 _1144_
rlabel metal2 47544 34832 47544 34832 0 _1145_
rlabel metal2 48328 35336 48328 35336 0 _1146_
rlabel metal3 48384 36232 48384 36232 0 _1147_
rlabel metal2 47096 44184 47096 44184 0 _1148_
rlabel metal2 47880 44184 47880 44184 0 _1149_
rlabel metal2 47768 25200 47768 25200 0 _1150_
rlabel metal2 48888 35000 48888 35000 0 _1151_
rlabel metal2 49168 41272 49168 41272 0 _1152_
rlabel metal3 43904 42504 43904 42504 0 _1153_
rlabel metal2 48720 43624 48720 43624 0 _1154_
rlabel metal2 49112 44072 49112 44072 0 _1155_
rlabel metal2 49448 43624 49448 43624 0 _1156_
rlabel metal2 49560 42224 49560 42224 0 _1157_
rlabel metal3 47880 27888 47880 27888 0 _1158_
rlabel metal2 48160 24136 48160 24136 0 _1159_
rlabel metal2 48664 24080 48664 24080 0 _1160_
rlabel metal2 51352 36848 51352 36848 0 _1161_
rlabel metal2 52696 36120 52696 36120 0 _1162_
rlabel metal2 52808 36904 52808 36904 0 _1163_
rlabel metal3 46704 45752 46704 45752 0 _1164_
rlabel metal3 52528 45640 52528 45640 0 _1165_
rlabel metal3 53816 43624 53816 43624 0 _1166_
rlabel metal2 50456 42952 50456 42952 0 _1167_
rlabel metal2 52080 40376 52080 40376 0 _1168_
rlabel metal2 19544 36512 19544 36512 0 _1169_
rlabel metal2 53032 42560 53032 42560 0 _1170_
rlabel metal3 54880 40600 54880 40600 0 _1171_
rlabel metal2 52920 33544 52920 33544 0 _1172_
rlabel metal2 52920 34048 52920 34048 0 _1173_
rlabel metal2 52920 38724 52920 38724 0 _1174_
rlabel metal2 53312 39032 53312 39032 0 _1175_
rlabel metal3 52080 32536 52080 32536 0 _1176_
rlabel metal2 52584 33208 52584 33208 0 _1177_
rlabel metal2 51016 35280 51016 35280 0 _1178_
rlabel metal2 51688 36568 51688 36568 0 _1179_
rlabel metal2 51408 34888 51408 34888 0 _1180_
rlabel metal2 51800 36736 51800 36736 0 _1181_
rlabel metal2 50960 44408 50960 44408 0 _1182_
rlabel metal2 51688 44968 51688 44968 0 _1183_
rlabel metal3 50148 43288 50148 43288 0 _1184_
rlabel metal2 51800 41160 51800 41160 0 _1185_
rlabel metal2 51352 42672 51352 42672 0 _1186_
rlabel metal2 51576 41496 51576 41496 0 _1187_
rlabel metal3 52528 33432 52528 33432 0 _1188_
rlabel metal3 52248 34888 52248 34888 0 _1189_
rlabel metal2 52696 35336 52696 35336 0 _1190_
rlabel metal2 52248 39312 52248 39312 0 _1191_
rlabel metal3 40040 34664 40040 34664 0 _1192_
rlabel metal2 39256 34832 39256 34832 0 _1193_
rlabel metal2 39816 37016 39816 37016 0 _1194_
rlabel metal2 40152 37520 40152 37520 0 _1195_
rlabel metal3 40208 37128 40208 37128 0 _1196_
rlabel metal2 39480 37856 39480 37856 0 _1197_
rlabel metal2 40264 43904 40264 43904 0 _1198_
rlabel metal2 40152 43008 40152 43008 0 _1199_
rlabel metal2 40488 40600 40488 40600 0 _1200_
rlabel metal2 39704 35056 39704 35056 0 _1201_
rlabel metal2 18760 40712 18760 40712 0 _1202_
rlabel metal3 39928 36456 39928 36456 0 _1203_
rlabel metal2 39872 40600 39872 40600 0 _1204_
rlabel metal2 39368 43568 39368 43568 0 _1205_
rlabel metal2 39032 43008 39032 43008 0 _1206_
rlabel metal2 39256 42000 39256 42000 0 _1207_
rlabel metal2 26712 42784 26712 42784 0 _1208_
rlabel metal2 26264 45136 26264 45136 0 _1209_
rlabel metal4 26712 41384 26712 41384 0 _1210_
rlabel metal2 26712 41832 26712 41832 0 _1211_
rlabel metal2 26936 41160 26936 41160 0 _1212_
rlabel metal2 27832 30856 27832 30856 0 _1213_
rlabel metal3 38724 34664 38724 34664 0 _1214_
rlabel metal2 28336 35672 28336 35672 0 _1215_
rlabel metal2 26544 40264 26544 40264 0 _1216_
rlabel metal2 29904 35000 29904 35000 0 _1217_
rlabel metal2 30296 35000 30296 35000 0 _1218_
rlabel metal2 30240 35784 30240 35784 0 _1219_
rlabel metal2 27272 44520 27272 44520 0 _1220_
rlabel metal3 28504 43624 28504 43624 0 _1221_
rlabel metal2 29736 39592 29736 39592 0 _1222_
rlabel metal2 24360 42784 24360 42784 0 _1223_
rlabel metal2 14504 43904 14504 43904 0 _1224_
rlabel metal2 25648 39032 25648 39032 0 _1225_
rlabel metal2 25704 40936 25704 40936 0 _1226_
rlabel metal2 25928 39592 25928 39592 0 _1227_
rlabel metal2 23016 31416 23016 31416 0 _1228_
rlabel metal2 23576 36960 23576 36960 0 _1229_
rlabel metal2 25480 35952 25480 35952 0 _1230_
rlabel metal2 25592 36904 25592 36904 0 _1231_
rlabel metal2 25480 38668 25480 38668 0 _1232_
rlabel metal2 22232 30296 22232 30296 0 _1233_
rlabel metal2 23912 35896 23912 35896 0 _1234_
rlabel metal2 24360 38360 24360 38360 0 _1235_
rlabel metal3 26824 43400 26824 43400 0 _1236_
rlabel metal2 28168 43008 28168 43008 0 _1237_
rlabel metal2 28616 40264 28616 40264 0 _1238_
rlabel metal2 18088 31472 18088 31472 0 _1239_
rlabel metal2 21336 37184 21336 37184 0 _1240_
rlabel metal2 19824 36456 19824 36456 0 _1241_
rlabel metal2 20272 36456 20272 36456 0 _1242_
rlabel metal3 18648 42616 18648 42616 0 _1243_
rlabel metal2 19544 41832 19544 41832 0 _1244_
rlabel metal2 19432 40544 19432 40544 0 _1245_
rlabel metal2 19544 39452 19544 39452 0 _1246_
rlabel metal2 19096 40656 19096 40656 0 _1247_
rlabel metal3 26544 39480 26544 39480 0 _1248_
rlabel metal2 16856 32928 16856 32928 0 _1249_
rlabel metal3 27664 34776 27664 34776 0 _1250_
rlabel metal2 31920 34888 31920 34888 0 _1251_
rlabel metal2 32984 35280 32984 35280 0 _1252_
rlabel metal2 34552 39312 34552 39312 0 _1253_
rlabel metal2 6384 38584 6384 38584 0 _1254_
rlabel metal2 5880 38612 5880 38612 0 _1255_
rlabel metal2 8232 41440 8232 41440 0 _1256_
rlabel metal3 8176 42616 8176 42616 0 _1257_
rlabel metal2 7672 41832 7672 41832 0 _1258_
rlabel metal2 6216 42448 6216 42448 0 _1259_
rlabel metal2 5432 42616 5432 42616 0 _1260_
rlabel metal2 7112 42112 7112 42112 0 _1261_
rlabel metal2 3976 42336 3976 42336 0 _1262_
rlabel metal2 4088 43120 4088 43120 0 _1263_
rlabel metal2 4984 42616 4984 42616 0 _1264_
rlabel metal2 6216 41552 6216 41552 0 _1265_
rlabel metal2 6552 40320 6552 40320 0 _1266_
rlabel metal3 5992 38248 5992 38248 0 _1267_
rlabel metal2 6384 37464 6384 37464 0 _1268_
rlabel metal2 5936 38808 5936 38808 0 _1269_
rlabel metal2 6552 37632 6552 37632 0 _1270_
rlabel metal2 12040 43288 12040 43288 0 _1271_
rlabel metal2 12096 39816 12096 39816 0 _1272_
rlabel metal3 12936 41944 12936 41944 0 _1273_
rlabel metal2 16968 50120 16968 50120 0 _1274_
rlabel metal2 17192 51128 17192 51128 0 _1275_
rlabel metal2 23352 53144 23352 53144 0 _1276_
rlabel metal2 14728 49896 14728 49896 0 _1277_
rlabel metal3 15008 45080 15008 45080 0 _1278_
rlabel metal2 14392 45416 14392 45416 0 _1279_
rlabel metal2 14840 46984 14840 46984 0 _1280_
rlabel metal2 39928 49000 39928 49000 0 _1281_
rlabel metal2 39816 49672 39816 49672 0 _1282_
rlabel metal2 41496 49672 41496 49672 0 _1283_
rlabel metal2 40264 51156 40264 51156 0 _1284_
rlabel metal3 15512 49000 15512 49000 0 _1285_
rlabel metal2 13888 48776 13888 48776 0 _1286_
rlabel metal2 12600 42336 12600 42336 0 _1287_
rlabel metal2 13048 40488 13048 40488 0 _1288_
rlabel metal3 12096 11480 12096 11480 0 _1289_
rlabel metal2 12712 20832 12712 20832 0 _1290_
rlabel metal2 15960 25592 15960 25592 0 _1291_
rlabel metal3 13048 39032 13048 39032 0 _1292_
rlabel metal2 13384 37184 13384 37184 0 _1293_
rlabel metal3 12320 44072 12320 44072 0 _1294_
rlabel metal3 21504 21784 21504 21784 0 _1295_
rlabel metal2 21112 24024 21112 24024 0 _1296_
rlabel metal2 15064 46648 15064 46648 0 _1297_
rlabel metal3 19544 17080 19544 17080 0 _1298_
rlabel metal3 21448 20776 21448 20776 0 _1299_
rlabel metal2 25368 22176 25368 22176 0 _1300_
rlabel metal2 21112 22008 21112 22008 0 _1301_
rlabel metal2 25256 19264 25256 19264 0 _1302_
rlabel metal2 22288 20888 22288 20888 0 _1303_
rlabel metal2 22008 17248 22008 17248 0 _1304_
rlabel metal2 22232 19152 22232 19152 0 _1305_
rlabel metal3 21896 16072 21896 16072 0 _1306_
rlabel metal2 22120 15484 22120 15484 0 _1307_
rlabel metal2 26712 9408 26712 9408 0 _1308_
rlabel metal2 26824 9352 26824 9352 0 _1309_
rlabel metal2 23800 9856 23800 9856 0 _1310_
rlabel metal2 28840 12488 28840 12488 0 _1311_
rlabel metal2 26264 9128 26264 9128 0 _1312_
rlabel metal2 35112 9352 35112 9352 0 _1313_
rlabel metal2 28616 9352 28616 9352 0 _1314_
rlabel metal2 14952 50176 14952 50176 0 _1315_
rlabel metal3 52332 13832 52332 13832 0 _1316_
rlabel metal2 43512 10248 43512 10248 0 _1317_
rlabel metal2 38696 9128 38696 9128 0 _1318_
rlabel metal2 34832 6552 34832 6552 0 _1319_
rlabel metal2 25480 17136 25480 17136 0 _1320_
rlabel metal2 46536 13776 46536 13776 0 _1321_
rlabel metal2 39592 8736 39592 8736 0 _1322_
rlabel metal2 38360 8624 38360 8624 0 _1323_
rlabel metal3 42728 9576 42728 9576 0 _1324_
rlabel metal2 41384 7728 41384 7728 0 _1325_
rlabel metal2 43624 8960 43624 8960 0 _1326_
rlabel metal2 49784 15848 49784 15848 0 _1327_
rlabel metal2 45808 16072 45808 16072 0 _1328_
rlabel metal2 46984 13272 46984 13272 0 _1329_
rlabel metal2 53424 15960 53424 15960 0 _1330_
rlabel metal2 50792 13888 50792 13888 0 _1331_
rlabel metal2 50904 15792 50904 15792 0 _1332_
rlabel metal2 51464 17752 51464 17752 0 _1333_
rlabel metal2 55384 23016 55384 23016 0 _1334_
rlabel metal2 53480 18144 53480 18144 0 _1335_
rlabel metal2 55608 25480 55608 25480 0 _1336_
rlabel metal3 55384 21448 55384 21448 0 _1337_
rlabel metal3 56112 23016 56112 23016 0 _1338_
rlabel metal3 55664 24584 55664 24584 0 _1339_
rlabel metal2 54376 26432 54376 26432 0 _1340_
rlabel metal2 55160 26572 55160 26572 0 _1341_
rlabel metal3 56056 26152 56056 26152 0 _1342_
rlabel metal2 42728 31360 42728 31360 0 _1343_
rlabel metal3 54488 30072 54488 30072 0 _1344_
rlabel metal2 55552 28728 55552 28728 0 _1345_
rlabel metal2 53032 31416 53032 31416 0 _1346_
rlabel metal3 55160 30968 55160 30968 0 _1347_
rlabel metal2 54432 31864 54432 31864 0 _1348_
rlabel metal2 22120 53256 22120 53256 0 _1349_
rlabel metal2 25536 34216 25536 34216 0 _1350_
rlabel metal2 41832 31864 41832 31864 0 _1351_
rlabel metal2 21672 53144 21672 53144 0 _1352_
rlabel metal2 25928 32592 25928 32592 0 _1353_
rlabel metal2 31752 32984 31752 32984 0 _1354_
rlabel metal3 29176 32760 29176 32760 0 _1355_
rlabel metal3 24388 32648 24388 32648 0 _1356_
rlabel metal3 25032 32760 25032 32760 0 _1357_
rlabel metal2 17304 43456 17304 43456 0 _1358_
rlabel metal3 18144 33992 18144 33992 0 _1359_
rlabel metal3 16072 50568 16072 50568 0 _1360_
rlabel metal2 16296 34944 16296 34944 0 _1361_
rlabel metal3 12600 33096 12600 33096 0 _1362_
rlabel metal2 14280 34104 14280 34104 0 _1363_
rlabel metal2 14952 43932 14952 43932 0 _1364_
rlabel metal2 16352 44184 16352 44184 0 _1365_
rlabel metal2 15960 44576 15960 44576 0 _1366_
rlabel metal2 16520 47824 16520 47824 0 _1367_
rlabel metal2 14896 31640 14896 31640 0 _1368_
rlabel metal2 51464 24248 51464 24248 0 _1369_
rlabel metal3 53480 24136 53480 24136 0 _1370_
rlabel metal2 50456 23464 50456 23464 0 _1371_
rlabel metal3 52808 21672 52808 21672 0 _1372_
rlabel metal3 52360 22232 52360 22232 0 _1373_
rlabel metal2 51576 21280 51576 21280 0 _1374_
rlabel metal2 52696 22176 52696 22176 0 _1375_
rlabel metal2 52136 25144 52136 25144 0 _1376_
rlabel metal2 51912 25592 51912 25592 0 _1377_
rlabel metal2 51240 26264 51240 26264 0 _1378_
rlabel metal3 50372 25368 50372 25368 0 _1379_
rlabel metal2 51240 25592 51240 25592 0 _1380_
rlabel metal2 51520 26488 51520 26488 0 _1381_
rlabel metal2 53032 27216 53032 27216 0 _1382_
rlabel metal2 54152 27944 54152 27944 0 _1383_
rlabel metal2 53928 28448 53928 28448 0 _1384_
rlabel metal2 53592 27720 53592 27720 0 _1385_
rlabel metal2 52248 28728 52248 28728 0 _1386_
rlabel metal2 55440 29512 55440 29512 0 _1387_
rlabel metal2 55160 29456 55160 29456 0 _1388_
rlabel metal2 52024 29344 52024 29344 0 _1389_
rlabel metal2 52584 29232 52584 29232 0 _1390_
rlabel metal2 51576 31808 51576 31808 0 _1391_
rlabel metal2 53144 31192 53144 31192 0 _1392_
rlabel metal2 53592 30576 53592 30576 0 _1393_
rlabel metal2 36344 30352 36344 30352 0 _1394_
rlabel metal3 29176 19208 29176 19208 0 _1395_
rlabel metal2 29400 19544 29400 19544 0 _1396_
rlabel metal2 27720 23408 27720 23408 0 _1397_
rlabel metal2 28896 23240 28896 23240 0 _1398_
rlabel metal3 24584 25480 24584 25480 0 _1399_
rlabel metal2 27720 24696 27720 24696 0 _1400_
rlabel metal2 28728 23072 28728 23072 0 _1401_
rlabel metal3 27720 21672 27720 21672 0 _1402_
rlabel metal2 26712 20328 26712 20328 0 _1403_
rlabel metal2 28728 22064 28728 22064 0 _1404_
rlabel metal2 29512 19712 29512 19712 0 _1405_
rlabel metal2 30800 11256 30800 11256 0 _1406_
rlabel metal3 28448 12152 28448 12152 0 _1407_
rlabel metal2 28168 12656 28168 12656 0 _1408_
rlabel metal3 29344 17640 29344 17640 0 _1409_
rlabel metal3 26152 15960 26152 15960 0 _1410_
rlabel metal3 28448 15400 28448 15400 0 _1411_
rlabel metal2 29400 15176 29400 15176 0 _1412_
rlabel metal2 39480 14168 39480 14168 0 _1413_
rlabel metal3 30744 11256 30744 11256 0 _1414_
rlabel metal2 29064 12264 29064 12264 0 _1415_
rlabel metal2 27496 14056 27496 14056 0 _1416_
rlabel metal2 28056 13832 28056 13832 0 _1417_
rlabel metal2 25872 16296 25872 16296 0 _1418_
rlabel metal2 27608 13832 27608 13832 0 _1419_
rlabel metal3 28784 12936 28784 12936 0 _1420_
rlabel metal2 39592 14168 39592 14168 0 _1421_
rlabel metal2 47320 17304 47320 17304 0 _1422_
rlabel metal3 45920 16296 45920 16296 0 _1423_
rlabel metal3 4774 55160 4774 55160 0 clk
rlabel metal2 48776 52304 48776 52304 0 clknet_0_clk
rlabel metal2 1848 10584 1848 10584 0 clknet_4_0_0_clk
rlabel metal2 48888 29456 48888 29456 0 clknet_4_10_0_clk
rlabel metal3 47096 40376 47096 40376 0 clknet_4_11_0_clk
rlabel metal2 25816 40936 25816 40936 0 clknet_4_12_0_clk
rlabel metal2 25704 51688 25704 51688 0 clknet_4_13_0_clk
rlabel metal2 42392 41888 42392 41888 0 clknet_4_14_0_clk
rlabel metal2 44968 52528 44968 52528 0 clknet_4_15_0_clk
rlabel metal2 1848 29400 1848 29400 0 clknet_4_1_0_clk
rlabel via2 22904 17640 22904 17640 0 clknet_4_2_0_clk
rlabel metal3 16576 25256 16576 25256 0 clknet_4_3_0_clk
rlabel metal2 7672 39648 7672 39648 0 clknet_4_4_0_clk
rlabel metal2 8232 45080 8232 45080 0 clknet_4_5_0_clk
rlabel metal2 20776 44744 20776 44744 0 clknet_4_6_0_clk
rlabel metal2 21448 50512 21448 50512 0 clknet_4_7_0_clk
rlabel metal2 44968 20048 44968 20048 0 clknet_4_8_0_clk
rlabel metal2 51688 14560 51688 14560 0 clknet_4_9_0_clk
rlabel metal2 2072 41216 2072 41216 0 net1
rlabel metal2 2520 46760 2520 46760 0 net10
rlabel metal2 44240 38136 44240 38136 0 net100
rlabel metal2 41720 41384 41720 41384 0 net101
rlabel metal2 28616 45192 28616 45192 0 net102
rlabel metal2 33432 44520 33432 44520 0 net103
rlabel metal2 24024 56336 24024 56336 0 net104
rlabel metal2 30072 50232 30072 50232 0 net105
rlabel metal2 32144 44408 32144 44408 0 net106
rlabel metal2 18088 37352 18088 37352 0 net107
rlabel metal2 46424 56056 46424 56056 0 net108
rlabel metal2 30352 46536 30352 46536 0 net109
rlabel metal2 2128 42168 2128 42168 0 net11
rlabel metal2 24752 54488 24752 54488 0 net110
rlabel metal3 26040 48216 26040 48216 0 net111
rlabel metal2 27216 48104 27216 48104 0 net112
rlabel metal2 48776 40544 48776 40544 0 net113
rlabel metal2 40040 34104 40040 34104 0 net114
rlabel metal3 39928 50792 39928 50792 0 net115
rlabel metal2 3808 44072 3808 44072 0 net116
rlabel metal2 7112 39648 7112 39648 0 net117
rlabel metal2 8120 43064 8120 43064 0 net118
rlabel metal3 2856 47208 2856 47208 0 net12
rlabel metal2 2744 36456 2744 36456 0 net13
rlabel metal2 5264 38808 5264 38808 0 net14
rlabel metal2 2072 40320 2072 40320 0 net15
rlabel metal3 3248 43848 3248 43848 0 net16
rlabel metal1 2688 46424 2688 46424 0 net17
rlabel metal2 4872 43120 4872 43120 0 net18
rlabel metal2 33152 21448 33152 21448 0 net19
rlabel metal2 6888 43120 6888 43120 0 net2
rlabel metal3 37856 14504 37856 14504 0 net20
rlabel metal2 36232 13608 36232 13608 0 net21
rlabel metal2 37128 17640 37128 17640 0 net22
rlabel metal2 46424 17976 46424 17976 0 net23
rlabel metal2 40488 18256 40488 18256 0 net24
rlabel metal2 40040 18704 40040 18704 0 net25
rlabel metal2 41496 22904 41496 22904 0 net26
rlabel metal2 41944 22736 41944 22736 0 net27
rlabel metal2 43176 24584 43176 24584 0 net28
rlabel metal3 42952 23352 42952 23352 0 net29
rlabel metal2 5656 38528 5656 38528 0 net3
rlabel metal2 33880 21448 33880 21448 0 net30
rlabel metal2 41160 25984 41160 25984 0 net31
rlabel metal2 40376 26040 40376 26040 0 net32
rlabel metal2 41888 26488 41888 26488 0 net33
rlabel metal2 41944 29120 41944 29120 0 net34
rlabel metal2 37240 26656 37240 26656 0 net35
rlabel metal2 57848 26656 57848 26656 0 net36
rlabel metal2 35336 27216 35336 27216 0 net37
rlabel metal2 24976 25256 24976 25256 0 net38
rlabel metal2 22456 27384 22456 27384 0 net39
rlabel metal2 5992 39536 5992 39536 0 net4
rlabel metal2 2072 27104 2072 27104 0 net40
rlabel metal3 34888 21840 34888 21840 0 net41
rlabel metal2 19152 25592 19152 25592 0 net42
rlabel metal2 18760 24976 18760 24976 0 net43
rlabel metal2 49000 18172 49000 18172 0 net44
rlabel metal2 32648 10024 32648 10024 0 net45
rlabel metal2 33320 7224 33320 7224 0 net46
rlabel metal3 32704 15400 32704 15400 0 net47
rlabel metal2 31192 14224 31192 14224 0 net48
rlabel metal2 35448 13944 35448 13944 0 net49
rlabel metal3 3360 38920 3360 38920 0 net5
rlabel metal2 35056 15288 35056 15288 0 net50
rlabel metal2 8008 30296 8008 30296 0 net51
rlabel metal2 2408 22008 2408 22008 0 net52
rlabel metal2 2968 20720 2968 20720 0 net53
rlabel metal2 6104 19152 6104 19152 0 net54
rlabel metal2 2072 18200 2072 18200 0 net55
rlabel metal2 2744 16632 2744 16632 0 net56
rlabel metal3 2072 15288 2072 15288 0 net57
rlabel metal2 7000 12824 7000 12824 0 net58
rlabel metal2 2072 12432 2072 12432 0 net59
rlabel metal3 4424 45192 4424 45192 0 net6
rlabel metal2 2072 11200 2072 11200 0 net60
rlabel metal2 2744 13272 2744 13272 0 net61
rlabel metal3 2072 31416 2072 31416 0 net62
rlabel metal2 2072 14560 2072 14560 0 net63
rlabel metal2 2744 14504 2744 14504 0 net64
rlabel metal2 14056 15204 14056 15204 0 net65
rlabel metal2 2744 11088 2744 11088 0 net66
rlabel metal2 2072 16800 2072 16800 0 net67
rlabel metal2 15288 15848 15288 15848 0 net68
rlabel metal2 17360 13608 17360 13608 0 net69
rlabel metal3 3752 44520 3752 44520 0 net7
rlabel metal2 18088 3584 18088 3584 0 net70
rlabel metal2 18424 3696 18424 3696 0 net71
rlabel metal2 15512 18760 15512 18760 0 net72
rlabel metal2 2744 30912 2744 30912 0 net73
rlabel metal2 2968 21896 2968 21896 0 net74
rlabel metal2 2744 27048 2744 27048 0 net75
rlabel metal2 8456 31024 8456 31024 0 net76
rlabel metal2 7000 29512 7000 29512 0 net77
rlabel metal2 2072 27832 2072 27832 0 net78
rlabel metal2 2296 25648 2296 25648 0 net79
rlabel metal3 4032 48328 4032 48328 0 net8
rlabel metal2 2072 25704 2072 25704 0 net80
rlabel metal2 8176 20776 8176 20776 0 net81
rlabel metal2 8512 20776 8512 20776 0 net82
rlabel metal2 2744 41440 2744 41440 0 net83
rlabel metal2 20664 51464 20664 51464 0 net84
rlabel metal3 50008 56056 50008 56056 0 net85
rlabel metal3 39928 51128 39928 51128 0 net86
rlabel metal2 45528 35728 45528 35728 0 net87
rlabel metal2 44296 39984 44296 39984 0 net88
rlabel metal2 49672 43792 49672 43792 0 net89
rlabel metal3 3024 49896 3024 49896 0 net9
rlabel metal2 48104 40208 48104 40208 0 net90
rlabel metal2 51688 38864 51688 38864 0 net91
rlabel metal2 51296 41272 51296 41272 0 net92
rlabel metal2 51688 37856 51688 37856 0 net93
rlabel metal3 53088 40264 53088 40264 0 net94
rlabel metal2 33544 42336 33544 42336 0 net95
rlabel metal2 56616 36904 56616 36904 0 net96
rlabel metal2 53256 40432 53256 40432 0 net97
rlabel metal2 55944 39648 55944 39648 0 net98
rlabel metal2 55664 40264 55664 40264 0 net99
rlabel metal2 20216 57946 20216 57946 0 pcpi_div_rd[0]
rlabel metal2 38360 57610 38360 57610 0 pcpi_div_rd[10]
rlabel metal2 42168 55328 42168 55328 0 pcpi_div_rd[11]
rlabel metal2 57960 34664 57960 34664 0 pcpi_div_rd[12]
rlabel metal2 55272 40824 55272 40824 0 pcpi_div_rd[13]
rlabel metal2 54936 45192 54936 45192 0 pcpi_div_rd[14]
rlabel metal2 55384 42504 55384 42504 0 pcpi_div_rd[15]
rlabel metal3 58338 38360 58338 38360 0 pcpi_div_rd[16]
rlabel metal2 55048 43736 55048 43736 0 pcpi_div_rd[17]
rlabel metal2 55384 35224 55384 35224 0 pcpi_div_rd[18]
rlabel metal2 57736 44184 57736 44184 0 pcpi_div_rd[19]
rlabel metal2 33656 57218 33656 57218 0 pcpi_div_rd[1]
rlabel metal2 55048 36344 55048 36344 0 pcpi_div_rd[20]
rlabel metal3 58058 41048 58058 41048 0 pcpi_div_rd[21]
rlabel metal3 58618 37688 58618 37688 0 pcpi_div_rd[22]
rlabel metal2 57848 42392 57848 42392 0 pcpi_div_rd[23]
rlabel metal2 55384 37800 55384 37800 0 pcpi_div_rd[24]
rlabel metal2 57960 45640 57960 45640 0 pcpi_div_rd[25]
rlabel metal2 28952 57554 28952 57554 0 pcpi_div_rd[26]
rlabel metal2 32312 56378 32312 56378 0 pcpi_div_rd[27]
rlabel metal2 23016 55552 23016 55552 0 pcpi_div_rd[28]
rlabel metal2 30296 55818 30296 55818 0 pcpi_div_rd[29]
rlabel metal2 31640 57778 31640 57778 0 pcpi_div_rd[2]
rlabel metal3 1358 35000 1358 35000 0 pcpi_div_rd[30]
rlabel metal2 43848 55664 43848 55664 0 pcpi_div_rd[31]
rlabel metal2 30968 57610 30968 57610 0 pcpi_div_rd[3]
rlabel metal2 23632 57400 23632 57400 0 pcpi_div_rd[4]
rlabel metal3 26320 52360 26320 52360 0 pcpi_div_rd[5]
rlabel metal2 26824 55608 26824 55608 0 pcpi_div_rd[6]
rlabel metal2 55048 40152 55048 40152 0 pcpi_div_rd[7]
rlabel metal2 58016 33544 58016 33544 0 pcpi_div_rd[8]
rlabel metal2 42504 53088 42504 53088 0 pcpi_div_rd[9]
rlabel metal3 1358 49784 1358 49784 0 pcpi_div_ready
rlabel metal2 1848 40768 1848 40768 0 pcpi_div_valid
rlabel metal3 1358 39704 1358 39704 0 pcpi_div_wait
rlabel metal3 1358 43736 1358 43736 0 pcpi_div_wr
rlabel metal2 1736 43288 1736 43288 0 pcpi_insn[0]
rlabel metal2 1736 37128 1736 37128 0 pcpi_insn[12]
rlabel metal2 1736 37800 1736 37800 0 pcpi_insn[13]
rlabel metal2 1736 38584 1736 38584 0 pcpi_insn[14]
rlabel metal2 1736 44744 1736 44744 0 pcpi_insn[1]
rlabel metal2 1848 45472 1848 45472 0 pcpi_insn[25]
rlabel metal2 1736 47992 1736 47992 0 pcpi_insn[26]
rlabel metal2 1736 49448 1736 49448 0 pcpi_insn[27]
rlabel metal2 1736 48664 1736 48664 0 pcpi_insn[28]
rlabel metal2 1736 41832 1736 41832 0 pcpi_insn[29]
rlabel metal2 1736 47208 1736 47208 0 pcpi_insn[2]
rlabel metal3 1582 36344 1582 36344 0 pcpi_insn[30]
rlabel metal2 1736 36008 1736 36008 0 pcpi_insn[31]
rlabel metal2 1736 39704 1736 39704 0 pcpi_insn[3]
rlabel metal3 1582 45752 1582 45752 0 pcpi_insn[4]
rlabel metal2 1736 46536 1736 46536 0 pcpi_insn[5]
rlabel metal2 1736 42504 1736 42504 0 pcpi_insn[6]
rlabel metal2 29736 2296 29736 2296 0 pcpi_rs1[0]
rlabel metal2 38416 3304 38416 3304 0 pcpi_rs1[10]
rlabel metal3 36960 3528 36960 3528 0 pcpi_rs1[11]
rlabel metal1 37632 2408 37632 2408 0 pcpi_rs1[12]
rlabel metal2 39032 3864 39032 3864 0 pcpi_rs1[13]
rlabel metal2 39704 2856 39704 2856 0 pcpi_rs1[14]
rlabel metal2 39816 2744 39816 2744 0 pcpi_rs1[15]
rlabel metal2 57512 23352 57512 23352 0 pcpi_rs1[16]
rlabel metal2 58184 22008 58184 22008 0 pcpi_rs1[17]
rlabel metal3 58394 24920 58394 24920 0 pcpi_rs1[18]
rlabel metal2 58184 23744 58184 23744 0 pcpi_rs1[19]
rlabel metal2 33544 3864 33544 3864 0 pcpi_rs1[1]
rlabel metal2 58184 25032 58184 25032 0 pcpi_rs1[20]
rlabel metal3 58394 26264 58394 26264 0 pcpi_rs1[21]
rlabel metal3 58730 29624 58730 29624 0 pcpi_rs1[22]
rlabel metal2 57512 29176 57512 29176 0 pcpi_rs1[23]
rlabel metal2 58184 27720 58184 27720 0 pcpi_rs1[24]
rlabel metal2 58072 26096 58072 26096 0 pcpi_rs1[25]
rlabel metal2 58184 28448 58184 28448 0 pcpi_rs1[26]
rlabel metal2 24416 3416 24416 3416 0 pcpi_rs1[27]
rlabel metal2 2408 29176 2408 29176 0 pcpi_rs1[28]
rlabel metal2 1736 27216 1736 27216 0 pcpi_rs1[29]
rlabel metal2 35000 2968 35000 2968 0 pcpi_rs1[2]
rlabel metal2 2576 27832 2576 27832 0 pcpi_rs1[30]
rlabel metal2 2408 24472 2408 24472 0 pcpi_rs1[31]
rlabel metal2 34048 2520 34048 2520 0 pcpi_rs1[3]
rlabel metal2 31640 1246 31640 1246 0 pcpi_rs1[4]
rlabel metal2 32592 2520 32592 2520 0 pcpi_rs1[5]
rlabel metal2 30296 2058 30296 2058 0 pcpi_rs1[6]
rlabel metal2 31080 3528 31080 3528 0 pcpi_rs1[7]
rlabel metal2 35112 2856 35112 2856 0 pcpi_rs1[8]
rlabel metal1 36288 2520 36288 2520 0 pcpi_rs1[9]
rlabel metal2 3080 30632 3080 30632 0 pcpi_rs2[0]
rlabel metal2 1736 22792 1736 22792 0 pcpi_rs2[10]
rlabel metal2 2744 20104 2744 20104 0 pcpi_rs2[11]
rlabel metal2 2408 18984 2408 18984 0 pcpi_rs2[12]
rlabel metal2 1736 18088 1736 18088 0 pcpi_rs2[13]
rlabel metal3 1582 16856 1582 16856 0 pcpi_rs2[14]
rlabel metal2 1736 15792 1736 15792 0 pcpi_rs2[15]
rlabel metal2 3080 10360 3080 10360 0 pcpi_rs2[16]
rlabel metal3 1246 12152 1246 12152 0 pcpi_rs2[17]
rlabel metal2 1736 11088 1736 11088 0 pcpi_rs2[18]
rlabel metal3 1582 12824 1582 12824 0 pcpi_rs2[19]
rlabel metal2 1792 33992 1792 33992 0 pcpi_rs2[1]
rlabel metal2 1736 14784 1736 14784 0 pcpi_rs2[20]
rlabel metal3 854 14168 854 14168 0 pcpi_rs2[21]
rlabel metal2 1736 13160 1736 13160 0 pcpi_rs2[22]
rlabel metal2 2408 10752 2408 10752 0 pcpi_rs2[23]
rlabel metal2 3024 14616 3024 14616 0 pcpi_rs2[24]
rlabel metal2 2408 15456 2408 15456 0 pcpi_rs2[25]
rlabel metal2 16688 3416 16688 3416 0 pcpi_rs2[26]
rlabel metal2 17640 3304 17640 3304 0 pcpi_rs2[27]
rlabel metal2 18648 3864 18648 3864 0 pcpi_rs2[28]
rlabel metal3 1246 19544 1246 19544 0 pcpi_rs2[29]
rlabel metal3 1582 30968 1582 30968 0 pcpi_rs2[2]
rlabel metal3 3038 21560 3038 21560 0 pcpi_rs2[30]
rlabel metal2 2520 26992 2520 26992 0 pcpi_rs2[31]
rlabel metal2 1848 31080 1848 31080 0 pcpi_rs2[3]
rlabel metal3 2464 29400 2464 29400 0 pcpi_rs2[4]
rlabel metal2 1736 28168 1736 28168 0 pcpi_rs2[5]
rlabel metal2 1736 25536 1736 25536 0 pcpi_rs2[6]
rlabel metal2 1736 24360 1736 24360 0 pcpi_rs2[7]
rlabel metal2 1736 22008 1736 22008 0 pcpi_rs2[8]
rlabel metal2 1736 20384 1736 20384 0 pcpi_rs2[9]
rlabel metal2 26712 24808 26712 24808 0 picorv32_pcpi_div_inst_0.dividend\[0\]
rlabel metal2 40656 23688 40656 23688 0 picorv32_pcpi_div_inst_0.dividend\[10\]
rlabel metal2 43400 11424 43400 11424 0 picorv32_pcpi_div_inst_0.dividend\[11\]
rlabel metal3 42560 22344 42560 22344 0 picorv32_pcpi_div_inst_0.dividend\[12\]
rlabel metal2 42504 16184 42504 16184 0 picorv32_pcpi_div_inst_0.dividend\[13\]
rlabel metal2 47656 16576 47656 16576 0 picorv32_pcpi_div_inst_0.dividend\[14\]
rlabel metal2 48216 19152 48216 19152 0 picorv32_pcpi_div_inst_0.dividend\[15\]
rlabel metal2 48216 21616 48216 21616 0 picorv32_pcpi_div_inst_0.dividend\[16\]
rlabel metal3 50008 21560 50008 21560 0 picorv32_pcpi_div_inst_0.dividend\[17\]
rlabel metal2 48888 26208 48888 26208 0 picorv32_pcpi_div_inst_0.dividend\[18\]
rlabel metal2 49448 24976 49448 24976 0 picorv32_pcpi_div_inst_0.dividend\[19\]
rlabel metal2 25704 23968 25704 23968 0 picorv32_pcpi_div_inst_0.dividend\[1\]
rlabel metal2 52248 35952 52248 35952 0 picorv32_pcpi_div_inst_0.dividend\[20\]
rlabel metal2 47768 33488 47768 33488 0 picorv32_pcpi_div_inst_0.dividend\[21\]
rlabel metal2 50344 32144 50344 32144 0 picorv32_pcpi_div_inst_0.dividend\[22\]
rlabel metal2 47880 30632 47880 30632 0 picorv32_pcpi_div_inst_0.dividend\[23\]
rlabel metal2 38920 32536 38920 32536 0 picorv32_pcpi_div_inst_0.dividend\[24\]
rlabel metal2 39704 30632 39704 30632 0 picorv32_pcpi_div_inst_0.dividend\[25\]
rlabel metal2 30408 30464 30408 30464 0 picorv32_pcpi_div_inst_0.dividend\[26\]
rlabel metal2 30968 29456 30968 29456 0 picorv32_pcpi_div_inst_0.dividend\[27\]
rlabel metal2 22344 33656 22344 33656 0 picorv32_pcpi_div_inst_0.dividend\[28\]
rlabel metal3 19488 30968 19488 30968 0 picorv32_pcpi_div_inst_0.dividend\[29\]
rlabel metal2 26264 22680 26264 22680 0 picorv32_pcpi_div_inst_0.dividend\[2\]
rlabel metal3 15400 30856 15400 30856 0 picorv32_pcpi_div_inst_0.dividend\[30\]
rlabel metal2 18200 26768 18200 26768 0 picorv32_pcpi_div_inst_0.dividend\[31\]
rlabel metal2 26656 20888 26656 20888 0 picorv32_pcpi_div_inst_0.dividend\[3\]
rlabel metal2 24360 16520 24360 16520 0 picorv32_pcpi_div_inst_0.dividend\[4\]
rlabel metal3 25872 14840 25872 14840 0 picorv32_pcpi_div_inst_0.dividend\[5\]
rlabel metal2 25368 11424 25368 11424 0 picorv32_pcpi_div_inst_0.dividend\[6\]
rlabel metal2 30072 10640 30072 10640 0 picorv32_pcpi_div_inst_0.dividend\[7\]
rlabel metal2 34552 9464 34552 9464 0 picorv32_pcpi_div_inst_0.dividend\[8\]
rlabel metal2 37296 16744 37296 16744 0 picorv32_pcpi_div_inst_0.dividend\[9\]
rlabel metal2 22232 24248 22232 24248 0 picorv32_pcpi_div_inst_0.divisor\[0\]
rlabel metal3 40544 9016 40544 9016 0 picorv32_pcpi_div_inst_0.divisor\[10\]
rlabel metal2 45192 9240 45192 9240 0 picorv32_pcpi_div_inst_0.divisor\[11\]
rlabel metal2 42952 16128 42952 16128 0 picorv32_pcpi_div_inst_0.divisor\[12\]
rlabel metal2 48888 14560 48888 14560 0 picorv32_pcpi_div_inst_0.divisor\[13\]
rlabel metal3 48384 16072 48384 16072 0 picorv32_pcpi_div_inst_0.divisor\[14\]
rlabel metal2 49448 16800 49448 16800 0 picorv32_pcpi_div_inst_0.divisor\[15\]
rlabel metal2 52360 17976 52360 17976 0 picorv32_pcpi_div_inst_0.divisor\[16\]
rlabel metal2 54040 21224 54040 21224 0 picorv32_pcpi_div_inst_0.divisor\[17\]
rlabel metal2 53592 24640 53592 24640 0 picorv32_pcpi_div_inst_0.divisor\[18\]
rlabel metal2 50232 24752 50232 24752 0 picorv32_pcpi_div_inst_0.divisor\[19\]
rlabel metal2 22008 23128 22008 23128 0 picorv32_pcpi_div_inst_0.divisor\[1\]
rlabel metal2 55496 25928 55496 25928 0 picorv32_pcpi_div_inst_0.divisor\[20\]
rlabel metal2 55720 27496 55720 27496 0 picorv32_pcpi_div_inst_0.divisor\[21\]
rlabel metal2 54488 30240 54488 30240 0 picorv32_pcpi_div_inst_0.divisor\[22\]
rlabel metal2 50120 30856 50120 30856 0 picorv32_pcpi_div_inst_0.divisor\[23\]
rlabel metal2 44632 32312 44632 32312 0 picorv32_pcpi_div_inst_0.divisor\[24\]
rlabel metal2 40152 30632 40152 30632 0 picorv32_pcpi_div_inst_0.divisor\[25\]
rlabel metal2 30744 31080 30744 31080 0 picorv32_pcpi_div_inst_0.divisor\[26\]
rlabel metal2 25704 32816 25704 32816 0 picorv32_pcpi_div_inst_0.divisor\[27\]
rlabel metal2 21112 32984 21112 32984 0 picorv32_pcpi_div_inst_0.divisor\[28\]
rlabel metal2 19880 31836 19880 31836 0 picorv32_pcpi_div_inst_0.divisor\[29\]
rlabel metal2 26040 21504 26040 21504 0 picorv32_pcpi_div_inst_0.divisor\[2\]
rlabel metal2 15512 34048 15512 34048 0 picorv32_pcpi_div_inst_0.divisor\[30\]
rlabel metal2 13384 32256 13384 32256 0 picorv32_pcpi_div_inst_0.divisor\[31\]
rlabel metal3 10976 33432 10976 33432 0 picorv32_pcpi_div_inst_0.divisor\[32\]
rlabel metal2 7000 32592 7000 32592 0 picorv32_pcpi_div_inst_0.divisor\[33\]
rlabel metal2 5320 32256 5320 32256 0 picorv32_pcpi_div_inst_0.divisor\[34\]
rlabel metal2 4648 32536 4648 32536 0 picorv32_pcpi_div_inst_0.divisor\[35\]
rlabel metal2 5096 25928 5096 25928 0 picorv32_pcpi_div_inst_0.divisor\[36\]
rlabel metal2 5264 26040 5264 26040 0 picorv32_pcpi_div_inst_0.divisor\[37\]
rlabel metal3 5040 26152 5040 26152 0 picorv32_pcpi_div_inst_0.divisor\[38\]
rlabel metal3 11256 24024 11256 24024 0 picorv32_pcpi_div_inst_0.divisor\[39\]
rlabel metal2 25704 19600 25704 19600 0 picorv32_pcpi_div_inst_0.divisor\[3\]
rlabel metal2 9240 23800 9240 23800 0 picorv32_pcpi_div_inst_0.divisor\[40\]
rlabel metal2 5320 23072 5320 23072 0 picorv32_pcpi_div_inst_0.divisor\[41\]
rlabel metal2 4872 23240 4872 23240 0 picorv32_pcpi_div_inst_0.divisor\[42\]
rlabel metal2 4648 20888 4648 20888 0 picorv32_pcpi_div_inst_0.divisor\[43\]
rlabel metal2 4648 17696 4648 17696 0 picorv32_pcpi_div_inst_0.divisor\[44\]
rlabel metal2 4032 16856 4032 16856 0 picorv32_pcpi_div_inst_0.divisor\[45\]
rlabel metal2 4200 16016 4200 16016 0 picorv32_pcpi_div_inst_0.divisor\[46\]
rlabel metal2 5320 14280 5320 14280 0 picorv32_pcpi_div_inst_0.divisor\[47\]
rlabel metal2 5992 10976 5992 10976 0 picorv32_pcpi_div_inst_0.divisor\[48\]
rlabel metal3 8064 10584 8064 10584 0 picorv32_pcpi_div_inst_0.divisor\[49\]
rlabel metal3 23352 16072 23352 16072 0 picorv32_pcpi_div_inst_0.divisor\[4\]
rlabel metal2 9520 11368 9520 11368 0 picorv32_pcpi_div_inst_0.divisor\[50\]
rlabel metal2 11984 9800 11984 9800 0 picorv32_pcpi_div_inst_0.divisor\[51\]
rlabel metal2 13832 10808 13832 10808 0 picorv32_pcpi_div_inst_0.divisor\[52\]
rlabel metal2 12712 9520 12712 9520 0 picorv32_pcpi_div_inst_0.divisor\[53\]
rlabel metal2 14504 6888 14504 6888 0 picorv32_pcpi_div_inst_0.divisor\[54\]
rlabel metal2 15400 11200 15400 11200 0 picorv32_pcpi_div_inst_0.divisor\[55\]
rlabel metal2 16072 9688 16072 9688 0 picorv32_pcpi_div_inst_0.divisor\[56\]
rlabel metal2 16632 10976 16632 10976 0 picorv32_pcpi_div_inst_0.divisor\[57\]
rlabel metal2 20776 10920 20776 10920 0 picorv32_pcpi_div_inst_0.divisor\[58\]
rlabel metal2 19320 11760 19320 11760 0 picorv32_pcpi_div_inst_0.divisor\[59\]
rlabel metal3 23856 15288 23856 15288 0 picorv32_pcpi_div_inst_0.divisor\[5\]
rlabel metal2 18872 16912 18872 16912 0 picorv32_pcpi_div_inst_0.divisor\[60\]
rlabel metal2 18200 21112 18200 21112 0 picorv32_pcpi_div_inst_0.divisor\[61\]
rlabel metal2 18424 21000 18424 21000 0 picorv32_pcpi_div_inst_0.divisor\[62\]
rlabel metal2 27608 9744 27608 9744 0 picorv32_pcpi_div_inst_0.divisor\[6\]
rlabel metal2 30296 8176 30296 8176 0 picorv32_pcpi_div_inst_0.divisor\[7\]
rlabel metal2 36008 8624 36008 8624 0 picorv32_pcpi_div_inst_0.divisor\[8\]
rlabel metal2 38920 8624 38920 8624 0 picorv32_pcpi_div_inst_0.divisor\[9\]
rlabel metal2 11592 28112 11592 28112 0 picorv32_pcpi_div_inst_0.instr_div
rlabel metal2 11592 37968 11592 37968 0 picorv32_pcpi_div_inst_0.instr_divu
rlabel metal2 8008 35672 8008 35672 0 picorv32_pcpi_div_inst_0.instr_rem
rlabel metal2 7448 40376 7448 40376 0 picorv32_pcpi_div_inst_0.instr_remu
rlabel metal2 18760 38304 18760 38304 0 picorv32_pcpi_div_inst_0.outsign
rlabel metal2 12712 40264 12712 40264 0 picorv32_pcpi_div_inst_0.pcpi_wait_q
rlabel metal2 20552 45920 20552 45920 0 picorv32_pcpi_div_inst_0.quotient\[0\]
rlabel metal2 33544 53536 33544 53536 0 picorv32_pcpi_div_inst_0.quotient\[10\]
rlabel metal3 34496 50456 34496 50456 0 picorv32_pcpi_div_inst_0.quotient\[11\]
rlabel metal2 39872 52920 39872 52920 0 picorv32_pcpi_div_inst_0.quotient\[12\]
rlabel metal2 40096 51352 40096 51352 0 picorv32_pcpi_div_inst_0.quotient\[13\]
rlabel metal2 44296 47880 44296 47880 0 picorv32_pcpi_div_inst_0.quotient\[14\]
rlabel metal2 44520 45752 44520 45752 0 picorv32_pcpi_div_inst_0.quotient\[15\]
rlabel metal2 47544 45528 47544 45528 0 picorv32_pcpi_div_inst_0.quotient\[16\]
rlabel metal3 47600 46088 47600 46088 0 picorv32_pcpi_div_inst_0.quotient\[17\]
rlabel metal2 47992 51688 47992 51688 0 picorv32_pcpi_div_inst_0.quotient\[18\]
rlabel metal2 48720 45864 48720 45864 0 picorv32_pcpi_div_inst_0.quotient\[19\]
rlabel metal2 20328 47488 20328 47488 0 picorv32_pcpi_div_inst_0.quotient\[1\]
rlabel metal2 55608 51072 55608 51072 0 picorv32_pcpi_div_inst_0.quotient\[20\]
rlabel metal2 53312 51352 53312 51352 0 picorv32_pcpi_div_inst_0.quotient\[21\]
rlabel metal2 52136 45864 52136 45864 0 picorv32_pcpi_div_inst_0.quotient\[22\]
rlabel metal2 50568 47320 50568 47320 0 picorv32_pcpi_div_inst_0.quotient\[23\]
rlabel metal2 39032 45472 39032 45472 0 picorv32_pcpi_div_inst_0.quotient\[24\]
rlabel metal2 39928 47600 39928 47600 0 picorv32_pcpi_div_inst_0.quotient\[25\]
rlabel metal2 26040 45528 26040 45528 0 picorv32_pcpi_div_inst_0.quotient\[26\]
rlabel metal2 25816 48720 25816 48720 0 picorv32_pcpi_div_inst_0.quotient\[27\]
rlabel metal2 17864 43400 17864 43400 0 picorv32_pcpi_div_inst_0.quotient\[28\]
rlabel metal2 13496 43288 13496 43288 0 picorv32_pcpi_div_inst_0.quotient\[29\]
rlabel metal2 19992 45752 19992 45752 0 picorv32_pcpi_div_inst_0.quotient\[2\]
rlabel via2 16408 40376 16408 40376 0 picorv32_pcpi_div_inst_0.quotient\[30\]
rlabel metal2 16856 39928 16856 39928 0 picorv32_pcpi_div_inst_0.quotient\[31\]
rlabel metal2 20552 50904 20552 50904 0 picorv32_pcpi_div_inst_0.quotient\[3\]
rlabel metal2 22456 48048 22456 48048 0 picorv32_pcpi_div_inst_0.quotient\[4\]
rlabel metal2 24248 50540 24248 50540 0 picorv32_pcpi_div_inst_0.quotient\[5\]
rlabel metal2 23576 52472 23576 52472 0 picorv32_pcpi_div_inst_0.quotient\[6\]
rlabel metal2 33992 46536 33992 46536 0 picorv32_pcpi_div_inst_0.quotient\[7\]
rlabel metal3 31864 49784 31864 49784 0 picorv32_pcpi_div_inst_0.quotient\[8\]
rlabel metal2 32536 50904 32536 50904 0 picorv32_pcpi_div_inst_0.quotient\[9\]
rlabel metal2 16072 46704 16072 46704 0 picorv32_pcpi_div_inst_0.quotient_msk\[0\]
rlabel via2 30520 53704 30520 53704 0 picorv32_pcpi_div_inst_0.quotient_msk\[10\]
rlabel metal2 38808 53256 38808 53256 0 picorv32_pcpi_div_inst_0.quotient_msk\[11\]
rlabel metal2 39592 52528 39592 52528 0 picorv32_pcpi_div_inst_0.quotient_msk\[12\]
rlabel metal2 39816 51800 39816 51800 0 picorv32_pcpi_div_inst_0.quotient_msk\[13\]
rlabel metal2 41160 53256 41160 53256 0 picorv32_pcpi_div_inst_0.quotient_msk\[14\]
rlabel metal2 44072 53256 44072 53256 0 picorv32_pcpi_div_inst_0.quotient_msk\[15\]
rlabel metal2 46144 54712 46144 54712 0 picorv32_pcpi_div_inst_0.quotient_msk\[16\]
rlabel metal2 46424 52472 46424 52472 0 picorv32_pcpi_div_inst_0.quotient_msk\[17\]
rlabel metal2 46984 50904 46984 50904 0 picorv32_pcpi_div_inst_0.quotient_msk\[18\]
rlabel metal2 49672 54544 49672 54544 0 picorv32_pcpi_div_inst_0.quotient_msk\[19\]
rlabel metal2 15064 49616 15064 49616 0 picorv32_pcpi_div_inst_0.quotient_msk\[1\]
rlabel metal2 52640 51352 52640 51352 0 picorv32_pcpi_div_inst_0.quotient_msk\[20\]
rlabel metal2 51184 52024 51184 52024 0 picorv32_pcpi_div_inst_0.quotient_msk\[21\]
rlabel metal2 50232 51184 50232 51184 0 picorv32_pcpi_div_inst_0.quotient_msk\[22\]
rlabel metal2 49336 51352 49336 51352 0 picorv32_pcpi_div_inst_0.quotient_msk\[23\]
rlabel metal2 36624 49784 36624 49784 0 picorv32_pcpi_div_inst_0.quotient_msk\[24\]
rlabel metal2 26768 51240 26768 51240 0 picorv32_pcpi_div_inst_0.quotient_msk\[25\]
rlabel metal2 26824 49336 26824 49336 0 picorv32_pcpi_div_inst_0.quotient_msk\[26\]
rlabel metal2 12936 47936 12936 47936 0 picorv32_pcpi_div_inst_0.quotient_msk\[27\]
rlabel metal2 13720 45696 13720 45696 0 picorv32_pcpi_div_inst_0.quotient_msk\[28\]
rlabel metal3 12880 45752 12880 45752 0 picorv32_pcpi_div_inst_0.quotient_msk\[29\]
rlabel metal2 16072 51912 16072 51912 0 picorv32_pcpi_div_inst_0.quotient_msk\[2\]
rlabel metal2 14336 45976 14336 45976 0 picorv32_pcpi_div_inst_0.quotient_msk\[30\]
rlabel metal2 15400 43064 15400 43064 0 picorv32_pcpi_div_inst_0.quotient_msk\[31\]
rlabel metal3 17864 52080 17864 52080 0 picorv32_pcpi_div_inst_0.quotient_msk\[3\]
rlabel metal2 17976 51912 17976 51912 0 picorv32_pcpi_div_inst_0.quotient_msk\[4\]
rlabel metal2 21784 54152 21784 54152 0 picorv32_pcpi_div_inst_0.quotient_msk\[5\]
rlabel metal2 22008 53256 22008 53256 0 picorv32_pcpi_div_inst_0.quotient_msk\[6\]
rlabel metal2 24248 52752 24248 52752 0 picorv32_pcpi_div_inst_0.quotient_msk\[7\]
rlabel metal2 26600 53256 26600 53256 0 picorv32_pcpi_div_inst_0.quotient_msk\[8\]
rlabel metal2 26656 54488 26656 54488 0 picorv32_pcpi_div_inst_0.quotient_msk\[9\]
rlabel metal2 14952 44912 14952 44912 0 picorv32_pcpi_div_inst_0.running
rlabel metal3 1582 41048 1582 41048 0 resetn
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>

magic
tech gf180mcuD
magscale 1 5
timestamp 1702206232
<< metal1 >>
rect 672 23141 24304 23158
rect 672 23115 2239 23141
rect 2265 23115 2291 23141
rect 2317 23115 2343 23141
rect 2369 23115 17599 23141
rect 17625 23115 17651 23141
rect 17677 23115 17703 23141
rect 17729 23115 24304 23141
rect 672 23098 24304 23115
rect 672 22749 24304 22766
rect 672 22723 9919 22749
rect 9945 22723 9971 22749
rect 9997 22723 10023 22749
rect 10049 22723 24304 22749
rect 672 22706 24304 22723
rect 672 22357 24304 22374
rect 672 22331 2239 22357
rect 2265 22331 2291 22357
rect 2317 22331 2343 22357
rect 2369 22331 17599 22357
rect 17625 22331 17651 22357
rect 17677 22331 17703 22357
rect 17729 22331 24304 22357
rect 672 22314 24304 22331
rect 672 21965 24304 21982
rect 672 21939 9919 21965
rect 9945 21939 9971 21965
rect 9997 21939 10023 21965
rect 10049 21939 24304 21965
rect 672 21922 24304 21939
rect 672 21573 24304 21590
rect 672 21547 2239 21573
rect 2265 21547 2291 21573
rect 2317 21547 2343 21573
rect 2369 21547 17599 21573
rect 17625 21547 17651 21573
rect 17677 21547 17703 21573
rect 17729 21547 24304 21573
rect 672 21530 24304 21547
rect 672 21181 24304 21198
rect 672 21155 9919 21181
rect 9945 21155 9971 21181
rect 9997 21155 10023 21181
rect 10049 21155 24304 21181
rect 672 21138 24304 21155
rect 672 20789 24304 20806
rect 672 20763 2239 20789
rect 2265 20763 2291 20789
rect 2317 20763 2343 20789
rect 2369 20763 17599 20789
rect 17625 20763 17651 20789
rect 17677 20763 17703 20789
rect 17729 20763 24304 20789
rect 672 20746 24304 20763
rect 672 20397 24304 20414
rect 672 20371 9919 20397
rect 9945 20371 9971 20397
rect 9997 20371 10023 20397
rect 10049 20371 24304 20397
rect 672 20354 24304 20371
rect 672 20005 24304 20022
rect 672 19979 2239 20005
rect 2265 19979 2291 20005
rect 2317 19979 2343 20005
rect 2369 19979 17599 20005
rect 17625 19979 17651 20005
rect 17677 19979 17703 20005
rect 17729 19979 24304 20005
rect 672 19962 24304 19979
rect 672 19613 24304 19630
rect 672 19587 9919 19613
rect 9945 19587 9971 19613
rect 9997 19587 10023 19613
rect 10049 19587 24304 19613
rect 672 19570 24304 19587
rect 672 19221 24304 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 24304 19221
rect 672 19178 24304 19195
rect 672 18829 24304 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 24304 18829
rect 672 18786 24304 18803
rect 672 18437 24304 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 24304 18437
rect 672 18394 24304 18411
rect 672 18045 24304 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 24304 18045
rect 672 18002 24304 18019
rect 672 17653 24304 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 24304 17653
rect 672 17610 24304 17627
rect 672 17261 24304 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 24304 17261
rect 672 17218 24304 17235
rect 672 16869 24304 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 24304 16869
rect 672 16826 24304 16843
rect 672 16477 24304 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 24304 16477
rect 672 16434 24304 16451
rect 672 16085 24304 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 24304 16085
rect 672 16042 24304 16059
rect 672 15693 24304 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 24304 15693
rect 672 15650 24304 15667
rect 672 15301 24304 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 24304 15301
rect 672 15258 24304 15275
rect 672 14909 24304 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 24304 14909
rect 672 14866 24304 14883
rect 672 14517 24304 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 24304 14517
rect 672 14474 24304 14491
rect 672 14125 24304 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 24304 14125
rect 672 14082 24304 14099
rect 672 13733 24304 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 24304 13733
rect 672 13690 24304 13707
rect 12049 13511 12055 13537
rect 12081 13511 12087 13537
rect 13169 13511 13175 13537
rect 13201 13511 13207 13537
rect 13505 13511 13511 13537
rect 13537 13511 13543 13537
rect 11607 13425 11633 13431
rect 11607 13393 11633 13399
rect 672 13341 24304 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 24304 13341
rect 672 13298 24304 13315
rect 24095 13033 24121 13039
rect 24095 13001 24121 13007
rect 672 12949 24304 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 24304 12949
rect 672 12906 24304 12923
rect 23983 12809 24009 12815
rect 23983 12777 24009 12783
rect 11601 12727 11607 12753
rect 11633 12727 11639 12753
rect 11881 12727 11887 12753
rect 11913 12727 11919 12753
rect 13001 12727 13007 12753
rect 13033 12727 13039 12753
rect 22801 12727 22807 12753
rect 22833 12727 22839 12753
rect 13791 12697 13817 12703
rect 13791 12665 13817 12671
rect 22639 12641 22665 12647
rect 13505 12615 13511 12641
rect 13537 12615 13543 12641
rect 22639 12609 22665 12615
rect 672 12557 24304 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 24304 12557
rect 672 12514 24304 12531
rect 12335 12473 12361 12479
rect 12335 12441 12361 12447
rect 12783 12473 12809 12479
rect 12783 12441 12809 12447
rect 14345 12391 14351 12417
rect 14377 12391 14383 12417
rect 10537 12335 10543 12361
rect 10569 12335 10575 12361
rect 10761 12335 10767 12361
rect 10793 12335 10799 12361
rect 11825 12335 11831 12361
rect 11857 12335 11863 12361
rect 12945 12335 12951 12361
rect 12977 12335 12983 12361
rect 13393 12335 13399 12361
rect 13425 12335 13431 12361
rect 22857 12335 22863 12361
rect 22889 12335 22895 12361
rect 22639 12305 22665 12311
rect 13113 12279 13119 12305
rect 13145 12279 13151 12305
rect 22639 12273 22665 12279
rect 23983 12249 24009 12255
rect 23983 12217 24009 12223
rect 672 12165 24304 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 24304 12165
rect 672 12122 24304 12139
rect 11551 12025 11577 12031
rect 23815 12025 23841 12031
rect 13393 11999 13399 12025
rect 13425 11999 13431 12025
rect 11551 11993 11577 11999
rect 23815 11993 23841 11999
rect 11657 11943 11663 11969
rect 11689 11943 11695 11969
rect 23703 11857 23729 11863
rect 23703 11825 23729 11831
rect 24095 11857 24121 11863
rect 24095 11825 24121 11831
rect 672 11773 24304 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 24304 11773
rect 672 11730 24304 11747
rect 12167 11689 12193 11695
rect 12167 11657 12193 11663
rect 12615 11689 12641 11695
rect 12615 11657 12641 11663
rect 11831 11633 11857 11639
rect 11831 11601 11857 11607
rect 12279 11633 12305 11639
rect 12279 11601 12305 11607
rect 13113 11551 13119 11577
rect 13145 11551 13151 11577
rect 14177 11551 14183 11577
rect 14209 11551 14215 11577
rect 14401 11551 14407 11577
rect 14433 11551 14439 11577
rect 12335 11465 12361 11471
rect 12335 11433 12361 11439
rect 672 11381 24304 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 24304 11381
rect 672 11338 24304 11355
rect 13281 11159 13287 11185
rect 13313 11159 13319 11185
rect 11433 11103 11439 11129
rect 11465 11103 11471 11129
rect 672 10989 24304 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 24304 10989
rect 672 10946 24304 10963
rect 672 10597 24304 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 24304 10597
rect 672 10554 24304 10571
rect 13337 10487 13343 10513
rect 13369 10487 13375 10513
rect 11433 10375 11439 10401
rect 11465 10375 11471 10401
rect 11769 10375 11775 10401
rect 11801 10375 11807 10401
rect 12889 10375 12895 10401
rect 12921 10375 12927 10401
rect 672 10205 24304 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 24304 10205
rect 672 10162 24304 10179
rect 672 9813 24304 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 24304 9813
rect 672 9770 24304 9787
rect 672 9421 24304 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 24304 9421
rect 672 9378 24304 9395
rect 672 9029 24304 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 24304 9029
rect 672 8986 24304 9003
rect 672 8637 24304 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 24304 8637
rect 672 8594 24304 8611
rect 672 8245 24304 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 24304 8245
rect 672 8202 24304 8219
rect 672 7853 24304 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 24304 7853
rect 672 7810 24304 7827
rect 672 7461 24304 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 24304 7461
rect 672 7418 24304 7435
rect 672 7069 24304 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 24304 7069
rect 672 7026 24304 7043
rect 672 6677 24304 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 24304 6677
rect 672 6634 24304 6651
rect 672 6285 24304 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 24304 6285
rect 672 6242 24304 6259
rect 672 5893 24304 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 24304 5893
rect 672 5850 24304 5867
rect 672 5501 24304 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 24304 5501
rect 672 5458 24304 5475
rect 672 5109 24304 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 24304 5109
rect 672 5066 24304 5083
rect 672 4717 24304 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 24304 4717
rect 672 4674 24304 4691
rect 672 4325 24304 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 24304 4325
rect 672 4282 24304 4299
rect 672 3933 24304 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 24304 3933
rect 672 3890 24304 3907
rect 672 3541 24304 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 24304 3541
rect 672 3498 24304 3515
rect 672 3149 24304 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 24304 3149
rect 672 3106 24304 3123
rect 672 2757 24304 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 24304 2757
rect 672 2714 24304 2731
rect 672 2365 24304 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 24304 2365
rect 672 2322 24304 2339
rect 672 1973 24304 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 24304 1973
rect 672 1930 24304 1947
rect 12559 1833 12585 1839
rect 12559 1801 12585 1807
rect 12279 1665 12305 1671
rect 12279 1633 12305 1639
rect 12895 1665 12921 1671
rect 12895 1633 12921 1639
rect 672 1581 24304 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 24304 1581
rect 672 1538 24304 1555
<< via1 >>
rect 2239 23115 2265 23141
rect 2291 23115 2317 23141
rect 2343 23115 2369 23141
rect 17599 23115 17625 23141
rect 17651 23115 17677 23141
rect 17703 23115 17729 23141
rect 9919 22723 9945 22749
rect 9971 22723 9997 22749
rect 10023 22723 10049 22749
rect 2239 22331 2265 22357
rect 2291 22331 2317 22357
rect 2343 22331 2369 22357
rect 17599 22331 17625 22357
rect 17651 22331 17677 22357
rect 17703 22331 17729 22357
rect 9919 21939 9945 21965
rect 9971 21939 9997 21965
rect 10023 21939 10049 21965
rect 2239 21547 2265 21573
rect 2291 21547 2317 21573
rect 2343 21547 2369 21573
rect 17599 21547 17625 21573
rect 17651 21547 17677 21573
rect 17703 21547 17729 21573
rect 9919 21155 9945 21181
rect 9971 21155 9997 21181
rect 10023 21155 10049 21181
rect 2239 20763 2265 20789
rect 2291 20763 2317 20789
rect 2343 20763 2369 20789
rect 17599 20763 17625 20789
rect 17651 20763 17677 20789
rect 17703 20763 17729 20789
rect 9919 20371 9945 20397
rect 9971 20371 9997 20397
rect 10023 20371 10049 20397
rect 2239 19979 2265 20005
rect 2291 19979 2317 20005
rect 2343 19979 2369 20005
rect 17599 19979 17625 20005
rect 17651 19979 17677 20005
rect 17703 19979 17729 20005
rect 9919 19587 9945 19613
rect 9971 19587 9997 19613
rect 10023 19587 10049 19613
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 12055 13511 12081 13537
rect 13175 13511 13201 13537
rect 13511 13511 13537 13537
rect 11607 13399 11633 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 24095 13007 24121 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 23983 12783 24009 12809
rect 11607 12727 11633 12753
rect 11887 12727 11913 12753
rect 13007 12727 13033 12753
rect 22807 12727 22833 12753
rect 13791 12671 13817 12697
rect 13511 12615 13537 12641
rect 22639 12615 22665 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 12335 12447 12361 12473
rect 12783 12447 12809 12473
rect 14351 12391 14377 12417
rect 10543 12335 10569 12361
rect 10767 12335 10793 12361
rect 11831 12335 11857 12361
rect 12951 12335 12977 12361
rect 13399 12335 13425 12361
rect 22863 12335 22889 12361
rect 13119 12279 13145 12305
rect 22639 12279 22665 12305
rect 23983 12223 24009 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 11551 11999 11577 12025
rect 13399 11999 13425 12025
rect 23815 11999 23841 12025
rect 11663 11943 11689 11969
rect 23703 11831 23729 11857
rect 24095 11831 24121 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 12167 11663 12193 11689
rect 12615 11663 12641 11689
rect 11831 11607 11857 11633
rect 12279 11607 12305 11633
rect 13119 11551 13145 11577
rect 14183 11551 14209 11577
rect 14407 11551 14433 11577
rect 12335 11439 12361 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 13287 11159 13313 11185
rect 11439 11103 11465 11129
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 13343 10487 13369 10513
rect 11439 10375 11465 10401
rect 11775 10375 11801 10401
rect 12895 10375 12921 10401
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 12559 1807 12585 1833
rect 12279 1639 12305 1665
rect 12895 1639 12921 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 2238 23142 2370 23147
rect 2266 23114 2290 23142
rect 2318 23114 2342 23142
rect 2238 23109 2370 23114
rect 17598 23142 17730 23147
rect 17626 23114 17650 23142
rect 17678 23114 17702 23142
rect 17598 23109 17730 23114
rect 9918 22750 10050 22755
rect 9946 22722 9970 22750
rect 9998 22722 10022 22750
rect 9918 22717 10050 22722
rect 2238 22358 2370 22363
rect 2266 22330 2290 22358
rect 2318 22330 2342 22358
rect 2238 22325 2370 22330
rect 17598 22358 17730 22363
rect 17626 22330 17650 22358
rect 17678 22330 17702 22358
rect 17598 22325 17730 22330
rect 9918 21966 10050 21971
rect 9946 21938 9970 21966
rect 9998 21938 10022 21966
rect 9918 21933 10050 21938
rect 2238 21574 2370 21579
rect 2266 21546 2290 21574
rect 2318 21546 2342 21574
rect 2238 21541 2370 21546
rect 17598 21574 17730 21579
rect 17626 21546 17650 21574
rect 17678 21546 17702 21574
rect 17598 21541 17730 21546
rect 9918 21182 10050 21187
rect 9946 21154 9970 21182
rect 9998 21154 10022 21182
rect 9918 21149 10050 21154
rect 2238 20790 2370 20795
rect 2266 20762 2290 20790
rect 2318 20762 2342 20790
rect 2238 20757 2370 20762
rect 17598 20790 17730 20795
rect 17626 20762 17650 20790
rect 17678 20762 17702 20790
rect 17598 20757 17730 20762
rect 9918 20398 10050 20403
rect 9946 20370 9970 20398
rect 9998 20370 10022 20398
rect 9918 20365 10050 20370
rect 2238 20006 2370 20011
rect 2266 19978 2290 20006
rect 2318 19978 2342 20006
rect 2238 19973 2370 19978
rect 17598 20006 17730 20011
rect 17626 19978 17650 20006
rect 17678 19978 17702 20006
rect 17598 19973 17730 19978
rect 9918 19614 10050 19619
rect 9946 19586 9970 19614
rect 9998 19586 10022 19614
rect 9918 19581 10050 19586
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 12054 13538 12082 13543
rect 13174 13538 13202 13543
rect 11830 13537 12082 13538
rect 11830 13511 12055 13537
rect 12081 13511 12082 13537
rect 11830 13510 12082 13511
rect 10766 13426 10794 13431
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10542 12362 10570 12367
rect 10542 12315 10570 12334
rect 10766 12361 10794 13398
rect 11606 13426 11634 13431
rect 11606 13379 11634 13398
rect 11606 12754 11634 12759
rect 11494 12753 11634 12754
rect 11494 12727 11607 12753
rect 11633 12727 11634 12753
rect 11494 12726 11634 12727
rect 10766 12335 10767 12361
rect 10793 12335 10794 12361
rect 10766 12329 10794 12335
rect 11438 12362 11466 12367
rect 11494 12362 11522 12726
rect 11606 12721 11634 12726
rect 11466 12334 11522 12362
rect 11550 12474 11578 12479
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 11438 11129 11466 12334
rect 11550 12026 11578 12446
rect 11830 12362 11858 13510
rect 12054 13505 12082 13510
rect 12614 13537 13202 13538
rect 12614 13511 13175 13537
rect 13201 13511 13202 13537
rect 12614 13510 13202 13511
rect 11886 12754 11914 12759
rect 11886 12753 12362 12754
rect 11886 12727 11887 12753
rect 11913 12727 12362 12753
rect 11886 12726 12362 12727
rect 11886 12721 11914 12726
rect 12334 12473 12362 12726
rect 12334 12447 12335 12473
rect 12361 12447 12362 12473
rect 12334 12441 12362 12447
rect 11830 12315 11858 12334
rect 12278 12306 12306 12311
rect 11550 12025 11690 12026
rect 11550 11999 11551 12025
rect 11577 11999 11690 12025
rect 11550 11998 11690 11999
rect 11550 11993 11578 11998
rect 11662 11969 11690 11998
rect 11662 11943 11663 11969
rect 11689 11943 11690 11969
rect 11662 11937 11690 11943
rect 12166 11690 12194 11695
rect 12278 11690 12306 12278
rect 12166 11689 12306 11690
rect 12166 11663 12167 11689
rect 12193 11663 12306 11689
rect 12166 11662 12306 11663
rect 12166 11657 12194 11662
rect 11830 11634 11858 11639
rect 11438 11103 11439 11129
rect 11465 11103 11466 11129
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 11438 10401 11466 11103
rect 11438 10375 11439 10401
rect 11465 10375 11466 10401
rect 11438 10369 11466 10375
rect 11774 11633 11858 11634
rect 11774 11607 11831 11633
rect 11857 11607 11858 11633
rect 11774 11606 11858 11607
rect 11774 10401 11802 11606
rect 11830 11601 11858 11606
rect 12278 11633 12306 11662
rect 12614 11689 12642 13510
rect 13174 13505 13202 13510
rect 13510 13537 13538 13543
rect 13510 13511 13511 13537
rect 13537 13511 13538 13537
rect 13006 12753 13034 12759
rect 13006 12727 13007 12753
rect 13033 12727 13034 12753
rect 13006 12698 13034 12727
rect 13510 12754 13538 13511
rect 24094 13033 24122 13039
rect 24094 13007 24095 13033
rect 24121 13007 24122 13033
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 23982 12809 24010 12815
rect 23982 12783 23983 12809
rect 24009 12783 24010 12809
rect 13510 12721 13538 12726
rect 14350 12754 14378 12759
rect 12950 12670 13006 12698
rect 12782 12474 12810 12479
rect 12950 12474 12978 12670
rect 13006 12665 13034 12670
rect 13790 12698 13818 12703
rect 13790 12651 13818 12670
rect 12782 12473 12978 12474
rect 12782 12447 12783 12473
rect 12809 12447 12978 12473
rect 12782 12446 12978 12447
rect 12782 12441 12810 12446
rect 12950 12361 12978 12446
rect 13510 12641 13538 12647
rect 13510 12615 13511 12641
rect 13537 12615 13538 12641
rect 12950 12335 12951 12361
rect 12977 12335 12978 12361
rect 12950 12329 12978 12335
rect 13118 12362 13146 12367
rect 12614 11663 12615 11689
rect 12641 11663 12642 11689
rect 12614 11657 12642 11663
rect 13118 12305 13146 12334
rect 13118 12279 13119 12305
rect 13145 12279 13146 12305
rect 12278 11607 12279 11633
rect 12305 11607 12306 11633
rect 12278 11601 12306 11607
rect 13118 11578 13146 12279
rect 12894 11577 13146 11578
rect 12894 11551 13119 11577
rect 13145 11551 13146 11577
rect 12894 11550 13146 11551
rect 12334 11466 12362 11471
rect 12334 11419 12362 11438
rect 11774 10375 11775 10401
rect 11801 10375 11802 10401
rect 11774 10369 11802 10375
rect 12894 10401 12922 11550
rect 13118 11545 13146 11550
rect 13398 12361 13426 12367
rect 13398 12335 13399 12361
rect 13425 12335 13426 12361
rect 13398 12025 13426 12335
rect 13510 12306 13538 12615
rect 14350 12418 14378 12726
rect 22806 12753 22834 12759
rect 22806 12727 22807 12753
rect 22833 12727 22834 12753
rect 22638 12642 22666 12647
rect 22806 12642 22834 12727
rect 22582 12641 22834 12642
rect 22582 12615 22639 12641
rect 22665 12615 22834 12641
rect 22582 12614 22834 12615
rect 23814 12698 23842 12703
rect 14350 12417 14434 12418
rect 14350 12391 14351 12417
rect 14377 12391 14434 12417
rect 14350 12390 14434 12391
rect 14350 12385 14378 12390
rect 13510 12273 13538 12278
rect 13398 11999 13399 12025
rect 13425 11999 13426 12025
rect 13286 11186 13314 11191
rect 13398 11186 13426 11999
rect 13286 11185 13426 11186
rect 13286 11159 13287 11185
rect 13313 11159 13426 11185
rect 13286 11158 13426 11159
rect 14182 11577 14210 11583
rect 14182 11551 14183 11577
rect 14209 11551 14210 11577
rect 13286 11153 13314 11158
rect 13342 10962 13370 10967
rect 13342 10513 13370 10934
rect 14182 10962 14210 11551
rect 14406 11577 14434 12390
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 14406 11551 14407 11577
rect 14433 11551 14434 11577
rect 14406 11545 14434 11551
rect 22526 11466 22554 11471
rect 22582 11466 22610 12614
rect 22638 12609 22666 12614
rect 22862 12361 22890 12367
rect 22862 12335 22863 12361
rect 22889 12335 22890 12361
rect 22638 12306 22666 12311
rect 22638 12259 22666 12278
rect 22862 12306 22890 12335
rect 22862 12273 22890 12278
rect 23814 12025 23842 12670
rect 23982 12474 24010 12783
rect 24094 12810 24122 13007
rect 24094 12777 24122 12782
rect 23982 12441 24010 12446
rect 23982 12249 24010 12255
rect 23982 12223 23983 12249
rect 24009 12223 24010 12249
rect 23982 12138 24010 12223
rect 23982 12105 24010 12110
rect 23814 11999 23815 12025
rect 23841 11999 23842 12025
rect 23814 11993 23842 11999
rect 23702 11857 23730 11863
rect 23702 11831 23703 11857
rect 23729 11831 23730 11857
rect 23702 11802 23730 11831
rect 23702 11769 23730 11774
rect 24094 11857 24122 11863
rect 24094 11831 24095 11857
rect 24121 11831 24122 11857
rect 24094 11802 24122 11831
rect 24094 11769 24122 11774
rect 22554 11438 22610 11466
rect 22526 11433 22554 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 14182 10929 14210 10934
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 13342 10487 13343 10513
rect 13369 10487 13370 10513
rect 13342 10481 13370 10487
rect 12894 10375 12895 10401
rect 12921 10375 12922 10401
rect 12894 10369 12922 10375
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12558 1834 12586 1839
rect 12446 1833 12586 1834
rect 12446 1807 12559 1833
rect 12585 1807 12586 1833
rect 12446 1806 12586 1807
rect 12278 1666 12306 1671
rect 12110 1665 12306 1666
rect 12110 1639 12279 1665
rect 12305 1639 12306 1665
rect 12110 1638 12306 1639
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 12110 400 12138 1638
rect 12278 1633 12306 1638
rect 12446 400 12474 1806
rect 12558 1801 12586 1806
rect 12894 1666 12922 1671
rect 12782 1665 12922 1666
rect 12782 1639 12895 1665
rect 12921 1639 12922 1665
rect 12782 1638 12922 1639
rect 12782 400 12810 1638
rect 12894 1633 12922 1638
rect 12096 0 12152 400
rect 12432 0 12488 400
rect 12768 0 12824 400
<< via2 >>
rect 2238 23141 2266 23142
rect 2238 23115 2239 23141
rect 2239 23115 2265 23141
rect 2265 23115 2266 23141
rect 2238 23114 2266 23115
rect 2290 23141 2318 23142
rect 2290 23115 2291 23141
rect 2291 23115 2317 23141
rect 2317 23115 2318 23141
rect 2290 23114 2318 23115
rect 2342 23141 2370 23142
rect 2342 23115 2343 23141
rect 2343 23115 2369 23141
rect 2369 23115 2370 23141
rect 2342 23114 2370 23115
rect 17598 23141 17626 23142
rect 17598 23115 17599 23141
rect 17599 23115 17625 23141
rect 17625 23115 17626 23141
rect 17598 23114 17626 23115
rect 17650 23141 17678 23142
rect 17650 23115 17651 23141
rect 17651 23115 17677 23141
rect 17677 23115 17678 23141
rect 17650 23114 17678 23115
rect 17702 23141 17730 23142
rect 17702 23115 17703 23141
rect 17703 23115 17729 23141
rect 17729 23115 17730 23141
rect 17702 23114 17730 23115
rect 9918 22749 9946 22750
rect 9918 22723 9919 22749
rect 9919 22723 9945 22749
rect 9945 22723 9946 22749
rect 9918 22722 9946 22723
rect 9970 22749 9998 22750
rect 9970 22723 9971 22749
rect 9971 22723 9997 22749
rect 9997 22723 9998 22749
rect 9970 22722 9998 22723
rect 10022 22749 10050 22750
rect 10022 22723 10023 22749
rect 10023 22723 10049 22749
rect 10049 22723 10050 22749
rect 10022 22722 10050 22723
rect 2238 22357 2266 22358
rect 2238 22331 2239 22357
rect 2239 22331 2265 22357
rect 2265 22331 2266 22357
rect 2238 22330 2266 22331
rect 2290 22357 2318 22358
rect 2290 22331 2291 22357
rect 2291 22331 2317 22357
rect 2317 22331 2318 22357
rect 2290 22330 2318 22331
rect 2342 22357 2370 22358
rect 2342 22331 2343 22357
rect 2343 22331 2369 22357
rect 2369 22331 2370 22357
rect 2342 22330 2370 22331
rect 17598 22357 17626 22358
rect 17598 22331 17599 22357
rect 17599 22331 17625 22357
rect 17625 22331 17626 22357
rect 17598 22330 17626 22331
rect 17650 22357 17678 22358
rect 17650 22331 17651 22357
rect 17651 22331 17677 22357
rect 17677 22331 17678 22357
rect 17650 22330 17678 22331
rect 17702 22357 17730 22358
rect 17702 22331 17703 22357
rect 17703 22331 17729 22357
rect 17729 22331 17730 22357
rect 17702 22330 17730 22331
rect 9918 21965 9946 21966
rect 9918 21939 9919 21965
rect 9919 21939 9945 21965
rect 9945 21939 9946 21965
rect 9918 21938 9946 21939
rect 9970 21965 9998 21966
rect 9970 21939 9971 21965
rect 9971 21939 9997 21965
rect 9997 21939 9998 21965
rect 9970 21938 9998 21939
rect 10022 21965 10050 21966
rect 10022 21939 10023 21965
rect 10023 21939 10049 21965
rect 10049 21939 10050 21965
rect 10022 21938 10050 21939
rect 2238 21573 2266 21574
rect 2238 21547 2239 21573
rect 2239 21547 2265 21573
rect 2265 21547 2266 21573
rect 2238 21546 2266 21547
rect 2290 21573 2318 21574
rect 2290 21547 2291 21573
rect 2291 21547 2317 21573
rect 2317 21547 2318 21573
rect 2290 21546 2318 21547
rect 2342 21573 2370 21574
rect 2342 21547 2343 21573
rect 2343 21547 2369 21573
rect 2369 21547 2370 21573
rect 2342 21546 2370 21547
rect 17598 21573 17626 21574
rect 17598 21547 17599 21573
rect 17599 21547 17625 21573
rect 17625 21547 17626 21573
rect 17598 21546 17626 21547
rect 17650 21573 17678 21574
rect 17650 21547 17651 21573
rect 17651 21547 17677 21573
rect 17677 21547 17678 21573
rect 17650 21546 17678 21547
rect 17702 21573 17730 21574
rect 17702 21547 17703 21573
rect 17703 21547 17729 21573
rect 17729 21547 17730 21573
rect 17702 21546 17730 21547
rect 9918 21181 9946 21182
rect 9918 21155 9919 21181
rect 9919 21155 9945 21181
rect 9945 21155 9946 21181
rect 9918 21154 9946 21155
rect 9970 21181 9998 21182
rect 9970 21155 9971 21181
rect 9971 21155 9997 21181
rect 9997 21155 9998 21181
rect 9970 21154 9998 21155
rect 10022 21181 10050 21182
rect 10022 21155 10023 21181
rect 10023 21155 10049 21181
rect 10049 21155 10050 21181
rect 10022 21154 10050 21155
rect 2238 20789 2266 20790
rect 2238 20763 2239 20789
rect 2239 20763 2265 20789
rect 2265 20763 2266 20789
rect 2238 20762 2266 20763
rect 2290 20789 2318 20790
rect 2290 20763 2291 20789
rect 2291 20763 2317 20789
rect 2317 20763 2318 20789
rect 2290 20762 2318 20763
rect 2342 20789 2370 20790
rect 2342 20763 2343 20789
rect 2343 20763 2369 20789
rect 2369 20763 2370 20789
rect 2342 20762 2370 20763
rect 17598 20789 17626 20790
rect 17598 20763 17599 20789
rect 17599 20763 17625 20789
rect 17625 20763 17626 20789
rect 17598 20762 17626 20763
rect 17650 20789 17678 20790
rect 17650 20763 17651 20789
rect 17651 20763 17677 20789
rect 17677 20763 17678 20789
rect 17650 20762 17678 20763
rect 17702 20789 17730 20790
rect 17702 20763 17703 20789
rect 17703 20763 17729 20789
rect 17729 20763 17730 20789
rect 17702 20762 17730 20763
rect 9918 20397 9946 20398
rect 9918 20371 9919 20397
rect 9919 20371 9945 20397
rect 9945 20371 9946 20397
rect 9918 20370 9946 20371
rect 9970 20397 9998 20398
rect 9970 20371 9971 20397
rect 9971 20371 9997 20397
rect 9997 20371 9998 20397
rect 9970 20370 9998 20371
rect 10022 20397 10050 20398
rect 10022 20371 10023 20397
rect 10023 20371 10049 20397
rect 10049 20371 10050 20397
rect 10022 20370 10050 20371
rect 2238 20005 2266 20006
rect 2238 19979 2239 20005
rect 2239 19979 2265 20005
rect 2265 19979 2266 20005
rect 2238 19978 2266 19979
rect 2290 20005 2318 20006
rect 2290 19979 2291 20005
rect 2291 19979 2317 20005
rect 2317 19979 2318 20005
rect 2290 19978 2318 19979
rect 2342 20005 2370 20006
rect 2342 19979 2343 20005
rect 2343 19979 2369 20005
rect 2369 19979 2370 20005
rect 2342 19978 2370 19979
rect 17598 20005 17626 20006
rect 17598 19979 17599 20005
rect 17599 19979 17625 20005
rect 17625 19979 17626 20005
rect 17598 19978 17626 19979
rect 17650 20005 17678 20006
rect 17650 19979 17651 20005
rect 17651 19979 17677 20005
rect 17677 19979 17678 20005
rect 17650 19978 17678 19979
rect 17702 20005 17730 20006
rect 17702 19979 17703 20005
rect 17703 19979 17729 20005
rect 17729 19979 17730 20005
rect 17702 19978 17730 19979
rect 9918 19613 9946 19614
rect 9918 19587 9919 19613
rect 9919 19587 9945 19613
rect 9945 19587 9946 19613
rect 9918 19586 9946 19587
rect 9970 19613 9998 19614
rect 9970 19587 9971 19613
rect 9971 19587 9997 19613
rect 9997 19587 9998 19613
rect 9970 19586 9998 19587
rect 10022 19613 10050 19614
rect 10022 19587 10023 19613
rect 10023 19587 10049 19613
rect 10049 19587 10050 19613
rect 10022 19586 10050 19587
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 10766 13398 10794 13426
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10542 12361 10570 12362
rect 10542 12335 10543 12361
rect 10543 12335 10569 12361
rect 10569 12335 10570 12361
rect 10542 12334 10570 12335
rect 11606 13425 11634 13426
rect 11606 13399 11607 13425
rect 11607 13399 11633 13425
rect 11633 13399 11634 13425
rect 11606 13398 11634 13399
rect 11438 12334 11466 12362
rect 11550 12446 11578 12474
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 11830 12361 11858 12362
rect 11830 12335 11831 12361
rect 11831 12335 11857 12361
rect 11857 12335 11858 12361
rect 11830 12334 11858 12335
rect 12278 12278 12306 12306
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 13510 12726 13538 12754
rect 14350 12726 14378 12754
rect 13006 12670 13034 12698
rect 13790 12697 13818 12698
rect 13790 12671 13791 12697
rect 13791 12671 13817 12697
rect 13817 12671 13818 12697
rect 13790 12670 13818 12671
rect 13118 12334 13146 12362
rect 12334 11465 12362 11466
rect 12334 11439 12335 11465
rect 12335 11439 12361 11465
rect 12361 11439 12362 11465
rect 12334 11438 12362 11439
rect 23814 12670 23842 12698
rect 13510 12278 13538 12306
rect 13342 10934 13370 10962
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 22638 12305 22666 12306
rect 22638 12279 22639 12305
rect 22639 12279 22665 12305
rect 22665 12279 22666 12305
rect 22638 12278 22666 12279
rect 22862 12278 22890 12306
rect 24094 12782 24122 12810
rect 23982 12446 24010 12474
rect 23982 12110 24010 12138
rect 23702 11774 23730 11802
rect 24094 11774 24122 11802
rect 22526 11438 22554 11466
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 14182 10934 14210 10962
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
<< metal3 >>
rect 2233 23114 2238 23142
rect 2266 23114 2290 23142
rect 2318 23114 2342 23142
rect 2370 23114 2375 23142
rect 17593 23114 17598 23142
rect 17626 23114 17650 23142
rect 17678 23114 17702 23142
rect 17730 23114 17735 23142
rect 9913 22722 9918 22750
rect 9946 22722 9970 22750
rect 9998 22722 10022 22750
rect 10050 22722 10055 22750
rect 2233 22330 2238 22358
rect 2266 22330 2290 22358
rect 2318 22330 2342 22358
rect 2370 22330 2375 22358
rect 17593 22330 17598 22358
rect 17626 22330 17650 22358
rect 17678 22330 17702 22358
rect 17730 22330 17735 22358
rect 9913 21938 9918 21966
rect 9946 21938 9970 21966
rect 9998 21938 10022 21966
rect 10050 21938 10055 21966
rect 2233 21546 2238 21574
rect 2266 21546 2290 21574
rect 2318 21546 2342 21574
rect 2370 21546 2375 21574
rect 17593 21546 17598 21574
rect 17626 21546 17650 21574
rect 17678 21546 17702 21574
rect 17730 21546 17735 21574
rect 9913 21154 9918 21182
rect 9946 21154 9970 21182
rect 9998 21154 10022 21182
rect 10050 21154 10055 21182
rect 2233 20762 2238 20790
rect 2266 20762 2290 20790
rect 2318 20762 2342 20790
rect 2370 20762 2375 20790
rect 17593 20762 17598 20790
rect 17626 20762 17650 20790
rect 17678 20762 17702 20790
rect 17730 20762 17735 20790
rect 9913 20370 9918 20398
rect 9946 20370 9970 20398
rect 9998 20370 10022 20398
rect 10050 20370 10055 20398
rect 2233 19978 2238 20006
rect 2266 19978 2290 20006
rect 2318 19978 2342 20006
rect 2370 19978 2375 20006
rect 17593 19978 17598 20006
rect 17626 19978 17650 20006
rect 17678 19978 17702 20006
rect 17730 19978 17735 20006
rect 9913 19586 9918 19614
rect 9946 19586 9970 19614
rect 9998 19586 10022 19614
rect 10050 19586 10055 19614
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 10761 13398 10766 13426
rect 10794 13398 11606 13426
rect 11634 13398 11639 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 24600 12810 25000 12824
rect 24089 12782 24094 12810
rect 24122 12782 25000 12810
rect 24600 12768 25000 12782
rect 13505 12726 13510 12754
rect 13538 12726 14350 12754
rect 14378 12726 14383 12754
rect 13001 12670 13006 12698
rect 13034 12670 13790 12698
rect 13818 12670 23814 12698
rect 23842 12670 23847 12698
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 0 12474 400 12488
rect 24600 12474 25000 12488
rect 0 12446 11550 12474
rect 11578 12446 11583 12474
rect 23977 12446 23982 12474
rect 24010 12446 25000 12474
rect 0 12432 400 12446
rect 24600 12432 25000 12446
rect 10537 12334 10542 12362
rect 10570 12334 11438 12362
rect 11466 12334 11471 12362
rect 11825 12334 11830 12362
rect 11858 12334 13118 12362
rect 13146 12334 13151 12362
rect 12273 12278 12278 12306
rect 12306 12278 13510 12306
rect 13538 12278 22638 12306
rect 22666 12278 22862 12306
rect 22890 12278 22895 12306
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 24600 12138 25000 12152
rect 23977 12110 23982 12138
rect 24010 12110 25000 12138
rect 24600 12096 25000 12110
rect 24600 11802 25000 11816
rect 23697 11774 23702 11802
rect 23730 11774 24094 11802
rect 24122 11774 25000 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 24600 11760 25000 11774
rect 12329 11438 12334 11466
rect 12362 11438 22526 11466
rect 22554 11438 22559 11466
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 13337 10934 13342 10962
rect 13370 10934 14182 10962
rect 14210 10934 14215 10962
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 23114 2266 23142
rect 2290 23114 2318 23142
rect 2342 23114 2370 23142
rect 17598 23114 17626 23142
rect 17650 23114 17678 23142
rect 17702 23114 17730 23142
rect 9918 22722 9946 22750
rect 9970 22722 9998 22750
rect 10022 22722 10050 22750
rect 2238 22330 2266 22358
rect 2290 22330 2318 22358
rect 2342 22330 2370 22358
rect 17598 22330 17626 22358
rect 17650 22330 17678 22358
rect 17702 22330 17730 22358
rect 9918 21938 9946 21966
rect 9970 21938 9998 21966
rect 10022 21938 10050 21966
rect 2238 21546 2266 21574
rect 2290 21546 2318 21574
rect 2342 21546 2370 21574
rect 17598 21546 17626 21574
rect 17650 21546 17678 21574
rect 17702 21546 17730 21574
rect 9918 21154 9946 21182
rect 9970 21154 9998 21182
rect 10022 21154 10050 21182
rect 2238 20762 2266 20790
rect 2290 20762 2318 20790
rect 2342 20762 2370 20790
rect 17598 20762 17626 20790
rect 17650 20762 17678 20790
rect 17702 20762 17730 20790
rect 9918 20370 9946 20398
rect 9970 20370 9998 20398
rect 10022 20370 10050 20398
rect 2238 19978 2266 20006
rect 2290 19978 2318 20006
rect 2342 19978 2370 20006
rect 17598 19978 17626 20006
rect 17650 19978 17678 20006
rect 17702 19978 17730 20006
rect 9918 19586 9946 19614
rect 9970 19586 9998 19614
rect 10022 19586 10050 19614
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 23142 2384 23158
rect 2224 23114 2238 23142
rect 2266 23114 2290 23142
rect 2318 23114 2342 23142
rect 2370 23114 2384 23142
rect 2224 22358 2384 23114
rect 2224 22330 2238 22358
rect 2266 22330 2290 22358
rect 2318 22330 2342 22358
rect 2370 22330 2384 22358
rect 2224 21574 2384 22330
rect 2224 21546 2238 21574
rect 2266 21546 2290 21574
rect 2318 21546 2342 21574
rect 2370 21546 2384 21574
rect 2224 20790 2384 21546
rect 2224 20762 2238 20790
rect 2266 20762 2290 20790
rect 2318 20762 2342 20790
rect 2370 20762 2384 20790
rect 2224 20006 2384 20762
rect 2224 19978 2238 20006
rect 2266 19978 2290 20006
rect 2318 19978 2342 20006
rect 2370 19978 2384 20006
rect 2224 19222 2384 19978
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 22750 10064 23158
rect 9904 22722 9918 22750
rect 9946 22722 9970 22750
rect 9998 22722 10022 22750
rect 10050 22722 10064 22750
rect 9904 21966 10064 22722
rect 9904 21938 9918 21966
rect 9946 21938 9970 21966
rect 9998 21938 10022 21966
rect 10050 21938 10064 21966
rect 9904 21182 10064 21938
rect 9904 21154 9918 21182
rect 9946 21154 9970 21182
rect 9998 21154 10022 21182
rect 10050 21154 10064 21182
rect 9904 20398 10064 21154
rect 9904 20370 9918 20398
rect 9946 20370 9970 20398
rect 9998 20370 10022 20398
rect 10050 20370 10064 20398
rect 9904 19614 10064 20370
rect 9904 19586 9918 19614
rect 9946 19586 9970 19614
rect 9998 19586 10022 19614
rect 10050 19586 10064 19614
rect 9904 18830 10064 19586
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 23142 17744 23158
rect 17584 23114 17598 23142
rect 17626 23114 17650 23142
rect 17678 23114 17702 23142
rect 17730 23114 17744 23142
rect 17584 22358 17744 23114
rect 17584 22330 17598 22358
rect 17626 22330 17650 22358
rect 17678 22330 17702 22358
rect 17730 22330 17744 22358
rect 17584 21574 17744 22330
rect 17584 21546 17598 21574
rect 17626 21546 17650 21574
rect 17678 21546 17702 21574
rect 17730 21546 17744 21574
rect 17584 20790 17744 21546
rect 17584 20762 17598 20790
rect 17626 20762 17650 20790
rect 17678 20762 17702 20790
rect 17730 20762 17744 20790
rect 17584 20006 17744 20762
rect 17584 19978 17598 20006
rect 17626 19978 17650 20006
rect 17678 19978 17702 20006
rect 17730 19978 17744 20006
rect 17584 19222 17744 19978
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _01_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12208 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  _02__6 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11984 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _02_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11424 0 1 10192
box -43 -43 2059 435
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _03_
timestamp 1698431365
transform -1 0 14560 0 -1 11760
box -43 -43 2059 435
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _04_
timestamp 1698431365
transform -1 0 13552 0 1 13328
box -43 -43 2059 435
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _05_
timestamp 1698431365
transform 1 0 10416 0 -1 12544
box -43 -43 2059 435
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_2  _06_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11536 0 1 12544
box -43 -43 2171 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__01__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12208 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__06__SETN
timestamp 1698431365
transform 1 0 13776 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_ctrl_in[0]_I
timestamp 1698431365
transform -1 0 11592 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout1_I
timestamp 1698431365
transform -1 0 12824 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 23744 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output2_I
timestamp 1698431365
transform 1 0 22624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output3_I
timestamp 1698431365
transform 1 0 22624 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_ctrl_in[0] dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11592 0 1 11760
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_ctrl_in[0]
timestamp 1698431365
transform -1 0 13384 0 1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_ctrl_in[0]
timestamp 1698431365
transform 1 0 13272 0 -1 12544
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ctrl_4
timestamp 1698431365
transform -1 0 13048 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ctrl_5
timestamp 1698431365
transform -1 0 12432 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tieh  ctrl_7 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23968 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tieh  ctrl_8
timestamp 1698431365
transform -1 0 12712 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12824 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 8400 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 10304 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12432 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_215 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_221 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13048 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 13944 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 19824 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698431365
transform 1 0 21728 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_410 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23632 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_418
timestamp 1698431365
transform 1 0 24080 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 8624 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 12208 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 20048 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698431365
transform 1 0 20384 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698431365
transform 1 0 23968 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 18424 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 22008 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_387
timestamp 1698431365
transform 1 0 22344 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_419
timestamp 1698431365
transform 1 0 24136 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 20048 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 20384 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 23968 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 18424 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 22008 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_387
timestamp 1698431365
transform 1 0 22344 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_419
timestamp 1698431365
transform 1 0 24136 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 20048 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698431365
transform 1 0 20384 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698431365
transform 1 0 23968 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 18424 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698431365
transform 1 0 22008 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_387
timestamp 1698431365
transform 1 0 22344 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_419
timestamp 1698431365
transform 1 0 24136 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 20048 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698431365
transform 1 0 20384 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698431365
transform 1 0 23968 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 18424 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698431365
transform 1 0 22008 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_387
timestamp 1698431365
transform 1 0 22344 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_419
timestamp 1698431365
transform 1 0 24136 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 20048 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1698431365
transform 1 0 20384 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698431365
transform 1 0 23968 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698431365
transform 1 0 18424 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698431365
transform 1 0 22008 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_387
timestamp 1698431365
transform 1 0 22344 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_419
timestamp 1698431365
transform 1 0 24136 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698431365
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698431365
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1698431365
transform 1 0 20048 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1698431365
transform 1 0 20384 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698431365
transform 1 0 23968 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698431365
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698431365
transform 1 0 18424 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1698431365
transform 1 0 22008 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_387
timestamp 1698431365
transform 1 0 22344 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_419
timestamp 1698431365
transform 1 0 24136 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698431365
transform 1 0 8624 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 12208 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698431365
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698431365
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698431365
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1698431365
transform 1 0 20048 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698431365
transform 1 0 20384 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698431365
transform 1 0 23968 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698431365
transform 1 0 6664 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698431365
transform 1 0 10248 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698431365
transform 1 0 10584 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698431365
transform 1 0 14168 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698431365
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698431365
transform 1 0 18424 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698431365
transform 1 0 22008 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_387
timestamp 1698431365
transform 1 0 22344 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_419
timestamp 1698431365
transform 1 0 24136 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 4704 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 8288 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698431365
transform 1 0 8624 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698431365
transform 1 0 12208 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698431365
transform 1 0 12544 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698431365
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698431365
transform 1 0 20048 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698431365
transform 1 0 20384 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698431365
transform 1 0 23968 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698431365
transform 1 0 6664 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698431365
transform 1 0 10248 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698431365
transform 1 0 10584 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698431365
transform 1 0 14168 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698431365
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698431365
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698431365
transform 1 0 18424 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698431365
transform 1 0 22008 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_387
timestamp 1698431365
transform 1 0 22344 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_419
timestamp 1698431365
transform 1 0 24136 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698431365
transform 1 0 4704 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 8288 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698431365
transform 1 0 8624 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698431365
transform 1 0 12208 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698431365
transform 1 0 12544 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698431365
transform 1 0 16128 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698431365
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1698431365
transform 1 0 20048 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698431365
transform 1 0 20384 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698431365
transform 1 0 23968 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698431365
transform 1 0 6664 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698431365
transform 1 0 10248 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698431365
transform 1 0 10584 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 14168 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698431365
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_317
timestamp 1698431365
transform 1 0 18424 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698431365
transform 1 0 22008 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_387
timestamp 1698431365
transform 1 0 22344 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_419
timestamp 1698431365
transform 1 0 24136 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 4704 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698431365
transform 1 0 8288 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698431365
transform 1 0 8624 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698431365
transform 1 0 12208 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698431365
transform 1 0 12544 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698431365
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698431365
transform 1 0 20048 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698431365
transform 1 0 20384 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698431365
transform 1 0 23968 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698431365
transform 1 0 6664 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 10248 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698431365
transform 1 0 10584 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 14168 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698431365
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_317
timestamp 1698431365
transform 1 0 18424 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_381
timestamp 1698431365
transform 1 0 22008 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_387
timestamp 1698431365
transform 1 0 22344 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_419
timestamp 1698431365
transform 1 0 24136 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698431365
transform 1 0 4704 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 8288 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_142
timestamp 1698431365
transform 1 0 8624 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698431365
transform 1 0 12208 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698431365
transform 1 0 12544 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 16128 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698431365
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_346
timestamp 1698431365
transform 1 0 20048 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_352
timestamp 1698431365
transform 1 0 20384 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_416
timestamp 1698431365
transform 1 0 23968 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698431365
transform 1 0 6664 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 10248 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_177
timestamp 1698431365
transform 1 0 10584 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_185
timestamp 1698431365
transform 1 0 11032 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_189
timestamp 1698431365
transform 1 0 11256 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_191
timestamp 1698431365
transform 1 0 11368 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_228
timestamp 1698431365
transform 1 0 13440 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698431365
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_317
timestamp 1698431365
transform 1 0 18424 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_381
timestamp 1698431365
transform 1 0 22008 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_387
timestamp 1698431365
transform 1 0 22344 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_419
timestamp 1698431365
transform 1 0 24136 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698431365
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 4704 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 8288 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698431365
transform 1 0 8624 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 12208 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698431365
transform 1 0 12544 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 16128 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698431365
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_346
timestamp 1698431365
transform 1 0 20048 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_352
timestamp 1698431365
transform 1 0 20384 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_416
timestamp 1698431365
transform 1 0 23968 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 6664 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 10248 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_227
timestamp 1698431365
transform 1 0 13384 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698431365
transform 1 0 14280 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698431365
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_317
timestamp 1698431365
transform 1 0 18424 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_381
timestamp 1698431365
transform 1 0 22008 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_387
timestamp 1698431365
transform 1 0 22344 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_419
timestamp 1698431365
transform 1 0 24136 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698431365
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698431365
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 4704 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 8288 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_142
timestamp 1698431365
transform 1 0 8624 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_174
timestamp 1698431365
transform 1 0 10416 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_190
timestamp 1698431365
transform 1 0 11312 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_202
timestamp 1698431365
transform 1 0 11984 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_248
timestamp 1698431365
transform 1 0 14560 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698431365
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_346
timestamp 1698431365
transform 1 0 20048 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_352
timestamp 1698431365
transform 1 0 20384 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698431365
transform 1 0 23968 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_107
timestamp 1698431365
transform 1 0 6664 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 10248 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_177
timestamp 1698431365
transform 1 0 10584 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698431365
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_317
timestamp 1698431365
transform 1 0 18424 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_381
timestamp 1698431365
transform 1 0 22008 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_387
timestamp 1698431365
transform 1 0 22344 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_403
timestamp 1698431365
transform 1 0 23240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_407
timestamp 1698431365
transform 1 0 23464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_409
timestamp 1698431365
transform 1 0 23576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698431365
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698431365
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 4704 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_142
timestamp 1698431365
transform 1 0 8624 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698431365
transform 1 0 12544 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_214
timestamp 1698431365
transform 1 0 12656 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_275
timestamp 1698431365
transform 1 0 16072 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698431365
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_346
timestamp 1698431365
transform 1 0 20048 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_352
timestamp 1698431365
transform 1 0 20384 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_384
timestamp 1698431365
transform 1 0 22176 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698431365
transform 1 0 6664 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 10248 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_177
timestamp 1698431365
transform 1 0 10584 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_193
timestamp 1698431365
transform 1 0 11480 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_232
timestamp 1698431365
transform 1 0 13664 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_236
timestamp 1698431365
transform 1 0 13888 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698431365
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698431365
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_317
timestamp 1698431365
transform 1 0 18424 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_381
timestamp 1698431365
transform 1 0 22008 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_387
timestamp 1698431365
transform 1 0 22344 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_391
timestamp 1698431365
transform 1 0 22568 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698431365
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698431365
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 4704 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 8288 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698431365
transform 1 0 8624 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 12208 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 12544 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 16128 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698431365
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_346
timestamp 1698431365
transform 1 0 20048 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_352
timestamp 1698431365
transform 1 0 20384 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 6664 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 10248 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_177
timestamp 1698431365
transform 1 0 10584 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_193
timestamp 1698431365
transform 1 0 11480 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_230
timestamp 1698431365
transform 1 0 13552 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698431365
transform 1 0 14000 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_317
timestamp 1698431365
transform 1 0 18424 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_381
timestamp 1698431365
transform 1 0 22008 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_387
timestamp 1698431365
transform 1 0 22344 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_419
timestamp 1698431365
transform 1 0 24136 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698431365
transform 1 0 8624 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 12208 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698431365
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698431365
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_346
timestamp 1698431365
transform 1 0 20048 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_352
timestamp 1698431365
transform 1 0 20384 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698431365
transform 1 0 23968 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_317
timestamp 1698431365
transform 1 0 18424 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_381
timestamp 1698431365
transform 1 0 22008 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_387
timestamp 1698431365
transform 1 0 22344 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_419
timestamp 1698431365
transform 1 0 24136 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698431365
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698431365
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_346
timestamp 1698431365
transform 1 0 20048 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_352
timestamp 1698431365
transform 1 0 20384 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_416
timestamp 1698431365
transform 1 0 23968 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_317
timestamp 1698431365
transform 1 0 18424 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_381
timestamp 1698431365
transform 1 0 22008 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_387
timestamp 1698431365
transform 1 0 22344 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_419
timestamp 1698431365
transform 1 0 24136 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698431365
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698431365
transform 1 0 20048 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_352
timestamp 1698431365
transform 1 0 20384 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_416
timestamp 1698431365
transform 1 0 23968 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_317
timestamp 1698431365
transform 1 0 18424 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_381
timestamp 1698431365
transform 1 0 22008 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_387
timestamp 1698431365
transform 1 0 22344 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_419
timestamp 1698431365
transform 1 0 24136 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698431365
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698431365
transform 1 0 20048 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_352
timestamp 1698431365
transform 1 0 20384 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_416
timestamp 1698431365
transform 1 0 23968 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_317
timestamp 1698431365
transform 1 0 18424 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_381
timestamp 1698431365
transform 1 0 22008 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_387
timestamp 1698431365
transform 1 0 22344 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_419
timestamp 1698431365
transform 1 0 24136 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698431365
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_346
timestamp 1698431365
transform 1 0 20048 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_352
timestamp 1698431365
transform 1 0 20384 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_416
timestamp 1698431365
transform 1 0 23968 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_317
timestamp 1698431365
transform 1 0 18424 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_381
timestamp 1698431365
transform 1 0 22008 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_387
timestamp 1698431365
transform 1 0 22344 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_419
timestamp 1698431365
transform 1 0 24136 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 20048 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_352
timestamp 1698431365
transform 1 0 20384 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698431365
transform 1 0 23968 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698431365
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698431365
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_317
timestamp 1698431365
transform 1 0 18424 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_381
timestamp 1698431365
transform 1 0 22008 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_387
timestamp 1698431365
transform 1 0 22344 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_419
timestamp 1698431365
transform 1 0 24136 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698431365
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 8624 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 12208 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698431365
transform 1 0 12544 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 16128 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698431365
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_346
timestamp 1698431365
transform 1 0 20048 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_352
timestamp 1698431365
transform 1 0 20384 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1698431365
transform 1 0 23968 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 2576 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 2744 0 1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 6328 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 6664 0 1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 10248 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 10584 0 1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 14168 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 14504 0 1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 18088 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_317
timestamp 1698431365
transform 1 0 18424 0 1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_381
timestamp 1698431365
transform 1 0 22008 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_387
timestamp 1698431365
transform 1 0 22344 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_419
timestamp 1698431365
transform 1 0 24136 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 784 0 -1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 4368 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 4704 0 -1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 8288 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 8624 0 -1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 12208 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 12544 0 -1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 16128 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_282
timestamp 1698431365
transform 1 0 16464 0 -1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698431365
transform 1 0 20048 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_352
timestamp 1698431365
transform 1 0 20384 0 -1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_416
timestamp 1698431365
transform 1 0 23968 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 784 0 1 19600
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 2576 0 1 19600
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 2744 0 1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 6328 0 1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 6664 0 1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 10248 0 1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 10584 0 1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 14168 0 1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 14504 0 1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 18088 0 1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_317
timestamp 1698431365
transform 1 0 18424 0 1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698431365
transform 1 0 22008 0 1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_387
timestamp 1698431365
transform 1 0 22344 0 1 19600
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_419
timestamp 1698431365
transform 1 0 24136 0 1 19600
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 784 0 -1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 4368 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 4704 0 -1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 8288 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 8624 0 -1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 12208 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 12544 0 -1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 16128 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_282
timestamp 1698431365
transform 1 0 16464 0 -1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698431365
transform 1 0 20048 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698431365
transform 1 0 20384 0 -1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 23968 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 784 0 1 20384
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 2576 0 1 20384
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 2744 0 1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 6328 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 6664 0 1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 10248 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 10584 0 1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 14168 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 14504 0 1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 18088 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698431365
transform 1 0 18424 0 1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 22008 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_387
timestamp 1698431365
transform 1 0 22344 0 1 20384
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_419
timestamp 1698431365
transform 1 0 24136 0 1 20384
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698431365
transform 1 0 784 0 -1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 4368 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698431365
transform 1 0 4704 0 -1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698431365
transform 1 0 8288 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698431365
transform 1 0 8624 0 -1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698431365
transform 1 0 12208 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_212
timestamp 1698431365
transform 1 0 12544 0 -1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698431365
transform 1 0 16128 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_282
timestamp 1698431365
transform 1 0 16464 0 -1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_346
timestamp 1698431365
transform 1 0 20048 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_352
timestamp 1698431365
transform 1 0 20384 0 -1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_416
timestamp 1698431365
transform 1 0 23968 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 784 0 1 21168
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 2576 0 1 21168
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 2744 0 1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 6328 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_107
timestamp 1698431365
transform 1 0 6664 0 1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_171
timestamp 1698431365
transform 1 0 10248 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_177
timestamp 1698431365
transform 1 0 10584 0 1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698431365
transform 1 0 14168 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_247
timestamp 1698431365
transform 1 0 14504 0 1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_311
timestamp 1698431365
transform 1 0 18088 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_317
timestamp 1698431365
transform 1 0 18424 0 1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 22008 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_387
timestamp 1698431365
transform 1 0 22344 0 1 21168
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_419
timestamp 1698431365
transform 1 0 24136 0 1 21168
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2
timestamp 1698431365
transform 1 0 784 0 -1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698431365
transform 1 0 4368 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_72
timestamp 1698431365
transform 1 0 4704 0 -1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 8288 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_142
timestamp 1698431365
transform 1 0 8624 0 -1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698431365
transform 1 0 12208 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_212
timestamp 1698431365
transform 1 0 12544 0 -1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_276
timestamp 1698431365
transform 1 0 16128 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_282
timestamp 1698431365
transform 1 0 16464 0 -1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_346
timestamp 1698431365
transform 1 0 20048 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_352
timestamp 1698431365
transform 1 0 20384 0 -1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_416
timestamp 1698431365
transform 1 0 23968 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 784 0 1 21952
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 2576 0 1 21952
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1698431365
transform 1 0 2744 0 1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698431365
transform 1 0 6328 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_107
timestamp 1698431365
transform 1 0 6664 0 1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_171
timestamp 1698431365
transform 1 0 10248 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_177
timestamp 1698431365
transform 1 0 10584 0 1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_241
timestamp 1698431365
transform 1 0 14168 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_247
timestamp 1698431365
transform 1 0 14504 0 1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_311
timestamp 1698431365
transform 1 0 18088 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_317
timestamp 1698431365
transform 1 0 18424 0 1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_381
timestamp 1698431365
transform 1 0 22008 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_387
timestamp 1698431365
transform 1 0 22344 0 1 21952
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_419
timestamp 1698431365
transform 1 0 24136 0 1 21952
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698431365
transform 1 0 784 0 -1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698431365
transform 1 0 4368 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_72
timestamp 1698431365
transform 1 0 4704 0 -1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1698431365
transform 1 0 8288 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_142
timestamp 1698431365
transform 1 0 8624 0 -1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_206
timestamp 1698431365
transform 1 0 12208 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_212
timestamp 1698431365
transform 1 0 12544 0 -1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_276
timestamp 1698431365
transform 1 0 16128 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_282
timestamp 1698431365
transform 1 0 16464 0 -1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_346
timestamp 1698431365
transform 1 0 20048 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_352
timestamp 1698431365
transform 1 0 20384 0 -1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_416
timestamp 1698431365
transform 1 0 23968 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 784 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_36
timestamp 1698431365
transform 1 0 2688 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_70
timestamp 1698431365
transform 1 0 4592 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_104
timestamp 1698431365
transform 1 0 6496 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_138
timestamp 1698431365
transform 1 0 8400 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_172
timestamp 1698431365
transform 1 0 10304 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_206
timestamp 1698431365
transform 1 0 12208 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_240
timestamp 1698431365
transform 1 0 14112 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_274
timestamp 1698431365
transform 1 0 16016 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_308
timestamp 1698431365
transform 1 0 17920 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_342
timestamp 1698431365
transform 1 0 19824 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_376
timestamp 1698431365
transform 1 0 21728 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_410
timestamp 1698431365
transform 1 0 23632 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_418
timestamp 1698431365
transform 1 0 24080 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input1
timestamp 1698431365
transform -1 0 24192 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22736 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698431365
transform 1 0 22736 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_55 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 24304 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_56
timestamp 1698431365
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 24304 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_57
timestamp 1698431365
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 24304 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_58
timestamp 1698431365
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 24304 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_59
timestamp 1698431365
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 24304 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_60
timestamp 1698431365
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 24304 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_61
timestamp 1698431365
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 24304 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_62
timestamp 1698431365
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 24304 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_63
timestamp 1698431365
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 24304 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_64
timestamp 1698431365
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 24304 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_65
timestamp 1698431365
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 24304 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_66
timestamp 1698431365
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 24304 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_67
timestamp 1698431365
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 24304 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_68
timestamp 1698431365
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 24304 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_69
timestamp 1698431365
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 24304 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_70
timestamp 1698431365
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 24304 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_71
timestamp 1698431365
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 24304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_72
timestamp 1698431365
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 24304 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_73
timestamp 1698431365
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 24304 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_74
timestamp 1698431365
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 24304 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_75
timestamp 1698431365
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 24304 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_76
timestamp 1698431365
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 24304 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_77
timestamp 1698431365
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 24304 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_78
timestamp 1698431365
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 24304 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_79
timestamp 1698431365
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 24304 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_80
timestamp 1698431365
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 24304 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_81
timestamp 1698431365
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 24304 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_82
timestamp 1698431365
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 24304 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_83
timestamp 1698431365
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 24304 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_84
timestamp 1698431365
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 24304 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_85
timestamp 1698431365
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 24304 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_86
timestamp 1698431365
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 24304 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_87
timestamp 1698431365
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 24304 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_88
timestamp 1698431365
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 24304 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_89
timestamp 1698431365
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 24304 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_90
timestamp 1698431365
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 24304 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_91
timestamp 1698431365
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 24304 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_92
timestamp 1698431365
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 24304 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_93
timestamp 1698431365
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 24304 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_94
timestamp 1698431365
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 24304 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_95
timestamp 1698431365
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 24304 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_96
timestamp 1698431365
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 24304 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_97
timestamp 1698431365
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 24304 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_98
timestamp 1698431365
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 24304 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_99
timestamp 1698431365
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 24304 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_100
timestamp 1698431365
transform 1 0 672 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 24304 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_101
timestamp 1698431365
transform 1 0 672 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 24304 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_102
timestamp 1698431365
transform 1 0 672 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 24304 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_103
timestamp 1698431365
transform 1 0 672 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 24304 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_104
timestamp 1698431365
transform 1 0 672 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 24304 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_105
timestamp 1698431365
transform 1 0 672 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 24304 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_106
timestamp 1698431365
transform 1 0 672 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 24304 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_107
timestamp 1698431365
transform 1 0 672 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 24304 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_108
timestamp 1698431365
transform 1 0 672 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 24304 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_109
timestamp 1698431365
transform 1 0 672 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 24304 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_118
timestamp 1698431365
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_119
timestamp 1698431365
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_120
timestamp 1698431365
transform 1 0 21616 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_121
timestamp 1698431365
transform 1 0 23520 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_122
timestamp 1698431365
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_123
timestamp 1698431365
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_124
timestamp 1698431365
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_125
timestamp 1698431365
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_126
timestamp 1698431365
transform 1 0 20272 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_128
timestamp 1698431365
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_129
timestamp 1698431365
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_130
timestamp 1698431365
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_131
timestamp 1698431365
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_132
timestamp 1698431365
transform 1 0 22232 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_133
timestamp 1698431365
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_134
timestamp 1698431365
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_135
timestamp 1698431365
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_136
timestamp 1698431365
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_137
timestamp 1698431365
transform 1 0 20272 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_138
timestamp 1698431365
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_139
timestamp 1698431365
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_140
timestamp 1698431365
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_141
timestamp 1698431365
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_142
timestamp 1698431365
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_143
timestamp 1698431365
transform 1 0 22232 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_144
timestamp 1698431365
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_145
timestamp 1698431365
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_146
timestamp 1698431365
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_147
timestamp 1698431365
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_148
timestamp 1698431365
transform 1 0 20272 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_149
timestamp 1698431365
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_150
timestamp 1698431365
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_151
timestamp 1698431365
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_152
timestamp 1698431365
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_153
timestamp 1698431365
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_154
timestamp 1698431365
transform 1 0 22232 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_155
timestamp 1698431365
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_156
timestamp 1698431365
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_157
timestamp 1698431365
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_158
timestamp 1698431365
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_159
timestamp 1698431365
transform 1 0 20272 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_160
timestamp 1698431365
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_161
timestamp 1698431365
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_162
timestamp 1698431365
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_163
timestamp 1698431365
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_164
timestamp 1698431365
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_165
timestamp 1698431365
transform 1 0 22232 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_166
timestamp 1698431365
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_167
timestamp 1698431365
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_168
timestamp 1698431365
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_169
timestamp 1698431365
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_170
timestamp 1698431365
transform 1 0 20272 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_171
timestamp 1698431365
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_172
timestamp 1698431365
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_173
timestamp 1698431365
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_174
timestamp 1698431365
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_175
timestamp 1698431365
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_176
timestamp 1698431365
transform 1 0 22232 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_177
timestamp 1698431365
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_178
timestamp 1698431365
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_179
timestamp 1698431365
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_180
timestamp 1698431365
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_181
timestamp 1698431365
transform 1 0 20272 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1698431365
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_183
timestamp 1698431365
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_184
timestamp 1698431365
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_185
timestamp 1698431365
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_186
timestamp 1698431365
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_187
timestamp 1698431365
transform 1 0 22232 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_188
timestamp 1698431365
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_189
timestamp 1698431365
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_190
timestamp 1698431365
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_191
timestamp 1698431365
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_192
timestamp 1698431365
transform 1 0 20272 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_193
timestamp 1698431365
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_194
timestamp 1698431365
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_195
timestamp 1698431365
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_196
timestamp 1698431365
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_197
timestamp 1698431365
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_198
timestamp 1698431365
transform 1 0 22232 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_199
timestamp 1698431365
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_200
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_201
timestamp 1698431365
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_202
timestamp 1698431365
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_203
timestamp 1698431365
transform 1 0 20272 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_204
timestamp 1698431365
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_205
timestamp 1698431365
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_206
timestamp 1698431365
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_207
timestamp 1698431365
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_208
timestamp 1698431365
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_209
timestamp 1698431365
transform 1 0 22232 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_210
timestamp 1698431365
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_211
timestamp 1698431365
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_212
timestamp 1698431365
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_213
timestamp 1698431365
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_214
timestamp 1698431365
transform 1 0 20272 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_215
timestamp 1698431365
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_216
timestamp 1698431365
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_217
timestamp 1698431365
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_218
timestamp 1698431365
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_219
timestamp 1698431365
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_220
timestamp 1698431365
transform 1 0 22232 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_221
timestamp 1698431365
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_222
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_223
timestamp 1698431365
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_224
timestamp 1698431365
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_225
timestamp 1698431365
transform 1 0 20272 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_226
timestamp 1698431365
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_227
timestamp 1698431365
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_228
timestamp 1698431365
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_229
timestamp 1698431365
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_230
timestamp 1698431365
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_231
timestamp 1698431365
transform 1 0 22232 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_232
timestamp 1698431365
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_233
timestamp 1698431365
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_234
timestamp 1698431365
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_235
timestamp 1698431365
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_236
timestamp 1698431365
transform 1 0 20272 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_237
timestamp 1698431365
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_238
timestamp 1698431365
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_239
timestamp 1698431365
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_240
timestamp 1698431365
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_241
timestamp 1698431365
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_242
timestamp 1698431365
transform 1 0 22232 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_243
timestamp 1698431365
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_244
timestamp 1698431365
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_245
timestamp 1698431365
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_246
timestamp 1698431365
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_247
timestamp 1698431365
transform 1 0 20272 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_248
timestamp 1698431365
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_249
timestamp 1698431365
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_250
timestamp 1698431365
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_251
timestamp 1698431365
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_252
timestamp 1698431365
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_253
timestamp 1698431365
transform 1 0 22232 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_254
timestamp 1698431365
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_255
timestamp 1698431365
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_256
timestamp 1698431365
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_257
timestamp 1698431365
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_258
timestamp 1698431365
transform 1 0 20272 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_259
timestamp 1698431365
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_260
timestamp 1698431365
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_261
timestamp 1698431365
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_262
timestamp 1698431365
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_263
timestamp 1698431365
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_264
timestamp 1698431365
transform 1 0 22232 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_265
timestamp 1698431365
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_266
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_267
timestamp 1698431365
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_268
timestamp 1698431365
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_269
timestamp 1698431365
transform 1 0 20272 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_270
timestamp 1698431365
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_271
timestamp 1698431365
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_272
timestamp 1698431365
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_273
timestamp 1698431365
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_274
timestamp 1698431365
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_275
timestamp 1698431365
transform 1 0 22232 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_276
timestamp 1698431365
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_277
timestamp 1698431365
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_278
timestamp 1698431365
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_279
timestamp 1698431365
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_280
timestamp 1698431365
transform 1 0 20272 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_281
timestamp 1698431365
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_282
timestamp 1698431365
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_283
timestamp 1698431365
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_284
timestamp 1698431365
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_285
timestamp 1698431365
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_286
timestamp 1698431365
transform 1 0 22232 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_287
timestamp 1698431365
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_288
timestamp 1698431365
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_289
timestamp 1698431365
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_290
timestamp 1698431365
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_291
timestamp 1698431365
transform 1 0 20272 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_292
timestamp 1698431365
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_293
timestamp 1698431365
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_294
timestamp 1698431365
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_295
timestamp 1698431365
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_296
timestamp 1698431365
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_297
timestamp 1698431365
transform 1 0 22232 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_298
timestamp 1698431365
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_299
timestamp 1698431365
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_300
timestamp 1698431365
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_301
timestamp 1698431365
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_302
timestamp 1698431365
transform 1 0 20272 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_303
timestamp 1698431365
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_304
timestamp 1698431365
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_305
timestamp 1698431365
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_306
timestamp 1698431365
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_307
timestamp 1698431365
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_308
timestamp 1698431365
transform 1 0 22232 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_309
timestamp 1698431365
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_310
timestamp 1698431365
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_311
timestamp 1698431365
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_312
timestamp 1698431365
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_313
timestamp 1698431365
transform 1 0 20272 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_314
timestamp 1698431365
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_315
timestamp 1698431365
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_316
timestamp 1698431365
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_317
timestamp 1698431365
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_318
timestamp 1698431365
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_319
timestamp 1698431365
transform 1 0 22232 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_320
timestamp 1698431365
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_321
timestamp 1698431365
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_322
timestamp 1698431365
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_323
timestamp 1698431365
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_324
timestamp 1698431365
transform 1 0 20272 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_325
timestamp 1698431365
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_326
timestamp 1698431365
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_327
timestamp 1698431365
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_328
timestamp 1698431365
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_329
timestamp 1698431365
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_330
timestamp 1698431365
transform 1 0 22232 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_331
timestamp 1698431365
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_332
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_333
timestamp 1698431365
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_334
timestamp 1698431365
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_335
timestamp 1698431365
transform 1 0 20272 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_336
timestamp 1698431365
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_337
timestamp 1698431365
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_338
timestamp 1698431365
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_339
timestamp 1698431365
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_340
timestamp 1698431365
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_341
timestamp 1698431365
transform 1 0 22232 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_342
timestamp 1698431365
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_343
timestamp 1698431365
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_344
timestamp 1698431365
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_345
timestamp 1698431365
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_346
timestamp 1698431365
transform 1 0 20272 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_347
timestamp 1698431365
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_348
timestamp 1698431365
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_349
timestamp 1698431365
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_350
timestamp 1698431365
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_351
timestamp 1698431365
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_352
timestamp 1698431365
transform 1 0 22232 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_353
timestamp 1698431365
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_354
timestamp 1698431365
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_355
timestamp 1698431365
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_356
timestamp 1698431365
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_357
timestamp 1698431365
transform 1 0 20272 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_358
timestamp 1698431365
transform 1 0 2632 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_359
timestamp 1698431365
transform 1 0 6552 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_360
timestamp 1698431365
transform 1 0 10472 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_361
timestamp 1698431365
transform 1 0 14392 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_362
timestamp 1698431365
transform 1 0 18312 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_363
timestamp 1698431365
transform 1 0 22232 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_364
timestamp 1698431365
transform 1 0 4592 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_365
timestamp 1698431365
transform 1 0 8512 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_366
timestamp 1698431365
transform 1 0 12432 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_367
timestamp 1698431365
transform 1 0 16352 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_368
timestamp 1698431365
transform 1 0 20272 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_369
timestamp 1698431365
transform 1 0 2632 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_370
timestamp 1698431365
transform 1 0 6552 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_371
timestamp 1698431365
transform 1 0 10472 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_372
timestamp 1698431365
transform 1 0 14392 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_373
timestamp 1698431365
transform 1 0 18312 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_374
timestamp 1698431365
transform 1 0 22232 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_375
timestamp 1698431365
transform 1 0 4592 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_376
timestamp 1698431365
transform 1 0 8512 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_377
timestamp 1698431365
transform 1 0 12432 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_378
timestamp 1698431365
transform 1 0 16352 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_379
timestamp 1698431365
transform 1 0 20272 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_380
timestamp 1698431365
transform 1 0 2632 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_381
timestamp 1698431365
transform 1 0 6552 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_382
timestamp 1698431365
transform 1 0 10472 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_383
timestamp 1698431365
transform 1 0 14392 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_384
timestamp 1698431365
transform 1 0 18312 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_385
timestamp 1698431365
transform 1 0 22232 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_386
timestamp 1698431365
transform 1 0 4592 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_387
timestamp 1698431365
transform 1 0 8512 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_388
timestamp 1698431365
transform 1 0 12432 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_389
timestamp 1698431365
transform 1 0 16352 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_390
timestamp 1698431365
transform 1 0 20272 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_391
timestamp 1698431365
transform 1 0 2632 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_392
timestamp 1698431365
transform 1 0 6552 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_393
timestamp 1698431365
transform 1 0 10472 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_394
timestamp 1698431365
transform 1 0 14392 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_395
timestamp 1698431365
transform 1 0 18312 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_396
timestamp 1698431365
transform 1 0 22232 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_397
timestamp 1698431365
transform 1 0 4592 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_398
timestamp 1698431365
transform 1 0 8512 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_399
timestamp 1698431365
transform 1 0 12432 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_400
timestamp 1698431365
transform 1 0 16352 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_401
timestamp 1698431365
transform 1 0 20272 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_402
timestamp 1698431365
transform 1 0 2632 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_403
timestamp 1698431365
transform 1 0 6552 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_404
timestamp 1698431365
transform 1 0 10472 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_405
timestamp 1698431365
transform 1 0 14392 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_406
timestamp 1698431365
transform 1 0 18312 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_407
timestamp 1698431365
transform 1 0 22232 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_408
timestamp 1698431365
transform 1 0 4592 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_409
timestamp 1698431365
transform 1 0 8512 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_410
timestamp 1698431365
transform 1 0 12432 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_411
timestamp 1698431365
transform 1 0 16352 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_412
timestamp 1698431365
transform 1 0 20272 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_413
timestamp 1698431365
transform 1 0 2576 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_414
timestamp 1698431365
transform 1 0 4480 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_415
timestamp 1698431365
transform 1 0 6384 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_416
timestamp 1698431365
transform 1 0 8288 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_417
timestamp 1698431365
transform 1 0 10192 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_418
timestamp 1698431365
transform 1 0 12096 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_419
timestamp 1698431365
transform 1 0 14000 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_420
timestamp 1698431365
transform 1 0 15904 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_421
timestamp 1698431365
transform 1 0 17808 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_422
timestamp 1698431365
transform 1 0 19712 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_423
timestamp 1698431365
transform 1 0 21616 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_424
timestamp 1698431365
transform 1 0 23520 0 1 22736
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 ctrl_in[0]
port 0 nsew signal input
flabel metal3 s 24600 11760 25000 11816 0 FreeSans 224 0 0 0 ctrl_in[1]
port 1 nsew signal input
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 ctrl_oeb[0]
port 2 nsew signal tristate
flabel metal3 s 24600 12768 25000 12824 0 FreeSans 224 0 0 0 ctrl_oeb[1]
port 3 nsew signal tristate
flabel metal2 s 12768 0 12824 400 0 FreeSans 224 90 0 0 ctrl_out[0]
port 4 nsew signal tristate
flabel metal2 s 12096 0 12152 400 0 FreeSans 224 90 0 0 ctrl_out[1]
port 5 nsew signal tristate
flabel metal3 s 24600 12096 25000 12152 0 FreeSans 224 0 0 0 reset
port 6 nsew signal tristate
flabel metal3 s 24600 12432 25000 12488 0 FreeSans 224 0 0 0 resetn
port 7 nsew signal tristate
flabel metal4 s 2224 1538 2384 23158 0 FreeSans 640 90 0 0 vdd
port 8 nsew power bidirectional
flabel metal4 s 17584 1538 17744 23158 0 FreeSans 640 90 0 0 vdd
port 8 nsew power bidirectional
flabel metal4 s 9904 1538 10064 23158 0 FreeSans 640 90 0 0 vss
port 9 nsew ground bidirectional
rlabel metal1 12488 23128 12488 23128 0 vdd
rlabel metal1 12488 22736 12488 22736 0 vss
rlabel metal2 13412 12180 13412 12180 0 clknet_0_ctrl_in[0]
rlabel metal2 11452 10752 11452 10752 0 clknet_1_0__leaf_ctrl_in[0]
rlabel metal2 14364 12572 14364 12572 0 clknet_1_1__leaf_ctrl_in[0]
rlabel metal2 11564 12236 11564 12236 0 ctrl_in[0]
rlabel metal2 24108 11816 24108 11816 0 ctrl_in[1]
rlabel metal2 13020 12712 13020 12712 0 net1
rlabel metal2 13524 12460 13524 12460 0 net2
rlabel metal2 22624 12628 22624 12628 0 net3
rlabel metal2 12796 1015 12796 1015 0 net4
rlabel metal2 12124 1015 12124 1015 0 net5
rlabel metal2 11788 11004 11788 11004 0 net6
rlabel metal2 24108 12908 24108 12908 0 net7
rlabel metal2 12460 1099 12460 1099 0 net8
rlabel metal2 11844 12936 11844 12936 0 net9
rlabel metal2 23996 12180 23996 12180 0 reset
rlabel metal2 23996 12628 23996 12628 0 resetn
rlabel metal2 13356 10724 13356 10724 0 rst_sync_0.sync_reg\[0\]
rlabel metal2 12628 12600 12628 12600 0 rst_sync_0.sync_reg\[1\]
rlabel metal2 10780 12880 10780 12880 0 rst_sync_0.sync_reg\[2\]
rlabel metal2 12348 12600 12348 12600 0 rst_sync_0.sync_reg\[3\]
<< properties >>
string FIXED_BBOX 0 0 25000 25000
<< end >>

* NGSPICE file created from pcpi_mul.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

.subckt pcpi_mul clk pcpi_insn[0] pcpi_insn[10] pcpi_insn[11] pcpi_insn[12] pcpi_insn[13]
+ pcpi_insn[14] pcpi_insn[15] pcpi_insn[16] pcpi_insn[17] pcpi_insn[18] pcpi_insn[19]
+ pcpi_insn[1] pcpi_insn[20] pcpi_insn[21] pcpi_insn[22] pcpi_insn[23] pcpi_insn[24]
+ pcpi_insn[25] pcpi_insn[26] pcpi_insn[27] pcpi_insn[28] pcpi_insn[29] pcpi_insn[2]
+ pcpi_insn[30] pcpi_insn[31] pcpi_insn[3] pcpi_insn[4] pcpi_insn[5] pcpi_insn[6]
+ pcpi_insn[7] pcpi_insn[8] pcpi_insn[9] pcpi_mul_rd[0] pcpi_mul_rd[10] pcpi_mul_rd[11]
+ pcpi_mul_rd[12] pcpi_mul_rd[13] pcpi_mul_rd[14] pcpi_mul_rd[15] pcpi_mul_rd[16]
+ pcpi_mul_rd[17] pcpi_mul_rd[18] pcpi_mul_rd[19] pcpi_mul_rd[1] pcpi_mul_rd[20] pcpi_mul_rd[21]
+ pcpi_mul_rd[22] pcpi_mul_rd[23] pcpi_mul_rd[24] pcpi_mul_rd[25] pcpi_mul_rd[26]
+ pcpi_mul_rd[27] pcpi_mul_rd[28] pcpi_mul_rd[29] pcpi_mul_rd[2] pcpi_mul_rd[30] pcpi_mul_rd[31]
+ pcpi_mul_rd[3] pcpi_mul_rd[4] pcpi_mul_rd[5] pcpi_mul_rd[6] pcpi_mul_rd[7] pcpi_mul_rd[8]
+ pcpi_mul_rd[9] pcpi_mul_ready pcpi_mul_valid pcpi_mul_wait pcpi_mul_wr pcpi_rs1[0]
+ pcpi_rs1[10] pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14] pcpi_rs1[15] pcpi_rs1[16]
+ pcpi_rs1[17] pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20] pcpi_rs1[21] pcpi_rs1[22]
+ pcpi_rs1[23] pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27] pcpi_rs1[28] pcpi_rs1[29]
+ pcpi_rs1[2] pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4] pcpi_rs1[5] pcpi_rs1[6]
+ pcpi_rs1[7] pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10] pcpi_rs2[11] pcpi_rs2[12]
+ pcpi_rs2[13] pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17] pcpi_rs2[18] pcpi_rs2[19]
+ pcpi_rs2[1] pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23] pcpi_rs2[24] pcpi_rs2[25]
+ pcpi_rs2[26] pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2] pcpi_rs2[30] pcpi_rs2[31]
+ pcpi_rs2[3] pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7] pcpi_rs2[8] pcpi_rs2[9]
+ resetn vdd vss
X_2106_ picorv32_pcpi_mul_inst_0.rd\[28\] picorv32_pcpi_mul_inst_0.rdx\[28\] _0485_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3086_ _0203_ clknet_leaf_11_clk picorv32_pcpi_mul_inst_0.next_rs1\[45\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2037_ picorv32_pcpi_mul_inst_0.rd\[21\] picorv32_pcpi_mul_inst_0.next_rs2\[22\]
+ _1427_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_37_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1454__A1 _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2246__A3 _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2174__B picorv32_pcpi_mul_inst_0.rd\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2939_ _0056_ clknet_leaf_26_clk picorv32_pcpi_mul_inst_0.next_rs2\[46\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input73_I pcpi_rs2[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2237__A3 _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1479__I _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2103__I _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1942__I _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2773__I net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1987__A2 _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3005__CLK clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2724_ net95 _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2655_ _0935_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1606_ _1211_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2586_ _0532_ picorv32_pcpi_mul_inst_0.next_rs1\[29\] picorv32_pcpi_mul_inst_0.next_rs1\[30\]
+ _0880_ _1158_ net42 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XANTENNA__2164__A2 _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1537_ _1190_ picorv32_pcpi_mul_inst_0.next_rs2\[8\] _1186_ picorv32_pcpi_mul_inst_0.next_rs2\[7\]
+ _1184_ net80 _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1468_ _1133_ _1135_ _1136_ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3069_ _0186_ clknet_leaf_3_clk picorv32_pcpi_mul_inst_0.next_rs1\[28\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1978__A2 picorv32_pcpi_mul_inst_0.rd\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2440_ _0779_ _0782_ _0780_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2371_ _0720_ _0724_ _1146_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_90_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2707_ _0888_ picorv32_pcpi_mul_inst_0.next_rs1\[61\] _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2638_ _0914_ picorv32_pcpi_mul_inst_0.next_rs1\[43\] _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2569_ _0868_ picorv32_pcpi_mul_inst_0.next_rs1\[22\] picorv32_pcpi_mul_inst_0.next_rs1\[23\]
+ _0873_ _0870_ net34 _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XANTENNA_input36_I pcpi_rs1[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2128__A2 _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2588__I _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2300__A2 _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1940_ _0306_ picorv32_pcpi_mul_inst_0.rd\[11\] _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1871_ picorv32_pcpi_mul_inst_0.rd\[5\] _0273_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_28_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2423_ _0770_ _1376_ _1437_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_50_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2354_ _0706_ _0708_ _0709_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2285_ _0637_ _0647_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_67_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1577__I _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_22_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_37_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2349__A2 _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2070_ picorv32_pcpi_mul_inst_0.next_rs2\[26\] _1410_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2781__I _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2972_ _0089_ clknet_leaf_40_clk picorv32_pcpi_mul_inst_0.rd\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1923_ picorv32_pcpi_mul_inst_0.next_rs2\[11\] _0320_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1854_ _0255_ _0257_ _0258_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_12_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1785_ _1249_ _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2406_ picorv32_pcpi_mul_inst_0.next_rs2\[59\] _1436_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2337_ _0686_ _0690_ _0687_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2268_ _0628_ _0630_ _0631_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2199_ _1260_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2503__A2 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2866__I net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1570_ _1213_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2122_ _0496_ _0498_ _0475_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2053_ _0433_ _0436_ _0429_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ _0072_ clknet_leaf_18_clk picorv32_pcpi_mul_inst_0.next_rs2\[62\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1906_ _0305_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2430__A1 _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2886_ _0005_ clknet_leaf_8_clk picorv32_pcpi_mul_inst_0.instr_mulh vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1837_ picorv32_pcpi_mul_inst_0.next_rs2\[3\] _1426_ _1430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1768_ _1370_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1699_ _1314_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output105_I net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput86 net86 pcpi_mul_rd[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput97 net97 pcpi_mul_rd[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2596__I _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2740_ _0982_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2671_ _0939_ picorv32_pcpi_mul_inst_0.next_rs1\[51\] _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1622_ picorv32_pcpi_mul_inst_0.instr_mulh _1244_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1553_ _1198_ _1200_ _1195_ picorv32_pcpi_mul_inst_0.next_rs2\[12\] _1201_ net54
+ _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_1_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1484_ _1141_ _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2191__A3 _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2105_ _0480_ _0482_ _0484_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3085_ _0202_ clknet_leaf_12_clk picorv32_pcpi_mul_inst_0.next_rs1\[44\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2036_ _0420_ _0421_ _0422_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_37_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2938_ _0055_ clknet_leaf_22_clk picorv32_pcpi_mul_inst_0.next_rs2\[45\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2403__A1 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2869_ _1102_ _1098_ _1103_ _1104_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input66_I pcpi_rs2[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2173__A3 _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_48_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2723_ _0977_ _0980_ _0984_ _0987_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2654_ _1393_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1605_ _1237_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2585_ _0883_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1536_ _1189_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1467_ _1124_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_66_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_93_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3068_ _0185_ clknet_leaf_3_clk picorv32_pcpi_mul_inst_0.next_rs1\[27\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2019_ picorv32_pcpi_mul_inst_0.rd\[20\] _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2394__A3 _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2370_ _0721_ _0723_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2024__I _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2706_ picorv32_pcpi_mul_inst_0.next_rs1\[60\] _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2385__A3 _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2637_ _1394_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2568_ _0858_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1519_ _1171_ picorv32_pcpi_mul_inst_0.next_rs2\[3\] _1175_ _1172_ _1176_ net73 _1178_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2499_ net117 _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input29_I pcpi_rs1[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2376__A3 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1584__A1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1887__A2 picorv32_pcpi_mul_inst_0.rd\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1948__I _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1870_ picorv32_pcpi_mul_inst_0.next_rs2\[6\] _0272_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2367__A3 _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2779__I net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1683__I _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2422_ picorv32_pcpi_mul_inst_0.rd\[60\] _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2353_ _0674_ _0703_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2284_ _0639_ _0644_ _0646_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1999_ _0378_ picorv32_pcpi_mul_inst_0.rd\[17\] _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2506__C2 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2809__A1 picorv32_pcpi_mul_inst_0.rd\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2971_ _0088_ clknet_leaf_43_clk picorv32_pcpi_mul_inst_0.rd\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2283__B _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1922_ _1423_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1853_ _1399_ picorv32_pcpi_mul_inst_0.rd\[3\] _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1796__A1 _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1784_ _1383_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2405_ picorv32_pcpi_mul_inst_0.rd\[58\] picorv32_pcpi_mul_inst_0.next_rs2\[59\]
+ _0651_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_4_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2336_ _0693_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_49_clk clknet_2_0__leaf_clk clknet_leaf_49_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2267_ picorv32_pcpi_mul_inst_0.next_rs2\[45\] _0592_ picorv32_pcpi_mul_inst_0.rd\[44\]
+ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_67_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2198_ _0561_ _0568_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2028__A2 _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_11_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_86_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2267__A2 _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_20_Left_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2121_ _0496_ _0498_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_21_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2052_ _0433_ _0436_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2258__A2 _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_36_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2954_ _0071_ clknet_leaf_19_clk picorv32_pcpi_mul_inst_0.next_rs2\[61\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1905_ _1160_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2885_ net117 clknet_leaf_8_clk picorv32_pcpi_mul_inst_0.pcpi_wait_q vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1836_ _1412_ _1425_ _1428_ _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1767_ _1358_ picorv32_pcpi_mul_inst_0.next_rs2\[59\] _1369_ _1370_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1698_ _1306_ picorv32_pcpi_mul_inst_0.next_rs2\[46\] _1313_ _1314_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2319_ _0666_ _0669_ _0677_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input11_I pcpi_insn[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1932__A1 picorv32_pcpi_mul_inst_0.rd\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput87 net87 pcpi_mul_rd[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput98 net98 pcpi_mul_rd[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_53_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2670_ _0935_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_81_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1621_ _1249_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_34_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1552_ _1183_ _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1483_ net4 net3 _1149_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1691__I _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I pcpi_insn[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2104_ _0483_ _0478_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3084_ _0201_ clknet_leaf_13_clk picorv32_pcpi_mul_inst_0.next_rs1\[43\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2035_ _0412_ picorv32_pcpi_mul_inst_0.rd\[21\] _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1454__A3 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2937_ _0054_ clknet_leaf_22_clk picorv32_pcpi_mul_inst_0.next_rs2\[44\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2868_ picorv32_pcpi_mul_inst_0.rd\[61\] _1095_ _0979_ _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1819_ _1407_ _1413_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2799_ _1045_ _1033_ _1046_ _1048_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1914__A1 picorv32_pcpi_mul_inst_0.rd\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input59_I pcpi_rs2[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2722_ _0511_ _1115_ _0986_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2653_ picorv32_pcpi_mul_inst_0.next_rs1\[46\] _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1604_ _1233_ _1235_ _1230_ picorv32_pcpi_mul_inst_0.next_rs2\[28\] _1236_ net71
+ _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2584_ _0532_ picorv32_pcpi_mul_inst_0.next_rs1\[28\] picorv32_pcpi_mul_inst_0.next_rs1\[29\]
+ _0880_ _1158_ net40 _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1535_ _1167_ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1466_ picorv32_pcpi_mul_inst_0.mul_counter\[3\] picorv32_pcpi_mul_inst_0.mul_counter\[4\]
+ picorv32_pcpi_mul_inst_0.mul_counter\[5\] _1134_ _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3136_ net116 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3067_ _0184_ clknet_leaf_3_clk picorv32_pcpi_mul_inst_0.next_rs1\[26\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2018_ _0404_ _0405_ _0406_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2312__A1 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2705_ _0967_ _0971_ _0969_ _0972_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2636_ picorv32_pcpi_mul_inst_0.next_rs1\[42\] _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2567_ _0872_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3136__I net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1518_ _1177_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2498_ _0822_ _0769_ _0826_ _0827_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1449_ net4 _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2196__B _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3119_ _0236_ clknet_leaf_35_clk net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_85_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2421_ picorv32_pcpi_mul_inst_0.rdx\[60\] _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2352_ _0595_ _0707_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2283_ _0639_ _0644_ _0645_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1998_ _0384_ _0386_ _0388_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2763__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2619_ _0898_ _0907_ _0900_ _0908_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_7_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input41_I pcpi_rs1[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2506__B2 _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2970_ _0087_ clknet_leaf_42_clk picorv32_pcpi_mul_inst_0.rd\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2037__A3 _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1921_ _0311_ _0313_ _0318_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1852_ _1147_ _0256_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1783_ _1375_ picorv32_pcpi_mul_inst_0.next_rs2\[62\] _1382_ _1383_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2404_ _0746_ _0749_ _0747_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_4_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2335_ _0685_ _0692_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2266_ _0629_ _1307_ _0590_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2197_ _0563_ _0566_ _0567_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1869__I _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2120_ picorv32_pcpi_mul_inst_0.rd\[30\] _0497_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2051_ _0434_ _0435_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2294__B _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1689__I _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2953_ _0070_ clknet_leaf_20_clk picorv32_pcpi_mul_inst_0.next_rs2\[60\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1904_ _0302_ _0303_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2884_ _0004_ clknet_leaf_6_clk picorv32_pcpi_mul_inst_0.mul_finish vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1835_ _1415_ picorv32_pcpi_mul_inst_0.next_rs2\[2\] _1427_ _1428_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1766_ _1367_ _1360_ _1368_ _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_40_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2194__A2 _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1697_ _1296_ _1308_ _1312_ _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2318_ _0667_ _1324_ _0601_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2249_ _0612_ _0614_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1599__I _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput88 net88 pcpi_mul_rd[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput99 net99 pcpi_mul_rd[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_74_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1999__A2 picorv32_pcpi_mul_inst_0.rd\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1620_ _1166_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1923__A2 _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1551_ picorv32_pcpi_mul_inst_0.next_rs2\[13\] _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1482_ net2 _1130_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2103_ _0446_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3083_ _0200_ clknet_leaf_13_clk picorv32_pcpi_mul_inst_0.next_rs1\[42\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2034_ _0417_ _0419_ _0388_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2100__A2 _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2936_ _0053_ clknet_leaf_22_clk picorv32_pcpi_mul_inst_0.next_rs2\[43\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2867_ picorv32_pcpi_mul_inst_0.rd\[29\] _1099_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2043__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1818_ _1152_ picorv32_pcpi_mul_inst_0.rd\[0\] _1409_ _1412_ _1413_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2798_ picorv32_pcpi_mul_inst_0.rd\[47\] _1047_ _1037_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1749_ _1354_ picorv32_pcpi_mul_inst_0.next_rs2\[55\] _1355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output110_I net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_20_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_35_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2330__A2 _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1841__A1 _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2721_ _0985_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2652_ _0932_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1603_ _1218_ _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2583_ _0882_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1534_ _1188_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1465_ picorv32_pcpi_mul_inst_0.mul_counter\[0\] picorv32_pcpi_mul_inst_0.mul_counter\[2\]
+ picorv32_pcpi_mul_inst_0.mul_counter\[1\] _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_3135_ _0252_ clknet_leaf_3_clk picorv32_pcpi_mul_inst_0.mul_counter\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3066_ _0183_ clknet_leaf_2_clk picorv32_pcpi_mul_inst_0.next_rs1\[25\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_93_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2017_ _0378_ picorv32_pcpi_mul_inst_0.rd\[19\] _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2919_ _0036_ clknet_leaf_43_clk picorv32_pcpi_mul_inst_0.next_rs2\[26\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input71_I pcpi_rs2[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1826__B _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2704_ _0888_ picorv32_pcpi_mul_inst_0.next_rs1\[60\] _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2635_ _0885_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2566_ _0868_ picorv32_pcpi_mul_inst_0.next_rs1\[21\] picorv32_pcpi_mul_inst_0.next_rs1\[22\]
+ _0866_ _0870_ net33 _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1517_ _1171_ _1172_ _1175_ picorv32_pcpi_mul_inst_0.next_rs2\[1\] _1176_ net62 _1177_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2497_ _0762_ _0765_ _0763_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1448_ _1119_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3118_ _0235_ clknet_leaf_35_clk net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3049_ _0166_ clknet_leaf_0_clk picorv32_pcpi_mul_inst_0.next_rs1\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1569__B1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_2__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2420_ _0766_ _0767_ _0768_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2351_ _0704_ _0705_ _0702_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2282_ _1140_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2460__A1 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1997_ _0286_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2618_ _0903_ picorv32_pcpi_mul_inst_0.next_rs1\[38\] _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2549_ _0845_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_7_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input34_I pcpi_rs1[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2203__A1 picorv32_pcpi_mul_inst_0.rd\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1920_ _0317_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1851_ _1438_ _1433_ _0254_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1782_ _1367_ _1377_ _1381_ _1382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_12_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2403_ _1250_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2334_ _0686_ _0690_ _0691_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2265_ picorv32_pcpi_mul_inst_0.rd\[44\] _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2196_ _0563_ _0566_ _1419_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1885__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2050_ picorv32_pcpi_mul_inst_0.next_rs2\[24\] _0331_ picorv32_pcpi_mul_inst_0.rd\[23\]
+ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2952_ _0069_ clknet_leaf_20_clk picorv32_pcpi_mul_inst_0.next_rs2\[59\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1903_ _1192_ _0263_ _0300_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_32_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2883_ _0003_ clknet_leaf_5_clk picorv32_pcpi_mul_inst_0.mul_counter\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1834_ _1426_ _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1765_ _1354_ picorv32_pcpi_mul_inst_0.next_rs2\[58\] _1368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1696_ _1301_ _1307_ _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2317_ _0636_ picorv32_pcpi_mul_inst_0.rd\[49\] _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2248_ _0609_ _0613_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2179_ _0519_ picorv32_pcpi_mul_inst_0.rd\[35\] _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1932__A3 _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput89 net89 pcpi_mul_rd[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_74_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_9_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1550_ _1199_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1481_ _1148_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2102_ _0443_ _0481_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3082_ _0199_ clknet_leaf_13_clk picorv32_pcpi_mul_inst_0.next_rs1\[41\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2033_ _0417_ _0419_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2935_ _0052_ clknet_leaf_15_clk picorv32_pcpi_mul_inst_0.next_rs2\[42\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2866_ net105 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1817_ picorv32_pcpi_mul_inst_0.rd\[0\] picorv32_pcpi_mul_inst_0.next_rs2\[1\] _1411_
+ _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2797_ _1029_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1748_ _1300_ _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1679_ _1296_ _1289_ _1297_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_88_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_17_Left_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2720_ _1118_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2651_ _1151_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1983__I _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1602_ picorv32_pcpi_mul_inst_0.next_rs2\[29\] _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2582_ _0532_ picorv32_pcpi_mul_inst_0.next_rs1\[27\] picorv32_pcpi_mul_inst_0.next_rs1\[28\]
+ _0880_ _0877_ net39 _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1533_ _1179_ picorv32_pcpi_mul_inst_0.next_rs2\[7\] _1186_ picorv32_pcpi_mul_inst_0.next_rs2\[6\]
+ _1184_ net79 _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XPHY_EDGE_ROW_26_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1464_ _1132_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3134_ _0251_ clknet_leaf_32_clk net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3065_ _0182_ clknet_leaf_2_clk picorv32_pcpi_mul_inst_0.next_rs1\[24\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_93_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2016_ _0400_ _0403_ _0388_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1832__A2 _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2918_ _0035_ clknet_leaf_37_clk picorv32_pcpi_mul_inst_0.next_rs2\[25\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_30_clk clknet_2_3__leaf_clk clknet_leaf_30_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2849_ picorv32_pcpi_mul_inst_0.rd\[57\] _1079_ _1085_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input64_I pcpi_rs2[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1823__A2 _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_clk clknet_2_3__leaf_clk clknet_leaf_21_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2067__A2 _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_12_clk clknet_2_2__leaf_clk clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2703_ picorv32_pcpi_mul_inst_0.next_rs1\[59\] _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2634_ _0909_ _0918_ _0911_ _0919_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2565_ _0871_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1516_ _1158_ _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2496_ _1140_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1447_ _1118_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3117_ _0234_ clknet_leaf_35_clk net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3048_ _0165_ clknet_leaf_1_clk picorv32_pcpi_mul_inst_0.next_rs1\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2058__A2 _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_34_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_49_clk_I clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2350_ _0702_ _0704_ _0705_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2281_ _0641_ _0643_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1799__A1 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1996_ _0384_ _0386_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1971__A1 picorv32_pcpi_mul_inst_0.rd\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2617_ picorv32_pcpi_mul_inst_0.next_rs1\[37\] _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2548_ _0860_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_58_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2479_ _1384_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input27_I pcpi_rs1[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output95_I net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1850_ _1438_ _1433_ _0254_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1781_ _1371_ _1376_ _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1953__A1 _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2402_ picorv32_pcpi_mul_inst_0.rd\[58\] _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2333_ _0686_ _0690_ _1146_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2264_ picorv32_pcpi_mul_inst_0.rdx\[44\] _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2195_ _0564_ _0565_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_9_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_63_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1979_ _0369_ _0370_ _0371_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2062__I _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1944__A1 _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1986__I _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2415__A2 _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2951_ _0068_ clknet_leaf_20_clk picorv32_pcpi_mul_inst_0.next_rs2\[58\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1902_ _1408_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2882_ _0002_ clknet_leaf_8_clk picorv32_pcpi_mul_inst_0.instr_mul vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1833_ _1422_ _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1764_ _1249_ _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1935__B picorv32_pcpi_mul_inst_0.rd\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1695_ _1311_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2316_ _0670_ _0672_ _0675_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2247_ picorv32_pcpi_mul_inst_0.next_rs2\[43\] _0574_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2178_ _0545_ _0548_ _0550_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_82_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1480_ picorv32_pcpi_mul_inst_0.mul_counter\[6\] _1147_ _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2101_ _1235_ _0375_ _0479_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3081_ _0198_ clknet_leaf_13_clk picorv32_pcpi_mul_inst_0.next_rs1\[40\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2032_ picorv32_pcpi_mul_inst_0.rd\[21\] _0418_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2934_ _0051_ clknet_leaf_21_clk picorv32_pcpi_mul_inst_0.next_rs2\[41\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2865_ _1097_ _1098_ _1100_ _1101_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1816_ _1410_ _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2796_ picorv32_pcpi_mul_inst_0.rd\[15\] _1035_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1747_ _1353_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1678_ _1283_ picorv32_pcpi_mul_inst_0.next_rs2\[42\] _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2315__A1 _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2650_ _0920_ _0930_ _0922_ _0931_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1601_ _1234_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2581_ _0881_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1532_ _1187_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1463_ picorv32_pcpi_mul_inst_0.mul_waiting _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I pcpi_insn[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3133_ _0250_ clknet_leaf_19_clk net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1504__I net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3064_ _0181_ clknet_leaf_2_clk picorv32_pcpi_mul_inst_0.next_rs1\[23\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2015_ _0400_ _0403_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2085__A3 _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2917_ _0034_ clknet_leaf_37_clk picorv32_pcpi_mul_inst_0.next_rs2\[24\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2793__A1 picorv32_pcpi_mul_inst_0.rd\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2848_ picorv32_pcpi_mul_inst_0.rd\[25\] _1083_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2779_ net87 _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input57_I pcpi_rs2[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_8_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2076__A3 _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2481__B1 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2702_ _0967_ _0968_ _0969_ _0970_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2633_ _0914_ picorv32_pcpi_mul_inst_0.next_rs1\[42\] _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2564_ _0868_ picorv32_pcpi_mul_inst_0.next_rs1\[20\] picorv32_pcpi_mul_inst_0.next_rs1\[21\]
+ _0866_ _0870_ net32 _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1515_ _1174_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2495_ _0822_ _0735_ _0820_ _0825_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1446_ _1117_ picorv32_pcpi_mul_inst_0.mul_finish _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3116_ _0233_ clknet_leaf_34_clk net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3047_ _0164_ clknet_leaf_46_clk picorv32_pcpi_mul_inst_0.next_rs1\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2766__A1 picorv32_pcpi_mul_inst_0.rd\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_45_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_69_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2049__A3 _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2280_ picorv32_pcpi_mul_inst_0.next_rs2\[46\] _0642_ picorv32_pcpi_mul_inst_0.rd\[45\]
+ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_72_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1995_ picorv32_pcpi_mul_inst_0.rd\[17\] _0385_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_27_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2616_ _0898_ _0905_ _0900_ _0906_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2547_ _0853_ picorv32_pcpi_mul_inst_0.next_rs1\[14\] picorv32_pcpi_mul_inst_0.next_rs1\[15\]
+ _0859_ _0855_ net25 _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XPHY_EDGE_ROW_81_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2478_ _0813_ _0814_ _0815_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_58_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_90_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2203__A3 _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1780_ _1380_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2401_ _0744_ _0751_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2332_ _0687_ _0689_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_33_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2263_ _0625_ _0626_ _0627_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2194_ picorv32_pcpi_mul_inst_0.next_rs2\[38\] _0527_ picorv32_pcpi_mul_inst_0.rd\[37\]
+ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_48_clk_I clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2433__A3 _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1978_ _0344_ picorv32_pcpi_mul_inst_0.rd\[15\] _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2188__A2 _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1935__A2 _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1871__A1 picorv32_pcpi_mul_inst_0.rd\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2950_ _0067_ clknet_leaf_20_clk picorv32_pcpi_mul_inst_0.next_rs2\[57\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1901_ _1192_ _1406_ _0300_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2881_ _0001_ clknet_leaf_8_clk picorv32_pcpi_mul_inst_0.instr_mulhsu vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1832_ _1172_ _1424_ picorv32_pcpi_mul_inst_0.rd\[1\] _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2179__A2 picorv32_pcpi_mul_inst_0.rd\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1763_ _1366_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1694_ _1306_ _1307_ _1310_ _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2315_ _0674_ _0667_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2246_ picorv32_pcpi_mul_inst_0.rd\[42\] picorv32_pcpi_mul_inst_0.next_rs2\[43\]
+ _0536_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2177_ _0474_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_23_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1917__A2 picorv32_pcpi_mul_inst_0.rd\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2801__I _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1853__A1 _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2100_ _1235_ _0263_ _0479_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3080_ _0197_ clknet_leaf_13_clk picorv32_pcpi_mul_inst_0.next_rs1\[39\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2031_ picorv32_pcpi_mul_inst_0.next_rs2\[22\] _1410_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2158__I _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1997__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2933_ _0050_ clknet_leaf_15_clk picorv32_pcpi_mul_inst_0.next_rs2\[40\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2864_ _0770_ _1095_ _0979_ _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1815_ _1401_ _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2795_ net90 _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1746_ _1341_ picorv32_pcpi_mul_inst_0.next_rs2\[55\] _1352_ _1353_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1677_ _1278_ _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2229_ _0595_ _0596_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2012__A1 picorv32_pcpi_mul_inst_0.rd\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2315__A2 _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1600_ _1233_ picorv32_pcpi_mul_inst_0.next_rs2\[28\] _1230_ picorv32_pcpi_mul_inst_0.next_rs2\[27\]
+ _1228_ net70 _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_81_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2580_ _0875_ picorv32_pcpi_mul_inst_0.next_rs1\[26\] picorv32_pcpi_mul_inst_0.next_rs1\[27\]
+ _0880_ _0877_ net38 _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1531_ _1179_ picorv32_pcpi_mul_inst_0.next_rs2\[6\] _1186_ _1181_ _1184_ net78 _1187_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1462_ net4 net3 _1131_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_38_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3132_ _0249_ clknet_leaf_32_clk net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3063_ _0180_ clknet_leaf_2_clk picorv32_pcpi_mul_inst_0.next_rs1\[22\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_93_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2014_ _0401_ _0402_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2916_ _0033_ clknet_leaf_37_clk picorv32_pcpi_mul_inst_0.next_rs2\[23\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2847_ net101 _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2778_ _1027_ _1016_ _1028_ _1031_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1729_ _1333_ _1326_ _1338_ _1339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2300__B picorv32_pcpi_mul_inst_0.rd\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2481__B2 _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2233__A1 _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2701_ _0961_ picorv32_pcpi_mul_inst_0.next_rs1\[59\] _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2632_ picorv32_pcpi_mul_inst_0.next_rs1\[41\] _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2563_ _1182_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1514_ _1173_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2494_ _0728_ _0731_ _0729_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1515__I _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1445_ net83 _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3115_ _0232_ clknet_leaf_33_clk net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3046_ _0163_ clknet_leaf_49_clk picorv32_pcpi_mul_inst_0.next_rs1\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2463__A1 _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_52_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1994_ picorv32_pcpi_mul_inst_0.next_rs2\[18\] _0272_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_7_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1971__A3 _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2615_ _0903_ picorv32_pcpi_mul_inst_0.next_rs1\[37\] _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2546_ _0858_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2477_ _0807_ picorv32_pcpi_mul_inst_0.rdx\[28\] _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1487__A2 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3029_ _0146_ clknet_leaf_36_clk picorv32_pcpi_mul_inst_0.rdx\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2427__A1 _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _0746_ _0749_ _0750_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2331_ _0684_ _0688_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2262_ _0598_ picorv32_pcpi_mul_inst_0.rd\[43\] _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2193_ picorv32_pcpi_mul_inst_0.rd\[37\] picorv32_pcpi_mul_inst_0.next_rs2\[38\]
+ _0525_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_27_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1977_ _0365_ _0368_ _0335_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2529_ _0839_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input32_I pcpi_rs1[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2534__I _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1613__I _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1900_ _0299_ picorv32_pcpi_mul_inst_0.rdx\[8\] _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2880_ _1112_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1831_ _1423_ _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1762_ _1358_ picorv32_pcpi_mul_inst_0.next_rs2\[58\] _1365_ _1366_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1693_ _1296_ _1308_ _1309_ _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2314_ _0673_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2245_ _0603_ _0606_ _0604_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2176_ _0545_ _0548_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1614__A2 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_74_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_32_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_47_clk_I clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2030_ _0414_ _0415_ _0416_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2932_ _0049_ clknet_leaf_15_clk picorv32_pcpi_mul_inst_0.next_rs2\[39\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_42_clk clknet_2_1__leaf_clk clknet_leaf_42_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_72_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2863_ _0478_ _1099_ _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1814_ _1408_ _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2794_ _1042_ _1033_ _1043_ _1044_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2021__A2 _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1745_ _1350_ _1343_ _1351_ _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1676_ _1295_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2228_ _0591_ _0593_ _0588_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2159_ picorv32_pcpi_mul_inst_0.rd\[34\] _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_36_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_33_clk clknet_2_1__leaf_clk clknet_leaf_33_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2208__B _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1530_ _1174_ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1461_ _1121_ _1131_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3131_ _0248_ clknet_leaf_32_clk net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3062_ _0179_ clknet_leaf_1_clk picorv32_pcpi_mul_inst_0.next_rs1\[21\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_93_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2013_ picorv32_pcpi_mul_inst_0.next_rs2\[20\] _0331_ picorv32_pcpi_mul_inst_0.rd\[19\]
+ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_clk clknet_2_2__leaf_clk clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2915_ _0032_ clknet_leaf_37_clk picorv32_pcpi_mul_inst_0.next_rs2\[22\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2846_ _1081_ _1082_ _1084_ _1086_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2777_ picorv32_pcpi_mul_inst_0.rd\[43\] _1030_ _1019_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1728_ _1337_ picorv32_pcpi_mul_inst_0.next_rs2\[51\] _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1659_ _1269_ picorv32_pcpi_mul_inst_0.next_rs2\[39\] _1281_ _1282_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2233__A2 picorv32_pcpi_mul_inst_0.rd\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1992__A1 _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2717__I _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2700_ _0935_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2631_ _0909_ _0916_ _0911_ _0917_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2562_ _0869_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1513_ _1139_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2493_ _0822_ _0702_ _0820_ _0824_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xclkbuf_leaf_4_clk clknet_2_0__leaf_clk clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1444_ _1116_ picorv32_pcpi_mul_inst_0.instr_any_mul vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2160__A1 _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3114_ _0231_ clknet_leaf_33_clk net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3045_ _0162_ clknet_leaf_49_clk picorv32_pcpi_mul_inst_0.next_rs1\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2829_ picorv32_pcpi_mul_inst_0.rd\[53\] _1063_ _1069_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input62_I pcpi_rs2[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1441__I _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1965__A1 picorv32_pcpi_mul_inst_0.rd\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_9_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2142__A1 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1993_ _0380_ _0382_ _0383_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1956__A1 picorv32_pcpi_mul_inst_0.rd\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2614_ picorv32_pcpi_mul_inst_0.next_rs1\[36\] _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1526__I _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2545_ _1173_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2381__A1 _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2476_ _0467_ _0472_ _0469_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3028_ _0145_ clknet_leaf_37_clk picorv32_pcpi_mul_inst_0.rdx\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1947__A1 _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2330_ picorv32_pcpi_mul_inst_0.next_rs2\[51\] _0574_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2261_ _0619_ _0624_ _0550_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2192_ _0553_ _0556_ _0562_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2177__I _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1976_ _0365_ _0368_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1929__A1 picorv32_pcpi_mul_inst_0.rd\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2528_ _0847_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2459_ _0796_ picorv32_pcpi_mul_inst_0.rdx\[8\] _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input25_I pcpi_rs1[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2087__I _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ _1422_ _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2584__A1 _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1761_ _1350_ _1360_ _1364_ _1365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1692_ _1301_ picorv32_pcpi_mul_inst_0.next_rs2\[44\] _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2313_ _1144_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2244_ _0569_ _0609_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2175_ _0546_ _0547_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_69_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1959_ _0344_ picorv32_pcpi_mul_inst_0.rd\[13\] _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_78_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2327__A1 _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_87_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_74_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2318__A1 _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1624__I _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2931_ _0048_ clknet_leaf_15_clk picorv32_pcpi_mul_inst_0.next_rs2\[38\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2862_ _0981_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1813_ _1145_ _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2793_ picorv32_pcpi_mul_inst_0.rd\[46\] _1030_ _1037_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1744_ _1337_ picorv32_pcpi_mul_inst_0.next_rs2\[54\] _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1675_ _1287_ picorv32_pcpi_mul_inst_0.next_rs2\[42\] _1294_ _1295_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2227_ _1408_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2088__A3 _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1835__A3 _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2493__B1 _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2158_ _1260_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2089_ _0330_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2796__A1 picorv32_pcpi_mul_inst_0.rd\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2012__A3 _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1460_ _1122_ _1130_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3130_ _0247_ clknet_leaf_31_clk net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3061_ _0178_ clknet_leaf_1_clk picorv32_pcpi_mul_inst_0.next_rs1\[20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_93_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2012_ picorv32_pcpi_mul_inst_0.rd\[19\] picorv32_pcpi_mul_inst_0.next_rs2\[20\]
+ _0328_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1817__A3 _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2914_ _0031_ clknet_leaf_37_clk picorv32_pcpi_mul_inst_0.next_rs2\[21\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2845_ _0736_ _1079_ _1085_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2776_ _1029_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1727_ _1300_ _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1658_ _1279_ _1271_ _1280_ _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1589_ _1226_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_31_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_46_clk_I clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_47_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2630_ _0914_ picorv32_pcpi_mul_inst_0.next_rs1\[41\] _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2561_ _0868_ picorv32_pcpi_mul_inst_0.next_rs1\[19\] picorv32_pcpi_mul_inst_0.next_rs1\[20\]
+ _0866_ _0863_ net31 _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1512_ picorv32_pcpi_mul_inst_0.next_rs2\[2\] _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2492_ _0694_ _0697_ _0695_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1735__A2 picorv32_pcpi_mul_inst_0.next_rs2\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1443_ picorv32_pcpi_mul_inst_0.instr_mul _1115_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3113_ _0230_ clknet_leaf_33_clk net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3044_ _0161_ clknet_leaf_49_clk picorv32_pcpi_mul_inst_0.next_rs1\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1974__A2 _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2828_ picorv32_pcpi_mul_inst_0.rd\[21\] _1067_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2759_ _0999_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input55_I pcpi_rs2[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_44_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2728__I net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1992_ _0372_ picorv32_pcpi_mul_inst_0.rdx\[16\] _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1807__I _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2613_ _0898_ _0902_ _0900_ _0904_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2544_ _0857_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2475_ _1141_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_50_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3027_ _0144_ clknet_leaf_40_clk picorv32_pcpi_mul_inst_0.rdx\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1571__B1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2260_ _0619_ _0624_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2191_ _0554_ _1270_ _1411_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1626__A1 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1975_ _0366_ _0367_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2527_ _0846_ picorv32_pcpi_mul_inst_0.next_rs1\[7\] picorv32_pcpi_mul_inst_0.next_rs1\[8\]
+ _0843_ _0840_ net49 _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_11_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2458_ _0292_ _0295_ _0293_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2389_ _1409_ _0740_ _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input18_I pcpi_mul_valid vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2290__A1 picorv32_pcpi_mul_inst_0.rd\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output86_I net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1760_ _1354_ _1359_ _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1691_ _1252_ _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2312_ _0595_ _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2243_ picorv32_pcpi_mul_inst_0.rd\[42\] _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2174_ picorv32_pcpi_mul_inst_0.next_rs2\[36\] _0470_ picorv32_pcpi_mul_inst_0.rd\[35\]
+ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1820__I _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2651__I _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1958_ _0349_ _0351_ _0335_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1889_ _1436_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_74_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1905__I _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2930_ _0047_ clknet_leaf_14_clk picorv32_pcpi_mul_inst_0.next_rs2\[37\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2861_ _1119_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1812_ picorv32_pcpi_mul_inst_0.next_rs2\[1\] _1406_ picorv32_pcpi_mul_inst_0.rd\[0\]
+ _1407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2792_ picorv32_pcpi_mul_inst_0.rd\[14\] _1035_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1743_ _1249_ _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1674_ _1279_ _1289_ _1293_ _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2309__A2 _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1517__B1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1815__I _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2226_ _0588_ _0591_ _0593_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2157_ _0521_ _0531_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2493__A1 _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2088_ picorv32_pcpi_mul_inst_0.rd\[27\] picorv32_pcpi_mul_inst_0.next_rs2\[28\]
+ _0468_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_48_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_5_clk_I clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2240__B _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3060_ _0177_ clknet_leaf_1_clk picorv32_pcpi_mul_inst_0.next_rs1\[19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2011_ _0393_ _0395_ _0399_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2466__I _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2913_ _0030_ clknet_leaf_39_clk picorv32_pcpi_mul_inst_0.next_rs2\[20\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2844_ _0978_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2775_ _1113_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1726_ _1336_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1657_ _1265_ picorv32_pcpi_mul_inst_0.next_rs2\[38\] _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1588_ _1225_ picorv32_pcpi_mul_inst_0.next_rs2\[24\] _1221_ picorv32_pcpi_mul_inst_0.next_rs2\[23\]
+ _1219_ net66 _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2209_ _0572_ _0577_ _0578_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_68_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2457__A1 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2286__I picorv32_pcpi_mul_inst_0.rd\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_2_0__f_clk clknet_0_clk clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_55_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2560_ _0845_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1511_ _1136_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2491_ _0822_ _0666_ _0820_ _0823_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1442_ _1114_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3112_ _0229_ clknet_leaf_32_clk net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3043_ _0160_ clknet_leaf_49_clk picorv32_pcpi_mul_inst_0.next_rs1\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2827_ net97 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2758_ net114 _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1709_ _1322_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2689_ _0925_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input48_I pcpi_rs1[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2151__A3 _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1991_ picorv32_pcpi_mul_inst_0.next_rs2\[17\] _0381_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2612_ _0903_ picorv32_pcpi_mul_inst_0.next_rs1\[36\] _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2543_ _0853_ picorv32_pcpi_mul_inst_0.next_rs1\[13\] picorv32_pcpi_mul_inst_0.next_rs1\[14\]
+ _0851_ _0855_ net24 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XANTENNA_clkbuf_leaf_45_clk_I clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2474_ _0803_ _0811_ _0812_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3026_ _0143_ clknet_leaf_43_clk picorv32_pcpi_mul_inst_0.rdx\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2060__A2 _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2739__I _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2190_ _1414_ picorv32_pcpi_mul_inst_0.rd\[37\] _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1874__A2 picorv32_pcpi_mul_inst_0.rd\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1974_ picorv32_pcpi_mul_inst_0.next_rs2\[16\] _0331_ picorv32_pcpi_mul_inst_0.rd\[15\]
+ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1929__A3 _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2526_ _0845_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2457_ _1150_ _0799_ _0800_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2388_ _0737_ _0738_ _0735_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3009_ _0126_ clknet_leaf_27_clk picorv32_pcpi_mul_inst_0.rd\[49\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2333__B _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_85_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2805__A1 _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1690_ picorv32_pcpi_mul_inst_0.next_rs2\[45\] _1307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2311_ _0668_ _0669_ _0666_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2242_ _0600_ _0608_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2173_ picorv32_pcpi_mul_inst_0.rd\[35\] picorv32_pcpi_mul_inst_0.next_rs2\[36\]
+ _0468_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_25_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2418__B _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_45_clk clknet_2_0__leaf_clk clknet_leaf_45_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1957_ _0349_ _0351_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1888_ _0285_ _0288_ _0289_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2509_ _0834_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input30_I pcpi_rs1[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_36_clk clknet_2_1__leaf_clk clknet_leaf_36_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_82_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2318__A3 _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2238__B picorv32_pcpi_mul_inst_0.rd\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_27_clk clknet_2_3__leaf_clk clknet_leaf_27_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2860_ net104 _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1811_ _1405_ _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2791_ net89 _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1742_ _1349_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1673_ _1283_ _1288_ _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1517__A1 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2199__I _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2190__A1 _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2225_ picorv32_pcpi_mul_inst_0.next_rs2\[41\] _0592_ picorv32_pcpi_mul_inst_0.rd\[40\]
+ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2156_ _0523_ _0529_ _0530_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2087_ _0282_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_18_clk clknet_2_2__leaf_clk clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2989_ _0106_ clknet_leaf_44_clk picorv32_pcpi_mul_inst_0.rd\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input78_I pcpi_rs2[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1995__A1 picorv32_pcpi_mul_inst_0.rd\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ picorv32_pcpi_mul_inst_0.rd\[18\] picorv32_pcpi_mul_inst_0.next_rs2\[19\]
+ _0363_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_93_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2912_ _0029_ clknet_leaf_39_clk picorv32_pcpi_mul_inst_0.next_rs2\[19\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2843_ _0440_ _1083_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2774_ picorv32_pcpi_mul_inst_0.rd\[11\] _1017_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1725_ _1323_ picorv32_pcpi_mul_inst_0.next_rs2\[51\] _1335_ _1336_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_7_clk clknet_2_2__leaf_clk clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1656_ _1278_ _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1587_ _1224_ _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2208_ _0572_ _0577_ _0541_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2139_ picorv32_pcpi_mul_inst_0.next_rs2\[33\] _0514_ picorv32_pcpi_mul_inst_0.rd\[32\]
+ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2218__A2 picorv32_pcpi_mul_inst_0.rd\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2393__A1 _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1646__I _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1510_ _1121_ _1149_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2490_ _0659_ _0662_ _0660_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1441_ _1113_ _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3111_ _0228_ clknet_leaf_32_clk net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3042_ _0159_ clknet_leaf_49_clk picorv32_pcpi_mul_inst_0.next_rs1\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_4_clk_I clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2826_ _1065_ _1066_ _1068_ _1070_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2757_ _1011_ _1000_ _1012_ _1014_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1708_ _1306_ picorv32_pcpi_mul_inst_0.next_rs2\[48\] _1321_ _1322_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2688_ picorv32_pcpi_mul_inst_0.next_rs1\[55\] _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1639_ _1242_ _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_44_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1990_ _1423_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2611_ _1388_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2542_ _0856_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2473_ _0807_ picorv32_pcpi_mul_inst_0.rdx\[24\] _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3025_ _0142_ clknet_leaf_47_clk picorv32_pcpi_mul_inst_0.rdx\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1892__A3 _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2809_ picorv32_pcpi_mul_inst_0.rd\[49\] _1047_ _1053_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input60_I pcpi_rs2[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1973_ picorv32_pcpi_mul_inst_0.rd\[15\] picorv32_pcpi_mul_inst_0.next_rs2\[16\]
+ _0328_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_71_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2339__A1 picorv32_pcpi_mul_inst_0.next_rs2\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2525_ _1124_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1834__I _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2456_ _0796_ picorv32_pcpi_mul_inst_0.rdx\[4\] _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2387_ _0735_ _0737_ _0738_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3008_ _0125_ clknet_leaf_27_clk picorv32_pcpi_mul_inst_0.rd\[48\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2290__A3 _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2750__A1 picorv32_pcpi_mul_inst_0.rd\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_44_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2310_ _0666_ _0668_ _0669_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2241_ _0603_ _0606_ _0607_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2172_ _0535_ _0540_ _0537_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_38_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1956_ picorv32_pcpi_mul_inst_0.rd\[13\] _0350_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_28_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1887_ _0266_ picorv32_pcpi_mul_inst_0.rd\[6\] _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1564__I _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2508_ _0830_ picorv32_pcpi_mul_inst_0.next_rs1\[1\] picorv32_pcpi_mul_inst_0.next_rs1\[2\]
+ _0826_ _0832_ net41 _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2439_ _0777_ _0785_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input23_I pcpi_rs1[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_56_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1810_ _1404_ _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2790_ _1039_ _1033_ _1040_ _1041_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1741_ _1341_ picorv32_pcpi_mul_inst_0.next_rs2\[54\] _1348_ _1349_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1672_ _1292_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2190__A2 picorv32_pcpi_mul_inst_0.rd\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2224_ _0524_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2155_ _0523_ _0529_ _1419_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2086_ _0460_ _0462_ _0466_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2988_ _0105_ clknet_leaf_43_clk picorv32_pcpi_mul_inst_0.rd\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1939_ _0327_ _0333_ _0335_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2911_ _0028_ clknet_leaf_39_clk picorv32_pcpi_mul_inst_0.next_rs2\[18\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2842_ _1034_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2773_ net86 _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1724_ _1333_ _1326_ _1334_ _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_79_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1655_ _1166_ _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1586_ _1124_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1910__A2 _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2207_ _0573_ _0576_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2138_ _0513_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2069_ _0449_ _0450_ _0451_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_76_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1901__A2 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1968__A2 picorv32_pcpi_mul_inst_0.rd\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1440_ picorv32_pcpi_mul_inst_0.instr_mulh picorv32_pcpi_mul_inst_0.instr_mulhu picorv32_pcpi_mul_inst_0.instr_mulhsu
+ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2758__I net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3110_ _0227_ clknet_leaf_45_clk net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3041_ _0158_ clknet_leaf_46_clk picorv32_pcpi_mul_inst_0.next_rs1\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1959__A2 picorv32_pcpi_mul_inst_0.rd\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2825_ _0703_ _1063_ _1069_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2756_ picorv32_pcpi_mul_inst_0.rd\[39\] _1013_ _1003_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1707_ _1315_ _1308_ _1320_ _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2687_ _0956_ _0957_ _0958_ _0959_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1592__C2 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1638_ _1264_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1569_ _1206_ picorv32_pcpi_mul_inst_0.next_rs2\[18\] _1212_ _1208_ _1209_ net59
+ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_39_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2127__A2 picorv32_pcpi_mul_inst_0.next_rs2\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2610_ picorv32_pcpi_mul_inst_0.next_rs1\[35\] _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2541_ _0853_ picorv32_pcpi_mul_inst_0.next_rs1\[12\] picorv32_pcpi_mul_inst_0.next_rs1\[13\]
+ _0851_ _0855_ net23 _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XANTENNA__1574__B1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2472_ _0433_ _0436_ _0434_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_50_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1877__A1 picorv32_pcpi_mul_inst_0.rd\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3024_ _0141_ clknet_leaf_46_clk picorv32_pcpi_mul_inst_0.rdx\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2437__B _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2808_ picorv32_pcpi_mul_inst_0.rd\[17\] _1051_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2739_ _0999_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input53_I pcpi_rs2[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_clk_I clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1972_ _0357_ _0359_ _0364_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_55_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2339__A2 _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2524_ _0844_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2455_ picorv32_pcpi_mul_inst_0.rd\[3\] _0798_ _0255_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2386_ picorv32_pcpi_mul_inst_0.next_rs2\[57\] _0525_ picorv32_pcpi_mul_inst_0.rd\[56\]
+ _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_3_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2275__A1 _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3007_ _0124_ clknet_leaf_23_clk picorv32_pcpi_mul_inst_0.rd\[47\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_46_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_85_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2266__A1 _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2591__I _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2240_ _0603_ _0606_ _1419_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2171_ _0544_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_76_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1480__A2 _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1955_ picorv32_pcpi_mul_inst_0.next_rs2\[14\] _0272_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1886_ _0281_ _0284_ _0287_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2507_ _0833_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2438_ _0779_ _0782_ _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2369_ _0718_ _0722_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input16_I pcpi_insn[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output84_I net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_73_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1740_ _1333_ _1343_ _1347_ _1348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1671_ _1287_ _1288_ _1291_ _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I pcpi_insn[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2478__A1 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2223_ _0589_ _1288_ _0590_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2154_ _0526_ _0528_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2085_ picorv32_pcpi_mul_inst_0.rd\[26\] picorv32_pcpi_mul_inst_0.next_rs2\[27\]
+ _0363_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_48_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2987_ _0104_ clknet_leaf_33_clk picorv32_pcpi_mul_inst_0.rd\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1938_ _0286_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1869_ _1422_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput80 pcpi_rs2[7] net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_43_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2910_ _0027_ clknet_leaf_39_clk picorv32_pcpi_mul_inst_0.next_rs2\[17\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2841_ _1119_ _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_75_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2772_ _1024_ _1016_ _1025_ _1026_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1723_ _1319_ picorv32_pcpi_mul_inst_0.next_rs2\[50\] _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1654_ _1277_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1585_ _1223_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2163__A3 _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2206_ _0570_ _0575_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2137_ _1401_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2068_ _0440_ picorv32_pcpi_mul_inst_0.rdx\[24\] _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_93_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input83_I resetn vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_30_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2090__A2 _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3040_ _0157_ clknet_leaf_47_clk picorv32_pcpi_mul_inst_0.rs1\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2824_ _0978_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2755_ _1114_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2686_ _0950_ picorv32_pcpi_mul_inst_0.next_rs1\[55\] _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1706_ _1319_ picorv32_pcpi_mul_inst_0.next_rs2\[47\] _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1637_ _1247_ picorv32_pcpi_mul_inst_0.next_rs2\[35\] _1263_ _1264_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2136__A3 _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1568_ _1211_ _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1499_ _1159_ _1161_ _1162_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2127__A3 _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2532__C2 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1938__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2540_ _0839_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2471_ _0803_ _0809_ _0810_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1574__A1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2769__I net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3023_ _0140_ clknet_leaf_5_clk picorv32_pcpi_mul_inst_0.rd\[63\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_66_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2807_ net92 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2738_ _1118_ _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2669_ picorv32_pcpi_mul_inst_0.next_rs1\[50\] _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input46_I pcpi_rs1[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2348__A3 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1493__I _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2808__A1 picorv32_pcpi_mul_inst_0.rd\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1971_ picorv32_pcpi_mul_inst_0.rd\[14\] picorv32_pcpi_mul_inst_0.next_rs2\[15\]
+ _0363_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_71_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1668__I _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2523_ _0837_ picorv32_pcpi_mul_inst_0.next_rs1\[6\] picorv32_pcpi_mul_inst_0.next_rs1\[7\]
+ _0843_ _0840_ net48 _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_11_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2454_ _0253_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2385_ _0736_ _1359_ _1437_ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_3_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput1 pcpi_insn[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_48_clk clknet_2_0__leaf_clk clknet_leaf_48_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3006_ _0123_ clknet_leaf_25_clk picorv32_pcpi_mul_inst_0.rd\[46\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1578__I _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_39_clk clknet_2_1__leaf_clk clknet_leaf_39_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_17_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2170_ _0534_ _0543_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_76_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1954_ _0346_ _0347_ _0348_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_28_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1885_ _0286_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2193__A1 picorv32_pcpi_mul_inst_0.rd\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2506_ _0830_ picorv32_pcpi_mul_inst_0.next_rs1\[0\] picorv32_pcpi_mul_inst_0.next_rs1\[1\]
+ _0826_ _0832_ net30 _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2437_ _0779_ _0782_ _0783_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2368_ picorv32_pcpi_mul_inst_0.next_rs2\[55\] _1436_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2299_ picorv32_pcpi_mul_inst_0.rd\[47\] picorv32_pcpi_mul_inst_0.next_rs2\[48\]
+ _0620_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_clkbuf_leaf_2_clk_I clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1670_ _1279_ _1289_ _1290_ _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_33_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2222_ _1404_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2153_ picorv32_pcpi_mul_inst_0.next_rs2\[34\] _0527_ picorv32_pcpi_mul_inst_0.rd\[33\]
+ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2084_ _0463_ _0464_ _0465_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2986_ _0103_ clknet_leaf_33_clk picorv32_pcpi_mul_inst_0.rd\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1937_ _0327_ _0333_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1868_ _0268_ _0269_ _0270_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput81 pcpi_rs2[8] net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput70 pcpi_rs2[27] net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1799_ _1171_ picorv32_pcpi_mul_inst_0.next_rs1\[62\] _1396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_87_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1591__I _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output115_I net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2371__B _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1904__A1 _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2840_ net100 _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2771_ picorv32_pcpi_mul_inst_0.rd\[42\] _1013_ _1019_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1722_ _1278_ _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1653_ _1269_ picorv32_pcpi_mul_inst_0.next_rs2\[38\] _1276_ _1277_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1584_ _1215_ picorv32_pcpi_mul_inst_0.next_rs2\[23\] _1221_ picorv32_pcpi_mul_inst_0.next_rs2\[22\]
+ _1219_ net65 _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2205_ picorv32_pcpi_mul_inst_0.next_rs2\[39\] _0574_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2320__A1 picorv32_pcpi_mul_inst_0.rd\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2136_ _0511_ _1248_ _1405_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_92_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2067_ picorv32_pcpi_mul_inst_0.next_rs2\[25\] _0381_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2969_ _0086_ clknet_leaf_42_clk picorv32_pcpi_mul_inst_0.rd\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1586__I _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input76_I pcpi_rs2[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_42_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2823_ _0407_ _1067_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2754_ picorv32_pcpi_mul_inst_0.rd\[7\] _1001_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1705_ _1300_ _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2685_ _0935_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1636_ _1261_ _1253_ _1262_ _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1567_ _1173_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1498_ picorv32_pcpi_mul_inst_0.mul_counter\[2\] _1156_ _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2119_ picorv32_pcpi_mul_inst_0.next_rs2\[31\] _1439_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3099_ _0216_ clknet_leaf_8_clk picorv32_pcpi_mul_inst_0.next_rs1\[58\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2470_ _0807_ picorv32_pcpi_mul_inst_0.rdx\[20\] _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2771__A1 picorv32_pcpi_mul_inst_0.rd\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1877__A3 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3022_ _0139_ clknet_leaf_18_clk picorv32_pcpi_mul_inst_0.rd\[62\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_66_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2806_ _1049_ _1050_ _1052_ _1054_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2737_ net110 _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2668_ _0932_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1619_ picorv32_pcpi_mul_inst_0.next_rs2\[33\] _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2599_ picorv32_pcpi_mul_inst_0.next_rs1\[32\] _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_6_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input39_I pcpi_rs1[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1774__I _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ _0330_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_71_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2522_ _0783_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2453_ _1150_ _0795_ _0797_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2384_ picorv32_pcpi_mul_inst_0.rd\[56\] _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_79_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput2 pcpi_insn[12] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3005_ _0122_ clknet_2_3__leaf_clk picorv32_pcpi_mul_inst_0.rd\[45\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2275__A3 _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1859__I _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2735__A1 picorv32_pcpi_mul_inst_0.rd\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2266__A3 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1953_ _0339_ picorv32_pcpi_mul_inst_0.rdx\[12\] _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1884_ _1145_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2505_ _1218_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1940__A2 picorv32_pcpi_mul_inst_0.rd\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2436_ _1173_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_16_Left_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2367_ picorv32_pcpi_mul_inst_0.rd\[54\] picorv32_pcpi_mul_inst_0.next_rs2\[55\]
+ _0651_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2298_ _0650_ _0655_ _0652_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2194__B picorv32_pcpi_mul_inst_0.rd\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2221_ picorv32_pcpi_mul_inst_0.rd\[40\] _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2152_ _0513_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2083_ _0447_ picorv32_pcpi_mul_inst_0.rd\[26\] _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2985_ _0102_ clknet_leaf_34_clk picorv32_pcpi_mul_inst_0.rd\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1936_ _0329_ _0332_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1867_ _0259_ picorv32_pcpi_mul_inst_0.rdx\[4\] _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput71 pcpi_rs2[28] net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput60 pcpi_rs2[18] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput82 pcpi_rs2[9] net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1798_ _1394_ _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1913__A2 _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2419_ _0742_ picorv32_pcpi_mul_inst_0.rd\[59\] _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input21_I pcpi_rs1[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output108_I net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2770_ picorv32_pcpi_mul_inst_0.rd\[10\] _1017_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_41_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1721_ _1332_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_1__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1652_ _1261_ _1271_ _1275_ _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_1_clk_I clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1583_ _1222_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2204_ _1403_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_49_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2135_ picorv32_pcpi_mul_inst_0.rd\[32\] _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_92_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2066_ picorv32_pcpi_mul_inst_0.rd\[24\] picorv32_pcpi_mul_inst_0.rdx\[24\] _0449_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2968_ _0085_ clknet_leaf_42_clk picorv32_pcpi_mul_inst_0.rd\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1919_ picorv32_pcpi_mul_inst_0.rd\[9\] picorv32_pcpi_mul_inst_0.next_rs2\[10\] _0278_
+ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2899_ _0016_ clknet_leaf_48_clk picorv32_pcpi_mul_inst_0.next_rs2\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input69_I pcpi_rs2[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1822__A1 _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2822_ _1034_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2753_ net113 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1704_ _1318_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2684_ picorv32_pcpi_mul_inst_0.next_rs1\[54\] _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1635_ _1243_ picorv32_pcpi_mul_inst_0.next_rs2\[34\] _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1566_ _1210_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1497_ _1160_ _1134_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_69_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2118_ _0488_ _0490_ _0495_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3098_ _0215_ clknet_leaf_9_clk picorv32_pcpi_mul_inst_0.next_rs1\[57\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2049_ picorv32_pcpi_mul_inst_0.rd\[23\] picorv32_pcpi_mul_inst_0.next_rs2\[24\]
+ _0328_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_49_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1804__A1 _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1970__I _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3021_ _0138_ clknet_leaf_18_clk picorv32_pcpi_mul_inst_0.rd\[61\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2287__A1 _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2805_ _0667_ _1047_ _1053_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2736_ _0994_ _0980_ _0995_ _0997_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2667_ _0933_ _0943_ _0936_ _0944_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1618_ _1168_ _1247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2598_ _0886_ _0891_ _1395_ _0893_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1880__I _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1549_ _1198_ picorv32_pcpi_mul_inst_0.next_rs2\[12\] _1195_ picorv32_pcpi_mul_inst_0.next_rs2\[11\]
+ _1193_ net53 _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XTAP_TAPCELL_ROW_6_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_41_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2521_ _0842_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2452_ _0796_ picorv32_pcpi_mul_inst_0.rd\[63\] _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2383_ picorv32_pcpi_mul_inst_0.rdx\[56\] _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_46_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput3 pcpi_insn[13] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3004_ _0121_ clknet_leaf_20_clk picorv32_pcpi_mul_inst_0.rd\[44\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_62_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2719_ picorv32_pcpi_mul_inst_0.rd\[0\] _0983_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input51_I pcpi_rs2[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1952_ picorv32_pcpi_mul_inst_0.next_rs2\[13\] _1424_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1883_ _0281_ _0284_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2504_ _0831_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2193__A3 _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2435_ _0780_ _0781_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2366_ _0712_ _0715_ _0713_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2297_ _0658_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_82_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2220_ picorv32_pcpi_mul_inst_0.rdx\[40\] _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2151_ picorv32_pcpi_mul_inst_0.rd\[33\] picorv32_pcpi_mul_inst_0.next_rs2\[34\]
+ _0525_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_17_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2082_ _0460_ _0462_ _0429_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2984_ _0101_ clknet_leaf_34_clk picorv32_pcpi_mul_inst_0.rd\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1935_ picorv32_pcpi_mul_inst_0.next_rs2\[12\] _0331_ picorv32_pcpi_mul_inst_0.rd\[11\]
+ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2314__I _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1866_ picorv32_pcpi_mul_inst_0.next_rs2\[5\] _1424_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput50 pcpi_rs1[9] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput72 pcpi_rs2[29] net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput61 pcpi_rs2[19] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1797_ _1393_ _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput83 resetn net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_87_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2418_ _0762_ _0765_ _0699_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2349_ picorv32_pcpi_mul_inst_0.next_rs2\[53\] _0592_ picorv32_pcpi_mul_inst_0.rd\[52\]
+ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_input14_I pcpi_insn[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_35_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1720_ _1323_ picorv32_pcpi_mul_inst_0.next_rs2\[50\] _1331_ _1332_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_44_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1651_ _1265_ _1270_ _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1582_ _1215_ picorv32_pcpi_mul_inst_0.next_rs2\[22\] _1221_ _1217_ _1219_ net64
+ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_0_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I pcpi_insn[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2203_ picorv32_pcpi_mul_inst_0.rd\[38\] picorv32_pcpi_mul_inst_0.next_rs2\[39\]
+ _0536_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_49_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2134_ picorv32_pcpi_mul_inst_0.rdx\[32\] _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_53_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_92_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2065_ _0442_ _0445_ _0448_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2967_ _0084_ clknet_leaf_47_clk picorv32_pcpi_mul_inst_0.rd\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1918_ _0314_ _0315_ _0316_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2898_ _0015_ clknet_leaf_49_clk picorv32_pcpi_mul_inst_0.next_rs2\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_62_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1849_ picorv32_pcpi_mul_inst_0.rd\[3\] _0253_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_71_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk clknet_leaf_20_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_46_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2821_ _1119_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2752_ _1008_ _1000_ _1009_ _1010_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1703_ _1306_ picorv32_pcpi_mul_inst_0.next_rs2\[47\] _1317_ _1318_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2683_ _0932_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1634_ _1260_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1565_ _1206_ _1208_ _1203_ picorv32_pcpi_mul_inst_0.next_rs2\[16\] _1209_ net58
+ _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1496_ _1144_ _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2117_ _0494_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3097_ _0214_ clknet_leaf_9_clk picorv32_pcpi_mul_inst_0.next_rs1\[56\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2048_ _0425_ _0427_ _0432_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input81_I pcpi_rs2[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2502__I _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_0_clk_I clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3020_ _0137_ clknet_leaf_19_clk picorv32_pcpi_mul_inst_0.rd\[60\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2804_ _0978_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_14_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2735_ picorv32_pcpi_mul_inst_0.rd\[35\] _0996_ _0986_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2666_ _0939_ picorv32_pcpi_mul_inst_0.next_rs1\[50\] _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1617_ _1245_ _1246_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2597_ _0892_ picorv32_pcpi_mul_inst_0.next_rs1\[32\] _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1548_ _1189_ _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_6_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1479_ _1146_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1961__A1 picorv32_pcpi_mul_inst_0.rd\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2520_ _0837_ picorv32_pcpi_mul_inst_0.next_rs1\[5\] picorv32_pcpi_mul_inst_0.next_rs1\[6\]
+ _0835_ _0840_ net47 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2451_ _0673_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2382_ _0732_ _0733_ _0734_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_79_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput4 pcpi_insn[14] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3003_ _0120_ clknet_leaf_23_clk picorv32_pcpi_mul_inst_0.rd\[43\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_2_1__f_clk clknet_0_clk clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_93_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_62_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2718_ _0982_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2649_ _0926_ picorv32_pcpi_mul_inst_0.next_rs1\[46\] _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input44_I pcpi_rs1[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2187__A1 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2137__I _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1951_ picorv32_pcpi_mul_inst_0.rd\[12\] picorv32_pcpi_mul_inst_0.rdx\[12\] _0346_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1882_ picorv32_pcpi_mul_inst_0.rd\[6\] _0283_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2503_ _0830_ _1406_ _1238_ picorv32_pcpi_mul_inst_0.next_rs1\[0\] _1236_ net19 _0831_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2434_ picorv32_pcpi_mul_inst_0.next_rs2\[62\] _1402_ picorv32_pcpi_mul_inst_0.rd\[61\]
+ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2365_ _1250_ _0718_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2296_ _0649_ _0657_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2102__A1 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_40_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2510__I _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1604__C2 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2150_ _0524_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2081_ _0460_ _0462_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_8_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2983_ _0100_ clknet_leaf_36_clk picorv32_pcpi_mul_inst_0.rd\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1934_ _0330_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1865_ picorv32_pcpi_mul_inst_0.rd\[4\] picorv32_pcpi_mul_inst_0.rdx\[4\] _0268_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput40 pcpi_rs1[29] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput73 pcpi_rs2[2] net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput62 pcpi_rs2[1] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput51 pcpi_rs2[0] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1796_ _1167_ _1392_ _1393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2417_ _0762_ _0765_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_87_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2348_ _0703_ _1342_ _0590_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2279_ _0513_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2505__I _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1650_ _1274_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1581_ _1211_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2202_ _0563_ _0566_ _0564_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2133_ _0507_ _0508_ _0509_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_49_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2064_ _0447_ _0440_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2966_ _0083_ clknet_leaf_47_clk picorv32_pcpi_mul_inst_0.rd\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1917_ _0306_ picorv32_pcpi_mul_inst_0.rd\[9\] _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2897_ _0014_ clknet_leaf_46_clk picorv32_pcpi_mul_inst_0.next_rs2\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1848_ picorv32_pcpi_mul_inst_0.next_rs2\[4\] _1439_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2792__A1 picorv32_pcpi_mul_inst_0.rd\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1779_ _1375_ _1376_ _1379_ _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output113_I net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2783__A1 _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2820_ net96 _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2751_ picorv32_pcpi_mul_inst_0.rd\[38\] _0996_ _1003_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1702_ _1315_ _1308_ _1316_ _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2774__A1 picorv32_pcpi_mul_inst_0.rd\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2682_ _0945_ _0954_ _0947_ _0955_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1633_ _1166_ _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1564_ _1183_ _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1495_ _1155_ _1156_ _1159_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2116_ picorv32_pcpi_mul_inst_0.rd\[29\] picorv32_pcpi_mul_inst_0.next_rs2\[30\]
+ _1427_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3096_ _0213_ clknet_leaf_9_clk picorv32_pcpi_mul_inst_0.next_rs1\[55\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2047_ picorv32_pcpi_mul_inst_0.rd\[22\] picorv32_pcpi_mul_inst_0.next_rs2\[23\]
+ _0363_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_49_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2949_ _0066_ clknet_leaf_28_clk picorv32_pcpi_mul_inst_0.next_rs2\[56\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input74_I pcpi_rs2[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2756__A1 picorv32_pcpi_mul_inst_0.rd\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2508__B2 _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2803_ _0372_ _1051_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2747__A1 picorv32_pcpi_mul_inst_0.rd\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2734_ _1114_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2665_ picorv32_pcpi_mul_inst_0.next_rs1\[49\] _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1616_ _1171_ picorv32_pcpi_mul_inst_0.next_rs2\[32\] _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2596_ _1388_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1547_ _1197_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1478_ _1145_ _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3079_ _0196_ clknet_leaf_13_clk picorv32_pcpi_mul_inst_0.next_rs1\[38\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2513__I _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1952__A2 _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2450_ picorv32_pcpi_mul_inst_0.rd\[63\] _0793_ _0794_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2381_ _0674_ picorv32_pcpi_mul_inst_0.rd\[55\] _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_79_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput5 pcpi_insn[1] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3002_ _0119_ clknet_leaf_21_clk picorv32_pcpi_mul_inst_0.rd\[42\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2717_ _0981_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2648_ picorv32_pcpi_mul_inst_0.next_rs1\[45\] _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2579_ _0858_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input37_I pcpi_rs1[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2423__A3 _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2243__I picorv32_pcpi_mul_inst_0.rd\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2399__B _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1950_ _0341_ _0343_ _0345_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2414__A3 _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1881_ picorv32_pcpi_mul_inst_0.next_rs2\[7\] _0282_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2502_ _1224_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_24_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2433_ picorv32_pcpi_mul_inst_0.rd\[61\] picorv32_pcpi_mul_inst_0.next_rs2\[62\]
+ _1422_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2364_ picorv32_pcpi_mul_inst_0.rd\[54\] _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2295_ _0650_ _0655_ _0656_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1861__A1 _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1456__A4 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2405__A3 _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2063__I _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1852__A1 _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1907__A2 _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2080_ picorv32_pcpi_mul_inst_0.rd\[26\] _0461_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2982_ _0099_ clknet_leaf_36_clk picorv32_pcpi_mul_inst_0.rd\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1933_ _1403_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1864_ _0261_ _0265_ _0267_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput30 pcpi_rs1[1] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 pcpi_rs2[10] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 pcpi_rs1[2] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput63 pcpi_rs2[20] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1795_ picorv32_pcpi_mul_inst_0.instr_mulh picorv32_pcpi_mul_inst_0.instr_mulhsu
+ _1132_ net43 _1392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2611__I _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput74 pcpi_rs2[30] net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2416_ _0763_ _0764_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_87_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2347_ picorv32_pcpi_mul_inst_0.rd\[52\] _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2278_ picorv32_pcpi_mul_inst_0.rd\[45\] picorv32_pcpi_mul_inst_0.next_rs2\[46\]
+ _0640_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_35_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1522__B1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1522__C2 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1580_ _1220_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2201_ _0569_ _0570_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2132_ _0483_ picorv32_pcpi_mul_inst_0.rd\[31\] _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2063_ _0446_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2965_ _0082_ clknet_leaf_48_clk picorv32_pcpi_mul_inst_0.rd\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1916_ _0311_ _0313_ _0287_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2896_ _0013_ clknet_leaf_4_clk picorv32_pcpi_mul_inst_0.next_rs2\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1847_ _1423_ _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1778_ _1367_ _1377_ _1378_ _1379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_67_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2516__I _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output106_I net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2299__A1 picorv32_pcpi_mul_inst_0.rd\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2471__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2750_ picorv32_pcpi_mul_inst_0.rd\[6\] _1001_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2223__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1701_ _1301_ picorv32_pcpi_mul_inst_0.next_rs2\[46\] _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2681_ _0950_ picorv32_pcpi_mul_inst_0.next_rs1\[54\] _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1632_ _1259_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1563_ picorv32_pcpi_mul_inst_0.next_rs2\[17\] _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_39_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1494_ _1158_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1505__I _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2115_ _0491_ _0492_ _0493_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3095_ _0212_ clknet_leaf_9_clk picorv32_pcpi_mul_inst_0.next_rs1\[54\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2046_ _0428_ _0430_ _0431_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2948_ _0065_ clknet_leaf_28_clk picorv32_pcpi_mul_inst_0.next_rs2\[55\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2879_ picorv32_pcpi_mul_inst_0.mul_counter\[5\] _1169_ _1111_ _1112_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input67_I pcpi_rs2[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2453__A1 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2802_ _1034_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_14_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2733_ picorv32_pcpi_mul_inst_0.rd\[3\] _0983_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2664_ _0933_ _0941_ _0936_ _0942_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1615_ _1243_ picorv32_pcpi_mul_inst_0.next_rs2\[31\] _1244_ _1152_ _1245_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2595_ picorv32_pcpi_mul_inst_0.next_rs1\[31\] _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1546_ _1190_ picorv32_pcpi_mul_inst_0.next_rs2\[11\] _1195_ picorv32_pcpi_mul_inst_0.next_rs2\[10\]
+ _1193_ net52 _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_1_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1477_ _1132_ _1144_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_65_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3078_ _0195_ clknet_leaf_13_clk picorv32_pcpi_mul_inst_0.next_rs1\[37\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2029_ _0407_ picorv32_pcpi_mul_inst_0.rdx\[20\] _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_59_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1961__A3 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_77_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_86_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_11_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2380_ _0728_ _0731_ _0699_ _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 pcpi_insn[25] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3001_ _0118_ clknet_leaf_21_clk picorv32_pcpi_mul_inst_0.rd\[41\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_19_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2716_ picorv32_pcpi_mul_inst_0.instr_mulh picorv32_pcpi_mul_inst_0.instr_mulhu picorv32_pcpi_mul_inst_0.instr_mulhsu
+ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2647_ _0920_ _0928_ _0922_ _0929_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2578_ _0879_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1529_ _1185_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1603__I _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1870__A2 _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1880_ _1426_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2501_ _0829_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2432_ _0769_ _0772_ _0778_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2363_ _0710_ _0717_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2294_ _0650_ _0655_ _0541_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_73_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2981_ _0098_ clknet_leaf_36_clk picorv32_pcpi_mul_inst_0.rd\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1932_ picorv32_pcpi_mul_inst_0.rd\[11\] picorv32_pcpi_mul_inst_0.next_rs2\[12\]
+ _0328_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xclkbuf_leaf_41_clk clknet_2_1__leaf_clk clknet_leaf_41_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1863_ _0266_ _0259_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput20 pcpi_rs1[10] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput31 pcpi_rs1[20] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 pcpi_rs2[11] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput64 pcpi_rs2[21] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput42 pcpi_rs1[30] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1794_ _1391_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput75 pcpi_rs2[31] net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2415_ picorv32_pcpi_mul_inst_0.next_rs2\[60\] _0290_ picorv32_pcpi_mul_inst_0.rd\[59\]
+ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_87_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1531__A1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2346_ picorv32_pcpi_mul_inst_0.rdx\[52\] _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2277_ _0524_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_32_clk clknet_2_1__leaf_clk clknet_leaf_32_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1522__A1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_23_clk clknet_2_3__leaf_clk clknet_leaf_23_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2712__I net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2200_ picorv32_pcpi_mul_inst_0.rd\[38\] _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2131_ _0503_ _0506_ _0475_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2062_ _1160_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_49_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_22_Left_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2964_ _0081_ clknet_leaf_46_clk picorv32_pcpi_mul_inst_0.rd\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_32_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1915_ _0311_ _0313_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_44_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_14_clk clknet_2_2__leaf_clk clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2895_ _0012_ clknet_leaf_4_clk picorv32_pcpi_mul_inst_0.next_rs2\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1846_ picorv32_pcpi_mul_inst_0.rd\[2\] picorv32_pcpi_mul_inst_0.next_rs2\[3\] _1437_
+ _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_71_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1777_ _1371_ picorv32_pcpi_mul_inst_0.next_rs2\[60\] _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_31_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2329_ picorv32_pcpi_mul_inst_0.rd\[50\] picorv32_pcpi_mul_inst_0.next_rs2\[51\]
+ _0651_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input12_I pcpi_insn[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_40_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2680_ picorv32_pcpi_mul_inst_0.next_rs1\[53\] _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1700_ _1278_ _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1631_ _1247_ picorv32_pcpi_mul_inst_0.next_rs2\[34\] _1258_ _1259_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1562_ _1207_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1493_ _1157_ _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input4_I pcpi_insn[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2114_ _0483_ picorv32_pcpi_mul_inst_0.rd\[29\] _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3094_ _0211_ clknet_leaf_9_clk picorv32_pcpi_mul_inst_0.next_rs1\[53\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1521__I _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2045_ _0412_ picorv32_pcpi_mul_inst_0.rd\[22\] _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2947_ _0064_ clknet_leaf_28_clk picorv32_pcpi_mul_inst_0.next_rs2\[54\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2214__A2 _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1973__A1 picorv32_pcpi_mul_inst_0.rd\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2878_ _1133_ _0982_ _1137_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1829_ picorv32_pcpi_mul_inst_0.rs1\[0\] _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2205__A2 _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2801_ _0999_ _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2732_ net109 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2663_ _0939_ picorv32_pcpi_mul_inst_0.next_rs1\[49\] _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1614_ _1132_ net75 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2594_ _0886_ _0887_ _0889_ _0890_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1545_ _1196_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1476_ net83 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3077_ _0194_ clknet_leaf_11_clk picorv32_pcpi_mul_inst_0.next_rs1\[36\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2028_ picorv32_pcpi_mul_inst_0.next_rs2\[21\] _0381_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2257__I _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 pcpi_insn[26] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3000_ _0117_ clknet_leaf_20_clk picorv32_pcpi_mul_inst_0.rd\[40\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2167__I _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2715_ _0979_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2646_ _0926_ picorv32_pcpi_mul_inst_0.next_rs1\[45\] _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2577_ _0875_ picorv32_pcpi_mul_inst_0.next_rs1\[25\] picorv32_pcpi_mul_inst_0.next_rs1\[26\]
+ _0873_ _0877_ net37 _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XANTENNA__2353__A1 _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1528_ _1179_ _1181_ _1175_ picorv32_pcpi_mul_inst_0.next_rs2\[4\] _1184_ net77 _1185_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1459_ _1126_ _1127_ _1129_ _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_2_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3129_ _0246_ clknet_leaf_30_clk net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1919__A1 picorv32_pcpi_mul_inst_0.rd\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2344__A1 _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1607__C2 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2500_ picorv32_pcpi_mul_inst_0.pcpi_wait_q _0828_ _1176_ _0826_ picorv32_pcpi_mul_inst_0.mul_counter\[6\]
+ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2431_ _0770_ _1376_ _1402_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2362_ _0712_ _0715_ _0716_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2293_ _0652_ _0654_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2629_ picorv32_pcpi_mul_inst_0.next_rs1\[40\] _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input42_I pcpi_rs1[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2317__A1 _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2980_ _0097_ clknet_leaf_37_clk picorv32_pcpi_mul_inst_0.rd\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1931_ _0282_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1862_ _1398_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput21 pcpi_rs1[11] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput10 pcpi_insn[29] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput54 pcpi_rs2[12] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 pcpi_rs1[21] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 pcpi_rs1[31] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1793_ _1375_ picorv32_pcpi_mul_inst_0.rs2\[63\] _1390_ _1391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput65 pcpi_rs2[22] net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput76 pcpi_rs2[3] net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2308__A1 _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2414_ picorv32_pcpi_mul_inst_0.rd\[59\] picorv32_pcpi_mul_inst_0.next_rs2\[60\]
+ _0536_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2345_ _0698_ _0700_ _0701_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2276_ _0628_ _0631_ _0638_ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_35_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1522__A2 picorv32_pcpi_mul_inst_0.next_rs2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2483__B1 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2214__B picorv32_pcpi_mul_inst_0.rd\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2130_ _0503_ _0506_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2061_ _0443_ _0444_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2963_ _0080_ clknet_leaf_46_clk picorv32_pcpi_mul_inst_0.rd\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_32_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1914_ picorv32_pcpi_mul_inst_0.rd\[9\] _0312_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2777__A1 picorv32_pcpi_mul_inst_0.rd\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2894_ _0011_ clknet_leaf_8_clk picorv32_pcpi_mul_inst_0.instr_mulhu vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1845_ _1436_ _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1776_ _1325_ _1377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2328_ _0678_ _0681_ _0679_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_79_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2259_ _0621_ _0623_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1991__A2 _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1873__B _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2299__A3 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2223__A3 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1982__A2 _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1630_ _1250_ _1253_ _1257_ _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_81_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1561_ _1206_ picorv32_pcpi_mul_inst_0.next_rs2\[16\] _1203_ picorv32_pcpi_mul_inst_0.next_rs2\[15\]
+ _1201_ net57 _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1492_ picorv32_pcpi_mul_inst_0.mul_waiting _1117_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2113_ _0488_ _0490_ _0475_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1802__I _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3093_ _0210_ clknet_leaf_9_clk picorv32_pcpi_mul_inst_0.next_rs1\[52\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2044_ _0425_ _0427_ _0429_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2946_ _0063_ clknet_leaf_28_clk picorv32_pcpi_mul_inst_0.next_rs2\[53\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2877_ _1108_ _1109_ _1110_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1828_ _1416_ _1421_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1759_ _1363_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1712__I _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output111_I net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1964__A2 _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2800_ net91 _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_14_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2731_ _0991_ _0980_ _0992_ _0993_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1955__A2 _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2662_ picorv32_pcpi_mul_inst_0.next_rs1\[48\] _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2593_ _1133_ net43 _1152_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1613_ _1242_ _1243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1544_ _1190_ picorv32_pcpi_mul_inst_0.next_rs2\[10\] _1195_ _1192_ _1193_ net82
+ _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_1_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1475_ _1143_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3076_ _0193_ clknet_leaf_11_clk picorv32_pcpi_mul_inst_0.next_rs1\[35\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2027_ picorv32_pcpi_mul_inst_0.rd\[20\] picorv32_pcpi_mul_inst_0.rdx\[20\] _0414_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_65_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2929_ _0046_ clknet_leaf_14_clk picorv32_pcpi_mul_inst_0.next_rs2\[36\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1946__A2 _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input72_I pcpi_rs2[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_5_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1882__A1 picorv32_pcpi_mul_inst_0.rd\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2273__I _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 pcpi_insn[27] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2714_ _0978_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1527__I _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2645_ picorv32_pcpi_mul_inst_0.next_rs1\[44\] _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2576_ _0878_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1527_ _1183_ _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1458_ net17 net7 _1128_ net9 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_TAPCELL_ROW_2_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3128_ _0245_ clknet_leaf_30_clk net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3059_ _0176_ clknet_leaf_2_clk picorv32_pcpi_mul_inst_0.next_rs1\[18\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1616__A1 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2093__I _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2430_ _1399_ picorv32_pcpi_mul_inst_0.rd\[61\] _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2361_ _0712_ _0715_ _0645_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2292_ _0648_ _0653_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1810__I _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2023__A1 _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2628_ _0909_ _0913_ _0911_ _0915_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2559_ _0867_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input35_I pcpi_rs1[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2317__A2 picorv32_pcpi_mul_inst_0.rd\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ _0319_ _0322_ _0326_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1861_ _1147_ _0264_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput22 pcpi_rs1[12] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2005__A1 picorv32_pcpi_mul_inst_0.rd\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput11 pcpi_insn[2] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput44 pcpi_rs1[3] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput55 pcpi_rs2[13] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput33 pcpi_rs1[22] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1792_ _1384_ _1377_ _1389_ _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput77 pcpi_rs2[4] net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput66 pcpi_rs2[23] net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2413_ _0754_ _0758_ _0755_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2344_ _0674_ picorv32_pcpi_mul_inst_0.rd\[51\] _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2275_ _0629_ _1307_ _0601_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_74_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1540__I _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2244__A1 _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2235__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2060_ _1227_ _0375_ _0441_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2474__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2962_ _0079_ clknet_leaf_4_clk picorv32_pcpi_mul_inst_0.rd\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1913_ picorv32_pcpi_mul_inst_0.next_rs2\[10\] _0272_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2893_ _0000_ clknet_leaf_44_clk net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1844_ _1403_ _1436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1775_ picorv32_pcpi_mul_inst_0.next_rs2\[61\] _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1535__I _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2327_ _0569_ _0684_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2258_ picorv32_pcpi_mul_inst_0.next_rs2\[44\] _0622_ picorv32_pcpi_mul_inst_0.rd\[43\]
+ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2189_ _0557_ _0559_ _0560_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1445__I net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2456__A1 _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1560_ _1189_ _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_34_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1491_ picorv32_pcpi_mul_inst_0.mul_counter\[1\] _1154_ _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2112_ _0488_ _0490_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3092_ _0209_ clknet_leaf_12_clk picorv32_pcpi_mul_inst_0.next_rs1\[51\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2043_ _0286_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2945_ _0062_ clknet_leaf_25_clk picorv32_pcpi_mul_inst_0.next_rs2\[52\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2876_ net108 _1098_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1973__A3 _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1974__B picorv32_pcpi_mul_inst_0.rd\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1827_ _1412_ _1418_ _1420_ _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1758_ _1358_ _1359_ _1362_ _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1689_ _1305_ _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1489__A2 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output104_I net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2730_ picorv32_pcpi_mul_inst_0.rd\[34\] _1115_ _0986_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2661_ _0933_ _0938_ _0936_ _0940_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1612_ _1241_ _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2592_ _0888_ picorv32_pcpi_mul_inst_0.next_rs1\[31\] _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1543_ _1174_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1474_ picorv32_pcpi_mul_inst_0.mul_counter\[6\] _1137_ _1142_ _1135_ _1143_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1813__I _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Left_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3075_ _0192_ clknet_leaf_17_clk picorv32_pcpi_mul_inst_0.next_rs1\[34\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2026_ _0409_ _0411_ _0413_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_65_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_28_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2928_ _0045_ clknet_leaf_14_clk picorv32_pcpi_mul_inst_0.next_rs2\[35\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2859_ _1093_ _1082_ _1094_ _1096_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input65_I pcpi_rs2[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_37_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_46_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1633__I _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 pcpi_insn[28] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1625__A2 picorv32_pcpi_mul_inst_0.next_rs2\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_27_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2050__A2 _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2713_ _1118_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2644_ _0920_ _0924_ _0922_ _0927_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2575_ _0875_ picorv32_pcpi_mul_inst_0.next_rs1\[24\] picorv32_pcpi_mul_inst_0.next_rs1\[25\]
+ _0873_ _0877_ net36 _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1526_ _1182_ _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1543__I _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1457_ net6 _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_2_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3127_ _0244_ clknet_leaf_33_clk net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3058_ _0175_ clknet_leaf_2_clk picorv32_pcpi_mul_inst_0.next_rs1\[17\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2009_ _0396_ _0397_ _0398_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2813__A1 picorv32_pcpi_mul_inst_0.rd\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1616__A2 picorv32_pcpi_mul_inst_0.next_rs2\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1919__A3 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2323__B _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1791__A1 _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ _0713_ _0714_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2291_ picorv32_pcpi_mul_inst_0.next_rs2\[47\] _0574_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_44_clk clknet_2_1__leaf_clk clknet_leaf_44_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2271__A2 _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput110 net110 pcpi_mul_rd[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_30_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2627_ _0914_ picorv32_pcpi_mul_inst_0.next_rs1\[40\] _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2558_ _0861_ picorv32_pcpi_mul_inst_0.next_rs1\[18\] picorv32_pcpi_mul_inst_0.next_rs1\[19\]
+ _0866_ _0863_ net29 _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1509_ _1169_ _1170_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2489_ _1384_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input28_I pcpi_rs1[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1837__A2 _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_35_clk clknet_2_1__leaf_clk clknet_leaf_35_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2262__A2 picorv32_pcpi_mul_inst_0.rd\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_26_clk clknet_2_3__leaf_clk clknet_leaf_26_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1860_ _1181_ _0263_ _0260_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput12 pcpi_insn[30] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1791_ _1388_ picorv32_pcpi_mul_inst_0.next_rs2\[63\] _1389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput23 pcpi_rs1[13] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput45 pcpi_rs1[4] net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput34 pcpi_rs1[23] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput78 pcpi_rs2[5] net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput56 pcpi_rs2[14] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput67 pcpi_rs2[24] net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2412_ _0761_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2308__A3 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2343_ _0694_ _0697_ _0699_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2274_ _0636_ picorv32_pcpi_mul_inst_0.rd\[45\] _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_17_clk clknet_2_2__leaf_clk clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1989_ picorv32_pcpi_mul_inst_0.rd\[16\] picorv32_pcpi_mul_inst_0.rdx\[16\] _0380_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_19_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1906__I _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2737__I net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2961_ _0078_ clknet_leaf_4_clk picorv32_pcpi_mul_inst_0.rd\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1912_ _0308_ _0309_ _0310_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_29_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1985__A1 _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2892_ picorv32_pcpi_mul_inst_0.instr_any_mul clknet_leaf_6_clk net117 vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1843_ _1432_ _1434_ _1435_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_40_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1774_ _1136_ _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1816__I _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_6_clk clknet_2_2__leaf_clk clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2326_ picorv32_pcpi_mul_inst_0.rd\[50\] _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2257_ _0330_ _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2188_ _0519_ _0554_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1900__A1 _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1490_ picorv32_pcpi_mul_inst_0.mul_counter\[1\] _1154_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2111_ picorv32_pcpi_mul_inst_0.rd\[29\] _0489_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_55_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3091_ _0208_ clknet_leaf_12_clk picorv32_pcpi_mul_inst_0.next_rs1\[50\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2042_ _0425_ _0427_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2944_ _0061_ clknet_leaf_26_clk picorv32_pcpi_mul_inst_0.next_rs2\[51\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2875_ picorv32_pcpi_mul_inst_0.rd\[63\] _1099_ _0000_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ _1412_ _1418_ _1419_ _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1757_ _1350_ _1360_ _1361_ _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1688_ _1167_ _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2309_ picorv32_pcpi_mul_inst_0.next_rs2\[49\] _0592_ picorv32_pcpi_mul_inst_0.rd\[48\]
+ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_input10_I pcpi_insn[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_51_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2660_ _0939_ picorv32_pcpi_mul_inst_0.next_rs1\[48\] _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1611_ _1138_ _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2365__A1 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2591_ _1242_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1542_ _1194_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1473_ picorv32_pcpi_mul_inst_0.mul_counter\[6\] _1141_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input2_I pcpi_insn[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3074_ _0191_ clknet_leaf_10_clk picorv32_pcpi_mul_inst_0.next_rs1\[33\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2025_ _0412_ _0407_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2927_ _0044_ clknet_leaf_7_clk picorv32_pcpi_mul_inst_0.next_rs2\[34\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2858_ picorv32_pcpi_mul_inst_0.rd\[59\] _1095_ _1085_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2789_ picorv32_pcpi_mul_inst_0.rd\[45\] _1030_ _1037_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1809_ _1403_ _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input58_I pcpi_rs2[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2745__I net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2586__A1 _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2712_ net84 _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2643_ _0926_ picorv32_pcpi_mul_inst_0.next_rs1\[44\] _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2574_ _1182_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1525_ _1157_ _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1456_ net8 net12 net10 net13 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_TAPCELL_ROW_2_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3126_ _0243_ clknet_leaf_30_clk net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3057_ _0174_ clknet_leaf_0_clk picorv32_pcpi_mul_inst_0.next_rs1\[16\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2008_ _0378_ picorv32_pcpi_mul_inst_0.rd\[18\] _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2390__I _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2329__A1 picorv32_pcpi_mul_inst_0.rd\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1644__I _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2290_ picorv32_pcpi_mul_inst_0.rd\[46\] picorv32_pcpi_mul_inst_0.next_rs2\[47\]
+ _0651_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_47_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1846__A3 _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2475__I _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput100 net100 pcpi_mul_rd[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_65_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2626_ _1388_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput111 net111 pcpi_mul_rd[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2557_ _0858_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1508_ picorv32_pcpi_mul_inst_0.mul_counter\[4\] _1164_ _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2488_ _0816_ _0628_ _0820_ _0821_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2495__B1 _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3109_ _0226_ clknet_leaf_45_clk net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_38_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2798__A1 picorv32_pcpi_mul_inst_0.rd\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_21_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_92_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_1_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1639__I _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 pcpi_insn[31] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1790_ _1241_ _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput24 pcpi_rs1[14] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 pcpi_rs1[5] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 pcpi_rs1[24] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput79 pcpi_rs2[6] net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput68 pcpi_rs2[25] net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput57 pcpi_rs2[15] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2411_ _0753_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2342_ _0474_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2273_ _1398_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1988_ _0374_ _0377_ _0379_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2609_ _0898_ _0899_ _0900_ _0901_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input40_I pcpi_rs1[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_2_2__f_clk clknet_0_clk clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__A3 _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1994__A2 _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2753__I net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2960_ _0077_ clknet_leaf_4_clk picorv32_pcpi_mul_inst_0.rd\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1911_ _0299_ picorv32_pcpi_mul_inst_0.rdx\[8\] _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2891_ _0010_ clknet_leaf_3_clk picorv32_pcpi_mul_inst_0.mul_counter\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1842_ _1399_ picorv32_pcpi_mul_inst_0.rd\[2\] _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1773_ _1374_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2325_ _0676_ _0683_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2256_ picorv32_pcpi_mul_inst_0.rd\[43\] picorv32_pcpi_mul_inst_0.next_rs2\[44\]
+ _0620_ _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2187_ _0443_ _0558_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2153__A2 _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2110_ picorv32_pcpi_mul_inst_0.next_rs2\[30\] _1410_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3090_ _0207_ clknet_leaf_12_clk picorv32_pcpi_mul_inst_0.next_rs1\[49\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2041_ picorv32_pcpi_mul_inst_0.rd\[22\] _0426_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2447__A3 _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2943_ _0060_ clknet_leaf_27_clk picorv32_pcpi_mul_inst_0.next_rs2\[50\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_18_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2874_ picorv32_pcpi_mul_inst_0.rd\[31\] _1114_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1825_ _1140_ _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1756_ _1354_ picorv32_pcpi_mul_inst_0.next_rs2\[56\] _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1687_ _1304_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2308_ _0667_ _1324_ _0590_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2239_ _0604_ _0605_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1949__A2 _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1610_ _1240_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2590_ picorv32_pcpi_mul_inst_0.next_rs1\[30\] _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1541_ _1190_ _1192_ _1186_ picorv32_pcpi_mul_inst_0.next_rs2\[8\] _1193_ net81 _1194_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_1_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1472_ _1140_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3073_ _0190_ clknet_leaf_7_clk picorv32_pcpi_mul_inst_0.next_rs1\[32\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2024_ _0305_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2926_ _0043_ clknet_leaf_17_clk picorv32_pcpi_mul_inst_0.next_rs2\[33\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2857_ _1113_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1808_ _1402_ _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2788_ picorv32_pcpi_mul_inst_0.rd\[13\] _1035_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1739_ _1337_ _1342_ _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1467__I _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2711_ _0967_ _0975_ _0969_ _0976_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_27_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2642_ _0925_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2573_ _0876_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2338__A2 picorv32_pcpi_mul_inst_0.next_rs2\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1524_ picorv32_pcpi_mul_inst_0.next_rs2\[5\] _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1455_ net14 net11 _1123_ _1125_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3125_ _0242_ clknet_leaf_30_clk net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3056_ _0173_ clknet_leaf_0_clk picorv32_pcpi_mul_inst_0.next_rs1\[15\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2007_ _0393_ _0395_ _0388_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2274__A1 _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2909_ _0026_ clknet_leaf_40_clk picorv32_pcpi_mul_inst_0.next_rs2\[16\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input70_I pcpi_rs2[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1528__B1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2256__A1 picorv32_pcpi_mul_inst_0.rd\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput101 net101 pcpi_mul_rd[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2625_ picorv32_pcpi_mul_inst_0.next_rs1\[39\] _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput112 net112 pcpi_mul_rd[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1519__B1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2556_ _0865_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1507_ _1133_ _1165_ _1168_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2487_ _0619_ _0624_ _0621_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2495__A1 _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3108_ _0225_ clknet_leaf_45_clk net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3039_ _0156_ clknet_leaf_6_clk picorv32_pcpi_mul_inst_0.mul_waiting vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_81_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput25 pcpi_rs1[15] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 pcpi_rs1[25] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput14 pcpi_insn[3] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput47 pcpi_rs1[6] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput69 pcpi_rs2[26] net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput58 pcpi_rs2[16] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2410_ _0754_ _0758_ _0759_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1655__I _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2341_ _0694_ _0697_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2272_ _0632_ _0634_ _0635_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2486__I _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2477__A1 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2229__A1 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1987_ _0378_ _0372_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2608_ _0892_ picorv32_pcpi_mul_inst_0.next_rs1\[35\] _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2539_ _0854_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_86_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input33_I pcpi_rs1[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2468__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2459__A1 _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1910_ picorv32_pcpi_mul_inst_0.next_rs2\[9\] _1424_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2890_ _0009_ clknet_leaf_3_clk picorv32_pcpi_mul_inst_0.mul_counter\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1841_ _1147_ _1433_ _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1772_ _1358_ picorv32_pcpi_mul_inst_0.next_rs2\[60\] _1373_ _1374_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2324_ _0678_ _0681_ _0682_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2255_ _0282_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2186_ _0555_ _0556_ _0553_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_54_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2040_ picorv32_pcpi_mul_inst_0.next_rs2\[23\] _0320_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2942_ _0059_ clknet_leaf_26_clk picorv32_pcpi_mul_inst_0.next_rs2\[49\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2873_ _1105_ _1098_ _1106_ _1107_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1824_ _1415_ _1417_ _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1755_ _1325_ _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1686_ _1287_ picorv32_pcpi_mul_inst_0.next_rs2\[44\] _1303_ _1304_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2307_ picorv32_pcpi_mul_inst_0.rd\[48\] _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2238_ picorv32_pcpi_mul_inst_0.next_rs2\[42\] _0527_ picorv32_pcpi_mul_inst_0.rd\[41\]
+ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_68_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2169_ _0535_ _0540_ _0542_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1582__A1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1753__I _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1540_ _1183_ _1193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2759__I _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1471_ _1139_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3072_ _0189_ clknet_leaf_7_clk picorv32_pcpi_mul_inst_0.next_rs1\[31\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2023_ _0302_ _0410_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2925_ _0042_ clknet_leaf_6_clk picorv32_pcpi_mul_inst_0.next_rs2\[32\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2856_ picorv32_pcpi_mul_inst_0.rd\[27\] _1083_ _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1807_ _1401_ _1402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2787_ net88 _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2356__A3 _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1738_ _1346_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1669_ _1283_ picorv32_pcpi_mul_inst_0.next_rs2\[40\] _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2816__A1 picorv32_pcpi_mul_inst_0.rd\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1748__I _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_17_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2710_ _0888_ picorv32_pcpi_mul_inst_0.next_rs1\[62\] _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2641_ _1241_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_10_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2572_ _0875_ picorv32_pcpi_mul_inst_0.next_rs1\[23\] picorv32_pcpi_mul_inst_0.next_rs1\[24\]
+ _0873_ _0870_ net35 _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XANTENNA__2338__A3 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1523_ _1180_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1454_ _1124_ net18 net1 net5 _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_10_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3124_ _0241_ clknet_leaf_30_clk net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3055_ _0172_ clknet_leaf_0_clk picorv32_pcpi_mul_inst_0.next_rs1\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_47_clk clknet_2_0__leaf_clk clknet_leaf_47_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2006_ _0393_ _0395_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2908_ _0025_ clknet_leaf_39_clk picorv32_pcpi_mul_inst_0.next_rs2\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2839_ _1077_ _1066_ _1078_ _1080_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input63_I pcpi_rs2[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2329__A3 _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_38_clk clknet_2_1__leaf_clk clknet_leaf_38_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_84_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2862__I _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2017__A2 picorv32_pcpi_mul_inst_0.rd\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1478__I _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1528__B2 picorv32_pcpi_mul_inst_0.next_rs2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1528__A1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2258__B picorv32_pcpi_mul_inst_0.rd\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_29_clk clknet_2_3__leaf_clk clknet_leaf_29_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2008__A2 picorv32_pcpi_mul_inst_0.rd\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2624_ _0909_ _0910_ _0911_ _0912_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput113 net113 pcpi_mul_rd[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1519__A1 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput102 net102 pcpi_mul_rd[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2555_ _0861_ picorv32_pcpi_mul_inst_0.next_rs1\[17\] picorv32_pcpi_mul_inst_0.next_rs1\[18\]
+ _0859_ _0863_ net28 _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_2486_ _1141_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1506_ _1167_ _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3107_ _0224_ clknet_leaf_44_clk net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2168__B _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3038_ _0155_ clknet_leaf_19_clk picorv32_pcpi_mul_inst_0.rdx\[60\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2247__A2 _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2183__A1 _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2857__I _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2238__A2 _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput26 pcpi_rs1[16] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput37 pcpi_rs1[26] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput15 pcpi_insn[4] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 pcpi_rs1[7] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput59 pcpi_rs2[17] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2340_ _0695_ _0696_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2271_ _0598_ _0629_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1986_ _0305_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_9_clk clknet_2_2__leaf_clk clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2607_ _1394_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2538_ _0853_ picorv32_pcpi_mul_inst_0.next_rs1\[11\] picorv32_pcpi_mul_inst_0.next_rs1\[12\]
+ _0851_ _0848_ net22 _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2469_ _0400_ _0403_ _0401_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input26_I pcpi_rs1[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2361__B _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1600__C2 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_7_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1840_ _1429_ _1431_ _1433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1771_ _1367_ _1360_ _1372_ _1373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1666__I _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2323_ _0678_ _0681_ _0645_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2254_ _0611_ _0615_ _0612_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2185_ _0553_ _0555_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1969_ _0360_ _0361_ _0362_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2200__I picorv32_pcpi_mul_inst_0.rd\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2870__I net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1486__I _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_89_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2941_ _0058_ clknet_leaf_22_clk picorv32_pcpi_mul_inst_0.next_rs2\[48\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2780__I _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2872_ picorv32_pcpi_mul_inst_0.rd\[62\] _1095_ _0979_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1823_ _1172_ _1404_ _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1754_ picorv32_pcpi_mul_inst_0.next_rs2\[57\] _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1685_ _1296_ _1289_ _1302_ _1303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2306_ picorv32_pcpi_mul_inst_0.rdx\[48\] _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2237_ picorv32_pcpi_mul_inst_0.rd\[41\] picorv32_pcpi_mul_inst_0.next_rs2\[42\]
+ _0525_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2168_ _0535_ _0540_ _0541_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2099_ _0478_ picorv32_pcpi_mul_inst_0.rdx\[28\] _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_0_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_59_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2770__A1 picorv32_pcpi_mul_inst_0.rd\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1470_ _1138_ _1117_ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2775__I _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3071_ _0188_ clknet_leaf_6_clk picorv32_pcpi_mul_inst_0.next_rs1\[30\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2022_ _1217_ _0375_ _0408_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2924_ _0041_ clknet_leaf_43_clk picorv32_pcpi_mul_inst_0.next_rs2\[31\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2855_ net103 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_13_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1806_ picorv32_pcpi_mul_inst_0.rs1\[0\] _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2786_ _1032_ _1033_ _1036_ _1038_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2761__A1 _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1737_ _1341_ _1342_ _1345_ _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1668_ _1252_ _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1599_ _1224_ _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2640_ picorv32_pcpi_mul_inst_0.next_rs1\[43\] _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2571_ _1260_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1522_ _1179_ picorv32_pcpi_mul_inst_0.next_rs2\[4\] _1175_ picorv32_pcpi_mul_inst_0.next_rs2\[3\]
+ _1176_ net76 _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XANTENNA__2743__A1 _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1453_ _1117_ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3123_ _0240_ clknet_leaf_30_clk net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3054_ _0171_ clknet_leaf_0_clk picorv32_pcpi_mul_inst_0.next_rs1\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2005_ picorv32_pcpi_mul_inst_0.rd\[18\] _0394_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1482__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2907_ _0024_ clknet_leaf_41_clk picorv32_pcpi_mul_inst_0.next_rs2\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2838_ picorv32_pcpi_mul_inst_0.rd\[55\] _1079_ _1069_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2769_ net85 _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input56_I pcpi_rs2[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2498__B1 _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2256__A3 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_25_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2623_ _0903_ picorv32_pcpi_mul_inst_0.next_rs1\[39\] _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2554_ _0864_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput114 net114 pcpi_mul_rd[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput103 net103 pcpi_mul_rd[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1505_ _1166_ _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2485_ _0816_ _0588_ _0813_ _0819_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_37_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3106_ _0223_ clknet_leaf_5_clk net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3037_ _0154_ clknet_leaf_31_clk picorv32_pcpi_mul_inst_0.rdx\[56\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_43_Left_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_2_0__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_16_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_52_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_89_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_61_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_72_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput27 pcpi_rs1[17] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput16 pcpi_insn[5] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput49 pcpi_rs1[8] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput38 pcpi_rs1[27] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_70_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2174__A2 _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2270_ _0595_ _0633_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1985_ _0302_ _0376_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2606_ picorv32_pcpi_mul_inst_0.next_rs1\[34\] _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2537_ _0845_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1862__I _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2468_ _0803_ _0806_ _0808_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2399_ _0746_ _0749_ _0645_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input19_I pcpi_rs1[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output87_I net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1903__A2 _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1770_ _1371_ picorv32_pcpi_mul_inst_0.next_rs2\[59\] _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1615__C _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2322_ _0679_ _0680_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_33_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2253_ _0618_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2184_ picorv32_pcpi_mul_inst_0.next_rs2\[37\] _0514_ picorv32_pcpi_mul_inst_0.rd\[36\]
+ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1968_ _0344_ picorv32_pcpi_mul_inst_0.rd\[14\] _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2386__A2 _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1899_ picorv32_pcpi_mul_inst_0.rd\[8\] _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2377__A2 _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2940_ _0057_ clknet_leaf_26_clk picorv32_pcpi_mul_inst_0.next_rs2\[47\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2871_ picorv32_pcpi_mul_inst_0.rd\[30\] _1099_ _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1822_ _1414_ _1415_ _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1753_ _1305_ _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1684_ _1301_ picorv32_pcpi_mul_inst_0.next_rs2\[43\] _1302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2305_ _0663_ _0664_ _0665_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2236_ _0588_ _0593_ _0602_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_45_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2167_ _0474_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2098_ picorv32_pcpi_mul_inst_0.rd\[28\] _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1587__I _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3070_ _0187_ clknet_leaf_3_clk picorv32_pcpi_mul_inst_0.next_rs1\[29\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2021_ _1217_ _0338_ _0408_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2923_ _0040_ clknet_leaf_43_clk picorv32_pcpi_mul_inst_0.next_rs2\[30\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2854_ _1090_ _1082_ _1091_ _1092_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_13_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1805_ _1397_ _1159_ _1400_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2785_ _0629_ _1030_ _1037_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1736_ _1333_ _1343_ _1344_ _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1667_ picorv32_pcpi_mul_inst_0.next_rs2\[41\] _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1598_ _1232_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2219_ _0585_ _0586_ _0587_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2201__A1 _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2570_ _0874_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1521_ _1136_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1452_ net15 net16 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3122_ _0239_ clknet_leaf_36_clk net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_78_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3053_ _0170_ clknet_leaf_0_clk picorv32_pcpi_mul_inst_0.next_rs1\[12\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2004_ picorv32_pcpi_mul_inst_0.next_rs2\[19\] _0320_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2906_ _0023_ clknet_leaf_41_clk picorv32_pcpi_mul_inst_0.next_rs2\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2837_ _1029_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2768_ _1021_ _1016_ _1022_ _1023_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2699_ picorv32_pcpi_mul_inst_0.next_rs1\[58\] _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1719_ _1315_ _1326_ _1330_ _1331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input49_I pcpi_rs1[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2498__A1 _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1473__A2 _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2380__B _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2622_ _1394_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2553_ _0861_ picorv32_pcpi_mul_inst_0.next_rs1\[16\] picorv32_pcpi_mul_inst_0.next_rs1\[17\]
+ _0859_ _0863_ net27 _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput115 net115 pcpi_mul_rd[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput104 net104 pcpi_mul_rd[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1504_ net83 _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2484_ _0581_ _0584_ _0582_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3105_ _0222_ clknet_leaf_6_clk net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3036_ _0153_ clknet_leaf_29_clk picorv32_pcpi_mul_inst_0.rdx\[52\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2183__A3 _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput28 pcpi_rs1[18] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput17 pcpi_insn[6] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput39 pcpi_rs1[28] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1984_ _1208_ _0375_ _0373_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_82_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2605_ _0885_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2536_ _0852_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2467_ _0807_ picorv32_pcpi_mul_inst_0.rdx\[16\] _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2398_ _0747_ _0748_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3019_ _0136_ clknet_leaf_31_clk picorv32_pcpi_mul_inst_0.rd\[59\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2147__A3 _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2321_ picorv32_pcpi_mul_inst_0.next_rs2\[50\] _0642_ picorv32_pcpi_mul_inst_0.rd\[49\]
+ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2252_ _0610_ _0617_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_leaf_15_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2183_ _0554_ _1270_ _1405_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_26_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _0357_ _0359_ _0335_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1898_ _0296_ _0297_ _0298_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2519_ _0841_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input31_I pcpi_rs1[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output118_I net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1812__A2 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2870_ net107 _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1821_ picorv32_pcpi_mul_inst_0.rd\[1\] _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_10_clk clknet_2_2__leaf_clk clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1752_ _1357_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1683_ _1300_ _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2304_ _0598_ picorv32_pcpi_mul_inst_0.rd\[47\] _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2235_ _0589_ _1288_ _0601_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2166_ _0537_ _0539_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2097_ _0473_ _0476_ _0477_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_51_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2999_ _0116_ clknet_leaf_15_clk picorv32_pcpi_mul_inst_0.rd\[39\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_71_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input79_I pcpi_rs2[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2020_ _0407_ picorv32_pcpi_mul_inst_0.rdx\[20\] _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1688__I _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2922_ _0039_ clknet_leaf_43_clk picorv32_pcpi_mul_inst_0.next_rs2\[29\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2853_ picorv32_pcpi_mul_inst_0.rd\[58\] _1079_ _1085_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1804_ _1399_ picorv32_pcpi_mul_inst_0.next_rs2\[1\] _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2784_ _0985_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1735_ _1337_ picorv32_pcpi_mul_inst_0.next_rs2\[52\] _1344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1666_ _1168_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1597_ _1225_ picorv32_pcpi_mul_inst_0.next_rs2\[27\] _1230_ picorv32_pcpi_mul_inst_0.next_rs2\[26\]
+ _1228_ net69 _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2218_ _0519_ picorv32_pcpi_mul_inst_0.rd\[39\] _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2149_ _1401_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2222__I _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_70_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1520_ _1178_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1451_ net2 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3121_ _0238_ clknet_leaf_35_clk net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_2_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3052_ _0169_ clknet_leaf_0_clk picorv32_pcpi_mul_inst_0.next_rs1\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2003_ _0384_ _0386_ _0392_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_18_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2905_ _0022_ clknet_leaf_41_clk picorv32_pcpi_mul_inst_0.next_rs2\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2836_ picorv32_pcpi_mul_inst_0.rd\[23\] _1067_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2767_ picorv32_pcpi_mul_inst_0.rd\[41\] _1013_ _1019_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2698_ _0932_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1718_ _1319_ _1324_ _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1649_ _1269_ _1270_ _1273_ _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_84_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2621_ picorv32_pcpi_mul_inst_0.next_rs1\[38\] _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2552_ _0839_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xoutput116 net116 pcpi_mul_ready vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput105 net105 pcpi_mul_rd[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_50_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1924__A1 picorv32_pcpi_mul_inst_0.rd\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1503_ picorv32_pcpi_mul_inst_0.mul_counter\[3\] picorv32_pcpi_mul_inst_0.mul_counter\[4\]
+ _1134_ _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2483_ _0816_ _0553_ _0813_ _0818_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3104_ _0221_ clknet_leaf_6_clk net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3035_ _0152_ clknet_leaf_25_clk picorv32_pcpi_mul_inst_0.rdx\[48\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1876__I _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2819_ _1061_ _1050_ _1062_ _1064_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input61_I pcpi_rs2[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput18 pcpi_mul_valid net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput29 pcpi_rs1[19] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1983_ _0290_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_82_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2604_ _0886_ _0896_ _1395_ _0897_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2535_ _0846_ picorv32_pcpi_mul_inst_0.next_rs1\[10\] picorv32_pcpi_mul_inst_0.next_rs1\[11\]
+ _0851_ _0848_ net21 _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2466_ _0673_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2397_ picorv32_pcpi_mul_inst_0.next_rs2\[58\] _0642_ picorv32_pcpi_mul_inst_0.rd\[57\]
+ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3018_ _0135_ clknet_leaf_31_clk picorv32_pcpi_mul_inst_0.rd\[58\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2389__A1 _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2230__I _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_40_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2320_ picorv32_pcpi_mul_inst_0.rd\[49\] picorv32_pcpi_mul_inst_0.next_rs2\[50\]
+ _0640_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2251_ _0611_ _0615_ _0616_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2182_ picorv32_pcpi_mul_inst_0.rd\[36\] _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1966_ _0357_ _0359_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1897_ _0266_ picorv32_pcpi_mul_inst_0.rd\[7\] _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2518_ _0837_ picorv32_pcpi_mul_inst_0.next_rs1\[4\] picorv32_pcpi_mul_inst_0.next_rs1\[5\]
+ _0835_ _0840_ net46 _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_11_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2449_ _0262_ picorv32_pcpi_mul_inst_0.rs2\[63\] _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input24_I pcpi_rs1[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_58_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_67_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1820_ _1398_ _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1751_ _1341_ picorv32_pcpi_mul_inst_0.next_rs2\[56\] _1356_ _1357_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1682_ _1138_ _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_76_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2303_ _0659_ _0662_ _0550_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2234_ _0513_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2165_ _0533_ _0538_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2096_ _0447_ picorv32_pcpi_mul_inst_0.rd\[27\] _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2998_ _0115_ clknet_leaf_15_clk picorv32_pcpi_mul_inst_0.rd\[38\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1949_ _0344_ _0339_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1884__I _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_67_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2047__A3 _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_29_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1730__A2 picorv32_pcpi_mul_inst_0.next_rs2\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2921_ _0038_ clknet_leaf_43_clk picorv32_pcpi_mul_inst_0.next_rs2\[28\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2852_ picorv32_pcpi_mul_inst_0.rd\[26\] _1083_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2783_ _0339_ _1035_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1803_ _1398_ _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2746__A1 picorv32_pcpi_mul_inst_0.rd\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1734_ _1325_ _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1665_ _1286_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1596_ _1231_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2217_ _0581_ _0584_ _0550_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2148_ _0510_ _0515_ _0522_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2079_ picorv32_pcpi_mul_inst_0.next_rs2\[27\] _1439_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1450_ _1120_ net3 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3120_ _0237_ clknet_leaf_35_clk net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_78_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3051_ _0168_ clknet_leaf_49_clk picorv32_pcpi_mul_inst_0.next_rs1\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2002_ _0391_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2904_ _0021_ clknet_leaf_41_clk picorv32_pcpi_mul_inst_0.next_rs2\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2835_ net99 _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2766_ picorv32_pcpi_mul_inst_0.rd\[9\] _1017_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2697_ _0956_ _0965_ _0958_ _0966_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1717_ _1329_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1648_ _1261_ _1271_ _1272_ _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1579_ _1215_ _1217_ _1212_ picorv32_pcpi_mul_inst_0.next_rs2\[20\] _1219_ net63
+ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_67_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1630__A1 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2110__A2 _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1468__B _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2143__I _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2620_ _0885_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2551_ _0862_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput106 net106 pcpi_mul_rd[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1502_ _1159_ _1163_ _1164_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput117 net117 pcpi_mul_wait vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2482_ _0545_ _0548_ _0546_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3103_ _0220_ clknet_leaf_18_clk net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3034_ _0151_ clknet_leaf_20_clk picorv32_pcpi_mul_inst_0.rdx\[44\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2101__A2 _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_12_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2818_ picorv32_pcpi_mul_inst_0.rd\[51\] _1063_ _1053_ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2749_ net112 _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input54_I pcpi_rs2[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Left_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput19 pcpi_rs1[0] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1842__A1 _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1982_ _1208_ _0338_ _0373_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2603_ _0892_ picorv32_pcpi_mul_inst_0.next_rs1\[34\] _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2534_ _0783_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2465_ _0365_ _0368_ _0366_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2396_ picorv32_pcpi_mul_inst_0.rd\[57\] picorv32_pcpi_mul_inst_0.next_rs2\[58\]
+ _0640_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3017_ _0134_ clknet_leaf_31_clk picorv32_pcpi_mul_inst_0.rd\[57\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1597__C2 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2010__A1 picorv32_pcpi_mul_inst_0.rd\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_57_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2001__A1 picorv32_pcpi_mul_inst_0.rd\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2250_ _0611_ _0615_ _0541_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2304__A2 picorv32_pcpi_mul_inst_0.rd\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2181_ picorv32_pcpi_mul_inst_0.rdx\[36\] _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_48_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1965_ picorv32_pcpi_mul_inst_0.rd\[14\] _0358_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1579__B1 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1896_ _0292_ _0295_ _0287_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2517_ _0839_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2448_ _0786_ _0788_ _0792_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2379_ _0728_ _0731_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input17_I pcpi_insn[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output85_I net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2470__A1 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1750_ _1350_ _1343_ _1355_ _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1681_ _1299_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2302_ _0659_ _0662_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input9_I pcpi_insn[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2233_ _1414_ picorv32_pcpi_mul_inst_0.rd\[41\] _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2164_ picorv32_pcpi_mul_inst_0.next_rs2\[35\] _1404_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2095_ _0467_ _0472_ _0475_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2326__I picorv32_pcpi_mul_inst_0.rd\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2997_ _0114_ clknet_leaf_14_clk picorv32_pcpi_mul_inst_0.rd\[37\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2213__A1 picorv32_pcpi_mul_inst_0.rd\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1948_ _0305_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1879_ _0271_ _0274_ _0280_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_43_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2452__A1 _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_3__f_clk clknet_0_clk clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2920_ _0037_ clknet_leaf_34_clk picorv32_pcpi_mul_inst_0.next_rs2\[27\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2851_ net102 _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1802_ _1160_ _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2782_ _1034_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1733_ picorv32_pcpi_mul_inst_0.next_rs2\[53\] _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1664_ _1269_ picorv32_pcpi_mul_inst_0.next_rs2\[40\] _1285_ _1286_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1595_ _1225_ picorv32_pcpi_mul_inst_0.next_rs2\[26\] _1230_ _1227_ _1228_ net68
+ _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2216_ _0581_ _0584_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2147_ _0511_ _1248_ _1411_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2078_ _0452_ _0454_ _0459_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_88_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_2_3__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3050_ _0167_ clknet_leaf_1_clk picorv32_pcpi_mul_inst_0.next_rs1\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2001_ picorv32_pcpi_mul_inst_0.rd\[17\] picorv32_pcpi_mul_inst_0.next_rs2\[18\]
+ _0278_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_26_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2903_ _0020_ clknet_leaf_41_clk picorv32_pcpi_mul_inst_0.next_rs2\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2834_ _1074_ _1066_ _1075_ _1076_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2765_ net115 _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2696_ _0961_ picorv32_pcpi_mul_inst_0.next_rs1\[58\] _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1716_ _1323_ _1324_ _1328_ _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1647_ _1265_ picorv32_pcpi_mul_inst_0.next_rs2\[36\] _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1578_ _1218_ _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_28_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2550_ _0861_ picorv32_pcpi_mul_inst_0.next_rs1\[15\] picorv32_pcpi_mul_inst_0.next_rs1\[16\]
+ _0859_ _0855_ net26 _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_50_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput107 net107 pcpi_mul_rd[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1501_ picorv32_pcpi_mul_inst_0.mul_counter\[3\] _1161_ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xoutput118 net118 pcpi_mul_wr vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2481_ _0816_ _0510_ _0813_ _0817_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_37_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3102_ _0219_ clknet_leaf_10_clk picorv32_pcpi_mul_inst_0.next_rs1\[61\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3033_ _0150_ clknet_leaf_21_clk picorv32_pcpi_mul_inst_0.rdx\[40\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1860__A2 _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2817_ _1029_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2748_ _1005_ _1000_ _1006_ _1007_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2679_ _0945_ _0952_ _0947_ _0953_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input47_I pcpi_rs1[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2876__A1 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1981_ _0372_ picorv32_pcpi_mul_inst_0.rdx\[16\] _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_clk clknet_2_1__leaf_clk clknet_leaf_40_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2602_ picorv32_pcpi_mul_inst_0.next_rs1\[33\] _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2533_ _0850_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2464_ _0803_ _0804_ _0805_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2395_ _0735_ _0738_ _0745_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3016_ _0133_ clknet_leaf_31_clk picorv32_pcpi_mul_inst_0.rd\[56\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_31_clk clknet_2_3__leaf_clk clknet_leaf_31_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2013__B picorv32_pcpi_mul_inst_0.rd\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_22_clk clknet_2_3__leaf_clk clknet_leaf_22_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_40_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2180_ _0549_ _0551_ _0552_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2149__I _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2593__B _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1579__A1 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1964_ picorv32_pcpi_mul_inst_0.next_rs2\[15\] _0320_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_13_clk clknet_2_2__leaf_clk clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1895_ _0292_ _0295_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2516_ _1157_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2447_ picorv32_pcpi_mul_inst_0.rd\[62\] picorv32_pcpi_mul_inst_0.next_rs2\[63\]
+ _1411_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2378_ _0729_ _0730_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2231__A2 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2522__I _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1680_ _1287_ picorv32_pcpi_mul_inst_0.next_rs2\[43\] _1298_ _1299_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1981__A1 _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2301_ _0660_ _0661_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2232_ _0594_ _0597_ _0599_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2163_ picorv32_pcpi_mul_inst_0.rd\[34\] picorv32_pcpi_mul_inst_0.next_rs2\[35\]
+ _0536_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2094_ _0474_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1511__I _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2996_ _0113_ clknet_leaf_16_clk picorv32_pcpi_mul_inst_0.rd\[36\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1947_ _0302_ _0342_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2342__I _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1878_ _0279_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output116_I net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2850_ _1087_ _1082_ _1088_ _1089_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1801_ net51 _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2781_ _0981_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1732_ _1305_ _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1663_ _1279_ _1271_ _1284_ _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_40_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1594_ _1211_ _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1506__I _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2215_ _0582_ _0583_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2146_ _1414_ picorv32_pcpi_mul_inst_0.rd\[33\] _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2077_ _0458_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2979_ _0096_ clknet_leaf_38_clk picorv32_pcpi_mul_inst_0.rd\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input77_I pcpi_rs2[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2000_ _0387_ _0389_ _0390_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_18_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2902_ _0019_ clknet_leaf_48_clk picorv32_pcpi_mul_inst_0.next_rs2\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2833_ picorv32_pcpi_mul_inst_0.rd\[54\] _1063_ _1069_ _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2764_ _1015_ _1016_ _1018_ _1020_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1715_ _1315_ _1326_ _1327_ _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2695_ picorv32_pcpi_mul_inst_0.next_rs1\[57\] _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1646_ _1252_ _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1577_ _1182_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2352__A1 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2129_ _0504_ _0505_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_68_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_24_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2582__A1 _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1500_ picorv32_pcpi_mul_inst_0.mul_counter\[3\] _1161_ _1163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2480_ _0503_ _0506_ _0504_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xoutput108 net108 pcpi_mul_rd[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput90 net90 pcpi_mul_rd[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_3101_ _0218_ clknet_leaf_10_clk picorv32_pcpi_mul_inst_0.next_rs1\[60\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3032_ _0149_ clknet_leaf_16_clk picorv32_pcpi_mul_inst_0.rdx\[36\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2816_ picorv32_pcpi_mul_inst_0.rd\[19\] _1051_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2747_ picorv32_pcpi_mul_inst_0.rd\[37\] _0996_ _1003_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2678_ _0950_ picorv32_pcpi_mul_inst_0.next_rs1\[53\] _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1629_ _1243_ _1248_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_89_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2525__I _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1980_ picorv32_pcpi_mul_inst_0.rd\[16\] _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_12_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2601_ _0886_ _0894_ _1395_ _0895_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2532_ _0846_ picorv32_pcpi_mul_inst_0.next_rs1\[9\] picorv32_pcpi_mul_inst_0.next_rs1\[10\]
+ _0843_ _0848_ net20 _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2463_ _0796_ picorv32_pcpi_mul_inst_0.rdx\[12\] _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_27_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2394_ _0736_ _1359_ _0527_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3015_ _0132_ clknet_leaf_30_clk picorv32_pcpi_mul_inst_0.rd\[55\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1818__B1 _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2491__B1 _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2010__A3 _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2255__I _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2785__A1 _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2001__A3 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ _0349_ _0351_ _0356_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_31_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1894_ _0293_ _0294_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2515_ _0838_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2446_ _0789_ _0790_ _0791_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2377_ picorv32_pcpi_mul_inst_0.next_rs2\[56\] _0622_ picorv32_pcpi_mul_inst_0.rd\[55\]
+ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2767__A1 picorv32_pcpi_mul_inst_0.rd\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Left_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_27_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2300_ picorv32_pcpi_mul_inst_0.next_rs2\[48\] _0622_ picorv32_pcpi_mul_inst_0.rd\[47\]
+ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2231_ _0598_ _0589_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1497__A1 _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2162_ _0514_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2093_ _1145_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2995_ _0112_ clknet_leaf_21_clk picorv32_pcpi_mul_inst_0.rd\[35\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1946_ _1200_ _0263_ _0340_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_71_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2213__A3 _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1877_ picorv32_pcpi_mul_inst_0.rd\[5\] picorv32_pcpi_mul_inst_0.next_rs2\[6\] _0278_
+ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_43_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2429_ _0773_ _0775_ _0776_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input22_I pcpi_rs1[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output109_I net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1800_ _1395_ _1396_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2780_ _0999_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1731_ _1340_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1662_ _1283_ picorv32_pcpi_mul_inst_0.next_rs2\[39\] _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1593_ _1229_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2214_ picorv32_pcpi_mul_inst_0.next_rs2\[40\] _0470_ picorv32_pcpi_mul_inst_0.rd\[39\]
+ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2145_ _0516_ _0518_ _0520_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1890__A1 picorv32_pcpi_mul_inst_0.rd\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2076_ picorv32_pcpi_mul_inst_0.rd\[25\] picorv32_pcpi_mul_inst_0.next_rs2\[26\]
+ _1427_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_64_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2978_ _0095_ clknet_leaf_38_clk picorv32_pcpi_mul_inst_0.rd\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1929_ picorv32_pcpi_mul_inst_0.rd\[10\] picorv32_pcpi_mul_inst_0.next_rs2\[11\]
+ _0290_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1945__A2 _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_78_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2901_ _0018_ clknet_leaf_48_clk picorv32_pcpi_mul_inst_0.next_rs2\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2832_ picorv32_pcpi_mul_inst_0.rd\[22\] _1067_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2763_ _0589_ _1013_ _1019_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1927__A2 picorv32_pcpi_mul_inst_0.rd\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1714_ _1319_ picorv32_pcpi_mul_inst_0.next_rs2\[48\] _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2694_ _0956_ _0963_ _0958_ _0964_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1645_ picorv32_pcpi_mul_inst_0.next_rs2\[37\] _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1576_ picorv32_pcpi_mul_inst_0.next_rs2\[21\] _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1458__A4 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2128_ picorv32_pcpi_mul_inst_0.next_rs2\[32\] _0470_ picorv32_pcpi_mul_inst_0.rd\[31\]
+ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2059_ _1408_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput109 net109 pcpi_mul_rd[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput91 net91 pcpi_mul_rd[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_3100_ _0217_ clknet_leaf_8_clk picorv32_pcpi_mul_inst_0.next_rs1\[59\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3031_ _0148_ clknet_leaf_16_clk picorv32_pcpi_mul_inst_0.rdx\[32\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2270__A1 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2815_ net94 _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2746_ picorv32_pcpi_mul_inst_0.rd\[5\] _1001_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2677_ picorv32_pcpi_mul_inst_0.next_rs1\[52\] _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1628_ _1256_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1559_ _1205_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1710__I _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1620__I _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2451__I _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2600_ _0892_ picorv32_pcpi_mul_inst_0.next_rs1\[33\] _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2531_ _0849_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2462_ _0327_ _0333_ _0329_ _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2393_ _0636_ picorv32_pcpi_mul_inst_0.rd\[57\] _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1818__A1 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3014_ _0131_ clknet_leaf_28_clk picorv32_pcpi_mul_inst_0.rd\[54\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1530__I _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2491__A1 _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2626__I _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2729_ picorv32_pcpi_mul_inst_0.rd\[2\] _0983_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input52_I pcpi_rs2[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1705__I _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_40_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2473__A1 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1962_ _0355_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_31_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1893_ picorv32_pcpi_mul_inst_0.next_rs2\[8\] _1437_ picorv32_pcpi_mul_inst_0.rd\[7\]
+ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2514_ _0837_ picorv32_pcpi_mul_inst_0.next_rs1\[3\] picorv32_pcpi_mul_inst_0.next_rs1\[4\]
+ _0835_ _0832_ net45 _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_11_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1525__I _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2445_ _0742_ picorv32_pcpi_mul_inst_0.rd\[62\] _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2376_ picorv32_pcpi_mul_inst_0.rd\[55\] picorv32_pcpi_mul_inst_0.next_rs2\[56\]
+ _0620_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2464__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_11_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_26_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2230_ _0446_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2161_ _0523_ _0529_ _0526_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2092_ _0467_ _0472_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2994_ _0111_ clknet_leaf_14_clk picorv32_pcpi_mul_inst_0.rd\[34\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1945_ _1200_ _0338_ _0340_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1876_ _1426_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2428_ _0742_ _0770_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1488__A2 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2359_ picorv32_pcpi_mul_inst_0.next_rs2\[54\] _0642_ picorv32_pcpi_mul_inst_0.rd\[53\]
+ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input15_I pcpi_insn[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2724__I net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1730_ _1323_ picorv32_pcpi_mul_inst_0.next_rs2\[52\] _1339_ _1340_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1661_ _1242_ _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1592_ _1225_ _1227_ _1221_ picorv32_pcpi_mul_inst_0.next_rs2\[24\] _1228_ net67
+ _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_0_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1803__I _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I pcpi_insn[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2213_ picorv32_pcpi_mul_inst_0.rd\[39\] picorv32_pcpi_mul_inst_0.next_rs2\[40\]
+ _0468_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2144_ _0519_ _0511_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2075_ _0455_ _0456_ _0457_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_64_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2977_ _0094_ clknet_leaf_38_clk picorv32_pcpi_mul_inst_0.rd\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1928_ _0323_ _0324_ _0325_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1859_ _0262_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_55_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1881__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_64_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_73_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1623__I _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_82_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2900_ _0017_ clknet_leaf_48_clk picorv32_pcpi_mul_inst_0.next_rs2\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2831_ net98 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2762_ _0985_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1713_ _1325_ _1326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_91_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2693_ _0961_ picorv32_pcpi_mul_inst_0.next_rs1\[57\] _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1644_ _1168_ _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1575_ _1216_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2127_ picorv32_pcpi_mul_inst_0.rd\[31\] picorv32_pcpi_mul_inst_0.next_rs2\[32\]
+ _0468_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2058_ _1227_ _0338_ _0441_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2812__A1 picorv32_pcpi_mul_inst_0.rd\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1615__A2 picorv32_pcpi_mul_inst_0.next_rs2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input82_I pcpi_rs2[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2040__A2 _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2500__B1 _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2803__A1 _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2031__A2 _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1618__I _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput92 net92 pcpi_mul_rd[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3030_ _0147_ clknet_leaf_44_clk picorv32_pcpi_mul_inst_0.rdx\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_43_clk clknet_2_1__leaf_clk clknet_leaf_43_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2814_ _1058_ _1050_ _1059_ _1060_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2022__A2 _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2745_ net111 _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2676_ _0945_ _0949_ _0947_ _0951_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1627_ _1247_ _1248_ _1255_ _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1533__A1 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1558_ _1198_ picorv32_pcpi_mul_inst_0.next_rs2\[15\] _1203_ picorv32_pcpi_mul_inst_0.next_rs2\[14\]
+ _1201_ net56 _1205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1489_ picorv32_pcpi_mul_inst_0.mul_counter\[0\] _1151_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2094__I _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_34_clk clknet_2_1__leaf_clk clknet_leaf_34_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_20_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2013__A2 _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_25_clk clknet_2_3__leaf_clk clknet_leaf_25_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2732__I net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2004__A2 _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2530_ _0846_ picorv32_pcpi_mul_inst_0.next_rs1\[8\] picorv32_pcpi_mul_inst_0.next_rs1\[9\]
+ _0843_ _0848_ net50 _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_23_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2461_ _1238_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2392_ _0739_ _0741_ _0743_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3013_ _0130_ clknet_leaf_29_clk picorv32_pcpi_mul_inst_0.rd\[53\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1811__I _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_16_clk clknet_2_2__leaf_clk clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_34_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2728_ net106 _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2659_ _0925_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input45_I pcpi_rs1[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2089__I _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1961_ picorv32_pcpi_mul_inst_0.rd\[13\] picorv32_pcpi_mul_inst_0.next_rs2\[14\]
+ _0278_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_31_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2225__A2 _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1892_ picorv32_pcpi_mul_inst_0.rd\[7\] picorv32_pcpi_mul_inst_0.next_rs2\[8\] _0262_
+ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2513_ _1224_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_5_clk clknet_2_0__leaf_clk clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2444_ _0786_ _0788_ _0699_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2375_ _0720_ _0724_ _0721_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2321__B picorv32_pcpi_mul_inst_0.rd\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1451__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2160_ _0532_ _0533_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2091_ _0469_ _0471_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2993_ _0110_ clknet_leaf_6_clk picorv32_pcpi_mul_inst_0.rd\[33\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1944_ _0339_ picorv32_pcpi_mul_inst_0.rdx\[12\] _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1875_ _0275_ _0276_ _0277_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2427_ _1409_ _0774_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2358_ picorv32_pcpi_mul_inst_0.rd\[53\] picorv32_pcpi_mul_inst_0.next_rs2\[54\]
+ _0640_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2289_ _0514_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_67_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1660_ _1282_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1591_ _1218_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2212_ _0572_ _0577_ _0573_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2143_ _0446_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1890__A3 _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2074_ _0447_ picorv32_pcpi_mul_inst_0.rd\[25\] _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2976_ _0093_ clknet_leaf_39_clk picorv32_pcpi_mul_inst_0.rd\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1927_ _0306_ picorv32_pcpi_mul_inst_0.rd\[10\] _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1858_ _1439_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_10_clk_I clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2355__A1 _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1789_ _1387_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_25_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output114_I net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2830_ _1071_ _1066_ _1072_ _1073_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2761_ _0299_ _1017_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2692_ picorv32_pcpi_mul_inst_0.next_rs1\[56\] _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1712_ _1251_ _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1643_ _1268_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1574_ _1215_ picorv32_pcpi_mul_inst_0.next_rs2\[20\] _1212_ picorv32_pcpi_mul_inst_0.next_rs2\[19\]
+ _1209_ net61 _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XTAP_TAPCELL_ROW_1_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2126_ _0496_ _0498_ _0502_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2057_ _0440_ picorv32_pcpi_mul_inst_0.rdx\[24\] _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2959_ _0076_ clknet_leaf_4_clk picorv32_pcpi_mul_inst_0.next_rs2\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input75_I pcpi_rs2[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1634__I _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput93 net93 pcpi_mul_rd[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2813_ picorv32_pcpi_mul_inst_0.rd\[50\] _1047_ _1053_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2744_ _0998_ _1000_ _1002_ _1004_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2675_ _0950_ picorv32_pcpi_mul_inst_0.next_rs1\[52\] _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1626_ _1250_ _1253_ _1254_ _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_78_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1557_ _1204_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1488_ picorv32_pcpi_mul_inst_0.mul_counter\[0\] _1150_ _1153_ _0006_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2109_ _0485_ _0486_ _0487_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_68_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3089_ _0206_ clknet_leaf_11_clk picorv32_pcpi_mul_inst_0.next_rs1\[48\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2485__B1 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2788__A1 picorv32_pcpi_mul_inst_0.rd\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2460_ _1150_ _0801_ _0802_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2391_ _0742_ _0736_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3012_ _0129_ clknet_leaf_29_clk picorv32_pcpi_mul_inst_0.rd\[52\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2409__B _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2727_ _0988_ _0980_ _0989_ _0990_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2658_ picorv32_pcpi_mul_inst_0.next_rs1\[47\] _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1609_ _1233_ picorv32_pcpi_mul_inst_0.next_rs2\[31\] _1238_ picorv32_pcpi_mul_inst_0.next_rs2\[30\]
+ _1236_ net74 _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2589_ _0885_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input38_I pcpi_rs1[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1960_ _0352_ _0353_ _0354_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_31_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1891_ _0281_ _0284_ _0291_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1984__A2 _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2512_ _0836_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2443_ _0786_ _0788_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2374_ _0727_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1732__I _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2563__I _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2090_ picorv32_pcpi_mul_inst_0.next_rs2\[28\] _0470_ picorv32_pcpi_mul_inst_0.rd\[27\]
+ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2992_ _0109_ clknet_leaf_17_clk picorv32_pcpi_mul_inst_0.rd\[32\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1943_ picorv32_pcpi_mul_inst_0.rd\[12\] _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1874_ _0266_ picorv32_pcpi_mul_inst_0.rd\[5\] _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2426_ _0771_ _0772_ _0769_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1552__I _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2357_ _0702_ _0705_ _0711_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2288_ _0639_ _0644_ _0641_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_67_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1727__I _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2125__A2 picorv32_pcpi_mul_inst_0.next_rs2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2061__A1 _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1590_ picorv32_pcpi_mul_inst_0.next_rs2\[25\] _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2211_ _0580_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2142_ _0443_ _0517_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2073_ _0452_ _0454_ _0429_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_64_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2975_ _0092_ clknet_leaf_40_clk picorv32_pcpi_mul_inst_0.rd\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1926_ _0319_ _0322_ _0287_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1857_ _1181_ _1406_ _0260_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1788_ _1375_ picorv32_pcpi_mul_inst_0.next_rs2\[63\] _1386_ _1387_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2107__A2 _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2409_ _0754_ _0758_ _1146_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input20_I pcpi_rs1[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output107_I net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2760_ _0982_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2691_ _0956_ _0960_ _0958_ _0962_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1711_ picorv32_pcpi_mul_inst_0.next_rs2\[49\] _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1642_ _1247_ picorv32_pcpi_mul_inst_0.next_rs2\[36\] _1267_ _1268_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1573_ _1189_ _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1848__A1 picorv32_pcpi_mul_inst_0.next_rs2\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1830__I _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2125_ picorv32_pcpi_mul_inst_0.rd\[30\] picorv32_pcpi_mul_inst_0.next_rs2\[31\]
+ _0262_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2056_ picorv32_pcpi_mul_inst_0.rd\[24\] _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2958_ _0075_ clknet_leaf_7_clk picorv32_pcpi_mul_inst_0.next_rs1\[62\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1909_ picorv32_pcpi_mul_inst_0.rd\[8\] picorv32_pcpi_mul_inst_0.rdx\[8\] _0308_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2889_ _0008_ clknet_leaf_4_clk picorv32_pcpi_mul_inst_0.mul_counter\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input68_I pcpi_rs2[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2571__I _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput94 net94 pcpi_mul_rd[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2812_ picorv32_pcpi_mul_inst_0.rd\[18\] _1051_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2743_ _0554_ _0996_ _1003_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_39_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2674_ _0925_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1625_ _1243_ picorv32_pcpi_mul_inst_0.next_rs2\[32\] _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1556_ _1198_ picorv32_pcpi_mul_inst_0.next_rs2\[14\] _1203_ _1200_ _1201_ net55
+ _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_1487_ picorv32_pcpi_mul_inst_0.mul_counter\[0\] _1152_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_6_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2108_ _0478_ picorv32_pcpi_mul_inst_0.rdx\[28\] _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_37_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3088_ _0205_ clknet_leaf_10_clk picorv32_pcpi_mul_inst_0.next_rs1\[47\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2039_ _0417_ _0419_ _0424_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2246__A1 picorv32_pcpi_mul_inst_0.rd\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2237__A1 picorv32_pcpi_mul_inst_0.rd\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2250__B _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2390_ _0673_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_79_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3011_ _0128_ clknet_leaf_29_clk picorv32_pcpi_mul_inst_0.rd\[51\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_88_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2726_ picorv32_pcpi_mul_inst_0.rd\[33\] _1115_ _0986_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1555__I _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2657_ _0933_ _0934_ _0936_ _0937_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1608_ _1239_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2588_ _1151_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1539_ picorv32_pcpi_mul_inst_0.next_rs2\[9\] _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2467__A1 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_56_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1890_ picorv32_pcpi_mul_inst_0.rd\[6\] picorv32_pcpi_mul_inst_0.next_rs2\[7\] _0290_
+ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_50_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2511_ _0830_ picorv32_pcpi_mul_inst_0.next_rs1\[2\] picorv32_pcpi_mul_inst_0.next_rs1\[3\]
+ _0835_ _0832_ net44 _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_11_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2442_ picorv32_pcpi_mul_inst_0.rd\[62\] _0787_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2373_ _0719_ _0726_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_75_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2449__A1 _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2155__B _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2709_ picorv32_pcpi_mul_inst_0.next_rs1\[61\] _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input50_I pcpi_rs1[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2991_ _0108_ clknet_leaf_44_clk picorv32_pcpi_mul_inst_0.rd\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1942_ _1405_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_61_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1873_ _0271_ _0274_ _1409_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1833__I _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2425_ _0769_ _0771_ _0772_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2356_ _0703_ _1342_ _0601_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1893__A2 _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2287_ _0569_ _0648_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_67_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2070__A2 _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2125__A3 _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2574__I _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2749__I net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2116__A3 _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2210_ _0571_ _0579_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2141_ _0512_ _0515_ _0510_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2072_ _0452_ _0454_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2974_ _0091_ clknet_leaf_39_clk picorv32_pcpi_mul_inst_0.rd\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1925_ _0319_ _0322_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1856_ _0259_ picorv32_pcpi_mul_inst_0.rdx\[4\] _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_15_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1787_ _1384_ _1377_ _1385_ _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2408_ _0755_ _0757_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_24_Left_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1866__A2 _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2339_ picorv32_pcpi_mul_inst_0.next_rs2\[52\] _0622_ picorv32_pcpi_mul_inst_0.rd\[51\]
+ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input13_I pcpi_insn[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2291__A2 _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2343__B _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Left_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2503__C2 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1857__A2 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1609__A2 picorv32_pcpi_mul_inst_0.next_rs2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1710_ _1305_ _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2690_ _0961_ picorv32_pcpi_mul_inst_0.next_rs1\[56\] _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1641_ _1261_ _1253_ _1266_ _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_34_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1572_ _1214_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_60_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input5_I pcpi_insn[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2124_ _0499_ _0500_ _0501_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_46_clk clknet_2_0__leaf_clk clknet_leaf_46_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2055_ _0437_ _0438_ _0439_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2957_ _0074_ clknet_leaf_18_clk picorv32_pcpi_mul_inst_0.rs2\[63\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1908_ _0301_ _0304_ _0307_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2888_ _0007_ clknet_leaf_4_clk picorv32_pcpi_mul_inst_0.mul_counter\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1839_ _1429_ _1431_ _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1507__B _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_37_clk clknet_2_1__leaf_clk clknet_leaf_37_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput84 net84 pcpi_mul_rd[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput95 net95 pcpi_mul_rd[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1931__I _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_28_clk clknet_2_3__leaf_clk clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2811_ net93 _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2742_ _0985_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2673_ picorv32_pcpi_mul_inst_0.next_rs1\[51\] _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1624_ _1252_ _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1555_ _1174_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2191__A1 _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1486_ _1151_ _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2107_ picorv32_pcpi_mul_inst_0.next_rs2\[29\] _0381_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk clknet_leaf_19_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3087_ _0204_ clknet_leaf_11_clk picorv32_pcpi_mul_inst_0.next_rs1\[46\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2038_ _0423_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_37_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input80_I pcpi_rs2[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2173__A1 picorv32_pcpi_mul_inst_0.rd\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1661__I _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3010_ _0127_ clknet_leaf_27_clk picorv32_pcpi_mul_inst_0.rd\[50\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_42_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2725_ _1415_ _0983_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_8_clk clknet_2_2__leaf_clk clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2656_ _0926_ picorv32_pcpi_mul_inst_0.next_rs1\[47\] _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1607_ _1233_ picorv32_pcpi_mul_inst_0.next_rs2\[30\] _1238_ _1235_ _1236_ net72
+ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
X_2587_ _0884_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1911__A1 _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1538_ _1191_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1469_ picorv32_pcpi_mul_inst_0.mul_waiting _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_23_clk_I clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_38_clk_I clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_31_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2510_ _0783_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2441_ picorv32_pcpi_mul_inst_0.next_rs2\[63\] _0524_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2146__A1 _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2372_ _0720_ _0724_ _0725_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2708_ _0967_ _0973_ _0969_ _0974_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2639_ _0920_ _0921_ _0922_ _0923_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input43_I pcpi_rs1[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2860__I net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1476__I net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2128__A1 picorv32_pcpi_mul_inst_0.next_rs2\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2990_ _0107_ clknet_leaf_44_clk picorv32_pcpi_mul_inst_0.rd\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1941_ _0334_ _0336_ _0337_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1872_ _0271_ _0274_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2119__A1 picorv32_pcpi_mul_inst_0.next_rs2\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2424_ picorv32_pcpi_mul_inst_0.next_rs2\[61\] _1402_ picorv32_pcpi_mul_inst_0.rd\[60\]
+ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2355_ _0636_ picorv32_pcpi_mul_inst_0.rd\[53\] _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2286_ picorv32_pcpi_mul_inst_0.rd\[46\] _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_67_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1934__I _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _0510_ _0512_ _0515_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2071_ picorv32_pcpi_mul_inst_0.rd\[25\] _0453_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2765__I net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2973_ _0090_ clknet_leaf_40_clk picorv32_pcpi_mul_inst_0.rd\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1924_ picorv32_pcpi_mul_inst_0.rd\[10\] _0321_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1855_ picorv32_pcpi_mul_inst_0.rd\[4\] _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_12_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1786_ _1371_ picorv32_pcpi_mul_inst_0.next_rs2\[62\] _1385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2407_ _0752_ _0756_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2338_ picorv32_pcpi_mul_inst_0.rd\[51\] picorv32_pcpi_mul_inst_0.next_rs2\[52\]
+ _0620_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2269_ _0630_ _0631_ _0628_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2751__A1 picorv32_pcpi_mul_inst_0.rd\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1640_ _1265_ picorv32_pcpi_mul_inst_0.next_rs2\[35\] _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1571_ _1206_ picorv32_pcpi_mul_inst_0.next_rs2\[19\] _1212_ picorv32_pcpi_mul_inst_0.next_rs2\[18\]
+ _1209_ net60 _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_67_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2123_ _0483_ picorv32_pcpi_mul_inst_0.rd\[30\] _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_77_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2054_ _0412_ picorv32_pcpi_mul_inst_0.rd\[23\] _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2444__B _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2956_ _0073_ clknet_leaf_18_clk picorv32_pcpi_mul_inst_0.next_rs2\[63\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1907_ _0306_ _0299_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2887_ _0006_ clknet_leaf_4_clk picorv32_pcpi_mul_inst_0.mul_counter\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1838_ picorv32_pcpi_mul_inst_0.rd\[2\] _1430_ _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_32_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1769_ _1241_ _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output112_I net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1484__I _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput85 net85 pcpi_mul_rd[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput96 net96 pcpi_mul_rd[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2488__B1 _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2810_ _1055_ _1050_ _1056_ _1057_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2741_ _0259_ _1001_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2672_ _0945_ _0946_ _0947_ _0948_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1623_ _1251_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1554_ _1202_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1485_ _1144_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
.ends


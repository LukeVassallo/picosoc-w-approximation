* NGSPICE file created from simple_interconnect.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

.subckt simple_interconnect clk gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[1] gpio_in[2] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6]
+ gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[14] gpio_oeb[15] gpio_oeb[2] gpio_oeb[3]
+ gpio_oeb[4] gpio_oeb[5] gpio_oeb[6] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10]
+ gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[1] gpio_out[2]
+ gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9]
+ mem_addr[0] mem_addr[10] mem_addr[11] mem_addr[12] mem_addr[13] mem_addr[14] mem_addr[15]
+ mem_addr[16] mem_addr[17] mem_addr[18] mem_addr[19] mem_addr[1] mem_addr[20] mem_addr[21]
+ mem_addr[22] mem_addr[23] mem_addr[24] mem_addr[25] mem_addr[26] mem_addr[27] mem_addr[28]
+ mem_addr[29] mem_addr[2] mem_addr[30] mem_addr[31] mem_addr[3] mem_addr[4] mem_addr[5]
+ mem_addr[6] mem_addr[7] mem_addr[8] mem_addr[9] mem_instr mem_rdata[0] mem_rdata[10]
+ mem_rdata[11] mem_rdata[12] mem_rdata[13] mem_rdata[14] mem_rdata[15] mem_rdata[16]
+ mem_rdata[17] mem_rdata[18] mem_rdata[19] mem_rdata[1] mem_rdata[20] mem_rdata[21]
+ mem_rdata[22] mem_rdata[23] mem_rdata[24] mem_rdata[25] mem_rdata[26] mem_rdata[27]
+ mem_rdata[28] mem_rdata[29] mem_rdata[2] mem_rdata[30] mem_rdata[31] mem_rdata[3]
+ mem_rdata[4] mem_rdata[5] mem_rdata[6] mem_rdata[7] mem_rdata[8] mem_rdata[9] mem_ready
+ mem_valid mem_wdata[0] mem_wdata[10] mem_wdata[11] mem_wdata[12] mem_wdata[13] mem_wdata[14]
+ mem_wdata[15] mem_wdata[16] mem_wdata[17] mem_wdata[18] mem_wdata[19] mem_wdata[1]
+ mem_wdata[20] mem_wdata[21] mem_wdata[22] mem_wdata[23] mem_wdata[24] mem_wdata[25]
+ mem_wdata[26] mem_wdata[27] mem_wdata[28] mem_wdata[29] mem_wdata[2] mem_wdata[30]
+ mem_wdata[31] mem_wdata[3] mem_wdata[4] mem_wdata[5] mem_wdata[6] mem_wdata[7] mem_wdata[8]
+ mem_wdata[9] mem_wstrb[0] mem_wstrb[1] mem_wstrb[2] mem_wstrb[3] ram_gwenb[0] ram_gwenb[1]
+ ram_gwenb[2] ram_gwenb[3] ram_rdata[0] ram_rdata[10] ram_rdata[11] ram_rdata[12]
+ ram_rdata[13] ram_rdata[14] ram_rdata[15] ram_rdata[16] ram_rdata[17] ram_rdata[18]
+ ram_rdata[19] ram_rdata[1] ram_rdata[20] ram_rdata[21] ram_rdata[22] ram_rdata[23]
+ ram_rdata[24] ram_rdata[25] ram_rdata[26] ram_rdata[27] ram_rdata[28] ram_rdata[29]
+ ram_rdata[2] ram_rdata[30] ram_rdata[31] ram_rdata[3] ram_rdata[4] ram_rdata[5]
+ ram_rdata[6] ram_rdata[7] ram_rdata[8] ram_rdata[9] ram_wenb[0] ram_wenb[10] ram_wenb[11]
+ ram_wenb[12] ram_wenb[13] ram_wenb[14] ram_wenb[15] ram_wenb[16] ram_wenb[17] ram_wenb[18]
+ ram_wenb[19] ram_wenb[1] ram_wenb[20] ram_wenb[21] ram_wenb[22] ram_wenb[23] ram_wenb[24]
+ ram_wenb[25] ram_wenb[26] ram_wenb[27] ram_wenb[28] ram_wenb[29] ram_wenb[2] ram_wenb[30]
+ ram_wenb[31] ram_wenb[3] ram_wenb[4] ram_wenb[5] ram_wenb[6] ram_wenb[7] ram_wenb[8]
+ ram_wenb[9] resetn simpleuart_dat_re simpleuart_dat_we simpleuart_div_we[0] simpleuart_div_we[1]
+ simpleuart_div_we[2] simpleuart_div_we[3] simpleuart_reg_dat_do[0] simpleuart_reg_dat_do[10]
+ simpleuart_reg_dat_do[11] simpleuart_reg_dat_do[12] simpleuart_reg_dat_do[13] simpleuart_reg_dat_do[14]
+ simpleuart_reg_dat_do[15] simpleuart_reg_dat_do[16] simpleuart_reg_dat_do[17] simpleuart_reg_dat_do[18]
+ simpleuart_reg_dat_do[19] simpleuart_reg_dat_do[1] simpleuart_reg_dat_do[20] simpleuart_reg_dat_do[21]
+ simpleuart_reg_dat_do[22] simpleuart_reg_dat_do[23] simpleuart_reg_dat_do[24] simpleuart_reg_dat_do[25]
+ simpleuart_reg_dat_do[26] simpleuart_reg_dat_do[27] simpleuart_reg_dat_do[28] simpleuart_reg_dat_do[29]
+ simpleuart_reg_dat_do[2] simpleuart_reg_dat_do[30] simpleuart_reg_dat_do[31] simpleuart_reg_dat_do[3]
+ simpleuart_reg_dat_do[4] simpleuart_reg_dat_do[5] simpleuart_reg_dat_do[6] simpleuart_reg_dat_do[7]
+ simpleuart_reg_dat_do[8] simpleuart_reg_dat_do[9] simpleuart_reg_dat_wait simpleuart_reg_div_do[0]
+ simpleuart_reg_div_do[10] simpleuart_reg_div_do[11] simpleuart_reg_div_do[12] simpleuart_reg_div_do[13]
+ simpleuart_reg_div_do[14] simpleuart_reg_div_do[15] simpleuart_reg_div_do[16] simpleuart_reg_div_do[17]
+ simpleuart_reg_div_do[18] simpleuart_reg_div_do[19] simpleuart_reg_div_do[1] simpleuart_reg_div_do[20]
+ simpleuart_reg_div_do[21] simpleuart_reg_div_do[22] simpleuart_reg_div_do[23] simpleuart_reg_div_do[24]
+ simpleuart_reg_div_do[25] simpleuart_reg_div_do[26] simpleuart_reg_div_do[27] simpleuart_reg_div_do[28]
+ simpleuart_reg_div_do[29] simpleuart_reg_div_do[2] simpleuart_reg_div_do[30] simpleuart_reg_div_do[31]
+ simpleuart_reg_div_do[3] simpleuart_reg_div_do[4] simpleuart_reg_div_do[5] simpleuart_reg_div_do[6]
+ simpleuart_reg_div_do[7] simpleuart_reg_div_do[8] simpleuart_reg_div_do[9] spimem_rdata[0]
+ spimem_rdata[10] spimem_rdata[11] spimem_rdata[12] spimem_rdata[13] spimem_rdata[14]
+ spimem_rdata[15] spimem_rdata[16] spimem_rdata[17] spimem_rdata[18] spimem_rdata[19]
+ spimem_rdata[1] spimem_rdata[20] spimem_rdata[21] spimem_rdata[22] spimem_rdata[23]
+ spimem_rdata[24] spimem_rdata[25] spimem_rdata[26] spimem_rdata[27] spimem_rdata[28]
+ spimem_rdata[29] spimem_rdata[2] spimem_rdata[30] spimem_rdata[31] spimem_rdata[3]
+ spimem_rdata[4] spimem_rdata[5] spimem_rdata[6] spimem_rdata[7] spimem_rdata[8]
+ spimem_rdata[9] spimem_ready spimem_valid spimemio_cfgreg_do[0] spimemio_cfgreg_do[10]
+ spimemio_cfgreg_do[11] spimemio_cfgreg_do[12] spimemio_cfgreg_do[13] spimemio_cfgreg_do[14]
+ spimemio_cfgreg_do[15] spimemio_cfgreg_do[16] spimemio_cfgreg_do[17] spimemio_cfgreg_do[18]
+ spimemio_cfgreg_do[19] spimemio_cfgreg_do[1] spimemio_cfgreg_do[20] spimemio_cfgreg_do[21]
+ spimemio_cfgreg_do[22] spimemio_cfgreg_do[23] spimemio_cfgreg_do[24] spimemio_cfgreg_do[25]
+ spimemio_cfgreg_do[26] spimemio_cfgreg_do[27] spimemio_cfgreg_do[28] spimemio_cfgreg_do[29]
+ spimemio_cfgreg_do[2] spimemio_cfgreg_do[30] spimemio_cfgreg_do[31] spimemio_cfgreg_do[3]
+ spimemio_cfgreg_do[4] spimemio_cfgreg_do[5] spimemio_cfgreg_do[6] spimemio_cfgreg_do[7]
+ spimemio_cfgreg_do[8] spimemio_cfgreg_do[9] spimemio_cfgreg_we[0] spimemio_cfgreg_we[1]
+ spimemio_cfgreg_we[2] spimemio_cfgreg_we[3] vdd vss gpio_oeb[13] gpio_oeb[1] gpio_oeb[12]
+ gpio_oeb[11] gpio_oeb[0] gpio_oeb[10] gpio_oeb[7]
XFILLER_0_92_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input108_I simpleuart_reg_dat_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input73_I ram_rdata[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output327_I net327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1270_ net243 _0079_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0985_ _0412_ _0438_ _0415_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_3_2__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1468_ net333 net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1399_ _0026_ clknet_3_3__leaf_clk iomem_rdata\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input225_I spimemio_cfgreg_do[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output277_I net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0770_ net125 _0239_ _0197_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1253_ gpio\[31\] _0657_ _0658_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1322_ gpio\[24\] _0111_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1184_ net39 _0606_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0968_ iomem_rdata\[17\] _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input175_I spimem_rdata[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput242 net242 gpio_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput286 net286 ram_wenb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_0899_ _0212_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_30_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput264 net264 mem_rdata[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput253 net253 mem_rdata[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput275 net275 mem_rdata[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput297 net297 ram_wenb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input36_I mem_wdata[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0822_ net164 _0262_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0753_ _0224_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0684_ _0149_ _0153_ _0157_ _0167_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1236_ _0651_ _0652_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1305_ _0423_ _0097_ _0101_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1098_ _0540_ _0542_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_35_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0746__I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1167_ net248 _0596_ _0598_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_49_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1021_ net214 _0446_ _0458_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_32_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0805_ _0226_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0736_ _0166_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0667_ net14 net13 net16 net15 _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input138_I simpleuart_reg_div_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1219_ _0638_ _0639_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1010__I net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1004_ _0404_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0719_ _0149_ _0153_ _0157_ _0165_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_79_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_43_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_91_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput186 spimem_rdata[26] net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput197 spimem_rdata[7] net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput175 spimem_rdata[16] net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput120 simpleuart_reg_dat_do[25] net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput131 simpleuart_reg_dat_do[6] net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_59_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput153 simpleuart_reg_div_do[25] net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput142 simpleuart_reg_div_do[15] net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1160__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput164 simpleuart_reg_div_do[6] net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_14_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1484_ net339 net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1151__A1 _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0717__A1 _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input66_I mem_wstrb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_39_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_48_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0984_ net79 _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_57_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0947__A1 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1467_ net333 net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_66_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1398_ _0025_ clknet_3_6__leaf_clk iomem_rdata\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1372__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input218_I spimemio_cfgreg_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input120_I simpleuart_reg_dat_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1363__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0929__A1 _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1252_ net58 _0655_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1354__A1 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1321_ _0098_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1183_ _0611_ _0612_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0967_ _0400_ _0402_ _0417_ _0422_ net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_6_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput243 net243 gpio_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input168_I spimem_rdata[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput298 net298 ram_wenb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_71_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput287 net287 ram_wenb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0898_ net139 _0357_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput276 net276 mem_rdata[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput265 net265 mem_rdata[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput254 net254 mem_rdata[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1345__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input29_I mem_addr[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_64_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0821_ net131 _0286_ _0249_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0752_ _0219_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0683_ net33 _0158_ _0164_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_10_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1166_ net65 _0592_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1235_ gpio\[26\] _0646_ _0647_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1304_ gpio\[17\] _0099_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1097_ _0507_ _0541_ _0509_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_35_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1020_ net149 _0456_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_32_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0735_ net103 _0180_ _0197_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_40_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0804_ _0224_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0666_ net17 _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_4_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input200_I spimem_ready vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1149_ _0182_ _0000_ net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1218_ gpio\[22\] _0632_ _0634_ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input96_I ram_rdata[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output252_I net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_82_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_20_Left_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1003_ net115 _0433_ _0443_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_1_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0718_ _0194_ net328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input150_I simpleuart_reg_div_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I mem_addr[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput110 simpleuart_reg_dat_do[16] net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput176 spimem_rdata[17] net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput198 spimem_rdata[8] net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput187 spimem_rdata[27] net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput121 simpleuart_reg_dat_do[26] net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput132 simpleuart_reg_dat_do[7] net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_59_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput154 simpleuart_reg_div_do[26] net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput143 simpleuart_reg_div_do[16] net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput165 simpleuart_reg_div_do[7] net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1483_ net339 net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input3_I mem_addr[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input198_I spimem_rdata[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input59_I mem_wdata[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0983_ _0434_ _0435_ _0436_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1466_ net334 net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0883__A1 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1397_ _0024_ clknet_3_4__leaf_clk gpio\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input113_I simpleuart_reg_dat_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_61_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1320_ _0096_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1251_ _0662_ _0066_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1182_ net237 _0608_ _0609_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1290__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0897_ _0208_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0966_ _0419_ net175 _0421_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_6_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput233 net233 gpio_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput244 net244 gpio_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput299 net299 ram_wenb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput288 net288 ram_wenb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput266 net266 mem_rdata[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput277 net277 mem_rdata[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput255 net255 mem_rdata[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input230_I spimemio_cfgreg_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1281__A1 _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_85_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_72_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1272__A1 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0820_ _0285_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0751_ _0215_ _0222_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0682_ _0149_ _0153_ _0157_ _0165_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_10_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1303_ _0400_ _0097_ _0100_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1096_ net89 _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1234_ net52 _0643_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1165_ _0593_ _0599_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input180_I spimem_rdata[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0949_ _0404_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input41_I mem_wdata[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0829__A1 _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_32_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0803_ _0266_ _0270_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0734_ _0205_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_24_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0665_ _0147_ _0148_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_12_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1148_ _0187_ _0000_ net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1079_ _0178_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1217_ net48 _0630_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input89_I ram_rdata[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0948__I _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output245_I net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1002_ _0401_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0717_ _0183_ _0190_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input143_I simpleuart_reg_div_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput122 simpleuart_reg_dat_do[27] net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput111 simpleuart_reg_dat_do[17] net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput133 simpleuart_reg_dat_do[8] net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput144 simpleuart_reg_div_do[17] net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput100 ram_rdata[8] net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0678__I _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput188 spimem_rdata[28] net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput177 spimem_rdata[18] net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput199 spimem_rdata[9] net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_59_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput155 simpleuart_reg_div_do[27] net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput166 simpleuart_reg_div_do[8] net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_14_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1482_ net339 net304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0892__A2 net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0982_ net210 _0393_ _0408_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1465_ net334 net317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1396_ _0023_ clknet_3_4__leaf_clk gpio\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input106_I simpleuart_reg_dat_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input71_I ram_rdata[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output325_I net325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1181_ net38 _0606_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1250_ gpio\[30\] _0657_ _0658_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput234 net234 gpio_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_0896_ net106 _0332_ _0343_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_30_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0965_ _0420_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput245 net245 gpio_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput289 net289 ram_wenb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_65_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput278 net278 mem_rdata[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput256 net256 mem_rdata[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput267 net267 mem_rdata[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input223_I spimemio_cfgreg_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1379_ _0006_ clknet_3_2__leaf_clk net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_73_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output275_I net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_72_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0750_ _0217_ _0218_ _0221_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0681_ _0163_ net23 _0164_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1233_ _0649_ _0650_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_9_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1302_ gpio\[16\] _0099_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_63_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1095_ _0536_ _0537_ _0539_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_35_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1164_ net247 _0596_ _0598_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0948_ _0166_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input173_I spimem_rdata[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0879_ _0331_ _0307_ _0339_ _0340_ net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input34_I mem_wdata[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0765__A1 _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1190__A1 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_32_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0802_ _0267_ _0268_ _0269_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0733_ _0204_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0664_ net21 net20 net19 net25 _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1216_ _0636_ _0637_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_48_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1147_ _0579_ _0546_ _0586_ _0587_ net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_1_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1078_ iomem_rdata\[26\] _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_35_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_93_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output238_I net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0986__A1 _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0738__A1 net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0910__A1 _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1001_ iomem_rdata\[20\] _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_16_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0729__A1 _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_5__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0716_ _0193_ net327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input136_I simpleuart_reg_div_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput178 spimem_rdata[19] net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput123 simpleuart_reg_dat_do[28] net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput112 simpleuart_reg_dat_do[18] net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput134 simpleuart_reg_dat_do[9] net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput156 simpleuart_reg_div_do[28] net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1145__A1 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput145 simpleuart_reg_div_do[18] net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput167 simpleuart_reg_div_do[9] net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput101 ram_rdata[9] net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput189 spimem_rdata[29] net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_59_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1481_ net341 net303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1127__A1 _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1366__A1 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0981_ net145 _0405_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_17_Left_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1357__A1 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1464_ net334 net316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_26_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1395_ _0022_ clknet_3_4__leaf_clk gpio\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_53_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input64_I mem_wdata[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1348__A1 net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1133__I net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_24_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1339__A1 _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1180_ _0607_ _0610_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0964_ _0204_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput235 net235 gpio_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput246 net246 gpio_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_30_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0895_ _0205_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput257 net257 mem_rdata[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput268 net268 mem_rdata[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_66_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput279 net279 mem_rdata[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1378_ _0005_ clknet_3_0__leaf_clk net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_input216_I spimemio_cfgreg_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output268_I net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0680_ net12 net1 net26 _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_10_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1232_ gpio\[25\] _0646_ _0647_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1301_ _0098_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_63_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1094_ net220 _0538_ _0504_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1163_ _0597_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0947_ net110 _0380_ _0390_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0878_ _0319_ net169 _0320_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_input166_I simpleuart_reg_div_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input27_I mem_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0697__I _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0801_ _0220_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0756__A2 net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0732_ _0172_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0663_ net24 net22 _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_12_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1146_ _0558_ net192 _0559_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_9_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1215_ gpio\[21\] _0632_ _0634_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0692__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1077_ _0515_ _0500_ _0522_ _0523_ net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_31_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1000_ _0442_ _0402_ _0451_ _0452_ net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_89_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout331_I net332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0715_ _0181_ _0190_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0729__A2 _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input129_I simpleuart_reg_dat_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1129_ net126 _0179_ _0535_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_51_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input94_I ram_rdata[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output250_I net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput135 simpleuart_reg_dat_wait net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput124 simpleuart_reg_dat_do[29] net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput179 spimem_rdata[1] net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput168 spimem_rdata[0] net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput113 simpleuart_reg_dat_do[19] net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_59_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput157 simpleuart_reg_div_do[29] net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput146 simpleuart_reg_div_do[19] net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput102 resetn net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1480_ net341 net302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1046__I net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1136__A2 net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0885__I _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1063__A1 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0877__A1 _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0980_ net112 _0433_ _0390_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_27_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1463_ net337 net315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0868__A1 _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input1_I mem_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1394_ _0021_ clknet_3_4__leaf_clk gpio\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input196_I spimem_rdata[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input57_I mem_wdata[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1036__A1 _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1284__A1 net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1275__A1 _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0963_ _0418_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0894_ iomem_rdata\[12\] _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__1027__A1 _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput236 net236 gpio_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput247 net247 gpio_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput269 net269 mem_rdata[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput258 net258 mem_rdata[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_66_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1377_ _0004_ clknet_3_0__leaf_clk net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_input209_I spimemio_cfgreg_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input111_I simpleuart_reg_dat_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1266__A1 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_54_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_63_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1231_ net51 _0643_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1162_ net102 _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_9_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1300_ _0069_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_72_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_63_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1093_ _0168_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0877_ _0336_ _0338_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0946_ _0401_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_81_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input159_I simpleuart_reg_div_do[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1429_ _0056_ clknet_3_5__leaf_clk iomem_rdata\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_90_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output280_I net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_77_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_6_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_32_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0731_ iomem_rdata\[0\] _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_24_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0800_ net96 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1145_ _0583_ _0585_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1214_ net47 _0630_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1076_ _0512_ net185 _0513_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_43_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0929_ _0384_ _0386_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_82_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0714_ _0192_ net326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1059_ _0411_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1128_ iomem_rdata\[30\] _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input87_I ram_rdata[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput169 spimem_rdata[10] net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output243_I net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput125 simpleuart_reg_dat_do[2] net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput114 simpleuart_reg_dat_do[1] net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput103 simpleuart_reg_dat_do[0] net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput136 simpleuart_reg_div_do[0] net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput147 simpleuart_reg_div_do[1] net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput158 simpleuart_reg_div_do[2] net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input141_I simpleuart_reg_div_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1462_ net337 net314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1393_ _0020_ clknet_3_4__leaf_clk gpio\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input189_I spimem_rdata[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_61_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_24_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0962_ _0219_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0893_ _0341_ _0307_ _0352_ _0353_ net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xoutput248 net248 gpio_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput237 net237 gpio_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_50_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput259 net259 mem_rdata[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_66_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1376_ _0003_ clknet_3_0__leaf_clk net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_92_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input104_I simpleuart_reg_dat_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_21_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1193__A1 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1092_ net155 _0502_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1161_ _0595_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1230_ _0644_ _0648_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_71_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0876_ _0314_ _0337_ _0316_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0945_ _0204_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1428_ _0055_ clknet_3_5__leaf_clk iomem_rdata\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input221_I spimemio_cfgreg_do[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1359_ _0123_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0998__A1 _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output273_I net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0730_ _0202_ net323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1213_ _0631_ _0635_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_48_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1144_ _0553_ _0584_ _0555_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1075_ _0519_ _0521_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_1_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input171_I spimem_rdata[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0928_ _0362_ _0385_ _0364_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0859_ iomem_rdata\[9\] _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_16_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input32_I mem_addr[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1148__A1 _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0938__B _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0713_ _0182_ _0190_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1139__A1 net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1058_ _0501_ _0503_ _0505_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1127_ _0561_ _0546_ _0568_ _0569_ net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_8_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput126 simpleuart_reg_dat_do[30] net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput115 simpleuart_reg_dat_do[20] net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput104 simpleuart_reg_dat_do[10] net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output236_I net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput159 simpleuart_reg_div_do[30] net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput148 simpleuart_reg_div_do[20] net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput137 simpleuart_reg_div_do[10] net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_42_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1369__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1343__I _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input134_I simpleuart_reg_dat_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1163__I _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_27_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1461_ net336 net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1392_ _0019_ clknet_3_4__leaf_clk gpio\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1073__I net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0961_ _0410_ _0416_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0892_ _0319_ net170 _0320_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput238 net238 gpio_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_49_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput249 net249 mem_rdata[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__0700__I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1375_ _0002_ clknet_3_0__leaf_clk net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_81_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0777__A2 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input62_I mem_wdata[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1091_ net122 _0525_ _0535_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1160_ net67 _0594_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_71_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0944_ iomem_rdata\[16\] _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_0875_ net71 _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_87_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1358_ _0134_ _0135_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1427_ _0054_ clknet_3_5__leaf_clk iomem_rdata\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input214_I spimemio_cfgreg_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1289_ _0072_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output266_I net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1212_ gpio\[20\] _0632_ _0634_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1143_ net94 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1074_ _0507_ _0520_ _0509_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0927_ net75 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_93_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0789_ _0225_ net193 _0227_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0858_ _0306_ _0307_ _0318_ _0321_ net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA_input164_I simpleuart_reg_div_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input25_I mem_addr[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0712_ _0191_ net325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_69_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1126_ _0558_ net189 _0559_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_0_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1057_ net217 _0492_ _0504_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1075__A1 _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_78_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput127 simpleuart_reg_dat_do[31] net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput116 simpleuart_reg_dat_do[21] net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput105 simpleuart_reg_dat_do[11] net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput149 simpleuart_reg_div_do[21] net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput138 simpleuart_reg_div_do[11] net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_87_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1057__A1 net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input127_I simpleuart_reg_dat_do[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1109_ _0411_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1296__A1 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1048__A1 _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input92_I ram_rdata[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1287__A1 _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1460_ net336 net312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1391_ _0018_ clknet_3_4__leaf_clk gpio\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0960_ _0412_ _0413_ _0415_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput239 net239 gpio_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0891_ _0349_ _0351_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1084__I net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1374_ _0001_ clknet_3_0__leaf_clk net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input194_I spimem_rdata[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input55_I mem_wdata[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_14_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_9_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1090_ _0195_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_41_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1079__I _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0874_ _0333_ _0334_ _0335_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0943_ _0389_ _0355_ _0398_ _0399_ net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_11_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1288_ _0070_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1357_ net242 _0127_ _0128_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1426_ _0053_ clknet_3_5__leaf_clk iomem_rdata\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input207_I spimemio_cfgreg_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output259_I net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1142_ _0580_ _0581_ _0582_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1211_ _0633_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1362__I net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1073_ net87 _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0857_ _0319_ net198 _0320_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0926_ _0381_ _0382_ _0383_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_3_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input157_I simpleuart_reg_div_do[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0788_ _0254_ _0256_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1409_ _0036_ clknet_3_3__leaf_clk iomem_rdata\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input18_I mem_addr[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0840__A2 net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0711_ _0187_ _0190_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1125_ _0565_ _0567_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_32_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1056_ _0407_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0909_ _0367_ net171 _0368_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_16_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput117 simpleuart_reg_dat_do[22] net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput106 simpleuart_reg_dat_do[12] net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput128 simpleuart_reg_dat_do[3] net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput139 simpleuart_reg_div_do[12] net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1066__A2 net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_90_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1108_ _0547_ _0549_ _0551_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1039_ iomem_rdata\[23\] _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input85_I ram_rdata[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output241_I net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0785__B _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0798__A1 _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1390_ _0017_ clknet_3_4__leaf_clk gpio\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0961__A1 _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_69_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0713__A1 _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_24_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0890_ _0314_ _0350_ _0316_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1373_ _0145_ _0146_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input187_I spimem_rdata[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0934__A1 net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input48_I mem_wdata[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0925__A1 net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0873_ net202 _0299_ _0311_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0942_ _0367_ net174 _0368_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_2_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1425_ _0052_ clknet_3_5__leaf_clk iomem_rdata\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1287_ _0341_ _0084_ _0089_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1356_ net59 _0124_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_34_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input102_I resetn vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_76_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1141_ net225 _0188_ _0550_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_48_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1072_ _0516_ _0517_ _0518_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1210_ net102 _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0925_ net206 _0347_ _0359_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0856_ _0226_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0787_ _0217_ _0255_ _0221_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1408_ _0035_ clknet_3_3__leaf_clk iomem_rdata\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_82_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1339_ _0579_ _0116_ _0121_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output271_I net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0710_ _0189_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1124_ _0553_ _0566_ _0555_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1055_ net152 _0502_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0908_ _0226_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0839_ _0301_ _0303_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput118 simpleuart_reg_dat_do[23] net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput107 simpleuart_reg_dat_do[13] net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput129 simpleuart_reg_dat_do[4] net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input30_I mem_addr[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1107_ net221 _0538_ _0550_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1038_ _0478_ _0454_ _0486_ _0487_ net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input78_I ram_rdata[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output234_I net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0789__A2 net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input132_I simpleuart_reg_dat_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1471__I net335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1372_ net246 _0138_ _0139_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0689__A1 net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0941_ _0395_ _0397_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0872_ net137 _0309_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_79_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1355_ _0132_ _0133_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1424_ _0051_ clknet_3_5__leaf_clk iomem_rdata\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1286_ net235 _0085_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input60_I mem_wdata[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1140_ net160 _0548_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1071_ net218 _0492_ _0504_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0924_ net141 _0357_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0855_ _0224_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0786_ net95 _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_93_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1407_ _0034_ clknet_3_2__leaf_clk iomem_rdata\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1338_ gpio\[31\] _0117_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input212_I spimemio_cfgreg_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1269_ _0072_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_19_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output264_I net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1069__A1 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_29_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1054_ _0404_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1123_ net91 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_38_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0807__A1 _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0907_ _0224_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput108 simpleuart_reg_dat_do[14] net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0769_ _0179_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0838_ _0267_ _0302_ _0269_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input162_I simpleuart_reg_div_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput119 simpleuart_reg_dat_do[24] net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input23_I mem_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_1__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_56_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1223__A1 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_90_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1106_ _0407_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1037_ _0466_ net182 _0467_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_44_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput90 ram_rdata[28] net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_10_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input125_I simpleuart_reg_dat_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input90_I ram_rdata[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_24_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1371_ net63 _0136_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0916__I net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0940_ _0362_ _0396_ _0364_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0871_ net104 _0332_ _0296_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_10_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_79_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1285_ _0331_ _0084_ _0088_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1354_ net241 _0127_ _0128_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1423_ _0050_ clknet_3_5__leaf_clk iomem_rdata\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0736__I _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input192_I spimem_rdata[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input53_I mem_wdata[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_76_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1070_ net153 _0502_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1087__A2 net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout338_I net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0923_ net108 _0380_ _0343_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0854_ _0313_ _0317_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_93_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0785_ _0250_ _0251_ _0253_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_23_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1268_ _0070_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1406_ _0033_ clknet_3_2__leaf_clk iomem_rdata\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_3_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1337_ _0570_ _0116_ _0120_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input205_I spimemio_cfgreg_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1199_ gpio\[17\] _0621_ _0622_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0761__A1 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output257_I net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0816__A2 net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1122_ _0562_ _0563_ _0564_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1053_ net119 _0479_ _0489_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_16_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0991__A1 net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0906_ _0361_ _0365_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0837_ net99 _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput109 simpleuart_reg_dat_do[15] net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input155_I simpleuart_reg_div_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0768_ iomem_rdata\[2\] _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_0699_ net68 _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input16_I mem_addr[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0982__A1 net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_58_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_90_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I mem_addr[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0725__A1 _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1150__A1 _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1105_ net156 _0548_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1036_ _0483_ _0485_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0744__I _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput91 ram_rdata[29] net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput80 ram_rdata[19] net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1141__A1 net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_75_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_84_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_69_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input118_I simpleuart_reg_dat_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1019_ net116 _0433_ _0443_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_24_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_93_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input83_I ram_rdata[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0937__A1 net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1370_ _0143_ _0144_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_66_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_37_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1335__A1 _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0689__A3 _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0870_ _0285_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1422_ _0049_ clknet_3_5__leaf_clk iomem_rdata\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1284_ net234 _0085_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1353_ net56 _0124_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_34_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input185_I spimem_rdata[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0999_ _0419_ net178 _0421_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_6_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input46_I mem_wdata[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1317__A1 _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0927__I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0837__I net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_48_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0922_ _0285_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0853_ _0314_ _0315_ _0316_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_93_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0784_ net226 _0252_ _0213_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1405_ _0032_ clknet_3_2__leaf_clk iomem_rdata\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1267_ _0248_ _0071_ _0077_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__0747__I net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1198_ net42 _0618_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput1 mem_addr[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1336_ gpio\[30\] _0117_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input100_I ram_rdata[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1121_ net222 _0538_ _0550_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1052_ _0401_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_28_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0836_ _0297_ _0298_ _0300_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0767_ _0229_ _0206_ _0236_ _0237_ net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_0905_ _0362_ _0363_ _0364_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0698_ _0179_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input148_I simpleuart_reg_div_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1319_ _0488_ _0104_ _0109_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_50_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0725__A2 _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1104_ _0404_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1035_ _0461_ _0484_ _0463_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0819_ _0178_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput92 ram_rdata[2] net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput81 ram_rdata[1] net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput70 ram_rdata[0] net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_55_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0891__A1 _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_69_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1018_ iomem_rdata\[21\] _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_72_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input76_I ram_rdata[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0873__A1 net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1050__A1 _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1041__A1 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0919__A2 net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input228_I spimemio_cfgreg_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input130_I simpleuart_reg_dat_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1280__A1 net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1032__A1 net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_71_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1271__A1 _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1421_ _0048_ clknet_3_6__leaf_clk iomem_rdata\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_79_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1283_ _0322_ _0084_ _0087_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1352_ _0130_ _0131_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1262__A1 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input178_I spimem_rdata[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0998_ _0448_ _0450_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input39_I mem_wdata[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0921_ iomem_rdata\[14\] _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0783_ _0188_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0852_ _0220_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1404_ _0031_ clknet_3_2__leaf_clk iomem_rdata\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1335_ _0561_ _0116_ _0119_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1266_ net242 _0073_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1197_ _0619_ _0623_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput2 mem_addr[10] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0763__I net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_81_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1226__A1 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_2_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1120_ net157 _0548_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1051_ iomem_rdata\[24\] _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_56_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0904_ _0220_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_16_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0835_ net230 _0299_ _0264_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0697_ _0178_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0766_ _0225_ net179 _0227_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_11_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1318_ gpio\[23\] _0105_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_16_Left_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input210_I spimemio_cfgreg_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1249_ net57 _0655_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output262_I net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1103_ net123 _0525_ _0535_ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1034_ net84 _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input160_I simpleuart_reg_div_do[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput93 ram_rdata[30] net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput82 ram_rdata[20] net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0818_ iomem_rdata\[6\] _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_0749_ _0220_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput60 mem_wdata[4] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput71 ram_rdata[10] net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_55_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input21_I mem_addr[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0951__I _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1017_ _0453_ _0454_ _0465_ _0468_ net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_8_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input69_I mem_wstrb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input123_I simpleuart_reg_dat_do[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_8_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1099__A2 net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1351_ net240 _0127_ _0128_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1420_ _0047_ clknet_3_3__leaf_clk iomem_rdata\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1282_ net248 _0085_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_34_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1210__I net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0997_ _0412_ _0449_ _0415_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0828__A2 net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_4__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0920_ _0370_ _0355_ _0377_ _0378_ net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_0782_ net161 _0209_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0851_ net100 _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1403_ _0030_ clknet_3_2__leaf_clk iomem_rdata\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1265_ _0238_ _0071_ _0076_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1334_ gpio\[29\] _0117_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_19_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput3 mem_addr[11] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1196_ gpio\[16\] _0621_ _0622_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input190_I spimem_rdata[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0994__A1 net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input51_I mem_wdata[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1050_ _0488_ _0454_ _0497_ _0498_ net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__0864__I net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout336_I net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0834_ _0188_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0903_ net73 _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_16_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0765_ _0233_ _0235_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0696_ _0161_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0900__A1 net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1248_ _0660_ _0661_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1317_ _0478_ _0104_ _0108_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input203_I spimemio_cfgreg_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0774__I net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1179_ net236 _0608_ _0609_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_50_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input99_I ram_rdata[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output255_I net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1135__A1 _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1102_ _0401_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_1033_ _0480_ _0481_ _0482_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0817_ _0275_ _0260_ _0282_ _0283_ net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_3_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput61 mem_wdata[5] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput50 mem_wdata[24] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput72 ram_rdata[11] net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput94 ram_rdata[31] net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input153_I simpleuart_reg_div_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput83 ram_rdata[21] net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0748_ _0219_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0679_ net33 _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_55_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input14_I mem_addr[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1117__A1 _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_35_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_44_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_53_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input6_I mem_addr[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_60_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1016_ _0466_ net180 _0467_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_62_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_71_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_68_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1123__I net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input116_I simpleuart_reg_dat_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1411__CLK clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input81_I ram_rdata[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0957__I net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1281_ _0306_ _0084_ _0086_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1350_ net45 _0124_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_8_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_34_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0996_ net80 _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1479_ net330 net301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output285_I net342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0850_ _0216_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0781_ net128 _0239_ _0249_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1402_ _0029_ clknet_3_2__leaf_clk iomem_rdata\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1264_ net241 _0073_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput4 mem_addr[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1333_ _0545_ _0116_ _0118_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1195_ _0597_ _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input183_I spimem_rdata[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0979_ _0285_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input44_I mem_wdata[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_2_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_44_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0833_ net165 _0262_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0902_ _0216_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__0976__A2 net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0695_ _0177_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0764_ _0217_ _0234_ _0221_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1247_ gpio\[29\] _0657_ _0658_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1178_ _0597_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1316_ gpio\[22\] _0105_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output248_I net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xsimple_interconnect_350 gpio_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_80_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1080__A1 net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1032_ net215 _0446_ _0458_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0875__I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1101_ iomem_rdata\[28\] _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_84_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0824__B _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1071__A1 net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0816_ _0272_ net195 _0273_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xinput84 ram_rdata[22] net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0747_ net200 _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput95 ram_rdata[3] net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput62 mem_wdata[6] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput40 mem_wdata[15] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput51 mem_wdata[25] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput73 ram_rdata[12] net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input146_I simpleuart_reg_div_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1126__A2 net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0678_ _0161_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_55_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1053__A1 net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1015_ _0420_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_60_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1044__A1 net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1292__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0858__A1 _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1283__A1 _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1340__S _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput230 spimemio_cfgreg_do[7] net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1274__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input109_I simpleuart_reg_dat_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_65_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input74_I ram_rdata[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1017__A1 _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output328_I net328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0973__I net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_71_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_79_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1280_ net247 _0085_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_8_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0995_ _0444_ _0445_ _0447_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_26_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input226_I spimemio_cfgreg_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1478_ net330 net300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output278_I net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_5_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0780_ _0196_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1401_ _0028_ clknet_3_3__leaf_clk iomem_rdata\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1263_ _0229_ _0071_ _0075_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput5 mem_addr[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1194_ _0620_ _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1332_ gpio\[28\] _0117_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_19_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input176_I spimem_rdata[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0978_ iomem_rdata\[18\] _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_14_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput320 net320 simpleuart_div_we[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input37_I mem_wdata[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1147__B1 _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_16_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0832_ net132 _0286_ _0296_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0901_ _0356_ _0358_ _0360_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0763_ net81 _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0694_ net18 net281 _0174_ _0176_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1315_ _0469_ _0104_ _0107_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1246_ net55 _0655_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1177_ _0595_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_50_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xsimple_interconnect_351 gpio_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_13_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1031_ net150 _0456_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_29_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1100_ _0534_ _0500_ _0543_ _0544_ net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout341_I net342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput85 ram_rdata[23] net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0815_ _0279_ _0281_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0746_ net70 _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput74 ram_rdata[13] net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput63 mem_wdata[7] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 mem_wdata[16] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 mem_wdata[26] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput30 mem_addr[7] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput96 ram_rdata[4] net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input139_I simpleuart_reg_div_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0677_ _0149_ _0153_ _0157_ _0160_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_55_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1229_ gpio\[24\] _0646_ _0647_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output260_I net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0867__A2 net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1014_ _0418_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_60_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0729_ _0183_ _0198_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput231 spimemio_cfgreg_do[8] net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput220 spimemio_cfgreg_do[27] net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1026__A2 net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0776__A1 _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input67_I mem_wstrb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1060__I net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0994_ net211 _0446_ _0408_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1477_ net330 net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input219_I spimemio_cfgreg_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input121_I simpleuart_reg_dat_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_68_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0984__I net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_77_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_86_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0988__A1 _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0912__A1 net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1400_ _0027_ clknet_3_6__leaf_clk iomem_rdata\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1331_ _0098_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_47_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1262_ net240 _0073_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1193_ net68 _0594_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput6 mem_addr[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput310 net310 ram_wenb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_30_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput321 net321 simpleuart_div_we[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0977_ _0423_ _0402_ _0430_ _0431_ net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA_input169_I spimem_rdata[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_2_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1156__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_92_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1147__A1 _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0900_ net204 _0347_ _0359_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_44_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0831_ _0196_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0762_ _0230_ _0231_ _0232_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0693_ _0151_ _0152_ _0154_ _0175_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_12_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0889__I net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1314_ gpio\[21\] _0105_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1176_ net37 _0606_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1245_ _0656_ _0659_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1129__A1 net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_13_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xsimple_interconnect_352 gpio_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_18_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1030_ net117 _0479_ _0443_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_29_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout334_I net335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0814_ _0267_ _0280_ _0269_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput31 mem_addr[8] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 mem_addr[27] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput86 ram_rdata[24] net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0745_ _0216_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput75 ram_rdata[14] net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0676_ net33 _0158_ net26 _0159_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xinput64 mem_wdata[8] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput42 mem_wdata[17] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 mem_wdata[27] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput97 ram_rdata[5] net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1243__I _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1228_ _0633_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1414__CLK clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input201_I spimemio_cfgreg_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_55_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1159_ _0589_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input97_I ram_rdata[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output253_I net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1013_ _0460_ _0464_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_22_Left_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_60_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input151_I simpleuart_reg_div_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0728_ _0201_ net322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_40_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input12_I mem_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_7__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput221 spimemio_cfgreg_do[28] net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput210 spimemio_cfgreg_do[18] net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput232 spimemio_cfgreg_do[9] net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I mem_addr[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input199_I spimem_rdata[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_8_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0993_ _0346_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1476_ net329 net298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0930__A2 net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input114_I simpleuart_reg_dat_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1261_ _0203_ _0071_ _0074_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1330_ _0096_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1192_ net41 _0618_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput7 mem_addr[15] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0976_ _0419_ net176 _0421_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xoutput300 net300 ram_wenb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput311 net311 ram_wenb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_30_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput322 net322 simpleuart_div_we[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input231_I spimemio_cfgreg_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1459_ net336 net311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output283_I net335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0830_ iomem_rdata\[7\] _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_16_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0761_ net212 _0189_ _0213_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_24_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0692_ net17 net3 _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_11_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1244_ gpio\[28\] _0657_ _0658_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1313_ _0453_ _0104_ _0106_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1175_ _0591_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input181_I spimem_rdata[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0821__A1 net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0959_ _0414_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input42_I mem_wdata[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xsimple_interconnect_353 gpio_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_78_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0879__A1 _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0803__A1 _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0813_ net97 _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput10 mem_addr[18] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 mem_wdata[18] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput54 mem_wdata[28] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 mem_addr[9] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 mem_addr[28] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput87 ram_rdata[25] net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__0849__B _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0744_ _0211_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput76 ram_rdata[15] net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput65 mem_wdata[9] net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0675_ net12 net1 _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput98 ram_rdata[6] net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_55_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1158_ net64 _0592_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1227_ _0645_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1089_ iomem_rdata\[27\] _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_90_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output246_I net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1286__A1 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1038__A1 _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1012_ _0461_ _0462_ _0463_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0727_ _0181_ _0198_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input144_I simpleuart_reg_div_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput211 spimemio_cfgreg_do[19] net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput200 spimem_ready net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput222 spimemio_cfgreg_do[29] net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_89_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0992_ net146 _0405_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0701__I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1475_ net329 net296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input107_I simpleuart_reg_dat_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0694__A2 net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input72_I ram_rdata[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output326_I net326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1260_ net233 _0073_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1191_ _0617_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput8 mem_addr[16] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0975_ _0427_ _0429_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput301 net301 ram_wenb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput312 net312 ram_wenb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput323 net323 simpleuart_div_we[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input224_I spimemio_cfgreg_do[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1458_ net336 net308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1389_ _0016_ clknet_3_3__leaf_clk gpio\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output276_I net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0760_ net147 _0209_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_16_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0691_ _0163_ _0170_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1347__I _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1174_ _0604_ _0605_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1243_ _0633_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1312_ gpio\[20\] _0105_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input174_I spimem_rdata[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0958_ _0219_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0889_ net72 _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input35_I mem_wdata[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xsimple_interconnect_354 gpio_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsimple_interconnect_343 gpio_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_92_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput88 ram_rdata[26] net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0743_ _0207_ _0210_ _0214_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0812_ _0276_ _0277_ _0278_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput77 ram_rdata[16] net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__0690__B _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput66 mem_wstrb[0] net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput44 mem_wdata[19] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput55 mem_wdata[29] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 mem_addr[29] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput33 mem_valid net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput11 mem_addr[19] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0674_ net23 _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xinput99 ram_rdata[7] net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1157_ _0591_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1226_ net69 _0594_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_90_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1088_ _0524_ _0500_ _0532_ _0533_ net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_70_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output239_I net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_26_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0797__A1 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1011_ _0414_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_60_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0788__A1 _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0726_ _0200_ net321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input137_I simpleuart_reg_div_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1209_ _0620_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_23_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput201 spimemio_cfgreg_do[0] net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput223 spimemio_cfgreg_do[2] net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput212 spimemio_cfgreg_do[1] net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_89_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1090__I _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0709_ _0188_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0991_ net113 _0433_ _0443_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1474_ net329 net295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Left_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_28_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input65_I mem_wdata[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_37_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0906__A1 _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 mem_addr[17] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1190_ net68 _0590_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0974_ _0412_ _0428_ _0415_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput324 net324 spimem_valid vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput302 net302 ram_wenb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_77_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput313 net313 ram_wenb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1457_ net338 net297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1417__CLK clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input217_I spimemio_cfgreg_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1388_ _0015_ clknet_3_3__leaf_clk gpio\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1313__A1 _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1077__B1 _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output269_I net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_44_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0690_ net135 _0162_ _0166_ _0173_ net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_51_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1311_ _0098_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1173_ net235 _0596_ _0598_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1242_ _0645_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0707__I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0888_ _0344_ _0345_ _0348_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0957_ net77 _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input167_I simpleuart_reg_div_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input28_I mem_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xsimple_interconnect_355 gpio_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsimple_interconnect_344 gpio_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_65_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0811_ net228 _0252_ _0264_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0742_ net201 _0189_ _0213_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xinput89 ram_rdata[27] net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput78 ram_rdata[17] net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput67 mem_wstrb[1] net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0673_ _0154_ _0155_ _0156_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xinput34 mem_wdata[0] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput56 mem_wdata[2] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput45 mem_wdata[1] net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 mem_addr[2] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput12 mem_addr[1] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1093__I _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1087_ _0512_ net186 _0513_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1225_ net50 _0643_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1156_ net67 _0590_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_63_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1178__I _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1010_ net82 _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout332_I net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0720__I _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0725_ _0182_ _0198_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1208_ net46 _0630_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1139_ net127 _0179_ _0196_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input95_I ram_rdata[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput213 spimemio_cfgreg_do[20] net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput224 spimemio_cfgreg_do[30] net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput202 spimemio_cfgreg_do[10] net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output251_I net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0942__A2 net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0708_ _0168_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I mem_addr[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0860__A1 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0990_ _0342_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1473_ net329 net294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input2_I mem_addr[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input197_I spimem_rdata[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input58_I mem_wdata[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_0__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1086__A1 _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput325 net325 spimemio_cfgreg_we[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput303 net303 ram_wenb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput314 net314 ram_wenb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_54_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1096__I net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0973_ net78 _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1456_ net338 net286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1387_ _0014_ clknet_3_1__leaf_clk gpio\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input112_I simpleuart_reg_dat_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0903__I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0815__A1 _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0813__I net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1241_ net54 _0655_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1310_ _0096_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1172_ net36 _0592_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0956_ _0411_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_65_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0887_ net203 _0347_ _0311_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_30_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_74_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1439_ _0065_ clknet_3_0__leaf_clk net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xsimple_interconnect_356 gpio_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsimple_interconnect_345 gpio_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_83_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output281_I net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_92_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0810_ net163 _0262_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_1_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput13 mem_addr[20] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0741_ _0212_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput79 ram_rdata[18] net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput24 mem_addr[30] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput68 mem_wstrb[2] net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0672_ net28 net27 net30 net29 _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput35 mem_wdata[10] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 mem_wdata[20] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput57 mem_wdata[30] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1224_ _0642_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_63_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1086_ _0529_ _0531_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1155_ _0589_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0939_ net76 _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input40_I mem_wdata[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0724_ _0199_ net320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_68_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1207_ _0617_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1069_ net120 _0479_ _0489_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1138_ iomem_rdata\[31\] _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_90_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input88_I ram_rdata[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput203 spimemio_cfgreg_do[11] net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput214 spimemio_cfgreg_do[21] net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput225 spimemio_cfgreg_do[31] net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output244_I net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0707_ net66 _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input142_I simpleuart_reg_div_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1472_ net331 net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0972_ _0424_ _0425_ _0426_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput326 net326 spimemio_cfgreg_we[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput304 net304 ram_wenb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput315 net315 ram_wenb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1386_ _0013_ clknet_3_1__leaf_clk gpio\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input105_I simpleuart_reg_dat_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input70_I ram_rdata[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0760__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output324_I net324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0751__A1 _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1171_ _0602_ _0603_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1240_ _0642_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0806__A2 net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0886_ _0346_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0955_ _0211_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0742__A1 net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input222_I spimemio_cfgreg_do[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1369_ net245 _0138_ _0139_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1438_ _0064_ clknet_3_0__leaf_clk net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xsimple_interconnect_357 gpio_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsimple_interconnect_346 gpio_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_21_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output274_I net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_57_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0740_ _0211_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput25 mem_addr[31] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput14 mem_addr[21] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 mem_wdata[11] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0671_ net32 net31 net3 net2 _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput69 mem_wstrb[3] net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput47 mem_wdata[21] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput58 mem_wdata[31] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1223_ net69 _0590_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1154_ _0169_ iomem_ready _0150_ _0174_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_90_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1085_ _0507_ _0530_ _0509_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input172_I spimem_rdata[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0938_ _0391_ _0392_ _0394_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0869_ iomem_rdata\[10\] _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0715__A1 _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input33_I mem_valid vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1131__A1 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0819__I _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_60_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0723_ _0187_ _0198_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_68_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1137_ _0570_ _0546_ _0577_ _0578_ net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_1206_ _0628_ _0629_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1068_ iomem_rdata\[25\] _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_31_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput215 spimemio_cfgreg_do[22] net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput204 spimemio_cfgreg_do[12] net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput226 spimemio_cfgreg_do[3] net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output237_I net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1113__A1 _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0918__A1 _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0706_ _0186_ net324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input135_I simpleuart_reg_dat_wait vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_70_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_78_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1471_ net335 net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1307__A1 _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_47_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0971_ net209 _0393_ _0408_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput327 net327 spimemio_cfgreg_we[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput305 net305 ram_wenb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_77_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput316 net316 ram_wenb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_22_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1385_ _0012_ clknet_3_1__leaf_clk gpio\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input63_I mem_wdata[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1170_ net234 _0596_ _0598_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0885_ _0168_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0954_ _0403_ _0406_ _0409_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1437_ _0063_ clknet_3_0__leaf_clk net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input215_I spimemio_cfgreg_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1430__CLK clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1368_ net62 _0136_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1299_ _0096_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xsimple_interconnect_358 gpio_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xsimple_interconnect_347 gpio_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_92_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output267_I net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout340 net341 net340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput37 mem_wdata[12] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput59 mem_wdata[3] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput15 mem_addr[22] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 mem_wdata[22] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 mem_addr[3] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0670_ net5 net4 net7 net6 _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1153_ _0588_ net319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1084_ net88 _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1222_ _0640_ _0641_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0937_ net207 _0393_ _0359_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_23_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0868_ _0322_ _0307_ _0329_ _0330_ net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_0799_ _0216_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input26_I mem_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input165_I simpleuart_reg_div_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_80_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0722_ _0197_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1136_ _0558_ net191 _0559_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1067_ _0499_ _0500_ _0511_ _0514_ net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_1205_ gpio\[19\] _0621_ _0622_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_31_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput216 spimemio_cfgreg_do[23] net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput205 spimemio_cfgreg_do[13] net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput227 spimemio_cfgreg_do[4] net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_89_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0705_ _0163_ _0169_ _0170_ _0176_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_input128_I simpleuart_reg_dat_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1119_ net124 _0525_ _0535_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0854__A1 _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input93_I ram_rdata[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0909__A2 net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1098__A1 _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1270__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1470_ net333 net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_33_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1013__A1 _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0827__A1 _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0970_ net144 _0405_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput328 net328 spimemio_cfgreg_we[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput306 net306 ram_wenb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_77_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput317 net317 ram_wenb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0809__A1 net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1384_ _0011_ clknet_3_1__leaf_clk gpio\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input195_I spimem_rdata[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input56_I mem_wdata[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_52_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_25_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0953_ net208 _0393_ _0408_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0884_ net138 _0309_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_34_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1367_ _0141_ _0142_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1436_ _0062_ clknet_3_0__leaf_clk net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input208_I spimemio_cfgreg_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input110_I simpleuart_reg_dat_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Left_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1298_ _0069_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xsimple_interconnect_348 gpio_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_46_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_52_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xfanout341 net342 net341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout330 net331 net330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_61_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_29_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_70_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput16 mem_addr[23] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput38 mem_wdata[13] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput49 mem_wdata[23] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 mem_addr[4] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1221_ gpio\[23\] _0632_ _0634_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1152_ _0187_ _0180_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1083_ _0526_ _0527_ _0528_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_90_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0936_ _0346_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0867_ _0319_ net199 _0320_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0798_ _0261_ _0263_ _0265_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input158_I simpleuart_reg_div_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1419_ _0046_ clknet_3_6__leaf_clk iomem_rdata\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_26_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input19_I mem_addr[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_5_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0851__I net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0721_ _0196_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1204_ net44 _0618_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1135_ _0574_ _0576_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_23_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1066_ _0512_ net184 _0513_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_31_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0919_ _0367_ net172 _0368_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_28_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput217 spimemio_cfgreg_do[24] net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput206 spimemio_cfgreg_do[14] net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput228 spimemio_cfgreg_do[5] net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_39_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_3__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0704_ _0185_ net318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_36_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1049_ _0466_ net183 _0467_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1118_ iomem_rdata\[29\] _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input86_I ram_rdata[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output242_I net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0666__I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_70_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0772__A1 net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input140_I simpleuart_reg_div_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1110__I net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_75_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput307 net307 ram_wenb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_50_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput318 net318 simpleuart_dat_re vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_50_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1383_ _0010_ clknet_3_1__leaf_clk gpio\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input188_I spimem_rdata[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input49_I mem_wdata[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1170__A1 net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0952_ _0407_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0883_ net105 _0332_ _0343_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0975__A1 _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0727__A1 _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1152__A1 _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1366_ net244 _0138_ _0139_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1435_ _0061_ clknet_3_0__leaf_clk net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_53_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input103_I simpleuart_reg_dat_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1297_ _0389_ _0090_ _0095_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xsimple_interconnect_349 gpio_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_58_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout331 net332 net331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0939__I net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout342 net285 net342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_29_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0674__I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput17 mem_addr[24] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput39 mem_wdata[14] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 mem_addr[5] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1151_ _0183_ _0177_ net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_20_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1220_ net49 _0630_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1082_ net219 _0492_ _0504_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0935_ net142 _0357_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0866_ _0326_ _0328_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0797_ net227 _0252_ _0264_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input220_I spimemio_cfgreg_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1125__A1 _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1349_ _0125_ _0129_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1418_ _0045_ clknet_3_3__leaf_clk iomem_rdata\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_62_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output272_I net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0720_ _0195_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1107__A1 net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1134_ _0553_ _0575_ _0555_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1203_ _0626_ _0627_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_23_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1065_ _0420_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input170_I spimem_rdata[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0849_ _0308_ _0310_ _0312_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0918_ _0374_ _0376_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput218 spimemio_cfgreg_do[25] net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput207 spimemio_cfgreg_do[15] net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput229 spimemio_cfgreg_do[6] net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input31_I mem_addr[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0901__B _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1337__A1 _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_73_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1023__I net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0703_ _0180_ _0184_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_88_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_36_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1117_ _0545_ _0546_ _0557_ _0560_ net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_75_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1048_ _0494_ _0496_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input79_I ram_rdata[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1319__A1 _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output235_I net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_78_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input133_I simpleuart_reg_dat_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput308 net308 ram_wenb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput319 net319 simpleuart_dat_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_35_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1382_ _0009_ clknet_3_1__leaf_clk gpio\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1211__I _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0690__A1 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_52_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0951_ _0211_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0882_ _0342_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0727__A2 _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1296_ net239 _0091_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1365_ net61 _0136_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1434_ _0060_ clknet_3_0__leaf_clk net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_92_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0966__A2 net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout332 net284 net332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input61_I mem_wdata[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0955__I _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput18 mem_addr[25] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput29 mem_addr[6] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1150_ _0181_ _0000_ net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1081_ net154 _0502_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__0893__A1 _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0934_ net109 _0380_ _0390_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0865_ _0314_ _0327_ _0316_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0796_ _0212_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1417_ _0044_ clknet_3_7__leaf_clk iomem_rdata\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input213_I spimemio_cfgreg_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1279_ _0072_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1348_ net233 _0127_ _0128_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output265_I net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1116__A2 net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1133_ net93 _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1064_ _0418_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1202_ gpio\[18\] _0621_ _0622_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__0866__A1 _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1291__A1 _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0848_ net231 _0299_ _0311_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_31_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0779_ iomem_rdata\[3\] _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_0917_ _0362_ _0375_ _0364_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput208 spimemio_cfgreg_do[16] net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput219 spimemio_cfgreg_do[26] net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input24_I mem_addr[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input163_I simpleuart_reg_div_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_49_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1282__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_58_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0848__A1 net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1273__A1 _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0702_ _0181_ _0182_ net66 _0183_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__1025__A1 _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_88_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1047_ _0461_ _0495_ _0463_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0839__A1 _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1116_ _0558_ net188 _0559_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1264__A1 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1255__A1 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1007__A1 net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1034__I net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_41_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input126_I simpleuart_reg_dat_do[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input91_I ram_rdata[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_75_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput309 net309 ram_wenb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1029__I _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1381_ _0008_ clknet_3_1__leaf_clk net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_1_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0681__A2 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0881_ _0195_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0950_ net143 _0405_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_15_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1137__B1 _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1433_ _0059_ clknet_3_0__leaf_clk net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_11_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1295_ _0379_ _0090_ _0094_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1364_ _0137_ _0140_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input193_I spimem_rdata[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout333 net334 net333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_21_Left_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input54_I mem_wdata[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput19 mem_addr[26] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1080_ net121 _0525_ _0489_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0881__I _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_28_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0933_ _0342_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0795_ net162 _0262_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0864_ net101 _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1347_ _0633_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1416_ _0043_ clknet_3_7__leaf_clk iomem_rdata\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input206_I spimemio_cfgreg_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1278_ _0070_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_62_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output258_I net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0915__B _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1201_ net43 _0618_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1132_ _0571_ _0572_ _0573_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1063_ _0506_ _0510_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_83_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0916_ net74 _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0847_ _0212_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_31_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0778_ _0238_ _0206_ _0246_ _0247_ net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_3_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput209 spimemio_cfgreg_do[17] net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input156_I simpleuart_reg_div_do[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0857__A2 net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0786__I net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input17_I mem_addr[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0793__A1 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0696__I _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0784__A1 net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0701_ net69 _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input9_I mem_addr[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1046_ net85 _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1115_ _0420_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1016__A2 net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_70_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1182__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input119_I simpleuart_reg_dat_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1029_ _0178_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input84_I ram_rdata[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output240_I net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1173__A1 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1380_ _0007_ clknet_3_1__leaf_clk net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1164__A1 net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0969__A1 net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0743__B _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0880_ iomem_rdata\[11\] _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1137__A1 _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1363_ net243 _0138_ _0139_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1432_ _0058_ clknet_3_0__leaf_clk net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1294_ net238 _0091_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input186_I spimem_rdata[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout334 net335 net334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input47_I mem_wdata[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1119__A1 net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0699__I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_6__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_28_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0932_ iomem_rdata\[15\] _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_23_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_93_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0794_ _0208_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0863_ _0323_ _0324_ _0325_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_2_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1346_ _0126_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1415_ _0042_ clknet_3_4__leaf_clk iomem_rdata\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_54_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1277_ _0295_ _0078_ _0083_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input101_I ram_rdata[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1143__I net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_25_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1200_ _0624_ _0625_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1131_ net224 _0538_ _0550_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1062_ _0507_ _0508_ _0509_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0915_ _0371_ _0372_ _0373_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0777_ _0225_ net190 _0227_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0846_ net166 _0309_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1228__I _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_67_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input149_I simpleuart_reg_div_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1329_ _0534_ _0110_ _0115_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_22_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output270_I net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput290 net290 ram_wenb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_69_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0926__B _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0700_ net67 _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1114_ _0418_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_64_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1045_ _0490_ _0491_ _0493_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0836__B _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0829_ _0284_ _0260_ _0293_ _0294_ net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_16_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0766__A2 net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_41_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1028_ iomem_rdata\[22\] _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_71_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input77_I ram_rdata[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output233_I net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0987__A2 net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input131_I simpleuart_reg_dat_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input229_I spimemio_cfgreg_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1091__A1 net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1146__A2 net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_43_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1082__A1 net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0896__A1 net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1293_ _0370_ _0090_ _0093_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1362_ net102 _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1431_ _0057_ clknet_3_5__leaf_clk iomem_ready vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput190 spimem_rdata[2] net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input179_I spimem_rdata[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout335 net283 net335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__0887__A1 net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0811__A1 net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0862_ net232 _0299_ _0311_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_36_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0931_ _0379_ _0355_ _0387_ _0388_ net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_0793_ net129 _0239_ _0249_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1276_ net246 _0079_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1345_ net66 _0589_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1414_ _0041_ clknet_3_7__leaf_clk iomem_rdata\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1294__A1 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1285__A1 _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_25_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1130_ net159 _0548_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_0_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1061_ _0414_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1276__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0914_ net205 _0347_ _0359_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0845_ _0208_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0776_ _0243_ _0245_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input211_I spimemio_cfgreg_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1259_ _0072_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1328_ gpio\[27\] _0111_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1019__A1 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_18_Left_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output263_I net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput291 net291 ram_wenb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput280 net280 mem_rdata[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_27_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_36_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_88_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1044_ net216 _0492_ _0458_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1113_ _0552_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_88_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_72_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0759_ net114 _0180_ _0197_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0828_ _0272_ net196 _0273_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_16_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input22_I mem_addr[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input161_I simpleuart_reg_div_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0762__B _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1100__B1 _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1027_ _0469_ _0454_ _0476_ _0477_ net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input124_I simpleuart_reg_dat_do[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1162__I net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1430_ _0000_ clknet_3_7__leaf_clk ram_ready vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput180 spimem_rdata[20] net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_91_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1292_ net237 _0091_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1361_ _0126_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput191 spimem_rdata[30] net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout336 net282 net336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0878__A2 net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0996__I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0930_ _0367_ net173 _0368_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0792_ _0205_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_0861_ net167 _0309_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1413_ _0040_ clknet_3_6__leaf_clk iomem_rdata\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1275_ _0284_ _0078_ _0082_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1344_ net34 _0124_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_62_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input191_I spimem_rdata[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input52_I mem_wdata[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1037__A2 net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1060_ net86 _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0844_ net133 _0286_ _0296_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0913_ net140 _0357_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0775_ _0217_ _0244_ _0221_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input204_I spimemio_cfgreg_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0711__A1 _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1258_ _0069_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1189_ _0615_ _0616_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1327_ _0524_ _0110_ _0114_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output256_I net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput270 net270 mem_rdata[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput292 net292 ram_wenb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__0702__A1 _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput281 net281 mem_ready vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0941__A1 _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1043_ _0346_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1112_ _0553_ _0554_ _0555_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_36_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0758_ iomem_rdata\[1\] _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_0827_ _0290_ _0292_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1185__A1 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input154_I simpleuart_reg_div_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0689_ net200 ram_ready _0168_ _0172_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA_input15_I mem_addr[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0923__A1 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_33_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1167__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0914__A1 net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I mem_addr[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0863__B _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1026_ _0466_ net181 _0467_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_8_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_55_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_64_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0773__B _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_73_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1149__A1 _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_82_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_46_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_91_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input117_I simpleuart_reg_dat_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1009_ _0411_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input82_I ram_rdata[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1416__CLK clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_43_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_15_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1360_ net60 _0136_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput181 spimem_rdata[21] net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput192 spimem_rdata[31] net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput170 spimem_rdata[11] net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1291_ _0354_ _0090_ _0092_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout337 net338 net337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0860_ net134 _0286_ _0296_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0791_ iomem_rdata\[4\] _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_3_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1412_ _0039_ clknet_3_6__leaf_clk iomem_rdata\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1343_ _0123_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1274_ net245 _0079_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input184_I spimem_rdata[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0989_ iomem_rdata\[19\] _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_14_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input45_I mem_wdata[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0800__I net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0912_ net107 _0332_ _0343_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0843_ _0205_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_0774_ net92 _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1326_ gpio\[26\] _0111_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1257_ _0070_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1188_ net239 _0608_ _0609_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput293 net293 ram_wenb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput282 net338 ram_gwenb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_42_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput271 net271 mem_rdata[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput260 net260 mem_rdata[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_output249_I net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0702__A2 _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1111_ _0414_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1042_ net151 _0456_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0757_ _0203_ _0206_ _0223_ _0228_ net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_0826_ _0267_ _0291_ _0269_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0688_ _0169_ _0170_ _0171_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_input147_I simpleuart_reg_div_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1309_ _0442_ _0097_ _0103_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0999__A2 net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1025_ _0473_ _0475_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0809_ net130 _0239_ _0249_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_4_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1094__A1 net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0832__A1 net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0874__B _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0823__A1 net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1008_ _0455_ _0457_ _0459_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input75_I ram_rdata[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput182 spimem_rdata[22] net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput171 spimem_rdata[12] net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput193 spimem_rdata[3] net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput160 simpleuart_reg_div_do[31] net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1290_ net236 _0091_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout338 net282 net338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_92_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input227_I spimemio_cfgreg_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output279_I net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0790_ _0248_ _0206_ _0257_ _0258_ net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_11_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1273_ _0275_ _0078_ _0081_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1411_ _0038_ clknet_3_7__leaf_clk iomem_rdata\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1342_ net66 _0594_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0708__I _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0988_ _0432_ _0402_ _0440_ _0441_ net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA_input177_I spimem_rdata[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input38_I mem_wdata[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0842_ iomem_rdata\[8\] _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_0911_ iomem_rdata\[13\] _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__1359__I _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0773_ _0240_ _0241_ _0242_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1256_ _0069_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1325_ _0515_ _0110_ _0113_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1187_ net40 _0606_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput294 net294 ram_wenb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput283 net335 ram_gwenb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput261 net261 mem_rdata[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput250 net250 mem_rdata[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput272 net272 mem_rdata[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__0702__A3 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_88_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1110_ net90 _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout342_I net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1041_ net118 _0479_ _0489_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0825_ net98 _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0756_ _0225_ net168 _0227_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0687_ _0163_ iomem_ready _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1239_ _0653_ _0654_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1308_ gpio\[19\] _0099_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output261_I net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1024_ _0461_ _0474_ _0463_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0808_ iomem_rdata\[5\] _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_0739_ ram_ready _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input20_I mem_addr[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_46_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1007_ net213 _0446_ _0458_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1076__A2 net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input68_I mem_wstrb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput172 spimem_rdata[13] net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput194 spimem_rdata[4] net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput183 spimem_rdata[23] net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_59_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput150 simpleuart_reg_div_do[22] net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput161 simpleuart_reg_div_do[3] net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1487_ net340 net310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout339 net341 net339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_6_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input122_I simpleuart_reg_dat_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1049__A2 net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0980__A1 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_56_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0971__A1 net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1410_ _0037_ clknet_3_6__leaf_clk iomem_rdata\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_79_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1272_ net244 _0079_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1341_ _0122_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0723__A1 _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_88_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_62_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0987_ _0419_ net177 _0421_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_13_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0953__A1 net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0772_ net223 _0189_ _0213_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_36_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0841_ _0295_ _0260_ _0304_ _0305_ net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_0910_ _0354_ _0355_ _0366_ _0369_ net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_3_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1121__A1 net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1255_ net102 _0589_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1186_ _0613_ _0614_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1324_ gpio\[25\] _0111_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1188__A1 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput240 net240 gpio_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput295 net295 ram_wenb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput284 net332 ram_gwenb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input50_I mem_wdata[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput251 net251 mem_rdata[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput262 net262 mem_rdata[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput273 net273 mem_rdata[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__0702__A4 _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1195__I _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1179__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1040_ _0342_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1103__A1 net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1351__A1 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout335_I net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0755_ _0226_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0824_ _0287_ _0288_ _0289_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0686_ _0147_ _0148_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1342__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input202_I spimemio_cfgreg_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1169_ net35 _0592_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1238_ gpio\[27\] _0646_ _0647_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1307_ _0432_ _0097_ _0102_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input98_I ram_rdata[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output254_I net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1333__A1 _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_77_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1023_ net83 _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_32_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0738_ net136 _0209_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0807_ _0259_ _0260_ _0271_ _0274_ net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_25_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0888__B _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_15_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input152_I simpleuart_reg_div_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1315__A1 _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0669_ net18 _0150_ _0151_ _0152_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_4_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input13_I mem_addr[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_33_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Left_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_85_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_51_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input5_I mem_addr[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1006_ _0407_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_17_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput151 simpleuart_reg_div_do[23] net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput140 simpleuart_reg_div_do[13] net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput162 simpleuart_reg_div_do[4] net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput184 spimem_rdata[24] net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput173 spimem_rdata[14] net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput195 spimem_rdata[5] net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout329 net331 net329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1486_ net340 net309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input115_I simpleuart_reg_dat_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input80_I ram_rdata[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1340_ iomem_ready _0590_ _0597_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1271_ _0259_ _0078_ _0080_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__0723__A2 _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0740__I _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0986_ _0437_ _0439_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1469_ net333 net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input232_I spimemio_cfgreg_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output284_I net332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0825__I net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0840_ _0272_ net197 _0273_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0771_ net158 _0209_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1323_ _0499_ _0110_ _0112_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1254_ _0067_ _0068_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1185_ net238 _0608_ _0609_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input182_I spimem_rdata[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput241 net241 gpio_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0969_ net111 _0380_ _0390_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_30_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput252 net252 mem_rdata[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_6_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput296 net296 ram_wenb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput285 net342 ram_gwenb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput274 net274 mem_rdata[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput263 net263 mem_rdata[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input43_I mem_wdata[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_38_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0871__A1 net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0862__A1 net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0823_ net229 _0252_ _0264_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0754_ _0204_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0685_ net18 _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_20_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1306_ gpio\[18\] _0099_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1099_ _0512_ net187 _0513_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1237_ net53 _0643_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1168_ _0600_ _0601_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1030__A1 net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output247_I net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0844__A1 net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1021__A1 net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0835__A1 net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1022_ _0470_ _0471_ _0472_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1260__A1 net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0806_ _0272_ net194 _0273_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0737_ _0208_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0668_ net9 net8 net11 net10 _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input145_I simpleuart_reg_div_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1003__A1 net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0817__A1 _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1005_ net148 _0456_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_51_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput185 spimem_rdata[25] net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput174 spimem_rdata[15] net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput196 spimem_rdata[6] net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_91_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput130 simpleuart_reg_dat_do[5] net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput152 simpleuart_reg_div_do[24] net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput141 simpleuart_reg_div_do[14] net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput163 simpleuart_reg_div_do[5] net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1485_ net339 net307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pcpi_approx_mul
  CLASS BLOCK ;
  FOREIGN pcpi_approx_mul ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 250.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END clk
  PIN pcpi_insn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 188.160 300.000 188.720 ;
    END
  END pcpi_insn[0]
  PIN pcpi_insn[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END pcpi_insn[10]
  PIN pcpi_insn[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END pcpi_insn[11]
  PIN pcpi_insn[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 246.000 141.680 250.000 ;
    END
  END pcpi_insn[12]
  PIN pcpi_insn[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 246.000 145.040 250.000 ;
    END
  END pcpi_insn[13]
  PIN pcpi_insn[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 246.000 148.400 250.000 ;
    END
  END pcpi_insn[14]
  PIN pcpi_insn[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 0.000 7.280 4.000 ;
    END
  END pcpi_insn[15]
  PIN pcpi_insn[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END pcpi_insn[16]
  PIN pcpi_insn[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END pcpi_insn[17]
  PIN pcpi_insn[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 4.000 ;
    END
  END pcpi_insn[18]
  PIN pcpi_insn[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 0.000 20.720 4.000 ;
    END
  END pcpi_insn[19]
  PIN pcpi_insn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 161.280 300.000 161.840 ;
    END
  END pcpi_insn[1]
  PIN pcpi_insn[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END pcpi_insn[20]
  PIN pcpi_insn[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END pcpi_insn[21]
  PIN pcpi_insn[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END pcpi_insn[22]
  PIN pcpi_insn[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END pcpi_insn[23]
  PIN pcpi_insn[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END pcpi_insn[24]
  PIN pcpi_insn[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 178.080 300.000 178.640 ;
    END
  END pcpi_insn[25]
  PIN pcpi_insn[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 154.560 300.000 155.120 ;
    END
  END pcpi_insn[26]
  PIN pcpi_insn[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 134.400 300.000 134.960 ;
    END
  END pcpi_insn[27]
  PIN pcpi_insn[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 151.200 300.000 151.760 ;
    END
  END pcpi_insn[28]
  PIN pcpi_insn[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 137.760 300.000 138.320 ;
    END
  END pcpi_insn[29]
  PIN pcpi_insn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 181.440 300.000 182.000 ;
    END
  END pcpi_insn[2]
  PIN pcpi_insn[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 164.640 300.000 165.200 ;
    END
  END pcpi_insn[30]
  PIN pcpi_insn[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 147.840 300.000 148.400 ;
    END
  END pcpi_insn[31]
  PIN pcpi_insn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 168.000 300.000 168.560 ;
    END
  END pcpi_insn[3]
  PIN pcpi_insn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 174.720 300.000 175.280 ;
    END
  END pcpi_insn[4]
  PIN pcpi_insn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 171.360 300.000 171.920 ;
    END
  END pcpi_insn[5]
  PIN pcpi_insn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 184.800 300.000 185.360 ;
    END
  END pcpi_insn[6]
  PIN pcpi_insn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 0.000 40.880 4.000 ;
    END
  END pcpi_insn[7]
  PIN pcpi_insn[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END pcpi_insn[8]
  PIN pcpi_insn[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 4.000 ;
    END
  END pcpi_insn[9]
  PIN pcpi_rd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 73.920 300.000 74.480 ;
    END
  END pcpi_rd[0]
  PIN pcpi_rd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 80.640 300.000 81.200 ;
    END
  END pcpi_rd[10]
  PIN pcpi_rd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 104.160 300.000 104.720 ;
    END
  END pcpi_rd[11]
  PIN pcpi_rd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 127.680 300.000 128.240 ;
    END
  END pcpi_rd[12]
  PIN pcpi_rd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 110.880 300.000 111.440 ;
    END
  END pcpi_rd[13]
  PIN pcpi_rd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 107.520 300.000 108.080 ;
    END
  END pcpi_rd[14]
  PIN pcpi_rd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END pcpi_rd[15]
  PIN pcpi_rd[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END pcpi_rd[16]
  PIN pcpi_rd[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END pcpi_rd[17]
  PIN pcpi_rd[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END pcpi_rd[18]
  PIN pcpi_rd[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END pcpi_rd[19]
  PIN pcpi_rd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 84.000 300.000 84.560 ;
    END
  END pcpi_rd[1]
  PIN pcpi_rd[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END pcpi_rd[20]
  PIN pcpi_rd[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 4.000 ;
    END
  END pcpi_rd[21]
  PIN pcpi_rd[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 246.000 134.960 250.000 ;
    END
  END pcpi_rd[22]
  PIN pcpi_rd[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 246.000 131.600 250.000 ;
    END
  END pcpi_rd[23]
  PIN pcpi_rd[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END pcpi_rd[24]
  PIN pcpi_rd[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END pcpi_rd[25]
  PIN pcpi_rd[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 141.120 300.000 141.680 ;
    END
  END pcpi_rd[26]
  PIN pcpi_rd[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 246.000 171.920 250.000 ;
    END
  END pcpi_rd[27]
  PIN pcpi_rd[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 144.480 300.000 145.040 ;
    END
  END pcpi_rd[28]
  PIN pcpi_rd[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 124.320 300.000 124.880 ;
    END
  END pcpi_rd[29]
  PIN pcpi_rd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 87.360 300.000 87.920 ;
    END
  END pcpi_rd[2]
  PIN pcpi_rd[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 120.960 300.000 121.520 ;
    END
  END pcpi_rd[30]
  PIN pcpi_rd[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 97.440 300.000 98.000 ;
    END
  END pcpi_rd[31]
  PIN pcpi_rd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 100.800 300.000 101.360 ;
    END
  END pcpi_rd[3]
  PIN pcpi_rd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 90.720 300.000 91.280 ;
    END
  END pcpi_rd[4]
  PIN pcpi_rd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 0.000 175.280 4.000 ;
    END
  END pcpi_rd[5]
  PIN pcpi_rd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END pcpi_rd[6]
  PIN pcpi_rd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 94.080 300.000 94.640 ;
    END
  END pcpi_rd[7]
  PIN pcpi_rd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 114.240 300.000 114.800 ;
    END
  END pcpi_rd[8]
  PIN pcpi_rd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 77.280 300.000 77.840 ;
    END
  END pcpi_rd[9]
  PIN pcpi_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 117.600 300.000 118.160 ;
    END
  END pcpi_ready
  PIN pcpi_rs1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END pcpi_rs1[0]
  PIN pcpi_rs1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.040 4.000 47.600 ;
    END
  END pcpi_rs1[10]
  PIN pcpi_rs1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 4.000 44.240 ;
    END
  END pcpi_rs1[11]
  PIN pcpi_rs1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.840 4.000 64.400 ;
    END
  END pcpi_rs1[12]
  PIN pcpi_rs1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.200 4.000 67.760 ;
    END
  END pcpi_rs1[13]
  PIN pcpi_rs1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 4.000 71.120 ;
    END
  END pcpi_rs1[14]
  PIN pcpi_rs1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.640 4.000 81.200 ;
    END
  END pcpi_rs1[15]
  PIN pcpi_rs1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 246.000 87.920 250.000 ;
    END
  END pcpi_rs1[16]
  PIN pcpi_rs1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 246.000 64.400 250.000 ;
    END
  END pcpi_rs1[17]
  PIN pcpi_rs1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 246.000 61.040 250.000 ;
    END
  END pcpi_rs1[18]
  PIN pcpi_rs1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 4.000 218.960 ;
    END
  END pcpi_rs1[19]
  PIN pcpi_rs1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END pcpi_rs1[1]
  PIN pcpi_rs1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 4.000 212.240 ;
    END
  END pcpi_rs1[20]
  PIN pcpi_rs1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 208.320 4.000 208.880 ;
    END
  END pcpi_rs1[21]
  PIN pcpi_rs1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END pcpi_rs1[22]
  PIN pcpi_rs1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END pcpi_rs1[23]
  PIN pcpi_rs1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 246.000 222.320 250.000 ;
    END
  END pcpi_rs1[24]
  PIN pcpi_rs1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 246.000 225.680 250.000 ;
    END
  END pcpi_rs1[25]
  PIN pcpi_rs1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 246.000 215.600 250.000 ;
    END
  END pcpi_rs1[26]
  PIN pcpi_rs1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 246.000 208.880 250.000 ;
    END
  END pcpi_rs1[27]
  PIN pcpi_rs1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 246.000 185.360 250.000 ;
    END
  END pcpi_rs1[28]
  PIN pcpi_rs1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 246.000 198.800 250.000 ;
    END
  END pcpi_rs1[29]
  PIN pcpi_rs1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 0.000 188.720 4.000 ;
    END
  END pcpi_rs1[2]
  PIN pcpi_rs1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 246.000 218.960 250.000 ;
    END
  END pcpi_rs1[30]
  PIN pcpi_rs1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 246.000 202.160 250.000 ;
    END
  END pcpi_rs1[31]
  PIN pcpi_rs1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END pcpi_rs1[3]
  PIN pcpi_rs1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END pcpi_rs1[4]
  PIN pcpi_rs1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END pcpi_rs1[5]
  PIN pcpi_rs1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 0.000 182.000 4.000 ;
    END
  END pcpi_rs1[6]
  PIN pcpi_rs1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END pcpi_rs1[7]
  PIN pcpi_rs1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 4.000 57.680 ;
    END
  END pcpi_rs1[8]
  PIN pcpi_rs1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 4.000 61.040 ;
    END
  END pcpi_rs1[9]
  PIN pcpi_rs2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END pcpi_rs2[0]
  PIN pcpi_rs2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END pcpi_rs2[10]
  PIN pcpi_rs2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END pcpi_rs2[11]
  PIN pcpi_rs2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END pcpi_rs2[12]
  PIN pcpi_rs2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.400 4.000 50.960 ;
    END
  END pcpi_rs2[13]
  PIN pcpi_rs2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.320 4.000 40.880 ;
    END
  END pcpi_rs2[14]
  PIN pcpi_rs2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END pcpi_rs2[15]
  PIN pcpi_rs2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.240 4.000 198.800 ;
    END
  END pcpi_rs2[16]
  PIN pcpi_rs2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END pcpi_rs2[17]
  PIN pcpi_rs2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 4.000 205.520 ;
    END
  END pcpi_rs2[18]
  PIN pcpi_rs2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 4.000 178.640 ;
    END
  END pcpi_rs2[19]
  PIN pcpi_rs2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 4.000 ;
    END
  END pcpi_rs2[1]
  PIN pcpi_rs2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 246.000 50.960 250.000 ;
    END
  END pcpi_rs2[20]
  PIN pcpi_rs2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 246.000 47.600 250.000 ;
    END
  END pcpi_rs2[21]
  PIN pcpi_rs2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 246.000 84.560 250.000 ;
    END
  END pcpi_rs2[22]
  PIN pcpi_rs2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 246.000 91.280 250.000 ;
    END
  END pcpi_rs2[23]
  PIN pcpi_rs2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 246.000 195.440 250.000 ;
    END
  END pcpi_rs2[24]
  PIN pcpi_rs2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 246.000 192.080 250.000 ;
    END
  END pcpi_rs2[25]
  PIN pcpi_rs2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 246.000 188.720 250.000 ;
    END
  END pcpi_rs2[26]
  PIN pcpi_rs2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 246.000 151.760 250.000 ;
    END
  END pcpi_rs2[27]
  PIN pcpi_rs2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 246.000 205.520 250.000 ;
    END
  END pcpi_rs2[28]
  PIN pcpi_rs2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 246.000 212.240 250.000 ;
    END
  END pcpi_rs2[29]
  PIN pcpi_rs2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 0.000 134.960 4.000 ;
    END
  END pcpi_rs2[2]
  PIN pcpi_rs2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 246.000 232.400 250.000 ;
    END
  END pcpi_rs2[30]
  PIN pcpi_rs2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 246.000 229.040 250.000 ;
    END
  END pcpi_rs2[31]
  PIN pcpi_rs2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 0.000 148.400 4.000 ;
    END
  END pcpi_rs2[3]
  PIN pcpi_rs2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END pcpi_rs2[4]
  PIN pcpi_rs2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END pcpi_rs2[5]
  PIN pcpi_rs2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 0.000 198.800 4.000 ;
    END
  END pcpi_rs2[6]
  PIN pcpi_rs2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 0.000 215.600 4.000 ;
    END
  END pcpi_rs2[7]
  PIN pcpi_rs2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.280 4.000 77.840 ;
    END
  END pcpi_rs2[8]
  PIN pcpi_rs2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.920 4.000 74.480 ;
    END
  END pcpi_rs2[9]
  PIN pcpi_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 157.920 300.000 158.480 ;
    END
  END pcpi_valid
  PIN pcpi_wait
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 4.000 ;
    END
  END pcpi_wait
  PIN pcpi_wr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 131.040 300.000 131.600 ;
    END
  END pcpi_wr
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END resetn
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 231.580 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 231.580 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 235.050 ;
      LAYER Metal2 ;
        RECT 7.980 245.700 46.740 246.000 ;
        RECT 47.900 245.700 50.100 246.000 ;
        RECT 51.260 245.700 60.180 246.000 ;
        RECT 61.340 245.700 63.540 246.000 ;
        RECT 64.700 245.700 83.700 246.000 ;
        RECT 84.860 245.700 87.060 246.000 ;
        RECT 88.220 245.700 90.420 246.000 ;
        RECT 91.580 245.700 130.740 246.000 ;
        RECT 131.900 245.700 134.100 246.000 ;
        RECT 135.260 245.700 140.820 246.000 ;
        RECT 141.980 245.700 144.180 246.000 ;
        RECT 145.340 245.700 147.540 246.000 ;
        RECT 148.700 245.700 150.900 246.000 ;
        RECT 152.060 245.700 171.060 246.000 ;
        RECT 172.220 245.700 184.500 246.000 ;
        RECT 185.660 245.700 187.860 246.000 ;
        RECT 189.020 245.700 191.220 246.000 ;
        RECT 192.380 245.700 194.580 246.000 ;
        RECT 195.740 245.700 197.940 246.000 ;
        RECT 199.100 245.700 201.300 246.000 ;
        RECT 202.460 245.700 204.660 246.000 ;
        RECT 205.820 245.700 208.020 246.000 ;
        RECT 209.180 245.700 211.380 246.000 ;
        RECT 212.540 245.700 214.740 246.000 ;
        RECT 215.900 245.700 218.100 246.000 ;
        RECT 219.260 245.700 221.460 246.000 ;
        RECT 222.620 245.700 224.820 246.000 ;
        RECT 225.980 245.700 228.180 246.000 ;
        RECT 229.340 245.700 231.540 246.000 ;
        RECT 232.700 245.700 292.180 246.000 ;
        RECT 7.980 4.300 292.180 245.700 ;
        RECT 7.980 3.500 9.780 4.300 ;
        RECT 10.940 3.500 13.140 4.300 ;
        RECT 14.300 3.500 16.500 4.300 ;
        RECT 17.660 3.500 19.860 4.300 ;
        RECT 21.020 3.500 23.220 4.300 ;
        RECT 24.380 3.500 26.580 4.300 ;
        RECT 27.740 3.500 29.940 4.300 ;
        RECT 31.100 3.500 33.300 4.300 ;
        RECT 34.460 3.500 36.660 4.300 ;
        RECT 37.820 3.500 40.020 4.300 ;
        RECT 41.180 3.500 43.380 4.300 ;
        RECT 44.540 3.500 46.740 4.300 ;
        RECT 47.900 3.500 50.100 4.300 ;
        RECT 51.260 3.500 70.260 4.300 ;
        RECT 71.420 3.500 107.220 4.300 ;
        RECT 108.380 3.500 127.380 4.300 ;
        RECT 128.540 3.500 130.740 4.300 ;
        RECT 131.900 3.500 134.100 4.300 ;
        RECT 135.260 3.500 137.460 4.300 ;
        RECT 138.620 3.500 140.820 4.300 ;
        RECT 141.980 3.500 144.180 4.300 ;
        RECT 145.340 3.500 147.540 4.300 ;
        RECT 148.700 3.500 150.900 4.300 ;
        RECT 152.060 3.500 154.260 4.300 ;
        RECT 155.420 3.500 157.620 4.300 ;
        RECT 158.780 3.500 160.980 4.300 ;
        RECT 162.140 3.500 164.340 4.300 ;
        RECT 165.500 3.500 167.700 4.300 ;
        RECT 168.860 3.500 171.060 4.300 ;
        RECT 172.220 3.500 174.420 4.300 ;
        RECT 175.580 3.500 177.780 4.300 ;
        RECT 178.940 3.500 181.140 4.300 ;
        RECT 182.300 3.500 184.500 4.300 ;
        RECT 185.660 3.500 187.860 4.300 ;
        RECT 189.020 3.500 197.940 4.300 ;
        RECT 199.100 3.500 214.740 4.300 ;
        RECT 215.900 3.500 292.180 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 219.260 296.000 234.500 ;
        RECT 4.300 218.100 296.000 219.260 ;
        RECT 4.000 212.540 296.000 218.100 ;
        RECT 4.300 211.380 296.000 212.540 ;
        RECT 4.000 209.180 296.000 211.380 ;
        RECT 4.300 208.020 296.000 209.180 ;
        RECT 4.000 205.820 296.000 208.020 ;
        RECT 4.300 204.660 296.000 205.820 ;
        RECT 4.000 202.460 296.000 204.660 ;
        RECT 4.300 201.300 296.000 202.460 ;
        RECT 4.000 199.100 296.000 201.300 ;
        RECT 4.300 197.940 296.000 199.100 ;
        RECT 4.000 195.740 296.000 197.940 ;
        RECT 4.300 194.580 296.000 195.740 ;
        RECT 4.000 189.020 296.000 194.580 ;
        RECT 4.000 187.860 295.700 189.020 ;
        RECT 4.000 185.660 296.000 187.860 ;
        RECT 4.000 184.500 295.700 185.660 ;
        RECT 4.000 182.300 296.000 184.500 ;
        RECT 4.000 181.140 295.700 182.300 ;
        RECT 4.000 178.940 296.000 181.140 ;
        RECT 4.300 177.780 295.700 178.940 ;
        RECT 4.000 175.580 296.000 177.780 ;
        RECT 4.000 174.420 295.700 175.580 ;
        RECT 4.000 172.220 296.000 174.420 ;
        RECT 4.000 171.060 295.700 172.220 ;
        RECT 4.000 168.860 296.000 171.060 ;
        RECT 4.300 167.700 295.700 168.860 ;
        RECT 4.000 165.500 296.000 167.700 ;
        RECT 4.000 164.340 295.700 165.500 ;
        RECT 4.000 162.140 296.000 164.340 ;
        RECT 4.000 160.980 295.700 162.140 ;
        RECT 4.000 158.780 296.000 160.980 ;
        RECT 4.000 157.620 295.700 158.780 ;
        RECT 4.000 155.420 296.000 157.620 ;
        RECT 4.000 154.260 295.700 155.420 ;
        RECT 4.000 152.060 296.000 154.260 ;
        RECT 4.000 150.900 295.700 152.060 ;
        RECT 4.000 148.700 296.000 150.900 ;
        RECT 4.000 147.540 295.700 148.700 ;
        RECT 4.000 145.340 296.000 147.540 ;
        RECT 4.000 144.180 295.700 145.340 ;
        RECT 4.000 141.980 296.000 144.180 ;
        RECT 4.300 140.820 295.700 141.980 ;
        RECT 4.000 138.620 296.000 140.820 ;
        RECT 4.000 137.460 295.700 138.620 ;
        RECT 4.000 135.260 296.000 137.460 ;
        RECT 4.300 134.100 295.700 135.260 ;
        RECT 4.000 131.900 296.000 134.100 ;
        RECT 4.300 130.740 295.700 131.900 ;
        RECT 4.000 128.540 296.000 130.740 ;
        RECT 4.300 127.380 295.700 128.540 ;
        RECT 4.000 125.180 296.000 127.380 ;
        RECT 4.300 124.020 295.700 125.180 ;
        RECT 4.000 121.820 296.000 124.020 ;
        RECT 4.300 120.660 295.700 121.820 ;
        RECT 4.000 118.460 296.000 120.660 ;
        RECT 4.300 117.300 295.700 118.460 ;
        RECT 4.000 115.100 296.000 117.300 ;
        RECT 4.000 113.940 295.700 115.100 ;
        RECT 4.000 111.740 296.000 113.940 ;
        RECT 4.000 110.580 295.700 111.740 ;
        RECT 4.000 108.380 296.000 110.580 ;
        RECT 4.000 107.220 295.700 108.380 ;
        RECT 4.000 105.020 296.000 107.220 ;
        RECT 4.000 103.860 295.700 105.020 ;
        RECT 4.000 101.660 296.000 103.860 ;
        RECT 4.000 100.500 295.700 101.660 ;
        RECT 4.000 98.300 296.000 100.500 ;
        RECT 4.000 97.140 295.700 98.300 ;
        RECT 4.000 94.940 296.000 97.140 ;
        RECT 4.300 93.780 295.700 94.940 ;
        RECT 4.000 91.580 296.000 93.780 ;
        RECT 4.000 90.420 295.700 91.580 ;
        RECT 4.000 88.220 296.000 90.420 ;
        RECT 4.300 87.060 295.700 88.220 ;
        RECT 4.000 84.860 296.000 87.060 ;
        RECT 4.000 83.700 295.700 84.860 ;
        RECT 4.000 81.500 296.000 83.700 ;
        RECT 4.300 80.340 295.700 81.500 ;
        RECT 4.000 78.140 296.000 80.340 ;
        RECT 4.300 76.980 295.700 78.140 ;
        RECT 4.000 74.780 296.000 76.980 ;
        RECT 4.300 73.620 295.700 74.780 ;
        RECT 4.000 71.420 296.000 73.620 ;
        RECT 4.300 70.260 296.000 71.420 ;
        RECT 4.000 68.060 296.000 70.260 ;
        RECT 4.300 66.900 296.000 68.060 ;
        RECT 4.000 64.700 296.000 66.900 ;
        RECT 4.300 63.540 296.000 64.700 ;
        RECT 4.000 61.340 296.000 63.540 ;
        RECT 4.300 60.180 296.000 61.340 ;
        RECT 4.000 57.980 296.000 60.180 ;
        RECT 4.300 56.820 296.000 57.980 ;
        RECT 4.000 54.620 296.000 56.820 ;
        RECT 4.300 53.460 296.000 54.620 ;
        RECT 4.000 51.260 296.000 53.460 ;
        RECT 4.300 50.100 296.000 51.260 ;
        RECT 4.000 47.900 296.000 50.100 ;
        RECT 4.300 46.740 296.000 47.900 ;
        RECT 4.000 44.540 296.000 46.740 ;
        RECT 4.300 43.380 296.000 44.540 ;
        RECT 4.000 41.180 296.000 43.380 ;
        RECT 4.300 40.020 296.000 41.180 ;
        RECT 4.000 15.260 296.000 40.020 ;
      LAYER Metal4 ;
        RECT 48.300 15.210 98.740 174.070 ;
        RECT 100.940 15.210 175.540 174.070 ;
        RECT 177.740 15.210 191.940 174.070 ;
  END
END pcpi_approx_mul
END LIBRARY


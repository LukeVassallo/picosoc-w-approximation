VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pcpi_exact_mul
  CLASS BLOCK ;
  FOREIGN pcpi_exact_mul ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 215.040 4.000 215.600 ;
    END
  END clk
  PIN pcpi_insn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END pcpi_insn[0]
  PIN pcpi_insn[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END pcpi_insn[10]
  PIN pcpi_insn[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END pcpi_insn[11]
  PIN pcpi_insn[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 296.000 124.880 300.000 ;
    END
  END pcpi_insn[12]
  PIN pcpi_insn[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 296.000 131.600 300.000 ;
    END
  END pcpi_insn[13]
  PIN pcpi_insn[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 296.000 141.680 300.000 ;
    END
  END pcpi_insn[14]
  PIN pcpi_insn[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 0.000 7.280 4.000 ;
    END
  END pcpi_insn[15]
  PIN pcpi_insn[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END pcpi_insn[16]
  PIN pcpi_insn[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END pcpi_insn[17]
  PIN pcpi_insn[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 4.000 ;
    END
  END pcpi_insn[18]
  PIN pcpi_insn[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 0.000 20.720 4.000 ;
    END
  END pcpi_insn[19]
  PIN pcpi_insn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END pcpi_insn[1]
  PIN pcpi_insn[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END pcpi_insn[20]
  PIN pcpi_insn[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END pcpi_insn[21]
  PIN pcpi_insn[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END pcpi_insn[22]
  PIN pcpi_insn[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END pcpi_insn[23]
  PIN pcpi_insn[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END pcpi_insn[24]
  PIN pcpi_insn[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END pcpi_insn[25]
  PIN pcpi_insn[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END pcpi_insn[26]
  PIN pcpi_insn[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END pcpi_insn[27]
  PIN pcpi_insn[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 4.000 218.960 ;
    END
  END pcpi_insn[28]
  PIN pcpi_insn[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END pcpi_insn[29]
  PIN pcpi_insn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 4.000 57.680 ;
    END
  END pcpi_insn[2]
  PIN pcpi_insn[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END pcpi_insn[30]
  PIN pcpi_insn[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END pcpi_insn[31]
  PIN pcpi_insn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 4.000 61.040 ;
    END
  END pcpi_insn[3]
  PIN pcpi_insn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END pcpi_insn[4]
  PIN pcpi_insn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END pcpi_insn[5]
  PIN pcpi_insn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END pcpi_insn[6]
  PIN pcpi_insn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 0.000 40.880 4.000 ;
    END
  END pcpi_insn[7]
  PIN pcpi_insn[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END pcpi_insn[8]
  PIN pcpi_insn[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 4.000 ;
    END
  END pcpi_insn[9]
  PIN pcpi_rd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END pcpi_rd[0]
  PIN pcpi_rd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 4.000 212.240 ;
    END
  END pcpi_rd[10]
  PIN pcpi_rd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 296.000 171.920 300.000 ;
    END
  END pcpi_rd[11]
  PIN pcpi_rd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END pcpi_rd[12]
  PIN pcpi_rd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 296.000 161.840 300.000 ;
    END
  END pcpi_rd[13]
  PIN pcpi_rd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END pcpi_rd[14]
  PIN pcpi_rd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 0.000 134.960 4.000 ;
    END
  END pcpi_rd[15]
  PIN pcpi_rd[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.920 4.000 74.480 ;
    END
  END pcpi_rd[16]
  PIN pcpi_rd[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END pcpi_rd[17]
  PIN pcpi_rd[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 124.320 300.000 124.880 ;
    END
  END pcpi_rd[18]
  PIN pcpi_rd[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END pcpi_rd[19]
  PIN pcpi_rd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END pcpi_rd[1]
  PIN pcpi_rd[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 120.960 300.000 121.520 ;
    END
  END pcpi_rd[20]
  PIN pcpi_rd[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END pcpi_rd[21]
  PIN pcpi_rd[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END pcpi_rd[22]
  PIN pcpi_rd[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END pcpi_rd[23]
  PIN pcpi_rd[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 296.000 165.200 300.000 ;
    END
  END pcpi_rd[24]
  PIN pcpi_rd[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 178.080 300.000 178.640 ;
    END
  END pcpi_rd[25]
  PIN pcpi_rd[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 296.000 178.640 300.000 ;
    END
  END pcpi_rd[26]
  PIN pcpi_rd[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 296.000 121.520 300.000 ;
    END
  END pcpi_rd[27]
  PIN pcpi_rd[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 161.280 300.000 161.840 ;
    END
  END pcpi_rd[28]
  PIN pcpi_rd[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 134.400 300.000 134.960 ;
    END
  END pcpi_rd[29]
  PIN pcpi_rd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END pcpi_rd[2]
  PIN pcpi_rd[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 141.120 300.000 141.680 ;
    END
  END pcpi_rd[30]
  PIN pcpi_rd[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 137.760 300.000 138.320 ;
    END
  END pcpi_rd[31]
  PIN pcpi_rd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.840 4.000 148.400 ;
    END
  END pcpi_rd[3]
  PIN pcpi_rd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 296.000 128.240 300.000 ;
    END
  END pcpi_rd[4]
  PIN pcpi_rd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.240 4.000 198.800 ;
    END
  END pcpi_rd[5]
  PIN pcpi_rd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 296.000 158.480 300.000 ;
    END
  END pcpi_rd[6]
  PIN pcpi_rd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 296.000 138.320 300.000 ;
    END
  END pcpi_rd[7]
  PIN pcpi_rd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END pcpi_rd[8]
  PIN pcpi_rd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END pcpi_rd[9]
  PIN pcpi_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 154.560 300.000 155.120 ;
    END
  END pcpi_ready
  PIN pcpi_rs1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END pcpi_rs1[0]
  PIN pcpi_rs1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END pcpi_rs1[10]
  PIN pcpi_rs1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 0.000 175.280 4.000 ;
    END
  END pcpi_rs1[11]
  PIN pcpi_rs1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 0.000 198.800 4.000 ;
    END
  END pcpi_rs1[12]
  PIN pcpi_rs1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 0.000 215.600 4.000 ;
    END
  END pcpi_rs1[13]
  PIN pcpi_rs1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 0.000 235.760 4.000 ;
    END
  END pcpi_rs1[14]
  PIN pcpi_rs1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 0.000 249.200 4.000 ;
    END
  END pcpi_rs1[15]
  PIN pcpi_rs1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 4.000 84.560 ;
    END
  END pcpi_rs1[16]
  PIN pcpi_rs1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END pcpi_rs1[17]
  PIN pcpi_rs1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.840 4.000 64.400 ;
    END
  END pcpi_rs1[18]
  PIN pcpi_rs1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 4.000 71.120 ;
    END
  END pcpi_rs1[19]
  PIN pcpi_rs1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END pcpi_rs1[1]
  PIN pcpi_rs1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.200 4.000 67.760 ;
    END
  END pcpi_rs1[20]
  PIN pcpi_rs1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.280 4.000 77.840 ;
    END
  END pcpi_rs1[21]
  PIN pcpi_rs1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.400 4.000 50.960 ;
    END
  END pcpi_rs1[22]
  PIN pcpi_rs1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 4.000 44.240 ;
    END
  END pcpi_rs1[23]
  PIN pcpi_rs1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 296.000 145.040 300.000 ;
    END
  END pcpi_rs1[24]
  PIN pcpi_rs1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 296.000 148.400 300.000 ;
    END
  END pcpi_rs1[25]
  PIN pcpi_rs1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 296.000 151.760 300.000 ;
    END
  END pcpi_rs1[26]
  PIN pcpi_rs1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 296.000 192.080 300.000 ;
    END
  END pcpi_rs1[27]
  PIN pcpi_rs1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 296.000 185.360 300.000 ;
    END
  END pcpi_rs1[28]
  PIN pcpi_rs1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 296.000 188.720 300.000 ;
    END
  END pcpi_rs1[29]
  PIN pcpi_rs1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.280 4.000 161.840 ;
    END
  END pcpi_rs1[2]
  PIN pcpi_rs1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 296.000 249.200 300.000 ;
    END
  END pcpi_rs1[30]
  PIN pcpi_rs1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 296.000 252.560 300.000 ;
    END
  END pcpi_rs1[31]
  PIN pcpi_rs1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 4.000 178.640 ;
    END
  END pcpi_rs1[3]
  PIN pcpi_rs1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 4.000 205.520 ;
    END
  END pcpi_rs1[4]
  PIN pcpi_rs1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.120 4.000 225.680 ;
    END
  END pcpi_rs1[5]
  PIN pcpi_rs1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END pcpi_rs1[6]
  PIN pcpi_rs1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 4.000 252.560 ;
    END
  END pcpi_rs1[7]
  PIN pcpi_rs1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END pcpi_rs1[8]
  PIN pcpi_rs1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END pcpi_rs1[9]
  PIN pcpi_rs2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.720 4.000 175.280 ;
    END
  END pcpi_rs2[0]
  PIN pcpi_rs2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 0.000 182.000 4.000 ;
    END
  END pcpi_rs2[10]
  PIN pcpi_rs2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 0.000 188.720 4.000 ;
    END
  END pcpi_rs2[11]
  PIN pcpi_rs2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 0.000 195.440 4.000 ;
    END
  END pcpi_rs2[12]
  PIN pcpi_rs2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END pcpi_rs2[13]
  PIN pcpi_rs2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 107.520 300.000 108.080 ;
    END
  END pcpi_rs2[14]
  PIN pcpi_rs2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 117.600 300.000 118.160 ;
    END
  END pcpi_rs2[15]
  PIN pcpi_rs2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END pcpi_rs2[16]
  PIN pcpi_rs2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.440 4.000 98.000 ;
    END
  END pcpi_rs2[17]
  PIN pcpi_rs2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END pcpi_rs2[18]
  PIN pcpi_rs2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.640 4.000 81.200 ;
    END
  END pcpi_rs2[19]
  PIN pcpi_rs2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END pcpi_rs2[1]
  PIN pcpi_rs2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END pcpi_rs2[20]
  PIN pcpi_rs2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END pcpi_rs2[21]
  PIN pcpi_rs2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END pcpi_rs2[22]
  PIN pcpi_rs2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END pcpi_rs2[23]
  PIN pcpi_rs2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 296.000 134.960 300.000 ;
    END
  END pcpi_rs2[24]
  PIN pcpi_rs2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 296.000 155.120 300.000 ;
    END
  END pcpi_rs2[25]
  PIN pcpi_rs2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 296.000 168.560 300.000 ;
    END
  END pcpi_rs2[26]
  PIN pcpi_rs2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 296.000 182.000 300.000 ;
    END
  END pcpi_rs2[27]
  PIN pcpi_rs2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 296.000 175.280 300.000 ;
    END
  END pcpi_rs2[28]
  PIN pcpi_rs2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 296.000 202.160 300.000 ;
    END
  END pcpi_rs2[29]
  PIN pcpi_rs2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.440 4.000 182.000 ;
    END
  END pcpi_rs2[2]
  PIN pcpi_rs2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 184.800 300.000 185.360 ;
    END
  END pcpi_rs2[30]
  PIN pcpi_rs2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 174.720 300.000 175.280 ;
    END
  END pcpi_rs2[31]
  PIN pcpi_rs2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 171.360 4.000 171.920 ;
    END
  END pcpi_rs2[3]
  PIN pcpi_rs2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 4.000 192.080 ;
    END
  END pcpi_rs2[4]
  PIN pcpi_rs2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 208.320 4.000 208.880 ;
    END
  END pcpi_rs2[5]
  PIN pcpi_rs2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END pcpi_rs2[6]
  PIN pcpi_rs2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 296.000 118.160 300.000 ;
    END
  END pcpi_rs2[7]
  PIN pcpi_rs2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END pcpi_rs2[8]
  PIN pcpi_rs2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END pcpi_rs2[9]
  PIN pcpi_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END pcpi_valid
  PIN pcpi_wait
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END pcpi_wait
  PIN pcpi_wr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 157.920 300.000 158.480 ;
    END
  END pcpi_wr
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END resetn
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 283.770 ;
      LAYER Metal2 ;
        RECT 6.300 295.700 117.300 296.660 ;
        RECT 118.460 295.700 120.660 296.660 ;
        RECT 121.820 295.700 124.020 296.660 ;
        RECT 125.180 295.700 127.380 296.660 ;
        RECT 128.540 295.700 130.740 296.660 ;
        RECT 131.900 295.700 134.100 296.660 ;
        RECT 135.260 295.700 137.460 296.660 ;
        RECT 138.620 295.700 140.820 296.660 ;
        RECT 141.980 295.700 144.180 296.660 ;
        RECT 145.340 295.700 147.540 296.660 ;
        RECT 148.700 295.700 150.900 296.660 ;
        RECT 152.060 295.700 154.260 296.660 ;
        RECT 155.420 295.700 157.620 296.660 ;
        RECT 158.780 295.700 160.980 296.660 ;
        RECT 162.140 295.700 164.340 296.660 ;
        RECT 165.500 295.700 167.700 296.660 ;
        RECT 168.860 295.700 171.060 296.660 ;
        RECT 172.220 295.700 174.420 296.660 ;
        RECT 175.580 295.700 177.780 296.660 ;
        RECT 178.940 295.700 181.140 296.660 ;
        RECT 182.300 295.700 184.500 296.660 ;
        RECT 185.660 295.700 187.860 296.660 ;
        RECT 189.020 295.700 191.220 296.660 ;
        RECT 192.380 295.700 201.300 296.660 ;
        RECT 202.460 295.700 248.340 296.660 ;
        RECT 249.500 295.700 251.700 296.660 ;
        RECT 252.860 295.700 291.620 296.660 ;
        RECT 6.300 4.300 291.620 295.700 ;
        RECT 6.300 4.000 6.420 4.300 ;
        RECT 7.580 4.000 9.780 4.300 ;
        RECT 10.940 4.000 13.140 4.300 ;
        RECT 14.300 4.000 16.500 4.300 ;
        RECT 17.660 4.000 19.860 4.300 ;
        RECT 21.020 4.000 23.220 4.300 ;
        RECT 24.380 4.000 26.580 4.300 ;
        RECT 27.740 4.000 29.940 4.300 ;
        RECT 31.100 4.000 33.300 4.300 ;
        RECT 34.460 4.000 36.660 4.300 ;
        RECT 37.820 4.000 40.020 4.300 ;
        RECT 41.180 4.000 43.380 4.300 ;
        RECT 44.540 4.000 46.740 4.300 ;
        RECT 47.900 4.000 50.100 4.300 ;
        RECT 51.260 4.000 97.140 4.300 ;
        RECT 98.300 4.000 110.580 4.300 ;
        RECT 111.740 4.000 124.020 4.300 ;
        RECT 125.180 4.000 134.100 4.300 ;
        RECT 135.260 4.000 140.820 4.300 ;
        RECT 141.980 4.000 144.180 4.300 ;
        RECT 145.340 4.000 150.900 4.300 ;
        RECT 152.060 4.000 154.260 4.300 ;
        RECT 155.420 4.000 157.620 4.300 ;
        RECT 158.780 4.000 160.980 4.300 ;
        RECT 162.140 4.000 164.340 4.300 ;
        RECT 165.500 4.000 167.700 4.300 ;
        RECT 168.860 4.000 171.060 4.300 ;
        RECT 172.220 4.000 174.420 4.300 ;
        RECT 175.580 4.000 177.780 4.300 ;
        RECT 178.940 4.000 181.140 4.300 ;
        RECT 182.300 4.000 184.500 4.300 ;
        RECT 185.660 4.000 187.860 4.300 ;
        RECT 189.020 4.000 191.220 4.300 ;
        RECT 192.380 4.000 194.580 4.300 ;
        RECT 195.740 4.000 197.940 4.300 ;
        RECT 199.100 4.000 214.740 4.300 ;
        RECT 215.900 4.000 234.900 4.300 ;
        RECT 236.060 4.000 248.340 4.300 ;
        RECT 249.500 4.000 291.620 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 252.860 296.000 282.380 ;
        RECT 4.300 251.700 296.000 252.860 ;
        RECT 4.000 225.980 296.000 251.700 ;
        RECT 4.300 224.820 296.000 225.980 ;
        RECT 4.000 222.620 296.000 224.820 ;
        RECT 4.300 221.460 296.000 222.620 ;
        RECT 4.000 219.260 296.000 221.460 ;
        RECT 4.300 218.100 296.000 219.260 ;
        RECT 4.000 215.900 296.000 218.100 ;
        RECT 4.300 214.740 296.000 215.900 ;
        RECT 4.000 212.540 296.000 214.740 ;
        RECT 4.300 211.380 296.000 212.540 ;
        RECT 4.000 209.180 296.000 211.380 ;
        RECT 4.300 208.020 296.000 209.180 ;
        RECT 4.000 205.820 296.000 208.020 ;
        RECT 4.300 204.660 296.000 205.820 ;
        RECT 4.000 202.460 296.000 204.660 ;
        RECT 4.300 201.300 296.000 202.460 ;
        RECT 4.000 199.100 296.000 201.300 ;
        RECT 4.300 197.940 296.000 199.100 ;
        RECT 4.000 195.740 296.000 197.940 ;
        RECT 4.300 194.580 296.000 195.740 ;
        RECT 4.000 192.380 296.000 194.580 ;
        RECT 4.300 191.220 296.000 192.380 ;
        RECT 4.000 189.020 296.000 191.220 ;
        RECT 4.300 187.860 296.000 189.020 ;
        RECT 4.000 185.660 296.000 187.860 ;
        RECT 4.300 184.500 295.700 185.660 ;
        RECT 4.000 182.300 296.000 184.500 ;
        RECT 4.300 181.140 296.000 182.300 ;
        RECT 4.000 178.940 296.000 181.140 ;
        RECT 4.300 177.780 295.700 178.940 ;
        RECT 4.000 175.580 296.000 177.780 ;
        RECT 4.300 174.420 295.700 175.580 ;
        RECT 4.000 172.220 296.000 174.420 ;
        RECT 4.300 171.060 296.000 172.220 ;
        RECT 4.000 168.860 296.000 171.060 ;
        RECT 4.300 167.700 296.000 168.860 ;
        RECT 4.000 165.500 296.000 167.700 ;
        RECT 4.300 164.340 296.000 165.500 ;
        RECT 4.000 162.140 296.000 164.340 ;
        RECT 4.300 160.980 295.700 162.140 ;
        RECT 4.000 158.780 296.000 160.980 ;
        RECT 4.300 157.620 295.700 158.780 ;
        RECT 4.000 155.420 296.000 157.620 ;
        RECT 4.300 154.260 295.700 155.420 ;
        RECT 4.000 152.060 296.000 154.260 ;
        RECT 4.300 150.900 296.000 152.060 ;
        RECT 4.000 148.700 296.000 150.900 ;
        RECT 4.300 147.540 296.000 148.700 ;
        RECT 4.000 145.340 296.000 147.540 ;
        RECT 4.300 144.180 296.000 145.340 ;
        RECT 4.000 141.980 296.000 144.180 ;
        RECT 4.300 140.820 295.700 141.980 ;
        RECT 4.000 138.620 296.000 140.820 ;
        RECT 4.300 137.460 295.700 138.620 ;
        RECT 4.000 135.260 296.000 137.460 ;
        RECT 4.300 134.100 295.700 135.260 ;
        RECT 4.000 131.900 296.000 134.100 ;
        RECT 4.300 130.740 296.000 131.900 ;
        RECT 4.000 128.540 296.000 130.740 ;
        RECT 4.300 127.380 296.000 128.540 ;
        RECT 4.000 125.180 296.000 127.380 ;
        RECT 4.300 124.020 295.700 125.180 ;
        RECT 4.000 121.820 296.000 124.020 ;
        RECT 4.300 120.660 295.700 121.820 ;
        RECT 4.000 118.460 296.000 120.660 ;
        RECT 4.300 117.300 295.700 118.460 ;
        RECT 4.000 115.100 296.000 117.300 ;
        RECT 4.300 113.940 296.000 115.100 ;
        RECT 4.000 111.740 296.000 113.940 ;
        RECT 4.300 110.580 296.000 111.740 ;
        RECT 4.000 108.380 296.000 110.580 ;
        RECT 4.300 107.220 295.700 108.380 ;
        RECT 4.000 105.020 296.000 107.220 ;
        RECT 4.300 103.860 296.000 105.020 ;
        RECT 4.000 101.660 296.000 103.860 ;
        RECT 4.300 100.500 296.000 101.660 ;
        RECT 4.000 98.300 296.000 100.500 ;
        RECT 4.300 97.140 296.000 98.300 ;
        RECT 4.000 94.940 296.000 97.140 ;
        RECT 4.300 93.780 296.000 94.940 ;
        RECT 4.000 91.580 296.000 93.780 ;
        RECT 4.300 90.420 296.000 91.580 ;
        RECT 4.000 88.220 296.000 90.420 ;
        RECT 4.300 87.060 296.000 88.220 ;
        RECT 4.000 84.860 296.000 87.060 ;
        RECT 4.300 83.700 296.000 84.860 ;
        RECT 4.000 81.500 296.000 83.700 ;
        RECT 4.300 80.340 296.000 81.500 ;
        RECT 4.000 78.140 296.000 80.340 ;
        RECT 4.300 76.980 296.000 78.140 ;
        RECT 4.000 74.780 296.000 76.980 ;
        RECT 4.300 73.620 296.000 74.780 ;
        RECT 4.000 71.420 296.000 73.620 ;
        RECT 4.300 70.260 296.000 71.420 ;
        RECT 4.000 68.060 296.000 70.260 ;
        RECT 4.300 66.900 296.000 68.060 ;
        RECT 4.000 64.700 296.000 66.900 ;
        RECT 4.300 63.540 296.000 64.700 ;
        RECT 4.000 61.340 296.000 63.540 ;
        RECT 4.300 60.180 296.000 61.340 ;
        RECT 4.000 57.980 296.000 60.180 ;
        RECT 4.300 56.820 296.000 57.980 ;
        RECT 4.000 54.620 296.000 56.820 ;
        RECT 4.300 53.460 296.000 54.620 ;
        RECT 4.000 51.260 296.000 53.460 ;
        RECT 4.300 50.100 296.000 51.260 ;
        RECT 4.000 44.540 296.000 50.100 ;
        RECT 4.300 43.380 296.000 44.540 ;
        RECT 4.000 12.460 296.000 43.380 ;
      LAYER Metal4 ;
        RECT 8.540 65.050 21.940 272.630 ;
        RECT 24.140 65.050 98.740 272.630 ;
        RECT 100.940 65.050 175.540 272.630 ;
        RECT 177.740 65.050 244.580 272.630 ;
  END
END pcpi_exact_mul
END LIBRARY


* NGSPICE file created from user_project_wrapper.ext - technology: gf180mcuD

* Black-box entry subcircuit for user_proj_example abstract view
.subckt user_proj_example io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12]
+ la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18]
+ la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23]
+ la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29]
+ la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34]
+ la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3]
+ la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45]
+ la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50]
+ la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56]
+ la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61]
+ la_data_in[62] la_data_in[63] la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9]
+ la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vdd vss wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for simple_interconnect abstract view
.subckt simple_interconnect clk gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[1] gpio_in[2] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6]
+ gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12]
+ gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[1] gpio_oeb[2] gpio_oeb[3] gpio_oeb[4]
+ gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10]
+ gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[1] gpio_out[2]
+ gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9]
+ mem_addr[0] mem_addr[10] mem_addr[11] mem_addr[12] mem_addr[13] mem_addr[14] mem_addr[15]
+ mem_addr[16] mem_addr[17] mem_addr[18] mem_addr[19] mem_addr[1] mem_addr[20] mem_addr[21]
+ mem_addr[22] mem_addr[23] mem_addr[24] mem_addr[25] mem_addr[26] mem_addr[27] mem_addr[28]
+ mem_addr[29] mem_addr[2] mem_addr[30] mem_addr[31] mem_addr[3] mem_addr[4] mem_addr[5]
+ mem_addr[6] mem_addr[7] mem_addr[8] mem_addr[9] mem_instr mem_rdata[0] mem_rdata[10]
+ mem_rdata[11] mem_rdata[12] mem_rdata[13] mem_rdata[14] mem_rdata[15] mem_rdata[16]
+ mem_rdata[17] mem_rdata[18] mem_rdata[19] mem_rdata[1] mem_rdata[20] mem_rdata[21]
+ mem_rdata[22] mem_rdata[23] mem_rdata[24] mem_rdata[25] mem_rdata[26] mem_rdata[27]
+ mem_rdata[28] mem_rdata[29] mem_rdata[2] mem_rdata[30] mem_rdata[31] mem_rdata[3]
+ mem_rdata[4] mem_rdata[5] mem_rdata[6] mem_rdata[7] mem_rdata[8] mem_rdata[9] mem_ready
+ mem_valid mem_wdata[0] mem_wdata[10] mem_wdata[11] mem_wdata[12] mem_wdata[13] mem_wdata[14]
+ mem_wdata[15] mem_wdata[16] mem_wdata[17] mem_wdata[18] mem_wdata[19] mem_wdata[1]
+ mem_wdata[20] mem_wdata[21] mem_wdata[22] mem_wdata[23] mem_wdata[24] mem_wdata[25]
+ mem_wdata[26] mem_wdata[27] mem_wdata[28] mem_wdata[29] mem_wdata[2] mem_wdata[30]
+ mem_wdata[31] mem_wdata[3] mem_wdata[4] mem_wdata[5] mem_wdata[6] mem_wdata[7] mem_wdata[8]
+ mem_wdata[9] mem_wstrb[0] mem_wstrb[1] mem_wstrb[2] mem_wstrb[3] ram_gwenb[0] ram_gwenb[1]
+ ram_gwenb[2] ram_gwenb[3] ram_rdata[0] ram_rdata[10] ram_rdata[11] ram_rdata[12]
+ ram_rdata[13] ram_rdata[14] ram_rdata[15] ram_rdata[16] ram_rdata[17] ram_rdata[18]
+ ram_rdata[19] ram_rdata[1] ram_rdata[20] ram_rdata[21] ram_rdata[22] ram_rdata[23]
+ ram_rdata[24] ram_rdata[25] ram_rdata[26] ram_rdata[27] ram_rdata[28] ram_rdata[29]
+ ram_rdata[2] ram_rdata[30] ram_rdata[31] ram_rdata[3] ram_rdata[4] ram_rdata[5]
+ ram_rdata[6] ram_rdata[7] ram_rdata[8] ram_rdata[9] ram_wenb[0] ram_wenb[10] ram_wenb[11]
+ ram_wenb[12] ram_wenb[13] ram_wenb[14] ram_wenb[15] ram_wenb[16] ram_wenb[17] ram_wenb[18]
+ ram_wenb[19] ram_wenb[1] ram_wenb[20] ram_wenb[21] ram_wenb[22] ram_wenb[23] ram_wenb[24]
+ ram_wenb[25] ram_wenb[26] ram_wenb[27] ram_wenb[28] ram_wenb[29] ram_wenb[2] ram_wenb[30]
+ ram_wenb[31] ram_wenb[3] ram_wenb[4] ram_wenb[5] ram_wenb[6] ram_wenb[7] ram_wenb[8]
+ ram_wenb[9] resetn simpleuart_dat_re simpleuart_dat_we simpleuart_div_we[0] simpleuart_div_we[1]
+ simpleuart_div_we[2] simpleuart_div_we[3] simpleuart_reg_dat_do[0] simpleuart_reg_dat_do[10]
+ simpleuart_reg_dat_do[11] simpleuart_reg_dat_do[12] simpleuart_reg_dat_do[13] simpleuart_reg_dat_do[14]
+ simpleuart_reg_dat_do[15] simpleuart_reg_dat_do[16] simpleuart_reg_dat_do[17] simpleuart_reg_dat_do[18]
+ simpleuart_reg_dat_do[19] simpleuart_reg_dat_do[1] simpleuart_reg_dat_do[20] simpleuart_reg_dat_do[21]
+ simpleuart_reg_dat_do[22] simpleuart_reg_dat_do[23] simpleuart_reg_dat_do[24] simpleuart_reg_dat_do[25]
+ simpleuart_reg_dat_do[26] simpleuart_reg_dat_do[27] simpleuart_reg_dat_do[28] simpleuart_reg_dat_do[29]
+ simpleuart_reg_dat_do[2] simpleuart_reg_dat_do[30] simpleuart_reg_dat_do[31] simpleuart_reg_dat_do[3]
+ simpleuart_reg_dat_do[4] simpleuart_reg_dat_do[5] simpleuart_reg_dat_do[6] simpleuart_reg_dat_do[7]
+ simpleuart_reg_dat_do[8] simpleuart_reg_dat_do[9] simpleuart_reg_dat_wait simpleuart_reg_div_do[0]
+ simpleuart_reg_div_do[10] simpleuart_reg_div_do[11] simpleuart_reg_div_do[12] simpleuart_reg_div_do[13]
+ simpleuart_reg_div_do[14] simpleuart_reg_div_do[15] simpleuart_reg_div_do[16] simpleuart_reg_div_do[17]
+ simpleuart_reg_div_do[18] simpleuart_reg_div_do[19] simpleuart_reg_div_do[1] simpleuart_reg_div_do[20]
+ simpleuart_reg_div_do[21] simpleuart_reg_div_do[22] simpleuart_reg_div_do[23] simpleuart_reg_div_do[24]
+ simpleuart_reg_div_do[25] simpleuart_reg_div_do[26] simpleuart_reg_div_do[27] simpleuart_reg_div_do[28]
+ simpleuart_reg_div_do[29] simpleuart_reg_div_do[2] simpleuart_reg_div_do[30] simpleuart_reg_div_do[31]
+ simpleuart_reg_div_do[3] simpleuart_reg_div_do[4] simpleuart_reg_div_do[5] simpleuart_reg_div_do[6]
+ simpleuart_reg_div_do[7] simpleuart_reg_div_do[8] simpleuart_reg_div_do[9] spimem_rdata[0]
+ spimem_rdata[10] spimem_rdata[11] spimem_rdata[12] spimem_rdata[13] spimem_rdata[14]
+ spimem_rdata[15] spimem_rdata[16] spimem_rdata[17] spimem_rdata[18] spimem_rdata[19]
+ spimem_rdata[1] spimem_rdata[20] spimem_rdata[21] spimem_rdata[22] spimem_rdata[23]
+ spimem_rdata[24] spimem_rdata[25] spimem_rdata[26] spimem_rdata[27] spimem_rdata[28]
+ spimem_rdata[29] spimem_rdata[2] spimem_rdata[30] spimem_rdata[31] spimem_rdata[3]
+ spimem_rdata[4] spimem_rdata[5] spimem_rdata[6] spimem_rdata[7] spimem_rdata[8]
+ spimem_rdata[9] spimem_ready spimem_valid spimemio_cfgreg_do[0] spimemio_cfgreg_do[10]
+ spimemio_cfgreg_do[11] spimemio_cfgreg_do[12] spimemio_cfgreg_do[13] spimemio_cfgreg_do[14]
+ spimemio_cfgreg_do[15] spimemio_cfgreg_do[16] spimemio_cfgreg_do[17] spimemio_cfgreg_do[18]
+ spimemio_cfgreg_do[19] spimemio_cfgreg_do[1] spimemio_cfgreg_do[20] spimemio_cfgreg_do[21]
+ spimemio_cfgreg_do[22] spimemio_cfgreg_do[23] spimemio_cfgreg_do[24] spimemio_cfgreg_do[25]
+ spimemio_cfgreg_do[26] spimemio_cfgreg_do[27] spimemio_cfgreg_do[28] spimemio_cfgreg_do[29]
+ spimemio_cfgreg_do[2] spimemio_cfgreg_do[30] spimemio_cfgreg_do[31] spimemio_cfgreg_do[3]
+ spimemio_cfgreg_do[4] spimemio_cfgreg_do[5] spimemio_cfgreg_do[6] spimemio_cfgreg_do[7]
+ spimemio_cfgreg_do[8] spimemio_cfgreg_do[9] spimemio_cfgreg_we[0] spimemio_cfgreg_we[1]
+ spimemio_cfgreg_we[2] spimemio_cfgreg_we[3] vdd vss
.ends

* Black-box entry subcircuit for gf180_ram_512x8x1 abstract view
.subckt gf180_ram_512x8x1 VDD VSS addr[0] addr[1] addr[2] addr[3] addr[4] addr[5]
+ addr[6] addr[7] addr[8] cen clk gwen rdata[0] rdata[1] rdata[2] rdata[3] rdata[4]
+ rdata[5] rdata[6] rdata[7] wdata[0] wdata[1] wdata[2] wdata[3] wdata[4] wdata[5]
+ wdata[6] wdata[7] wen[0] wen[1] wen[2] wen[3] wen[4] wen[5] wen[6] wen[7]
.ends

* Black-box entry subcircuit for pcpi_approx_mul abstract view
.subckt pcpi_approx_mul clk pcpi_insn[0] pcpi_insn[10] pcpi_insn[11] pcpi_insn[12]
+ pcpi_insn[13] pcpi_insn[14] pcpi_insn[15] pcpi_insn[16] pcpi_insn[17] pcpi_insn[18]
+ pcpi_insn[19] pcpi_insn[1] pcpi_insn[20] pcpi_insn[21] pcpi_insn[22] pcpi_insn[23]
+ pcpi_insn[24] pcpi_insn[25] pcpi_insn[26] pcpi_insn[27] pcpi_insn[28] pcpi_insn[29]
+ pcpi_insn[2] pcpi_insn[30] pcpi_insn[31] pcpi_insn[3] pcpi_insn[4] pcpi_insn[5]
+ pcpi_insn[6] pcpi_insn[7] pcpi_insn[8] pcpi_insn[9] pcpi_rd[0] pcpi_rd[10] pcpi_rd[11]
+ pcpi_rd[12] pcpi_rd[13] pcpi_rd[14] pcpi_rd[15] pcpi_rd[16] pcpi_rd[17] pcpi_rd[18]
+ pcpi_rd[19] pcpi_rd[1] pcpi_rd[20] pcpi_rd[21] pcpi_rd[22] pcpi_rd[23] pcpi_rd[24]
+ pcpi_rd[25] pcpi_rd[26] pcpi_rd[27] pcpi_rd[28] pcpi_rd[29] pcpi_rd[2] pcpi_rd[30]
+ pcpi_rd[31] pcpi_rd[3] pcpi_rd[4] pcpi_rd[5] pcpi_rd[6] pcpi_rd[7] pcpi_rd[8] pcpi_rd[9]
+ pcpi_ready pcpi_rs1[0] pcpi_rs1[10] pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14]
+ pcpi_rs1[15] pcpi_rs1[16] pcpi_rs1[17] pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20]
+ pcpi_rs1[21] pcpi_rs1[22] pcpi_rs1[23] pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27]
+ pcpi_rs1[28] pcpi_rs1[29] pcpi_rs1[2] pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4]
+ pcpi_rs1[5] pcpi_rs1[6] pcpi_rs1[7] pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10]
+ pcpi_rs2[11] pcpi_rs2[12] pcpi_rs2[13] pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17]
+ pcpi_rs2[18] pcpi_rs2[19] pcpi_rs2[1] pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23]
+ pcpi_rs2[24] pcpi_rs2[25] pcpi_rs2[26] pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2]
+ pcpi_rs2[30] pcpi_rs2[31] pcpi_rs2[3] pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7]
+ pcpi_rs2[8] pcpi_rs2[9] pcpi_valid pcpi_wait pcpi_wr resetn vdd vss
.ends

* Black-box entry subcircuit for pcpi_mul abstract view
.subckt pcpi_mul clk pcpi_insn[0] pcpi_insn[10] pcpi_insn[11] pcpi_insn[12] pcpi_insn[13]
+ pcpi_insn[14] pcpi_insn[15] pcpi_insn[16] pcpi_insn[17] pcpi_insn[18] pcpi_insn[19]
+ pcpi_insn[1] pcpi_insn[20] pcpi_insn[21] pcpi_insn[22] pcpi_insn[23] pcpi_insn[24]
+ pcpi_insn[25] pcpi_insn[26] pcpi_insn[27] pcpi_insn[28] pcpi_insn[29] pcpi_insn[2]
+ pcpi_insn[30] pcpi_insn[31] pcpi_insn[3] pcpi_insn[4] pcpi_insn[5] pcpi_insn[6]
+ pcpi_insn[7] pcpi_insn[8] pcpi_insn[9] pcpi_mul_rd[0] pcpi_mul_rd[10] pcpi_mul_rd[11]
+ pcpi_mul_rd[12] pcpi_mul_rd[13] pcpi_mul_rd[14] pcpi_mul_rd[15] pcpi_mul_rd[16]
+ pcpi_mul_rd[17] pcpi_mul_rd[18] pcpi_mul_rd[19] pcpi_mul_rd[1] pcpi_mul_rd[20] pcpi_mul_rd[21]
+ pcpi_mul_rd[22] pcpi_mul_rd[23] pcpi_mul_rd[24] pcpi_mul_rd[25] pcpi_mul_rd[26]
+ pcpi_mul_rd[27] pcpi_mul_rd[28] pcpi_mul_rd[29] pcpi_mul_rd[2] pcpi_mul_rd[30] pcpi_mul_rd[31]
+ pcpi_mul_rd[3] pcpi_mul_rd[4] pcpi_mul_rd[5] pcpi_mul_rd[6] pcpi_mul_rd[7] pcpi_mul_rd[8]
+ pcpi_mul_rd[9] pcpi_mul_ready pcpi_mul_valid pcpi_mul_wait pcpi_mul_wr pcpi_rs1[0]
+ pcpi_rs1[10] pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14] pcpi_rs1[15] pcpi_rs1[16]
+ pcpi_rs1[17] pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20] pcpi_rs1[21] pcpi_rs1[22]
+ pcpi_rs1[23] pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27] pcpi_rs1[28] pcpi_rs1[29]
+ pcpi_rs1[2] pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4] pcpi_rs1[5] pcpi_rs1[6]
+ pcpi_rs1[7] pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10] pcpi_rs2[11] pcpi_rs2[12]
+ pcpi_rs2[13] pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17] pcpi_rs2[18] pcpi_rs2[19]
+ pcpi_rs2[1] pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23] pcpi_rs2[24] pcpi_rs2[25]
+ pcpi_rs2[26] pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2] pcpi_rs2[30] pcpi_rs2[31]
+ pcpi_rs2[3] pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7] pcpi_rs2[8] pcpi_rs2[9]
+ resetn vdd vss
.ends

* Black-box entry subcircuit for ctrl abstract view
.subckt ctrl ctrl_in[0] ctrl_in[1] ctrl_oeb[0] ctrl_oeb[1] ctrl_out[0] ctrl_out[1]
+ reset resetn vdd vss
.ends

* Black-box entry subcircuit for cpu abstract view
.subckt cpu clk irq_in[0] irq_in[1] irq_in[2] irq_in[3] irq_oeb[0] irq_oeb[1] irq_oeb[2]
+ irq_oeb[3] irq_out[0] irq_out[1] irq_out[2] irq_out[3] mem_addr[0] mem_addr[10]
+ mem_addr[11] mem_addr[12] mem_addr[13] mem_addr[14] mem_addr[15] mem_addr[16] mem_addr[17]
+ mem_addr[18] mem_addr[19] mem_addr[1] mem_addr[20] mem_addr[21] mem_addr[22] mem_addr[23]
+ mem_addr[24] mem_addr[25] mem_addr[26] mem_addr[27] mem_addr[28] mem_addr[29] mem_addr[2]
+ mem_addr[30] mem_addr[31] mem_addr[3] mem_addr[4] mem_addr[5] mem_addr[6] mem_addr[7]
+ mem_addr[8] mem_addr[9] mem_instr mem_rdata[0] mem_rdata[10] mem_rdata[11] mem_rdata[12]
+ mem_rdata[13] mem_rdata[14] mem_rdata[15] mem_rdata[16] mem_rdata[17] mem_rdata[18]
+ mem_rdata[19] mem_rdata[1] mem_rdata[20] mem_rdata[21] mem_rdata[22] mem_rdata[23]
+ mem_rdata[24] mem_rdata[25] mem_rdata[26] mem_rdata[27] mem_rdata[28] mem_rdata[29]
+ mem_rdata[2] mem_rdata[30] mem_rdata[31] mem_rdata[3] mem_rdata[4] mem_rdata[5]
+ mem_rdata[6] mem_rdata[7] mem_rdata[8] mem_rdata[9] mem_ready mem_valid mem_wdata[0]
+ mem_wdata[10] mem_wdata[11] mem_wdata[12] mem_wdata[13] mem_wdata[14] mem_wdata[15]
+ mem_wdata[16] mem_wdata[17] mem_wdata[18] mem_wdata[19] mem_wdata[1] mem_wdata[20]
+ mem_wdata[21] mem_wdata[22] mem_wdata[23] mem_wdata[24] mem_wdata[25] mem_wdata[26]
+ mem_wdata[27] mem_wdata[28] mem_wdata[29] mem_wdata[2] mem_wdata[30] mem_wdata[31]
+ mem_wdata[3] mem_wdata[4] mem_wdata[5] mem_wdata[6] mem_wdata[7] mem_wdata[8] mem_wdata[9]
+ mem_wstrb[0] mem_wstrb[1] mem_wstrb[2] mem_wstrb[3] pcpi_approx_mul_rd[0] pcpi_approx_mul_rd[10]
+ pcpi_approx_mul_rd[11] pcpi_approx_mul_rd[12] pcpi_approx_mul_rd[13] pcpi_approx_mul_rd[14]
+ pcpi_approx_mul_rd[15] pcpi_approx_mul_rd[16] pcpi_approx_mul_rd[17] pcpi_approx_mul_rd[18]
+ pcpi_approx_mul_rd[19] pcpi_approx_mul_rd[1] pcpi_approx_mul_rd[20] pcpi_approx_mul_rd[21]
+ pcpi_approx_mul_rd[22] pcpi_approx_mul_rd[23] pcpi_approx_mul_rd[24] pcpi_approx_mul_rd[25]
+ pcpi_approx_mul_rd[26] pcpi_approx_mul_rd[27] pcpi_approx_mul_rd[28] pcpi_approx_mul_rd[29]
+ pcpi_approx_mul_rd[2] pcpi_approx_mul_rd[30] pcpi_approx_mul_rd[31] pcpi_approx_mul_rd[3]
+ pcpi_approx_mul_rd[4] pcpi_approx_mul_rd[5] pcpi_approx_mul_rd[6] pcpi_approx_mul_rd[7]
+ pcpi_approx_mul_rd[8] pcpi_approx_mul_rd[9] pcpi_approx_mul_ready pcpi_approx_mul_wait
+ pcpi_approx_mul_wr pcpi_div_rd[0] pcpi_div_rd[10] pcpi_div_rd[11] pcpi_div_rd[12]
+ pcpi_div_rd[13] pcpi_div_rd[14] pcpi_div_rd[15] pcpi_div_rd[16] pcpi_div_rd[17]
+ pcpi_div_rd[18] pcpi_div_rd[19] pcpi_div_rd[1] pcpi_div_rd[20] pcpi_div_rd[21] pcpi_div_rd[22]
+ pcpi_div_rd[23] pcpi_div_rd[24] pcpi_div_rd[25] pcpi_div_rd[26] pcpi_div_rd[27]
+ pcpi_div_rd[28] pcpi_div_rd[29] pcpi_div_rd[2] pcpi_div_rd[30] pcpi_div_rd[31] pcpi_div_rd[3]
+ pcpi_div_rd[4] pcpi_div_rd[5] pcpi_div_rd[6] pcpi_div_rd[7] pcpi_div_rd[8] pcpi_div_rd[9]
+ pcpi_div_ready pcpi_div_wait pcpi_div_wr pcpi_exact_mul_rd[0] pcpi_exact_mul_rd[10]
+ pcpi_exact_mul_rd[11] pcpi_exact_mul_rd[12] pcpi_exact_mul_rd[13] pcpi_exact_mul_rd[14]
+ pcpi_exact_mul_rd[15] pcpi_exact_mul_rd[16] pcpi_exact_mul_rd[17] pcpi_exact_mul_rd[18]
+ pcpi_exact_mul_rd[19] pcpi_exact_mul_rd[1] pcpi_exact_mul_rd[20] pcpi_exact_mul_rd[21]
+ pcpi_exact_mul_rd[22] pcpi_exact_mul_rd[23] pcpi_exact_mul_rd[24] pcpi_exact_mul_rd[25]
+ pcpi_exact_mul_rd[26] pcpi_exact_mul_rd[27] pcpi_exact_mul_rd[28] pcpi_exact_mul_rd[29]
+ pcpi_exact_mul_rd[2] pcpi_exact_mul_rd[30] pcpi_exact_mul_rd[31] pcpi_exact_mul_rd[3]
+ pcpi_exact_mul_rd[4] pcpi_exact_mul_rd[5] pcpi_exact_mul_rd[6] pcpi_exact_mul_rd[7]
+ pcpi_exact_mul_rd[8] pcpi_exact_mul_rd[9] pcpi_exact_mul_ready pcpi_exact_mul_wait
+ pcpi_exact_mul_wr pcpi_insn[0] pcpi_insn[10] pcpi_insn[11] pcpi_insn[12] pcpi_insn[13]
+ pcpi_insn[14] pcpi_insn[15] pcpi_insn[16] pcpi_insn[17] pcpi_insn[18] pcpi_insn[19]
+ pcpi_insn[1] pcpi_insn[20] pcpi_insn[21] pcpi_insn[22] pcpi_insn[23] pcpi_insn[24]
+ pcpi_insn[25] pcpi_insn[26] pcpi_insn[27] pcpi_insn[28] pcpi_insn[29] pcpi_insn[2]
+ pcpi_insn[30] pcpi_insn[31] pcpi_insn[3] pcpi_insn[4] pcpi_insn[5] pcpi_insn[6]
+ pcpi_insn[7] pcpi_insn[8] pcpi_insn[9] pcpi_mul_rd[0] pcpi_mul_rd[10] pcpi_mul_rd[11]
+ pcpi_mul_rd[12] pcpi_mul_rd[13] pcpi_mul_rd[14] pcpi_mul_rd[15] pcpi_mul_rd[16]
+ pcpi_mul_rd[17] pcpi_mul_rd[18] pcpi_mul_rd[19] pcpi_mul_rd[1] pcpi_mul_rd[20] pcpi_mul_rd[21]
+ pcpi_mul_rd[22] pcpi_mul_rd[23] pcpi_mul_rd[24] pcpi_mul_rd[25] pcpi_mul_rd[26]
+ pcpi_mul_rd[27] pcpi_mul_rd[28] pcpi_mul_rd[29] pcpi_mul_rd[2] pcpi_mul_rd[30] pcpi_mul_rd[31]
+ pcpi_mul_rd[3] pcpi_mul_rd[4] pcpi_mul_rd[5] pcpi_mul_rd[6] pcpi_mul_rd[7] pcpi_mul_rd[8]
+ pcpi_mul_rd[9] pcpi_mul_ready pcpi_mul_wait pcpi_mul_wr pcpi_rs1[0] pcpi_rs1[10]
+ pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14] pcpi_rs1[15] pcpi_rs1[16] pcpi_rs1[17]
+ pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20] pcpi_rs1[21] pcpi_rs1[22] pcpi_rs1[23]
+ pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27] pcpi_rs1[28] pcpi_rs1[29] pcpi_rs1[2]
+ pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4] pcpi_rs1[5] pcpi_rs1[6] pcpi_rs1[7]
+ pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10] pcpi_rs2[11] pcpi_rs2[12] pcpi_rs2[13]
+ pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17] pcpi_rs2[18] pcpi_rs2[19] pcpi_rs2[1]
+ pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23] pcpi_rs2[24] pcpi_rs2[25] pcpi_rs2[26]
+ pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2] pcpi_rs2[30] pcpi_rs2[31] pcpi_rs2[3]
+ pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7] pcpi_rs2[8] pcpi_rs2[9] pcpi_valid
+ resetn vdd vss
.ends

* Black-box entry subcircuit for pcpi_exact_mul abstract view
.subckt pcpi_exact_mul clk pcpi_insn[0] pcpi_insn[10] pcpi_insn[11] pcpi_insn[12]
+ pcpi_insn[13] pcpi_insn[14] pcpi_insn[15] pcpi_insn[16] pcpi_insn[17] pcpi_insn[18]
+ pcpi_insn[19] pcpi_insn[1] pcpi_insn[20] pcpi_insn[21] pcpi_insn[22] pcpi_insn[23]
+ pcpi_insn[24] pcpi_insn[25] pcpi_insn[26] pcpi_insn[27] pcpi_insn[28] pcpi_insn[29]
+ pcpi_insn[2] pcpi_insn[30] pcpi_insn[31] pcpi_insn[3] pcpi_insn[4] pcpi_insn[5]
+ pcpi_insn[6] pcpi_insn[7] pcpi_insn[8] pcpi_insn[9] pcpi_rd[0] pcpi_rd[10] pcpi_rd[11]
+ pcpi_rd[12] pcpi_rd[13] pcpi_rd[14] pcpi_rd[15] pcpi_rd[16] pcpi_rd[17] pcpi_rd[18]
+ pcpi_rd[19] pcpi_rd[1] pcpi_rd[20] pcpi_rd[21] pcpi_rd[22] pcpi_rd[23] pcpi_rd[24]
+ pcpi_rd[25] pcpi_rd[26] pcpi_rd[27] pcpi_rd[28] pcpi_rd[29] pcpi_rd[2] pcpi_rd[30]
+ pcpi_rd[31] pcpi_rd[3] pcpi_rd[4] pcpi_rd[5] pcpi_rd[6] pcpi_rd[7] pcpi_rd[8] pcpi_rd[9]
+ pcpi_ready pcpi_rs1[0] pcpi_rs1[10] pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14]
+ pcpi_rs1[15] pcpi_rs1[16] pcpi_rs1[17] pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20]
+ pcpi_rs1[21] pcpi_rs1[22] pcpi_rs1[23] pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27]
+ pcpi_rs1[28] pcpi_rs1[29] pcpi_rs1[2] pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4]
+ pcpi_rs1[5] pcpi_rs1[6] pcpi_rs1[7] pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10]
+ pcpi_rs2[11] pcpi_rs2[12] pcpi_rs2[13] pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17]
+ pcpi_rs2[18] pcpi_rs2[19] pcpi_rs2[1] pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23]
+ pcpi_rs2[24] pcpi_rs2[25] pcpi_rs2[26] pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2]
+ pcpi_rs2[30] pcpi_rs2[31] pcpi_rs2[3] pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7]
+ pcpi_rs2[8] pcpi_rs2[9] pcpi_valid pcpi_wait pcpi_wr resetn vdd vss
.ends

* Black-box entry subcircuit for spimemio abstract view
.subckt spimemio addr[0] addr[10] addr[11] addr[12] addr[13] addr[14] addr[15] addr[16]
+ addr[17] addr[18] addr[19] addr[1] addr[20] addr[21] addr[22] addr[23] addr[2] addr[3]
+ addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] cfgreg_di[0] cfgreg_di[10] cfgreg_di[11]
+ cfgreg_di[12] cfgreg_di[13] cfgreg_di[14] cfgreg_di[15] cfgreg_di[16] cfgreg_di[17]
+ cfgreg_di[18] cfgreg_di[19] cfgreg_di[1] cfgreg_di[20] cfgreg_di[21] cfgreg_di[22]
+ cfgreg_di[23] cfgreg_di[24] cfgreg_di[25] cfgreg_di[26] cfgreg_di[27] cfgreg_di[28]
+ cfgreg_di[29] cfgreg_di[2] cfgreg_di[30] cfgreg_di[31] cfgreg_di[3] cfgreg_di[4]
+ cfgreg_di[5] cfgreg_di[6] cfgreg_di[7] cfgreg_di[8] cfgreg_di[9] cfgreg_do[0] cfgreg_do[10]
+ cfgreg_do[11] cfgreg_do[12] cfgreg_do[13] cfgreg_do[14] cfgreg_do[15] cfgreg_do[16]
+ cfgreg_do[17] cfgreg_do[18] cfgreg_do[19] cfgreg_do[1] cfgreg_do[20] cfgreg_do[21]
+ cfgreg_do[22] cfgreg_do[23] cfgreg_do[24] cfgreg_do[25] cfgreg_do[26] cfgreg_do[27]
+ cfgreg_do[28] cfgreg_do[29] cfgreg_do[2] cfgreg_do[30] cfgreg_do[31] cfgreg_do[3]
+ cfgreg_do[4] cfgreg_do[5] cfgreg_do[6] cfgreg_do[7] cfgreg_do[8] cfgreg_do[9] cfgreg_we[0]
+ cfgreg_we[1] cfgreg_we[2] cfgreg_we[3] clk flash_in[0] flash_in[1] flash_in[2] flash_in[3]
+ flash_in[4] flash_in[5] flash_oeb[0] flash_oeb[1] flash_oeb[2] flash_oeb[3] flash_oeb[4]
+ flash_oeb[5] flash_out[0] flash_out[1] flash_out[2] flash_out[3] flash_out[4] flash_out[5]
+ rdata[0] rdata[10] rdata[11] rdata[12] rdata[13] rdata[14] rdata[15] rdata[16] rdata[17]
+ rdata[18] rdata[19] rdata[1] rdata[20] rdata[21] rdata[22] rdata[23] rdata[24] rdata[25]
+ rdata[26] rdata[27] rdata[28] rdata[29] rdata[2] rdata[30] rdata[31] rdata[3] rdata[4]
+ rdata[5] rdata[6] rdata[7] rdata[8] rdata[9] ready resetn valid vdd vss
.ends

* Black-box entry subcircuit for simpleuart abstract view
.subckt simpleuart clk reg_dat_di[0] reg_dat_di[10] reg_dat_di[11] reg_dat_di[12]
+ reg_dat_di[13] reg_dat_di[14] reg_dat_di[15] reg_dat_di[16] reg_dat_di[17] reg_dat_di[18]
+ reg_dat_di[19] reg_dat_di[1] reg_dat_di[20] reg_dat_di[21] reg_dat_di[22] reg_dat_di[23]
+ reg_dat_di[24] reg_dat_di[25] reg_dat_di[26] reg_dat_di[27] reg_dat_di[28] reg_dat_di[29]
+ reg_dat_di[2] reg_dat_di[30] reg_dat_di[31] reg_dat_di[3] reg_dat_di[4] reg_dat_di[5]
+ reg_dat_di[6] reg_dat_di[7] reg_dat_di[8] reg_dat_di[9] reg_dat_do[0] reg_dat_do[10]
+ reg_dat_do[11] reg_dat_do[12] reg_dat_do[13] reg_dat_do[14] reg_dat_do[15] reg_dat_do[16]
+ reg_dat_do[17] reg_dat_do[18] reg_dat_do[19] reg_dat_do[1] reg_dat_do[20] reg_dat_do[21]
+ reg_dat_do[22] reg_dat_do[23] reg_dat_do[24] reg_dat_do[25] reg_dat_do[26] reg_dat_do[27]
+ reg_dat_do[28] reg_dat_do[29] reg_dat_do[2] reg_dat_do[30] reg_dat_do[31] reg_dat_do[3]
+ reg_dat_do[4] reg_dat_do[5] reg_dat_do[6] reg_dat_do[7] reg_dat_do[8] reg_dat_do[9]
+ reg_dat_re reg_dat_wait reg_dat_we reg_div_di[0] reg_div_di[10] reg_div_di[11] reg_div_di[12]
+ reg_div_di[13] reg_div_di[14] reg_div_di[15] reg_div_di[16] reg_div_di[17] reg_div_di[18]
+ reg_div_di[19] reg_div_di[1] reg_div_di[20] reg_div_di[21] reg_div_di[22] reg_div_di[23]
+ reg_div_di[24] reg_div_di[25] reg_div_di[26] reg_div_di[27] reg_div_di[28] reg_div_di[29]
+ reg_div_di[2] reg_div_di[30] reg_div_di[31] reg_div_di[3] reg_div_di[4] reg_div_di[5]
+ reg_div_di[6] reg_div_di[7] reg_div_di[8] reg_div_di[9] reg_div_do[0] reg_div_do[10]
+ reg_div_do[11] reg_div_do[12] reg_div_do[13] reg_div_do[14] reg_div_do[15] reg_div_do[16]
+ reg_div_do[17] reg_div_do[18] reg_div_do[19] reg_div_do[1] reg_div_do[20] reg_div_do[21]
+ reg_div_do[22] reg_div_do[23] reg_div_do[24] reg_div_do[25] reg_div_do[26] reg_div_do[27]
+ reg_div_do[28] reg_div_do[29] reg_div_do[2] reg_div_do[30] reg_div_do[31] reg_div_do[3]
+ reg_div_do[4] reg_div_do[5] reg_div_do[6] reg_div_do[7] reg_div_do[8] reg_div_do[9]
+ reg_div_we[0] reg_div_we[1] reg_div_we[2] reg_div_we[3] resetn uart_in[0] uart_in[1]
+ uart_oeb[0] uart_oeb[1] uart_out[0] uart_out[1] vdd vss
.ends

* Black-box entry subcircuit for pcpi_div abstract view
.subckt pcpi_div clk pcpi_div_rd[0] pcpi_div_rd[10] pcpi_div_rd[11] pcpi_div_rd[12]
+ pcpi_div_rd[13] pcpi_div_rd[14] pcpi_div_rd[15] pcpi_div_rd[16] pcpi_div_rd[17]
+ pcpi_div_rd[18] pcpi_div_rd[19] pcpi_div_rd[1] pcpi_div_rd[20] pcpi_div_rd[21] pcpi_div_rd[22]
+ pcpi_div_rd[23] pcpi_div_rd[24] pcpi_div_rd[25] pcpi_div_rd[26] pcpi_div_rd[27]
+ pcpi_div_rd[28] pcpi_div_rd[29] pcpi_div_rd[2] pcpi_div_rd[30] pcpi_div_rd[31] pcpi_div_rd[3]
+ pcpi_div_rd[4] pcpi_div_rd[5] pcpi_div_rd[6] pcpi_div_rd[7] pcpi_div_rd[8] pcpi_div_rd[9]
+ pcpi_div_ready pcpi_div_valid pcpi_div_wait pcpi_div_wr pcpi_insn[0] pcpi_insn[10]
+ pcpi_insn[11] pcpi_insn[12] pcpi_insn[13] pcpi_insn[14] pcpi_insn[15] pcpi_insn[16]
+ pcpi_insn[17] pcpi_insn[18] pcpi_insn[19] pcpi_insn[1] pcpi_insn[20] pcpi_insn[21]
+ pcpi_insn[22] pcpi_insn[23] pcpi_insn[24] pcpi_insn[25] pcpi_insn[26] pcpi_insn[27]
+ pcpi_insn[28] pcpi_insn[29] pcpi_insn[2] pcpi_insn[30] pcpi_insn[31] pcpi_insn[3]
+ pcpi_insn[4] pcpi_insn[5] pcpi_insn[6] pcpi_insn[7] pcpi_insn[8] pcpi_insn[9] pcpi_rs1[0]
+ pcpi_rs1[10] pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14] pcpi_rs1[15] pcpi_rs1[16]
+ pcpi_rs1[17] pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20] pcpi_rs1[21] pcpi_rs1[22]
+ pcpi_rs1[23] pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27] pcpi_rs1[28] pcpi_rs1[29]
+ pcpi_rs1[2] pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4] pcpi_rs1[5] pcpi_rs1[6]
+ pcpi_rs1[7] pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10] pcpi_rs2[11] pcpi_rs2[12]
+ pcpi_rs2[13] pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17] pcpi_rs2[18] pcpi_rs2[19]
+ pcpi_rs2[1] pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23] pcpi_rs2[24] pcpi_rs2[25]
+ pcpi_rs2[26] pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2] pcpi_rs2[30] pcpi_rs2[31]
+ pcpi_rs2[3] pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7] pcpi_rs2[8] pcpi_rs2[9]
+ resetn vdd vss
.ends

.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xuser_proj_example_inst_0 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ user_irq[0] user_irq[1] user_irq[2] la_data_in[0] la_data_in[10] la_data_in[11]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33]
+ la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60]
+ la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[6] la_data_in[7] la_data_in[8]
+ la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] la_oenb[0] la_oenb[10]
+ la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i user_proj_example
Xsimple_interconnect_inst_0 io_in[8] io_in[22] io_in[32] io_in[33] io_in[34] io_in[35]
+ io_in[36] io_in[37] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28]
+ io_in[29] io_in[30] io_in[31] io_oeb[22] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[30] io_oeb[31] io_out[22] io_out[32] io_out[33] io_out[34] io_out[35]
+ io_out[36] io_out[37] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28]
+ io_out[29] io_out[30] io_out[31] mem_addr\[0\] mem_addr\[10\] mem_addr\[11\] mem_addr\[12\]
+ mem_addr\[13\] mem_addr\[14\] mem_addr\[15\] mem_addr\[16\] mem_addr\[17\] mem_addr\[18\]
+ mem_addr\[19\] mem_addr\[1\] mem_addr\[20\] mem_addr\[21\] mem_addr\[22\] mem_addr\[23\]
+ mem_addr\[24\] mem_addr\[25\] mem_addr\[26\] mem_addr\[27\] mem_addr\[28\] mem_addr\[29\]
+ mem_addr\[2\] mem_addr\[30\] mem_addr\[31\] mem_addr\[3\] mem_addr\[4\] mem_addr\[5\]
+ mem_addr\[6\] mem_addr\[7\] mem_addr\[8\] mem_addr\[9\] mem_instr mem_rdata\[0\]
+ mem_rdata\[10\] mem_rdata\[11\] mem_rdata\[12\] mem_rdata\[13\] mem_rdata\[14\]
+ mem_rdata\[15\] mem_rdata\[16\] mem_rdata\[17\] mem_rdata\[18\] mem_rdata\[19\]
+ mem_rdata\[1\] mem_rdata\[20\] mem_rdata\[21\] mem_rdata\[22\] mem_rdata\[23\] mem_rdata\[24\]
+ mem_rdata\[25\] mem_rdata\[26\] mem_rdata\[27\] mem_rdata\[28\] mem_rdata\[29\]
+ mem_rdata\[2\] mem_rdata\[30\] mem_rdata\[31\] mem_rdata\[3\] mem_rdata\[4\] mem_rdata\[5\]
+ mem_rdata\[6\] mem_rdata\[7\] mem_rdata\[8\] mem_rdata\[9\] mem_ready mem_valid
+ mem_wdata\[0\] mem_wdata\[10\] mem_wdata\[11\] mem_wdata\[12\] mem_wdata\[13\] mem_wdata\[14\]
+ mem_wdata\[15\] mem_wdata\[16\] mem_wdata\[17\] mem_wdata\[18\] mem_wdata\[19\]
+ mem_wdata\[1\] mem_wdata\[20\] mem_wdata\[21\] mem_wdata\[22\] mem_wdata\[23\] mem_wdata\[24\]
+ mem_wdata\[25\] mem_wdata\[26\] mem_wdata\[27\] mem_wdata\[28\] mem_wdata\[29\]
+ mem_wdata\[2\] mem_wdata\[30\] mem_wdata\[31\] mem_wdata\[3\] mem_wdata\[4\] mem_wdata\[5\]
+ mem_wdata\[6\] mem_wdata\[7\] mem_wdata\[8\] mem_wdata\[9\] mem_wstrb\[0\] mem_wstrb\[1\]
+ mem_wstrb\[2\] mem_wstrb\[3\] ram_gwenb\[0\] ram_gwenb\[1\] ram_gwenb\[2\] ram_gwenb\[3\]
+ ram_rdata\[0\] ram_rdata\[10\] ram_rdata\[11\] ram_rdata\[12\] ram_rdata\[13\] ram_rdata\[14\]
+ ram_rdata\[15\] ram_rdata\[16\] ram_rdata\[17\] ram_rdata\[18\] ram_rdata\[19\]
+ ram_rdata\[1\] ram_rdata\[20\] ram_rdata\[21\] ram_rdata\[22\] ram_rdata\[23\] ram_rdata\[24\]
+ ram_rdata\[25\] ram_rdata\[26\] ram_rdata\[27\] ram_rdata\[28\] ram_rdata\[29\]
+ ram_rdata\[2\] ram_rdata\[30\] ram_rdata\[31\] ram_rdata\[3\] ram_rdata\[4\] ram_rdata\[5\]
+ ram_rdata\[6\] ram_rdata\[7\] ram_rdata\[8\] ram_rdata\[9\] ram_wenb\[0\] ram_wenb\[10\]
+ ram_wenb\[11\] ram_wenb\[12\] ram_wenb\[13\] ram_wenb\[14\] ram_wenb\[15\] ram_wenb\[16\]
+ ram_wenb\[17\] ram_wenb\[18\] ram_wenb\[19\] ram_wenb\[1\] ram_wenb\[20\] ram_wenb\[21\]
+ ram_wenb\[22\] ram_wenb\[23\] ram_wenb\[24\] ram_wenb\[25\] ram_wenb\[26\] ram_wenb\[27\]
+ ram_wenb\[28\] ram_wenb\[29\] ram_wenb\[2\] ram_wenb\[30\] ram_wenb\[31\] ram_wenb\[3\]
+ ram_wenb\[4\] ram_wenb\[5\] ram_wenb\[6\] ram_wenb\[7\] ram_wenb\[8\] ram_wenb\[9\]
+ resetn simpleuart_dat_re simpleuart_dat_we simpleuart_div_we\[0\] simpleuart_div_we\[1\]
+ simpleuart_div_we\[2\] simpleuart_div_we\[3\] simpleuart_reg_dat_do\[0\] simpleuart_reg_dat_do\[10\]
+ simpleuart_reg_dat_do\[11\] simpleuart_reg_dat_do\[12\] simpleuart_reg_dat_do\[13\]
+ simpleuart_reg_dat_do\[14\] simpleuart_reg_dat_do\[15\] simpleuart_reg_dat_do\[16\]
+ simpleuart_reg_dat_do\[17\] simpleuart_reg_dat_do\[18\] simpleuart_reg_dat_do\[19\]
+ simpleuart_reg_dat_do\[1\] simpleuart_reg_dat_do\[20\] simpleuart_reg_dat_do\[21\]
+ simpleuart_reg_dat_do\[22\] simpleuart_reg_dat_do\[23\] simpleuart_reg_dat_do\[24\]
+ simpleuart_reg_dat_do\[25\] simpleuart_reg_dat_do\[26\] simpleuart_reg_dat_do\[27\]
+ simpleuart_reg_dat_do\[28\] simpleuart_reg_dat_do\[29\] simpleuart_reg_dat_do\[2\]
+ simpleuart_reg_dat_do\[30\] simpleuart_reg_dat_do\[31\] simpleuart_reg_dat_do\[3\]
+ simpleuart_reg_dat_do\[4\] simpleuart_reg_dat_do\[5\] simpleuart_reg_dat_do\[6\]
+ simpleuart_reg_dat_do\[7\] simpleuart_reg_dat_do\[8\] simpleuart_reg_dat_do\[9\]
+ simpleuart_reg_dat_wait simpleuart_reg_div_do\[0\] simpleuart_reg_div_do\[10\] simpleuart_reg_div_do\[11\]
+ simpleuart_reg_div_do\[12\] simpleuart_reg_div_do\[13\] simpleuart_reg_div_do\[14\]
+ simpleuart_reg_div_do\[15\] simpleuart_reg_div_do\[16\] simpleuart_reg_div_do\[17\]
+ simpleuart_reg_div_do\[18\] simpleuart_reg_div_do\[19\] simpleuart_reg_div_do\[1\]
+ simpleuart_reg_div_do\[20\] simpleuart_reg_div_do\[21\] simpleuart_reg_div_do\[22\]
+ simpleuart_reg_div_do\[23\] simpleuart_reg_div_do\[24\] simpleuart_reg_div_do\[25\]
+ simpleuart_reg_div_do\[26\] simpleuart_reg_div_do\[27\] simpleuart_reg_div_do\[28\]
+ simpleuart_reg_div_do\[29\] simpleuart_reg_div_do\[2\] simpleuart_reg_div_do\[30\]
+ simpleuart_reg_div_do\[31\] simpleuart_reg_div_do\[3\] simpleuart_reg_div_do\[4\]
+ simpleuart_reg_div_do\[5\] simpleuart_reg_div_do\[6\] simpleuart_reg_div_do\[7\]
+ simpleuart_reg_div_do\[8\] simpleuart_reg_div_do\[9\] spimem_rdata\[0\] spimem_rdata\[10\]
+ spimem_rdata\[11\] spimem_rdata\[12\] spimem_rdata\[13\] spimem_rdata\[14\] spimem_rdata\[15\]
+ spimem_rdata\[16\] spimem_rdata\[17\] spimem_rdata\[18\] spimem_rdata\[19\] spimem_rdata\[1\]
+ spimem_rdata\[20\] spimem_rdata\[21\] spimem_rdata\[22\] spimem_rdata\[23\] spimem_rdata\[24\]
+ spimem_rdata\[25\] spimem_rdata\[26\] spimem_rdata\[27\] spimem_rdata\[28\] spimem_rdata\[29\]
+ spimem_rdata\[2\] spimem_rdata\[30\] spimem_rdata\[31\] spimem_rdata\[3\] spimem_rdata\[4\]
+ spimem_rdata\[5\] spimem_rdata\[6\] spimem_rdata\[7\] spimem_rdata\[8\] spimem_rdata\[9\]
+ spimem_ready spimem_valid spimemio_cfgreg_do\[0\] spimemio_cfgreg_do\[10\] spimemio_cfgreg_do\[11\]
+ spimemio_cfgreg_do\[12\] spimemio_cfgreg_do\[13\] spimemio_cfgreg_do\[14\] spimemio_cfgreg_do\[15\]
+ spimemio_cfgreg_do\[16\] spimemio_cfgreg_do\[17\] spimemio_cfgreg_do\[18\] spimemio_cfgreg_do\[19\]
+ spimemio_cfgreg_do\[1\] spimemio_cfgreg_do\[20\] spimemio_cfgreg_do\[21\] spimemio_cfgreg_do\[22\]
+ spimemio_cfgreg_do\[23\] spimemio_cfgreg_do\[24\] spimemio_cfgreg_do\[25\] spimemio_cfgreg_do\[26\]
+ spimemio_cfgreg_do\[27\] spimemio_cfgreg_do\[28\] spimemio_cfgreg_do\[29\] spimemio_cfgreg_do\[2\]
+ spimemio_cfgreg_do\[30\] spimemio_cfgreg_do\[31\] spimemio_cfgreg_do\[3\] spimemio_cfgreg_do\[4\]
+ spimemio_cfgreg_do\[5\] spimemio_cfgreg_do\[6\] spimemio_cfgreg_do\[7\] spimemio_cfgreg_do\[8\]
+ spimemio_cfgreg_do\[9\] spimemio_cfgreg_we\[0\] spimemio_cfgreg_we\[1\] spimemio_cfgreg_we\[2\]
+ spimemio_cfgreg_we\[3\] vdd vss simple_interconnect
Xsram512x8_0 vdd vss mem_addr\[2\] mem_addr\[3\] mem_addr\[4\] mem_addr\[5\] mem_addr\[6\]
+ mem_addr\[7\] mem_addr\[8\] mem_addr\[9\] mem_addr\[10\] reset io_in[8] ram_gwenb\[0\]
+ ram_rdata\[0\] ram_rdata\[1\] ram_rdata\[2\] ram_rdata\[3\] ram_rdata\[4\] ram_rdata\[5\]
+ ram_rdata\[6\] ram_rdata\[7\] mem_wdata\[0\] mem_wdata\[1\] mem_wdata\[2\] mem_wdata\[3\]
+ mem_wdata\[4\] mem_wdata\[5\] mem_wdata\[6\] mem_wdata\[7\] ram_wenb\[0\] ram_wenb\[1\]
+ ram_wenb\[2\] ram_wenb\[3\] ram_wenb\[4\] ram_wenb\[5\] ram_wenb\[6\] ram_wenb\[7\]
+ gf180_ram_512x8x1
Xpcpi_approx_mul_inst_0 io_in[8] pcpi_insn\[0\] pcpi_insn\[10\] pcpi_insn\[11\] pcpi_insn\[12\]
+ pcpi_insn\[13\] pcpi_insn\[14\] pcpi_insn\[15\] pcpi_insn\[16\] pcpi_insn\[17\]
+ pcpi_insn\[18\] pcpi_insn\[19\] pcpi_insn\[1\] pcpi_insn\[20\] pcpi_insn\[21\] pcpi_insn\[22\]
+ pcpi_insn\[23\] pcpi_insn\[24\] pcpi_insn\[25\] pcpi_insn\[26\] pcpi_insn\[27\]
+ pcpi_insn\[28\] pcpi_insn\[29\] pcpi_insn\[2\] pcpi_insn\[30\] pcpi_insn\[31\] pcpi_insn\[3\]
+ pcpi_insn\[4\] pcpi_insn\[5\] pcpi_insn\[6\] pcpi_insn\[7\] pcpi_insn\[8\] pcpi_insn\[9\]
+ pcpi_approx_mul_rd\[0\] pcpi_approx_mul_rd\[10\] pcpi_approx_mul_rd\[11\] pcpi_approx_mul_rd\[12\]
+ pcpi_approx_mul_rd\[13\] pcpi_approx_mul_rd\[14\] pcpi_approx_mul_rd\[15\] pcpi_approx_mul_rd\[16\]
+ pcpi_approx_mul_rd\[17\] pcpi_approx_mul_rd\[18\] pcpi_approx_mul_rd\[19\] pcpi_approx_mul_rd\[1\]
+ pcpi_approx_mul_rd\[20\] pcpi_approx_mul_rd\[21\] pcpi_approx_mul_rd\[22\] pcpi_approx_mul_rd\[23\]
+ pcpi_approx_mul_rd\[24\] pcpi_approx_mul_rd\[25\] pcpi_approx_mul_rd\[26\] pcpi_approx_mul_rd\[27\]
+ pcpi_approx_mul_rd\[28\] pcpi_approx_mul_rd\[29\] pcpi_approx_mul_rd\[2\] pcpi_approx_mul_rd\[30\]
+ pcpi_approx_mul_rd\[31\] pcpi_approx_mul_rd\[3\] pcpi_approx_mul_rd\[4\] pcpi_approx_mul_rd\[5\]
+ pcpi_approx_mul_rd\[6\] pcpi_approx_mul_rd\[7\] pcpi_approx_mul_rd\[8\] pcpi_approx_mul_rd\[9\]
+ pcpi_approx_mul_ready pcpi_rs1\[0\] pcpi_rs1\[10\] pcpi_rs1\[11\] pcpi_rs1\[12\]
+ pcpi_rs1\[13\] pcpi_rs1\[14\] pcpi_rs1\[15\] pcpi_rs1\[16\] pcpi_rs1\[17\] pcpi_rs1\[18\]
+ pcpi_rs1\[19\] pcpi_rs1\[1\] pcpi_rs1\[20\] pcpi_rs1\[21\] pcpi_rs1\[22\] pcpi_rs1\[23\]
+ pcpi_rs1\[24\] pcpi_rs1\[25\] pcpi_rs1\[26\] pcpi_rs1\[27\] pcpi_rs1\[28\] pcpi_rs1\[29\]
+ pcpi_rs1\[2\] pcpi_rs1\[30\] pcpi_rs1\[31\] pcpi_rs1\[3\] pcpi_rs1\[4\] pcpi_rs1\[5\]
+ pcpi_rs1\[6\] pcpi_rs1\[7\] pcpi_rs1\[8\] pcpi_rs1\[9\] pcpi_rs2\[0\] pcpi_rs2\[10\]
+ pcpi_rs2\[11\] pcpi_rs2\[12\] pcpi_rs2\[13\] pcpi_rs2\[14\] pcpi_rs2\[15\] pcpi_rs2\[16\]
+ pcpi_rs2\[17\] pcpi_rs2\[18\] pcpi_rs2\[19\] pcpi_rs2\[1\] pcpi_rs2\[20\] pcpi_rs2\[21\]
+ pcpi_rs2\[22\] pcpi_rs2\[23\] pcpi_rs2\[24\] pcpi_rs2\[25\] pcpi_rs2\[26\] pcpi_rs2\[27\]
+ pcpi_rs2\[28\] pcpi_rs2\[29\] pcpi_rs2\[2\] pcpi_rs2\[30\] pcpi_rs2\[31\] pcpi_rs2\[3\]
+ pcpi_rs2\[4\] pcpi_rs2\[5\] pcpi_rs2\[6\] pcpi_rs2\[7\] pcpi_rs2\[8\] pcpi_rs2\[9\]
+ pcpi_valid pcpi_approx_mul_wait pcpi_approx_mul_wr resetn vdd vss pcpi_approx_mul
Xsram512x8_1 vdd vss mem_addr\[2\] mem_addr\[3\] mem_addr\[4\] mem_addr\[5\] mem_addr\[6\]
+ mem_addr\[7\] mem_addr\[8\] mem_addr\[9\] mem_addr\[10\] reset io_in[8] ram_gwenb\[1\]
+ ram_rdata\[8\] ram_rdata\[9\] ram_rdata\[10\] ram_rdata\[11\] ram_rdata\[12\] ram_rdata\[13\]
+ ram_rdata\[14\] ram_rdata\[15\] mem_wdata\[8\] mem_wdata\[9\] mem_wdata\[10\] mem_wdata\[11\]
+ mem_wdata\[12\] mem_wdata\[13\] mem_wdata\[14\] mem_wdata\[15\] ram_wenb\[8\] ram_wenb\[9\]
+ ram_wenb\[10\] ram_wenb\[11\] ram_wenb\[12\] ram_wenb\[13\] ram_wenb\[14\] ram_wenb\[15\]
+ gf180_ram_512x8x1
Xsram512x8_2 vdd vss mem_addr\[2\] mem_addr\[3\] mem_addr\[4\] mem_addr\[5\] mem_addr\[6\]
+ mem_addr\[7\] mem_addr\[8\] mem_addr\[9\] mem_addr\[10\] reset io_in[8] ram_gwenb\[2\]
+ ram_rdata\[16\] ram_rdata\[17\] ram_rdata\[18\] ram_rdata\[19\] ram_rdata\[20\]
+ ram_rdata\[21\] ram_rdata\[22\] ram_rdata\[23\] mem_wdata\[16\] mem_wdata\[17\]
+ mem_wdata\[18\] mem_wdata\[19\] mem_wdata\[20\] mem_wdata\[21\] mem_wdata\[22\]
+ mem_wdata\[23\] ram_wenb\[16\] ram_wenb\[17\] ram_wenb\[18\] ram_wenb\[19\] ram_wenb\[20\]
+ ram_wenb\[21\] ram_wenb\[22\] ram_wenb\[23\] gf180_ram_512x8x1
Xsram512x8_3 vdd vss mem_addr\[2\] mem_addr\[3\] mem_addr\[4\] mem_addr\[5\] mem_addr\[6\]
+ mem_addr\[7\] mem_addr\[8\] mem_addr\[9\] mem_addr\[10\] reset io_in[8] ram_gwenb\[3\]
+ ram_rdata\[24\] ram_rdata\[25\] ram_rdata\[26\] ram_rdata\[27\] ram_rdata\[28\]
+ ram_rdata\[29\] ram_rdata\[30\] ram_rdata\[31\] mem_wdata\[24\] mem_wdata\[25\]
+ mem_wdata\[26\] mem_wdata\[27\] mem_wdata\[28\] mem_wdata\[29\] mem_wdata\[30\]
+ mem_wdata\[31\] ram_wenb\[24\] ram_wenb\[25\] ram_wenb\[26\] ram_wenb\[27\] ram_wenb\[28\]
+ ram_wenb\[29\] ram_wenb\[30\] ram_wenb\[31\] gf180_ram_512x8x1
Xpcpi_mul_inst_0 io_in[8] pcpi_insn\[0\] pcpi_insn\[10\] pcpi_insn\[11\] pcpi_insn\[12\]
+ pcpi_insn\[13\] pcpi_insn\[14\] pcpi_insn\[15\] pcpi_insn\[16\] pcpi_insn\[17\]
+ pcpi_insn\[18\] pcpi_insn\[19\] pcpi_insn\[1\] pcpi_insn\[20\] pcpi_insn\[21\] pcpi_insn\[22\]
+ pcpi_insn\[23\] pcpi_insn\[24\] pcpi_insn\[25\] pcpi_insn\[26\] pcpi_insn\[27\]
+ pcpi_insn\[28\] pcpi_insn\[29\] pcpi_insn\[2\] pcpi_insn\[30\] pcpi_insn\[31\] pcpi_insn\[3\]
+ pcpi_insn\[4\] pcpi_insn\[5\] pcpi_insn\[6\] pcpi_insn\[7\] pcpi_insn\[8\] pcpi_insn\[9\]
+ pcpi_mul_rd\[0\] pcpi_mul_rd\[10\] pcpi_mul_rd\[11\] pcpi_mul_rd\[12\] pcpi_mul_rd\[13\]
+ pcpi_mul_rd\[14\] pcpi_mul_rd\[15\] pcpi_mul_rd\[16\] pcpi_mul_rd\[17\] pcpi_mul_rd\[18\]
+ pcpi_mul_rd\[19\] pcpi_mul_rd\[1\] pcpi_mul_rd\[20\] pcpi_mul_rd\[21\] pcpi_mul_rd\[22\]
+ pcpi_mul_rd\[23\] pcpi_mul_rd\[24\] pcpi_mul_rd\[25\] pcpi_mul_rd\[26\] pcpi_mul_rd\[27\]
+ pcpi_mul_rd\[28\] pcpi_mul_rd\[29\] pcpi_mul_rd\[2\] pcpi_mul_rd\[30\] pcpi_mul_rd\[31\]
+ pcpi_mul_rd\[3\] pcpi_mul_rd\[4\] pcpi_mul_rd\[5\] pcpi_mul_rd\[6\] pcpi_mul_rd\[7\]
+ pcpi_mul_rd\[8\] pcpi_mul_rd\[9\] pcpi_mul_ready pcpi_valid pcpi_mul_wait pcpi_mul_wr
+ pcpi_rs1\[0\] pcpi_rs1\[10\] pcpi_rs1\[11\] pcpi_rs1\[12\] pcpi_rs1\[13\] pcpi_rs1\[14\]
+ pcpi_rs1\[15\] pcpi_rs1\[16\] pcpi_rs1\[17\] pcpi_rs1\[18\] pcpi_rs1\[19\] pcpi_rs1\[1\]
+ pcpi_rs1\[20\] pcpi_rs1\[21\] pcpi_rs1\[22\] pcpi_rs1\[23\] pcpi_rs1\[24\] pcpi_rs1\[25\]
+ pcpi_rs1\[26\] pcpi_rs1\[27\] pcpi_rs1\[28\] pcpi_rs1\[29\] pcpi_rs1\[2\] pcpi_rs1\[30\]
+ pcpi_rs1\[31\] pcpi_rs1\[3\] pcpi_rs1\[4\] pcpi_rs1\[5\] pcpi_rs1\[6\] pcpi_rs1\[7\]
+ pcpi_rs1\[8\] pcpi_rs1\[9\] pcpi_rs2\[0\] pcpi_rs2\[10\] pcpi_rs2\[11\] pcpi_rs2\[12\]
+ pcpi_rs2\[13\] pcpi_rs2\[14\] pcpi_rs2\[15\] pcpi_rs2\[16\] pcpi_rs2\[17\] pcpi_rs2\[18\]
+ pcpi_rs2\[19\] pcpi_rs2\[1\] pcpi_rs2\[20\] pcpi_rs2\[21\] pcpi_rs2\[22\] pcpi_rs2\[23\]
+ pcpi_rs2\[24\] pcpi_rs2\[25\] pcpi_rs2\[26\] pcpi_rs2\[27\] pcpi_rs2\[28\] pcpi_rs2\[29\]
+ pcpi_rs2\[2\] pcpi_rs2\[30\] pcpi_rs2\[31\] pcpi_rs2\[3\] pcpi_rs2\[4\] pcpi_rs2\[5\]
+ pcpi_rs2\[6\] pcpi_rs2\[7\] pcpi_rs2\[8\] pcpi_rs2\[9\] resetn vdd vss pcpi_mul
Xctrl_inst_0 io_in[8] io_in[9] io_oeb[8] io_oeb[9] io_out[8] io_out[9] reset resetn
+ vdd vss ctrl
Xcpu_inst_0 io_in[8] io_in[18] io_in[19] io_in[20] io_in[21] io_oeb[18] io_oeb[19]
+ io_oeb[20] io_oeb[21] io_out[18] io_out[19] io_out[20] io_out[21] mem_addr\[0\]
+ mem_addr\[10\] mem_addr\[11\] mem_addr\[12\] mem_addr\[13\] mem_addr\[14\] mem_addr\[15\]
+ mem_addr\[16\] mem_addr\[17\] mem_addr\[18\] mem_addr\[19\] mem_addr\[1\] mem_addr\[20\]
+ mem_addr\[21\] mem_addr\[22\] mem_addr\[23\] mem_addr\[24\] mem_addr\[25\] mem_addr\[26\]
+ mem_addr\[27\] mem_addr\[28\] mem_addr\[29\] mem_addr\[2\] mem_addr\[30\] mem_addr\[31\]
+ mem_addr\[3\] mem_addr\[4\] mem_addr\[5\] mem_addr\[6\] mem_addr\[7\] mem_addr\[8\]
+ mem_addr\[9\] mem_instr mem_rdata\[0\] mem_rdata\[10\] mem_rdata\[11\] mem_rdata\[12\]
+ mem_rdata\[13\] mem_rdata\[14\] mem_rdata\[15\] mem_rdata\[16\] mem_rdata\[17\]
+ mem_rdata\[18\] mem_rdata\[19\] mem_rdata\[1\] mem_rdata\[20\] mem_rdata\[21\] mem_rdata\[22\]
+ mem_rdata\[23\] mem_rdata\[24\] mem_rdata\[25\] mem_rdata\[26\] mem_rdata\[27\]
+ mem_rdata\[28\] mem_rdata\[29\] mem_rdata\[2\] mem_rdata\[30\] mem_rdata\[31\] mem_rdata\[3\]
+ mem_rdata\[4\] mem_rdata\[5\] mem_rdata\[6\] mem_rdata\[7\] mem_rdata\[8\] mem_rdata\[9\]
+ mem_ready mem_valid mem_wdata\[0\] mem_wdata\[10\] mem_wdata\[11\] mem_wdata\[12\]
+ mem_wdata\[13\] mem_wdata\[14\] mem_wdata\[15\] mem_wdata\[16\] mem_wdata\[17\]
+ mem_wdata\[18\] mem_wdata\[19\] mem_wdata\[1\] mem_wdata\[20\] mem_wdata\[21\] mem_wdata\[22\]
+ mem_wdata\[23\] mem_wdata\[24\] mem_wdata\[25\] mem_wdata\[26\] mem_wdata\[27\]
+ mem_wdata\[28\] mem_wdata\[29\] mem_wdata\[2\] mem_wdata\[30\] mem_wdata\[31\] mem_wdata\[3\]
+ mem_wdata\[4\] mem_wdata\[5\] mem_wdata\[6\] mem_wdata\[7\] mem_wdata\[8\] mem_wdata\[9\]
+ mem_wstrb\[0\] mem_wstrb\[1\] mem_wstrb\[2\] mem_wstrb\[3\] pcpi_approx_mul_rd\[0\]
+ pcpi_approx_mul_rd\[10\] pcpi_approx_mul_rd\[11\] pcpi_approx_mul_rd\[12\] pcpi_approx_mul_rd\[13\]
+ pcpi_approx_mul_rd\[14\] pcpi_approx_mul_rd\[15\] pcpi_approx_mul_rd\[16\] pcpi_approx_mul_rd\[17\]
+ pcpi_approx_mul_rd\[18\] pcpi_approx_mul_rd\[19\] pcpi_approx_mul_rd\[1\] pcpi_approx_mul_rd\[20\]
+ pcpi_approx_mul_rd\[21\] pcpi_approx_mul_rd\[22\] pcpi_approx_mul_rd\[23\] pcpi_approx_mul_rd\[24\]
+ pcpi_approx_mul_rd\[25\] pcpi_approx_mul_rd\[26\] pcpi_approx_mul_rd\[27\] pcpi_approx_mul_rd\[28\]
+ pcpi_approx_mul_rd\[29\] pcpi_approx_mul_rd\[2\] pcpi_approx_mul_rd\[30\] pcpi_approx_mul_rd\[31\]
+ pcpi_approx_mul_rd\[3\] pcpi_approx_mul_rd\[4\] pcpi_approx_mul_rd\[5\] pcpi_approx_mul_rd\[6\]
+ pcpi_approx_mul_rd\[7\] pcpi_approx_mul_rd\[8\] pcpi_approx_mul_rd\[9\] pcpi_approx_mul_ready
+ pcpi_approx_mul_wait pcpi_approx_mul_wr pcpi_div_rd\[0\] pcpi_div_rd\[10\] pcpi_div_rd\[11\]
+ pcpi_div_rd\[12\] pcpi_div_rd\[13\] pcpi_div_rd\[14\] pcpi_div_rd\[15\] pcpi_div_rd\[16\]
+ pcpi_div_rd\[17\] pcpi_div_rd\[18\] pcpi_div_rd\[19\] pcpi_div_rd\[1\] pcpi_div_rd\[20\]
+ pcpi_div_rd\[21\] pcpi_div_rd\[22\] pcpi_div_rd\[23\] pcpi_div_rd\[24\] pcpi_div_rd\[25\]
+ pcpi_div_rd\[26\] pcpi_div_rd\[27\] pcpi_div_rd\[28\] pcpi_div_rd\[29\] pcpi_div_rd\[2\]
+ pcpi_div_rd\[30\] pcpi_div_rd\[31\] pcpi_div_rd\[3\] pcpi_div_rd\[4\] pcpi_div_rd\[5\]
+ pcpi_div_rd\[6\] pcpi_div_rd\[7\] pcpi_div_rd\[8\] pcpi_div_rd\[9\] pcpi_div_ready
+ pcpi_div_wait pcpi_div_wr pcpi_exact_mul_rd\[0\] pcpi_exact_mul_rd\[10\] pcpi_exact_mul_rd\[11\]
+ pcpi_exact_mul_rd\[12\] pcpi_exact_mul_rd\[13\] pcpi_exact_mul_rd\[14\] pcpi_exact_mul_rd\[15\]
+ pcpi_exact_mul_rd\[16\] pcpi_exact_mul_rd\[17\] pcpi_exact_mul_rd\[18\] pcpi_exact_mul_rd\[19\]
+ pcpi_exact_mul_rd\[1\] pcpi_exact_mul_rd\[20\] pcpi_exact_mul_rd\[21\] pcpi_exact_mul_rd\[22\]
+ pcpi_exact_mul_rd\[23\] pcpi_exact_mul_rd\[24\] pcpi_exact_mul_rd\[25\] pcpi_exact_mul_rd\[26\]
+ pcpi_exact_mul_rd\[27\] pcpi_exact_mul_rd\[28\] pcpi_exact_mul_rd\[29\] pcpi_exact_mul_rd\[2\]
+ pcpi_exact_mul_rd\[30\] pcpi_exact_mul_rd\[31\] pcpi_exact_mul_rd\[3\] pcpi_exact_mul_rd\[4\]
+ pcpi_exact_mul_rd\[5\] pcpi_exact_mul_rd\[6\] pcpi_exact_mul_rd\[7\] pcpi_exact_mul_rd\[8\]
+ pcpi_exact_mul_rd\[9\] pcpi_exact_mul_ready pcpi_exact_mul_wait pcpi_exact_mul_wr
+ pcpi_insn\[0\] pcpi_insn\[10\] pcpi_insn\[11\] pcpi_insn\[12\] pcpi_insn\[13\] pcpi_insn\[14\]
+ pcpi_insn\[15\] pcpi_insn\[16\] pcpi_insn\[17\] pcpi_insn\[18\] pcpi_insn\[19\]
+ pcpi_insn\[1\] pcpi_insn\[20\] pcpi_insn\[21\] pcpi_insn\[22\] pcpi_insn\[23\] pcpi_insn\[24\]
+ pcpi_insn\[25\] pcpi_insn\[26\] pcpi_insn\[27\] pcpi_insn\[28\] pcpi_insn\[29\]
+ pcpi_insn\[2\] pcpi_insn\[30\] pcpi_insn\[31\] pcpi_insn\[3\] pcpi_insn\[4\] pcpi_insn\[5\]
+ pcpi_insn\[6\] pcpi_insn\[7\] pcpi_insn\[8\] pcpi_insn\[9\] pcpi_mul_rd\[0\] pcpi_mul_rd\[10\]
+ pcpi_mul_rd\[11\] pcpi_mul_rd\[12\] pcpi_mul_rd\[13\] pcpi_mul_rd\[14\] pcpi_mul_rd\[15\]
+ pcpi_mul_rd\[16\] pcpi_mul_rd\[17\] pcpi_mul_rd\[18\] pcpi_mul_rd\[19\] pcpi_mul_rd\[1\]
+ pcpi_mul_rd\[20\] pcpi_mul_rd\[21\] pcpi_mul_rd\[22\] pcpi_mul_rd\[23\] pcpi_mul_rd\[24\]
+ pcpi_mul_rd\[25\] pcpi_mul_rd\[26\] pcpi_mul_rd\[27\] pcpi_mul_rd\[28\] pcpi_mul_rd\[29\]
+ pcpi_mul_rd\[2\] pcpi_mul_rd\[30\] pcpi_mul_rd\[31\] pcpi_mul_rd\[3\] pcpi_mul_rd\[4\]
+ pcpi_mul_rd\[5\] pcpi_mul_rd\[6\] pcpi_mul_rd\[7\] pcpi_mul_rd\[8\] pcpi_mul_rd\[9\]
+ pcpi_mul_ready pcpi_mul_wait pcpi_mul_wr pcpi_rs1\[0\] pcpi_rs1\[10\] pcpi_rs1\[11\]
+ pcpi_rs1\[12\] pcpi_rs1\[13\] pcpi_rs1\[14\] pcpi_rs1\[15\] pcpi_rs1\[16\] pcpi_rs1\[17\]
+ pcpi_rs1\[18\] pcpi_rs1\[19\] pcpi_rs1\[1\] pcpi_rs1\[20\] pcpi_rs1\[21\] pcpi_rs1\[22\]
+ pcpi_rs1\[23\] pcpi_rs1\[24\] pcpi_rs1\[25\] pcpi_rs1\[26\] pcpi_rs1\[27\] pcpi_rs1\[28\]
+ pcpi_rs1\[29\] pcpi_rs1\[2\] pcpi_rs1\[30\] pcpi_rs1\[31\] pcpi_rs1\[3\] pcpi_rs1\[4\]
+ pcpi_rs1\[5\] pcpi_rs1\[6\] pcpi_rs1\[7\] pcpi_rs1\[8\] pcpi_rs1\[9\] pcpi_rs2\[0\]
+ pcpi_rs2\[10\] pcpi_rs2\[11\] pcpi_rs2\[12\] pcpi_rs2\[13\] pcpi_rs2\[14\] pcpi_rs2\[15\]
+ pcpi_rs2\[16\] pcpi_rs2\[17\] pcpi_rs2\[18\] pcpi_rs2\[19\] pcpi_rs2\[1\] pcpi_rs2\[20\]
+ pcpi_rs2\[21\] pcpi_rs2\[22\] pcpi_rs2\[23\] pcpi_rs2\[24\] pcpi_rs2\[25\] pcpi_rs2\[26\]
+ pcpi_rs2\[27\] pcpi_rs2\[28\] pcpi_rs2\[29\] pcpi_rs2\[2\] pcpi_rs2\[30\] pcpi_rs2\[31\]
+ pcpi_rs2\[3\] pcpi_rs2\[4\] pcpi_rs2\[5\] pcpi_rs2\[6\] pcpi_rs2\[7\] pcpi_rs2\[8\]
+ pcpi_rs2\[9\] pcpi_valid resetn vdd vss cpu
Xpcpi_exact_mul_inst_0 io_in[8] pcpi_insn\[0\] pcpi_insn\[10\] pcpi_insn\[11\] pcpi_insn\[12\]
+ pcpi_insn\[13\] pcpi_insn\[14\] pcpi_insn\[15\] pcpi_insn\[16\] pcpi_insn\[17\]
+ pcpi_insn\[18\] pcpi_insn\[19\] pcpi_insn\[1\] pcpi_insn\[20\] pcpi_insn\[21\] pcpi_insn\[22\]
+ pcpi_insn\[23\] pcpi_insn\[24\] pcpi_insn\[25\] pcpi_insn\[26\] pcpi_insn\[27\]
+ pcpi_insn\[28\] pcpi_insn\[29\] pcpi_insn\[2\] pcpi_insn\[30\] pcpi_insn\[31\] pcpi_insn\[3\]
+ pcpi_insn\[4\] pcpi_insn\[5\] pcpi_insn\[6\] pcpi_insn\[7\] pcpi_insn\[8\] pcpi_insn\[9\]
+ pcpi_exact_mul_rd\[0\] pcpi_exact_mul_rd\[10\] pcpi_exact_mul_rd\[11\] pcpi_exact_mul_rd\[12\]
+ pcpi_exact_mul_rd\[13\] pcpi_exact_mul_rd\[14\] pcpi_exact_mul_rd\[15\] pcpi_exact_mul_rd\[16\]
+ pcpi_exact_mul_rd\[17\] pcpi_exact_mul_rd\[18\] pcpi_exact_mul_rd\[19\] pcpi_exact_mul_rd\[1\]
+ pcpi_exact_mul_rd\[20\] pcpi_exact_mul_rd\[21\] pcpi_exact_mul_rd\[22\] pcpi_exact_mul_rd\[23\]
+ pcpi_exact_mul_rd\[24\] pcpi_exact_mul_rd\[25\] pcpi_exact_mul_rd\[26\] pcpi_exact_mul_rd\[27\]
+ pcpi_exact_mul_rd\[28\] pcpi_exact_mul_rd\[29\] pcpi_exact_mul_rd\[2\] pcpi_exact_mul_rd\[30\]
+ pcpi_exact_mul_rd\[31\] pcpi_exact_mul_rd\[3\] pcpi_exact_mul_rd\[4\] pcpi_exact_mul_rd\[5\]
+ pcpi_exact_mul_rd\[6\] pcpi_exact_mul_rd\[7\] pcpi_exact_mul_rd\[8\] pcpi_exact_mul_rd\[9\]
+ pcpi_exact_mul_ready pcpi_rs1\[0\] pcpi_rs1\[10\] pcpi_rs1\[11\] pcpi_rs1\[12\]
+ pcpi_rs1\[13\] pcpi_rs1\[14\] pcpi_rs1\[15\] pcpi_rs1\[16\] pcpi_rs1\[17\] pcpi_rs1\[18\]
+ pcpi_rs1\[19\] pcpi_rs1\[1\] pcpi_rs1\[20\] pcpi_rs1\[21\] pcpi_rs1\[22\] pcpi_rs1\[23\]
+ pcpi_rs1\[24\] pcpi_rs1\[25\] pcpi_rs1\[26\] pcpi_rs1\[27\] pcpi_rs1\[28\] pcpi_rs1\[29\]
+ pcpi_rs1\[2\] pcpi_rs1\[30\] pcpi_rs1\[31\] pcpi_rs1\[3\] pcpi_rs1\[4\] pcpi_rs1\[5\]
+ pcpi_rs1\[6\] pcpi_rs1\[7\] pcpi_rs1\[8\] pcpi_rs1\[9\] pcpi_rs2\[0\] pcpi_rs2\[10\]
+ pcpi_rs2\[11\] pcpi_rs2\[12\] pcpi_rs2\[13\] pcpi_rs2\[14\] pcpi_rs2\[15\] pcpi_rs2\[16\]
+ pcpi_rs2\[17\] pcpi_rs2\[18\] pcpi_rs2\[19\] pcpi_rs2\[1\] pcpi_rs2\[20\] pcpi_rs2\[21\]
+ pcpi_rs2\[22\] pcpi_rs2\[23\] pcpi_rs2\[24\] pcpi_rs2\[25\] pcpi_rs2\[26\] pcpi_rs2\[27\]
+ pcpi_rs2\[28\] pcpi_rs2\[29\] pcpi_rs2\[2\] pcpi_rs2\[30\] pcpi_rs2\[31\] pcpi_rs2\[3\]
+ pcpi_rs2\[4\] pcpi_rs2\[5\] pcpi_rs2\[6\] pcpi_rs2\[7\] pcpi_rs2\[8\] pcpi_rs2\[9\]
+ pcpi_valid pcpi_exact_mul_wait pcpi_exact_mul_wr resetn vdd vss pcpi_exact_mul
Xspimemio mem_addr\[0\] mem_addr\[10\] mem_addr\[11\] mem_addr\[12\] mem_addr\[13\]
+ mem_addr\[14\] mem_addr\[15\] mem_addr\[16\] mem_addr\[17\] mem_addr\[18\] mem_addr\[19\]
+ mem_addr\[1\] mem_addr\[20\] mem_addr\[21\] mem_addr\[22\] mem_addr\[23\] mem_addr\[2\]
+ mem_addr\[3\] mem_addr\[4\] mem_addr\[5\] mem_addr\[6\] mem_addr\[7\] mem_addr\[8\]
+ mem_addr\[9\] mem_wdata\[0\] mem_wdata\[10\] mem_wdata\[11\] mem_wdata\[12\] mem_wdata\[13\]
+ mem_wdata\[14\] mem_wdata\[15\] mem_wdata\[16\] mem_wdata\[17\] mem_wdata\[18\]
+ mem_wdata\[19\] mem_wdata\[1\] mem_wdata\[20\] mem_wdata\[21\] mem_wdata\[22\] mem_wdata\[23\]
+ mem_wdata\[24\] mem_wdata\[25\] mem_wdata\[26\] mem_wdata\[27\] mem_wdata\[28\]
+ mem_wdata\[29\] mem_wdata\[2\] mem_wdata\[30\] mem_wdata\[31\] mem_wdata\[3\] mem_wdata\[4\]
+ mem_wdata\[5\] mem_wdata\[6\] mem_wdata\[7\] mem_wdata\[8\] mem_wdata\[9\] spimemio_cfgreg_do\[0\]
+ spimemio_cfgreg_do\[10\] spimemio_cfgreg_do\[11\] spimemio_cfgreg_do\[12\] spimemio_cfgreg_do\[13\]
+ spimemio_cfgreg_do\[14\] spimemio_cfgreg_do\[15\] spimemio_cfgreg_do\[16\] spimemio_cfgreg_do\[17\]
+ spimemio_cfgreg_do\[18\] spimemio_cfgreg_do\[19\] spimemio_cfgreg_do\[1\] spimemio_cfgreg_do\[20\]
+ spimemio_cfgreg_do\[21\] spimemio_cfgreg_do\[22\] spimemio_cfgreg_do\[23\] spimemio_cfgreg_do\[24\]
+ spimemio_cfgreg_do\[25\] spimemio_cfgreg_do\[26\] spimemio_cfgreg_do\[27\] spimemio_cfgreg_do\[28\]
+ spimemio_cfgreg_do\[29\] spimemio_cfgreg_do\[2\] spimemio_cfgreg_do\[30\] spimemio_cfgreg_do\[31\]
+ spimemio_cfgreg_do\[3\] spimemio_cfgreg_do\[4\] spimemio_cfgreg_do\[5\] spimemio_cfgreg_do\[6\]
+ spimemio_cfgreg_do\[7\] spimemio_cfgreg_do\[8\] spimemio_cfgreg_do\[9\] spimemio_cfgreg_we\[0\]
+ spimemio_cfgreg_we\[1\] spimemio_cfgreg_we\[2\] spimemio_cfgreg_we\[3\] io_in[8]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_oeb[10] io_oeb[11]
+ io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] spimem_rdata\[0\] spimem_rdata\[10\] spimem_rdata\[11\] spimem_rdata\[12\]
+ spimem_rdata\[13\] spimem_rdata\[14\] spimem_rdata\[15\] spimem_rdata\[16\] spimem_rdata\[17\]
+ spimem_rdata\[18\] spimem_rdata\[19\] spimem_rdata\[1\] spimem_rdata\[20\] spimem_rdata\[21\]
+ spimem_rdata\[22\] spimem_rdata\[23\] spimem_rdata\[24\] spimem_rdata\[25\] spimem_rdata\[26\]
+ spimem_rdata\[27\] spimem_rdata\[28\] spimem_rdata\[29\] spimem_rdata\[2\] spimem_rdata\[30\]
+ spimem_rdata\[31\] spimem_rdata\[3\] spimem_rdata\[4\] spimem_rdata\[5\] spimem_rdata\[6\]
+ spimem_rdata\[7\] spimem_rdata\[8\] spimem_rdata\[9\] spimem_ready resetn spimem_valid
+ vdd vss spimemio
Xsimpleuart io_in[8] mem_wdata\[0\] mem_wdata\[10\] mem_wdata\[11\] mem_wdata\[12\]
+ mem_wdata\[13\] mem_wdata\[14\] mem_wdata\[15\] mem_wdata\[16\] mem_wdata\[17\]
+ mem_wdata\[18\] mem_wdata\[19\] mem_wdata\[1\] mem_wdata\[20\] mem_wdata\[21\] mem_wdata\[22\]
+ mem_wdata\[23\] mem_wdata\[24\] mem_wdata\[25\] mem_wdata\[26\] mem_wdata\[27\]
+ mem_wdata\[28\] mem_wdata\[29\] mem_wdata\[2\] mem_wdata\[30\] mem_wdata\[31\] mem_wdata\[3\]
+ mem_wdata\[4\] mem_wdata\[5\] mem_wdata\[6\] mem_wdata\[7\] mem_wdata\[8\] mem_wdata\[9\]
+ simpleuart_reg_dat_do\[0\] simpleuart_reg_dat_do\[10\] simpleuart_reg_dat_do\[11\]
+ simpleuart_reg_dat_do\[12\] simpleuart_reg_dat_do\[13\] simpleuart_reg_dat_do\[14\]
+ simpleuart_reg_dat_do\[15\] simpleuart_reg_dat_do\[16\] simpleuart_reg_dat_do\[17\]
+ simpleuart_reg_dat_do\[18\] simpleuart_reg_dat_do\[19\] simpleuart_reg_dat_do\[1\]
+ simpleuart_reg_dat_do\[20\] simpleuart_reg_dat_do\[21\] simpleuart_reg_dat_do\[22\]
+ simpleuart_reg_dat_do\[23\] simpleuart_reg_dat_do\[24\] simpleuart_reg_dat_do\[25\]
+ simpleuart_reg_dat_do\[26\] simpleuart_reg_dat_do\[27\] simpleuart_reg_dat_do\[28\]
+ simpleuart_reg_dat_do\[29\] simpleuart_reg_dat_do\[2\] simpleuart_reg_dat_do\[30\]
+ simpleuart_reg_dat_do\[31\] simpleuart_reg_dat_do\[3\] simpleuart_reg_dat_do\[4\]
+ simpleuart_reg_dat_do\[5\] simpleuart_reg_dat_do\[6\] simpleuart_reg_dat_do\[7\]
+ simpleuart_reg_dat_do\[8\] simpleuart_reg_dat_do\[9\] simpleuart_dat_re simpleuart_reg_dat_wait
+ simpleuart_dat_we mem_wdata\[0\] mem_wdata\[10\] mem_wdata\[11\] mem_wdata\[12\]
+ mem_wdata\[13\] mem_wdata\[14\] mem_wdata\[15\] mem_wdata\[16\] mem_wdata\[17\]
+ mem_wdata\[18\] mem_wdata\[19\] mem_wdata\[1\] mem_wdata\[20\] mem_wdata\[21\] mem_wdata\[22\]
+ mem_wdata\[23\] mem_wdata\[24\] mem_wdata\[25\] mem_wdata\[26\] mem_wdata\[27\]
+ mem_wdata\[28\] mem_wdata\[29\] mem_wdata\[2\] mem_wdata\[30\] mem_wdata\[31\] mem_wdata\[3\]
+ mem_wdata\[4\] mem_wdata\[5\] mem_wdata\[6\] mem_wdata\[7\] mem_wdata\[8\] mem_wdata\[9\]
+ simpleuart_reg_div_do\[0\] simpleuart_reg_div_do\[10\] simpleuart_reg_div_do\[11\]
+ simpleuart_reg_div_do\[12\] simpleuart_reg_div_do\[13\] simpleuart_reg_div_do\[14\]
+ simpleuart_reg_div_do\[15\] simpleuart_reg_div_do\[16\] simpleuart_reg_div_do\[17\]
+ simpleuart_reg_div_do\[18\] simpleuart_reg_div_do\[19\] simpleuart_reg_div_do\[1\]
+ simpleuart_reg_div_do\[20\] simpleuart_reg_div_do\[21\] simpleuart_reg_div_do\[22\]
+ simpleuart_reg_div_do\[23\] simpleuart_reg_div_do\[24\] simpleuart_reg_div_do\[25\]
+ simpleuart_reg_div_do\[26\] simpleuart_reg_div_do\[27\] simpleuart_reg_div_do\[28\]
+ simpleuart_reg_div_do\[29\] simpleuart_reg_div_do\[2\] simpleuart_reg_div_do\[30\]
+ simpleuart_reg_div_do\[31\] simpleuart_reg_div_do\[3\] simpleuart_reg_div_do\[4\]
+ simpleuart_reg_div_do\[5\] simpleuart_reg_div_do\[6\] simpleuart_reg_div_do\[7\]
+ simpleuart_reg_div_do\[8\] simpleuart_reg_div_do\[9\] simpleuart_div_we\[0\] simpleuart_div_we\[1\]
+ simpleuart_div_we\[2\] simpleuart_div_we\[3\] resetn io_in[16] io_in[17] io_oeb[16]
+ io_oeb[17] io_out[16] io_out[17] vdd vss simpleuart
Xpcpi_div_inst_0 io_in[8] pcpi_div_rd\[0\] pcpi_div_rd\[10\] pcpi_div_rd\[11\] pcpi_div_rd\[12\]
+ pcpi_div_rd\[13\] pcpi_div_rd\[14\] pcpi_div_rd\[15\] pcpi_div_rd\[16\] pcpi_div_rd\[17\]
+ pcpi_div_rd\[18\] pcpi_div_rd\[19\] pcpi_div_rd\[1\] pcpi_div_rd\[20\] pcpi_div_rd\[21\]
+ pcpi_div_rd\[22\] pcpi_div_rd\[23\] pcpi_div_rd\[24\] pcpi_div_rd\[25\] pcpi_div_rd\[26\]
+ pcpi_div_rd\[27\] pcpi_div_rd\[28\] pcpi_div_rd\[29\] pcpi_div_rd\[2\] pcpi_div_rd\[30\]
+ pcpi_div_rd\[31\] pcpi_div_rd\[3\] pcpi_div_rd\[4\] pcpi_div_rd\[5\] pcpi_div_rd\[6\]
+ pcpi_div_rd\[7\] pcpi_div_rd\[8\] pcpi_div_rd\[9\] pcpi_div_ready pcpi_valid pcpi_div_wait
+ pcpi_div_wr pcpi_insn\[0\] pcpi_insn\[10\] pcpi_insn\[11\] pcpi_insn\[12\] pcpi_insn\[13\]
+ pcpi_insn\[14\] pcpi_insn\[15\] pcpi_insn\[16\] pcpi_insn\[17\] pcpi_insn\[18\]
+ pcpi_insn\[19\] pcpi_insn\[1\] pcpi_insn\[20\] pcpi_insn\[21\] pcpi_insn\[22\] pcpi_insn\[23\]
+ pcpi_insn\[24\] pcpi_insn\[25\] pcpi_insn\[26\] pcpi_insn\[27\] pcpi_insn\[28\]
+ pcpi_insn\[29\] pcpi_insn\[2\] pcpi_insn\[30\] pcpi_insn\[31\] pcpi_insn\[3\] pcpi_insn\[4\]
+ pcpi_insn\[5\] pcpi_insn\[6\] pcpi_insn\[7\] pcpi_insn\[8\] pcpi_insn\[9\] pcpi_rs1\[0\]
+ pcpi_rs1\[10\] pcpi_rs1\[11\] pcpi_rs1\[12\] pcpi_rs1\[13\] pcpi_rs1\[14\] pcpi_rs1\[15\]
+ pcpi_rs1\[16\] pcpi_rs1\[17\] pcpi_rs1\[18\] pcpi_rs1\[19\] pcpi_rs1\[1\] pcpi_rs1\[20\]
+ pcpi_rs1\[21\] pcpi_rs1\[22\] pcpi_rs1\[23\] pcpi_rs1\[24\] pcpi_rs1\[25\] pcpi_rs1\[26\]
+ pcpi_rs1\[27\] pcpi_rs1\[28\] pcpi_rs1\[29\] pcpi_rs1\[2\] pcpi_rs1\[30\] pcpi_rs1\[31\]
+ pcpi_rs1\[3\] pcpi_rs1\[4\] pcpi_rs1\[5\] pcpi_rs1\[6\] pcpi_rs1\[7\] pcpi_rs1\[8\]
+ pcpi_rs1\[9\] pcpi_rs2\[0\] pcpi_rs2\[10\] pcpi_rs2\[11\] pcpi_rs2\[12\] pcpi_rs2\[13\]
+ pcpi_rs2\[14\] pcpi_rs2\[15\] pcpi_rs2\[16\] pcpi_rs2\[17\] pcpi_rs2\[18\] pcpi_rs2\[19\]
+ pcpi_rs2\[1\] pcpi_rs2\[20\] pcpi_rs2\[21\] pcpi_rs2\[22\] pcpi_rs2\[23\] pcpi_rs2\[24\]
+ pcpi_rs2\[25\] pcpi_rs2\[26\] pcpi_rs2\[27\] pcpi_rs2\[28\] pcpi_rs2\[29\] pcpi_rs2\[2\]
+ pcpi_rs2\[30\] pcpi_rs2\[31\] pcpi_rs2\[3\] pcpi_rs2\[4\] pcpi_rs2\[5\] pcpi_rs2\[6\]
+ pcpi_rs2\[7\] pcpi_rs2\[8\] pcpi_rs2\[9\] resetn vdd vss pcpi_div
.ends


magic
tech gf180mcuD
magscale 1 10
timestamp 1702206252
<< nwell >>
rect 1258 25440 518646 26304
rect 1258 23872 518646 24736
rect 1258 22304 518646 23168
rect 1258 20736 518646 21600
rect 1258 19168 518646 20032
rect 1258 17600 518646 18464
rect 1258 16032 518646 16896
rect 1258 14464 518646 15328
rect 1258 12896 518646 13760
rect 1258 11328 518646 12192
rect 1258 9760 518646 10624
rect 1258 8192 518646 9056
rect 1258 7463 279000 7488
rect 1258 6649 518646 7463
rect 1258 6624 285048 6649
rect 1258 5895 210680 5920
rect 1258 5081 518646 5895
rect 1258 5056 213101 5081
rect 1258 4327 210680 4352
rect 1258 3513 518646 4327
rect 1258 3488 273422 3513
<< pwell >>
rect 1258 26304 518646 26742
rect 1258 24736 518646 25440
rect 1258 23168 518646 23872
rect 1258 21600 518646 22304
rect 1258 20032 518646 20736
rect 1258 18464 518646 19168
rect 1258 16896 518646 17600
rect 1258 15328 518646 16032
rect 1258 13760 518646 14464
rect 1258 12192 518646 12896
rect 1258 10624 518646 11328
rect 1258 9056 518646 9760
rect 1258 7488 518646 8192
rect 1258 5920 518646 6624
rect 1258 4352 518646 5056
rect 1258 3050 518646 3488
<< obsm1 >>
rect 1344 1710 518720 26716
<< metal2 >>
rect 24640 0 24752 800
rect 26208 0 26320 800
rect 27776 0 27888 800
rect 29344 0 29456 800
rect 30912 0 31024 800
rect 32480 0 32592 800
rect 34048 0 34160 800
rect 35616 0 35728 800
rect 37184 0 37296 800
rect 38752 0 38864 800
rect 40320 0 40432 800
rect 41888 0 42000 800
rect 43456 0 43568 800
rect 45024 0 45136 800
rect 46592 0 46704 800
rect 48160 0 48272 800
rect 49728 0 49840 800
rect 51296 0 51408 800
rect 52864 0 52976 800
rect 54432 0 54544 800
rect 56000 0 56112 800
rect 57568 0 57680 800
rect 59136 0 59248 800
rect 60704 0 60816 800
rect 62272 0 62384 800
rect 63840 0 63952 800
rect 65408 0 65520 800
rect 66976 0 67088 800
rect 68544 0 68656 800
rect 70112 0 70224 800
rect 71680 0 71792 800
rect 73248 0 73360 800
rect 74816 0 74928 800
rect 76384 0 76496 800
rect 77952 0 78064 800
rect 79520 0 79632 800
rect 81088 0 81200 800
rect 82656 0 82768 800
rect 84224 0 84336 800
rect 85792 0 85904 800
rect 87360 0 87472 800
rect 88928 0 89040 800
rect 90496 0 90608 800
rect 92064 0 92176 800
rect 93632 0 93744 800
rect 95200 0 95312 800
rect 96768 0 96880 800
rect 98336 0 98448 800
rect 99904 0 100016 800
rect 101472 0 101584 800
rect 103040 0 103152 800
rect 104608 0 104720 800
rect 106176 0 106288 800
rect 107744 0 107856 800
rect 109312 0 109424 800
rect 110880 0 110992 800
rect 112448 0 112560 800
rect 114016 0 114128 800
rect 115584 0 115696 800
rect 117152 0 117264 800
rect 118720 0 118832 800
rect 120288 0 120400 800
rect 121856 0 121968 800
rect 123424 0 123536 800
rect 124992 0 125104 800
rect 126560 0 126672 800
rect 128128 0 128240 800
rect 129696 0 129808 800
rect 131264 0 131376 800
rect 132832 0 132944 800
rect 134400 0 134512 800
rect 135968 0 136080 800
rect 137536 0 137648 800
rect 139104 0 139216 800
rect 140672 0 140784 800
rect 142240 0 142352 800
rect 143808 0 143920 800
rect 145376 0 145488 800
rect 146944 0 147056 800
rect 148512 0 148624 800
rect 150080 0 150192 800
rect 151648 0 151760 800
rect 153216 0 153328 800
rect 154784 0 154896 800
rect 156352 0 156464 800
rect 157920 0 158032 800
rect 159488 0 159600 800
rect 161056 0 161168 800
rect 162624 0 162736 800
rect 164192 0 164304 800
rect 165760 0 165872 800
rect 167328 0 167440 800
rect 168896 0 169008 800
rect 170464 0 170576 800
rect 172032 0 172144 800
rect 173600 0 173712 800
rect 175168 0 175280 800
rect 176736 0 176848 800
rect 178304 0 178416 800
rect 179872 0 179984 800
rect 181440 0 181552 800
rect 183008 0 183120 800
rect 184576 0 184688 800
rect 186144 0 186256 800
rect 187712 0 187824 800
rect 189280 0 189392 800
rect 190848 0 190960 800
rect 192416 0 192528 800
rect 193984 0 194096 800
rect 195552 0 195664 800
rect 197120 0 197232 800
rect 198688 0 198800 800
rect 200256 0 200368 800
rect 201824 0 201936 800
rect 203392 0 203504 800
rect 204960 0 205072 800
rect 206528 0 206640 800
rect 208096 0 208208 800
rect 209664 0 209776 800
rect 211232 0 211344 800
rect 212800 0 212912 800
rect 214368 0 214480 800
rect 215936 0 216048 800
rect 217504 0 217616 800
rect 219072 0 219184 800
rect 220640 0 220752 800
rect 222208 0 222320 800
rect 223776 0 223888 800
rect 225344 0 225456 800
rect 226912 0 227024 800
rect 228480 0 228592 800
rect 230048 0 230160 800
rect 231616 0 231728 800
rect 233184 0 233296 800
rect 234752 0 234864 800
rect 236320 0 236432 800
rect 237888 0 238000 800
rect 239456 0 239568 800
rect 241024 0 241136 800
rect 242592 0 242704 800
rect 244160 0 244272 800
rect 245728 0 245840 800
rect 247296 0 247408 800
rect 248864 0 248976 800
rect 250432 0 250544 800
rect 252000 0 252112 800
rect 253568 0 253680 800
rect 255136 0 255248 800
rect 256704 0 256816 800
rect 258272 0 258384 800
rect 259840 0 259952 800
rect 261408 0 261520 800
rect 262976 0 263088 800
rect 264544 0 264656 800
rect 266112 0 266224 800
rect 267680 0 267792 800
rect 269248 0 269360 800
rect 270816 0 270928 800
rect 272384 0 272496 800
rect 273952 0 274064 800
rect 275520 0 275632 800
rect 277088 0 277200 800
rect 278656 0 278768 800
rect 280224 0 280336 800
rect 281792 0 281904 800
rect 283360 0 283472 800
rect 284928 0 285040 800
rect 286496 0 286608 800
rect 288064 0 288176 800
rect 289632 0 289744 800
rect 291200 0 291312 800
rect 292768 0 292880 800
rect 294336 0 294448 800
rect 295904 0 296016 800
rect 297472 0 297584 800
rect 299040 0 299152 800
rect 300608 0 300720 800
rect 302176 0 302288 800
rect 303744 0 303856 800
rect 305312 0 305424 800
rect 306880 0 306992 800
rect 308448 0 308560 800
rect 310016 0 310128 800
rect 311584 0 311696 800
rect 313152 0 313264 800
rect 314720 0 314832 800
rect 316288 0 316400 800
rect 317856 0 317968 800
rect 319424 0 319536 800
rect 320992 0 321104 800
rect 322560 0 322672 800
rect 324128 0 324240 800
rect 325696 0 325808 800
rect 327264 0 327376 800
rect 328832 0 328944 800
rect 330400 0 330512 800
rect 331968 0 332080 800
rect 333536 0 333648 800
rect 335104 0 335216 800
rect 336672 0 336784 800
rect 338240 0 338352 800
rect 339808 0 339920 800
rect 341376 0 341488 800
rect 342944 0 343056 800
rect 344512 0 344624 800
rect 346080 0 346192 800
rect 347648 0 347760 800
rect 349216 0 349328 800
rect 350784 0 350896 800
rect 352352 0 352464 800
rect 353920 0 354032 800
rect 355488 0 355600 800
rect 357056 0 357168 800
rect 358624 0 358736 800
rect 360192 0 360304 800
rect 361760 0 361872 800
rect 363328 0 363440 800
rect 364896 0 365008 800
rect 366464 0 366576 800
rect 368032 0 368144 800
rect 369600 0 369712 800
rect 371168 0 371280 800
rect 372736 0 372848 800
rect 374304 0 374416 800
rect 375872 0 375984 800
rect 377440 0 377552 800
rect 379008 0 379120 800
rect 380576 0 380688 800
rect 382144 0 382256 800
rect 383712 0 383824 800
rect 385280 0 385392 800
rect 386848 0 386960 800
rect 388416 0 388528 800
rect 389984 0 390096 800
rect 391552 0 391664 800
rect 393120 0 393232 800
rect 394688 0 394800 800
rect 396256 0 396368 800
rect 397824 0 397936 800
rect 399392 0 399504 800
rect 400960 0 401072 800
rect 402528 0 402640 800
rect 404096 0 404208 800
rect 405664 0 405776 800
rect 407232 0 407344 800
rect 408800 0 408912 800
rect 410368 0 410480 800
rect 411936 0 412048 800
rect 413504 0 413616 800
rect 415072 0 415184 800
rect 416640 0 416752 800
rect 418208 0 418320 800
rect 419776 0 419888 800
rect 421344 0 421456 800
rect 422912 0 423024 800
rect 424480 0 424592 800
rect 426048 0 426160 800
rect 427616 0 427728 800
rect 429184 0 429296 800
rect 430752 0 430864 800
rect 432320 0 432432 800
rect 433888 0 434000 800
rect 435456 0 435568 800
rect 437024 0 437136 800
rect 438592 0 438704 800
rect 440160 0 440272 800
rect 441728 0 441840 800
rect 443296 0 443408 800
rect 444864 0 444976 800
rect 446432 0 446544 800
rect 448000 0 448112 800
rect 449568 0 449680 800
rect 451136 0 451248 800
rect 452704 0 452816 800
rect 454272 0 454384 800
rect 455840 0 455952 800
rect 457408 0 457520 800
rect 458976 0 459088 800
rect 460544 0 460656 800
rect 462112 0 462224 800
rect 463680 0 463792 800
rect 465248 0 465360 800
rect 466816 0 466928 800
rect 468384 0 468496 800
rect 469952 0 470064 800
rect 471520 0 471632 800
rect 473088 0 473200 800
rect 474656 0 474768 800
rect 476224 0 476336 800
rect 477792 0 477904 800
rect 479360 0 479472 800
rect 480928 0 481040 800
rect 482496 0 482608 800
rect 484064 0 484176 800
rect 485632 0 485744 800
rect 487200 0 487312 800
rect 488768 0 488880 800
rect 490336 0 490448 800
rect 491904 0 492016 800
rect 493472 0 493584 800
rect 495040 0 495152 800
<< obsm2 >>
rect 24668 860 518692 27870
rect 24812 700 26148 860
rect 26380 700 27716 860
rect 27948 700 29284 860
rect 29516 700 30852 860
rect 31084 700 32420 860
rect 32652 700 33988 860
rect 34220 700 35556 860
rect 35788 700 37124 860
rect 37356 700 38692 860
rect 38924 700 40260 860
rect 40492 700 41828 860
rect 42060 700 43396 860
rect 43628 700 44964 860
rect 45196 700 46532 860
rect 46764 700 48100 860
rect 48332 700 49668 860
rect 49900 700 51236 860
rect 51468 700 52804 860
rect 53036 700 54372 860
rect 54604 700 55940 860
rect 56172 700 57508 860
rect 57740 700 59076 860
rect 59308 700 60644 860
rect 60876 700 62212 860
rect 62444 700 63780 860
rect 64012 700 65348 860
rect 65580 700 66916 860
rect 67148 700 68484 860
rect 68716 700 70052 860
rect 70284 700 71620 860
rect 71852 700 73188 860
rect 73420 700 74756 860
rect 74988 700 76324 860
rect 76556 700 77892 860
rect 78124 700 79460 860
rect 79692 700 81028 860
rect 81260 700 82596 860
rect 82828 700 84164 860
rect 84396 700 85732 860
rect 85964 700 87300 860
rect 87532 700 88868 860
rect 89100 700 90436 860
rect 90668 700 92004 860
rect 92236 700 93572 860
rect 93804 700 95140 860
rect 95372 700 96708 860
rect 96940 700 98276 860
rect 98508 700 99844 860
rect 100076 700 101412 860
rect 101644 700 102980 860
rect 103212 700 104548 860
rect 104780 700 106116 860
rect 106348 700 107684 860
rect 107916 700 109252 860
rect 109484 700 110820 860
rect 111052 700 112388 860
rect 112620 700 113956 860
rect 114188 700 115524 860
rect 115756 700 117092 860
rect 117324 700 118660 860
rect 118892 700 120228 860
rect 120460 700 121796 860
rect 122028 700 123364 860
rect 123596 700 124932 860
rect 125164 700 126500 860
rect 126732 700 128068 860
rect 128300 700 129636 860
rect 129868 700 131204 860
rect 131436 700 132772 860
rect 133004 700 134340 860
rect 134572 700 135908 860
rect 136140 700 137476 860
rect 137708 700 139044 860
rect 139276 700 140612 860
rect 140844 700 142180 860
rect 142412 700 143748 860
rect 143980 700 145316 860
rect 145548 700 146884 860
rect 147116 700 148452 860
rect 148684 700 150020 860
rect 150252 700 151588 860
rect 151820 700 153156 860
rect 153388 700 154724 860
rect 154956 700 156292 860
rect 156524 700 157860 860
rect 158092 700 159428 860
rect 159660 700 160996 860
rect 161228 700 162564 860
rect 162796 700 164132 860
rect 164364 700 165700 860
rect 165932 700 167268 860
rect 167500 700 168836 860
rect 169068 700 170404 860
rect 170636 700 171972 860
rect 172204 700 173540 860
rect 173772 700 175108 860
rect 175340 700 176676 860
rect 176908 700 178244 860
rect 178476 700 179812 860
rect 180044 700 181380 860
rect 181612 700 182948 860
rect 183180 700 184516 860
rect 184748 700 186084 860
rect 186316 700 187652 860
rect 187884 700 189220 860
rect 189452 700 190788 860
rect 191020 700 192356 860
rect 192588 700 193924 860
rect 194156 700 195492 860
rect 195724 700 197060 860
rect 197292 700 198628 860
rect 198860 700 200196 860
rect 200428 700 201764 860
rect 201996 700 203332 860
rect 203564 700 204900 860
rect 205132 700 206468 860
rect 206700 700 208036 860
rect 208268 700 209604 860
rect 209836 700 211172 860
rect 211404 700 212740 860
rect 212972 700 214308 860
rect 214540 700 215876 860
rect 216108 700 217444 860
rect 217676 700 219012 860
rect 219244 700 220580 860
rect 220812 700 222148 860
rect 222380 700 223716 860
rect 223948 700 225284 860
rect 225516 700 226852 860
rect 227084 700 228420 860
rect 228652 700 229988 860
rect 230220 700 231556 860
rect 231788 700 233124 860
rect 233356 700 234692 860
rect 234924 700 236260 860
rect 236492 700 237828 860
rect 238060 700 239396 860
rect 239628 700 240964 860
rect 241196 700 242532 860
rect 242764 700 244100 860
rect 244332 700 245668 860
rect 245900 700 247236 860
rect 247468 700 248804 860
rect 249036 700 250372 860
rect 250604 700 251940 860
rect 252172 700 253508 860
rect 253740 700 255076 860
rect 255308 700 256644 860
rect 256876 700 258212 860
rect 258444 700 259780 860
rect 260012 700 261348 860
rect 261580 700 262916 860
rect 263148 700 264484 860
rect 264716 700 266052 860
rect 266284 700 267620 860
rect 267852 700 269188 860
rect 269420 700 270756 860
rect 270988 700 272324 860
rect 272556 700 273892 860
rect 274124 700 275460 860
rect 275692 700 277028 860
rect 277260 700 278596 860
rect 278828 700 280164 860
rect 280396 700 281732 860
rect 281964 700 283300 860
rect 283532 700 284868 860
rect 285100 700 286436 860
rect 286668 700 288004 860
rect 288236 700 289572 860
rect 289804 700 291140 860
rect 291372 700 292708 860
rect 292940 700 294276 860
rect 294508 700 295844 860
rect 296076 700 297412 860
rect 297644 700 298980 860
rect 299212 700 300548 860
rect 300780 700 302116 860
rect 302348 700 303684 860
rect 303916 700 305252 860
rect 305484 700 306820 860
rect 307052 700 308388 860
rect 308620 700 309956 860
rect 310188 700 311524 860
rect 311756 700 313092 860
rect 313324 700 314660 860
rect 314892 700 316228 860
rect 316460 700 317796 860
rect 318028 700 319364 860
rect 319596 700 320932 860
rect 321164 700 322500 860
rect 322732 700 324068 860
rect 324300 700 325636 860
rect 325868 700 327204 860
rect 327436 700 328772 860
rect 329004 700 330340 860
rect 330572 700 331908 860
rect 332140 700 333476 860
rect 333708 700 335044 860
rect 335276 700 336612 860
rect 336844 700 338180 860
rect 338412 700 339748 860
rect 339980 700 341316 860
rect 341548 700 342884 860
rect 343116 700 344452 860
rect 344684 700 346020 860
rect 346252 700 347588 860
rect 347820 700 349156 860
rect 349388 700 350724 860
rect 350956 700 352292 860
rect 352524 700 353860 860
rect 354092 700 355428 860
rect 355660 700 356996 860
rect 357228 700 358564 860
rect 358796 700 360132 860
rect 360364 700 361700 860
rect 361932 700 363268 860
rect 363500 700 364836 860
rect 365068 700 366404 860
rect 366636 700 367972 860
rect 368204 700 369540 860
rect 369772 700 371108 860
rect 371340 700 372676 860
rect 372908 700 374244 860
rect 374476 700 375812 860
rect 376044 700 377380 860
rect 377612 700 378948 860
rect 379180 700 380516 860
rect 380748 700 382084 860
rect 382316 700 383652 860
rect 383884 700 385220 860
rect 385452 700 386788 860
rect 387020 700 388356 860
rect 388588 700 389924 860
rect 390156 700 391492 860
rect 391724 700 393060 860
rect 393292 700 394628 860
rect 394860 700 396196 860
rect 396428 700 397764 860
rect 397996 700 399332 860
rect 399564 700 400900 860
rect 401132 700 402468 860
rect 402700 700 404036 860
rect 404268 700 405604 860
rect 405836 700 407172 860
rect 407404 700 408740 860
rect 408972 700 410308 860
rect 410540 700 411876 860
rect 412108 700 413444 860
rect 413676 700 415012 860
rect 415244 700 416580 860
rect 416812 700 418148 860
rect 418380 700 419716 860
rect 419948 700 421284 860
rect 421516 700 422852 860
rect 423084 700 424420 860
rect 424652 700 425988 860
rect 426220 700 427556 860
rect 427788 700 429124 860
rect 429356 700 430692 860
rect 430924 700 432260 860
rect 432492 700 433828 860
rect 434060 700 435396 860
rect 435628 700 436964 860
rect 437196 700 438532 860
rect 438764 700 440100 860
rect 440332 700 441668 860
rect 441900 700 443236 860
rect 443468 700 444804 860
rect 445036 700 446372 860
rect 446604 700 447940 860
rect 448172 700 449508 860
rect 449740 700 451076 860
rect 451308 700 452644 860
rect 452876 700 454212 860
rect 454444 700 455780 860
rect 456012 700 457348 860
rect 457580 700 458916 860
rect 459148 700 460484 860
rect 460716 700 462052 860
rect 462284 700 463620 860
rect 463852 700 465188 860
rect 465420 700 466756 860
rect 466988 700 468324 860
rect 468556 700 469892 860
rect 470124 700 471460 860
rect 471692 700 473028 860
rect 473260 700 474596 860
rect 474828 700 476164 860
rect 476396 700 477732 860
rect 477964 700 479300 860
rect 479532 700 480868 860
rect 481100 700 482436 860
rect 482668 700 484004 860
rect 484236 700 485572 860
rect 485804 700 487140 860
rect 487372 700 488708 860
rect 488940 700 490276 860
rect 490508 700 491844 860
rect 492076 700 493412 860
rect 493644 700 494980 860
rect 495212 700 518692 860
<< metal3 >>
rect 519200 27776 520000 27888
rect 519200 26656 520000 26768
rect 519200 25536 520000 25648
rect 519200 24416 520000 24528
rect 519200 23296 520000 23408
rect 519200 22176 520000 22288
rect 519200 21056 520000 21168
rect 519200 19936 520000 20048
rect 519200 18816 520000 18928
rect 519200 17696 520000 17808
rect 519200 16576 520000 16688
rect 519200 15456 520000 15568
rect 519200 14336 520000 14448
rect 519200 13216 520000 13328
rect 519200 12096 520000 12208
rect 519200 10976 520000 11088
rect 519200 9856 520000 9968
rect 519200 8736 520000 8848
rect 519200 7616 520000 7728
rect 519200 6496 520000 6608
rect 519200 5376 520000 5488
rect 519200 4256 520000 4368
rect 519200 3136 520000 3248
rect 519200 2016 520000 2128
<< obsm3 >>
rect 24658 27716 519140 27860
rect 24658 26828 519200 27716
rect 24658 26596 519140 26828
rect 24658 25708 519200 26596
rect 24658 25476 519140 25708
rect 24658 24588 519200 25476
rect 24658 24356 519140 24588
rect 24658 23468 519200 24356
rect 24658 23236 519140 23468
rect 24658 22348 519200 23236
rect 24658 22116 519140 22348
rect 24658 21228 519200 22116
rect 24658 20996 519140 21228
rect 24658 20108 519200 20996
rect 24658 19876 519140 20108
rect 24658 18988 519200 19876
rect 24658 18756 519140 18988
rect 24658 17868 519200 18756
rect 24658 17636 519140 17868
rect 24658 16748 519200 17636
rect 24658 16516 519140 16748
rect 24658 15628 519200 16516
rect 24658 15396 519140 15628
rect 24658 14508 519200 15396
rect 24658 14276 519140 14508
rect 24658 13388 519200 14276
rect 24658 13156 519140 13388
rect 24658 12268 519200 13156
rect 24658 12036 519140 12268
rect 24658 11148 519200 12036
rect 24658 10916 519140 11148
rect 24658 10028 519200 10916
rect 24658 9796 519140 10028
rect 24658 8908 519200 9796
rect 24658 8676 519140 8908
rect 24658 7788 519200 8676
rect 24658 7556 519140 7788
rect 24658 6668 519200 7556
rect 24658 6436 519140 6668
rect 24658 5548 519200 6436
rect 24658 5316 519140 5548
rect 24658 4428 519200 5316
rect 24658 4196 519140 4428
rect 24658 3308 519200 4196
rect 24658 3076 519140 3308
rect 24658 2188 519200 3076
rect 24658 1956 519140 2188
rect 24658 1036 519200 1956
<< metal4 >>
rect 65836 3076 66156 26716
rect 130488 3076 130808 26716
rect 195140 3076 195460 26716
rect 259792 3076 260112 26716
rect 324444 3076 324764 26716
rect 389096 3076 389416 26716
rect 453748 3076 454068 26716
rect 518400 3076 518720 26716
<< obsm4 >>
rect 286188 3602 286244 4014
<< labels >>
rlabel metal3 s 519200 2016 520000 2128 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 519200 5376 520000 5488 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 519200 8736 520000 8848 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 519200 12096 520000 12208 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 519200 15456 520000 15568 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 519200 18816 520000 18928 6 io_in[5]
port 6 nsew signal input
rlabel metal3 s 519200 22176 520000 22288 6 io_in[6]
port 7 nsew signal input
rlabel metal3 s 519200 25536 520000 25648 6 io_in[7]
port 8 nsew signal input
rlabel metal3 s 519200 4256 520000 4368 6 io_oeb[0]
port 9 nsew signal output
rlabel metal3 s 519200 7616 520000 7728 6 io_oeb[1]
port 10 nsew signal output
rlabel metal3 s 519200 10976 520000 11088 6 io_oeb[2]
port 11 nsew signal output
rlabel metal3 s 519200 14336 520000 14448 6 io_oeb[3]
port 12 nsew signal output
rlabel metal3 s 519200 17696 520000 17808 6 io_oeb[4]
port 13 nsew signal output
rlabel metal3 s 519200 21056 520000 21168 6 io_oeb[5]
port 14 nsew signal output
rlabel metal3 s 519200 24416 520000 24528 6 io_oeb[6]
port 15 nsew signal output
rlabel metal3 s 519200 27776 520000 27888 6 io_oeb[7]
port 16 nsew signal output
rlabel metal3 s 519200 3136 520000 3248 6 io_out[0]
port 17 nsew signal output
rlabel metal3 s 519200 6496 520000 6608 6 io_out[1]
port 18 nsew signal output
rlabel metal3 s 519200 9856 520000 9968 6 io_out[2]
port 19 nsew signal output
rlabel metal3 s 519200 13216 520000 13328 6 io_out[3]
port 20 nsew signal output
rlabel metal3 s 519200 16576 520000 16688 6 io_out[4]
port 21 nsew signal output
rlabel metal3 s 519200 19936 520000 20048 6 io_out[5]
port 22 nsew signal output
rlabel metal3 s 519200 23296 520000 23408 6 io_out[6]
port 23 nsew signal output
rlabel metal3 s 519200 26656 520000 26768 6 io_out[7]
port 24 nsew signal output
rlabel metal2 s 491904 0 492016 800 6 irq[0]
port 25 nsew signal output
rlabel metal2 s 493472 0 493584 800 6 irq[1]
port 26 nsew signal output
rlabel metal2 s 495040 0 495152 800 6 irq[2]
port 27 nsew signal output
rlabel metal2 s 190848 0 190960 800 6 la_data_in[0]
port 28 nsew signal input
rlabel metal2 s 237888 0 238000 800 6 la_data_in[10]
port 29 nsew signal input
rlabel metal2 s 242592 0 242704 800 6 la_data_in[11]
port 30 nsew signal input
rlabel metal2 s 247296 0 247408 800 6 la_data_in[12]
port 31 nsew signal input
rlabel metal2 s 252000 0 252112 800 6 la_data_in[13]
port 32 nsew signal input
rlabel metal2 s 256704 0 256816 800 6 la_data_in[14]
port 33 nsew signal input
rlabel metal2 s 261408 0 261520 800 6 la_data_in[15]
port 34 nsew signal input
rlabel metal2 s 266112 0 266224 800 6 la_data_in[16]
port 35 nsew signal input
rlabel metal2 s 270816 0 270928 800 6 la_data_in[17]
port 36 nsew signal input
rlabel metal2 s 275520 0 275632 800 6 la_data_in[18]
port 37 nsew signal input
rlabel metal2 s 280224 0 280336 800 6 la_data_in[19]
port 38 nsew signal input
rlabel metal2 s 195552 0 195664 800 6 la_data_in[1]
port 39 nsew signal input
rlabel metal2 s 284928 0 285040 800 6 la_data_in[20]
port 40 nsew signal input
rlabel metal2 s 289632 0 289744 800 6 la_data_in[21]
port 41 nsew signal input
rlabel metal2 s 294336 0 294448 800 6 la_data_in[22]
port 42 nsew signal input
rlabel metal2 s 299040 0 299152 800 6 la_data_in[23]
port 43 nsew signal input
rlabel metal2 s 303744 0 303856 800 6 la_data_in[24]
port 44 nsew signal input
rlabel metal2 s 308448 0 308560 800 6 la_data_in[25]
port 45 nsew signal input
rlabel metal2 s 313152 0 313264 800 6 la_data_in[26]
port 46 nsew signal input
rlabel metal2 s 317856 0 317968 800 6 la_data_in[27]
port 47 nsew signal input
rlabel metal2 s 322560 0 322672 800 6 la_data_in[28]
port 48 nsew signal input
rlabel metal2 s 327264 0 327376 800 6 la_data_in[29]
port 49 nsew signal input
rlabel metal2 s 200256 0 200368 800 6 la_data_in[2]
port 50 nsew signal input
rlabel metal2 s 331968 0 332080 800 6 la_data_in[30]
port 51 nsew signal input
rlabel metal2 s 336672 0 336784 800 6 la_data_in[31]
port 52 nsew signal input
rlabel metal2 s 341376 0 341488 800 6 la_data_in[32]
port 53 nsew signal input
rlabel metal2 s 346080 0 346192 800 6 la_data_in[33]
port 54 nsew signal input
rlabel metal2 s 350784 0 350896 800 6 la_data_in[34]
port 55 nsew signal input
rlabel metal2 s 355488 0 355600 800 6 la_data_in[35]
port 56 nsew signal input
rlabel metal2 s 360192 0 360304 800 6 la_data_in[36]
port 57 nsew signal input
rlabel metal2 s 364896 0 365008 800 6 la_data_in[37]
port 58 nsew signal input
rlabel metal2 s 369600 0 369712 800 6 la_data_in[38]
port 59 nsew signal input
rlabel metal2 s 374304 0 374416 800 6 la_data_in[39]
port 60 nsew signal input
rlabel metal2 s 204960 0 205072 800 6 la_data_in[3]
port 61 nsew signal input
rlabel metal2 s 379008 0 379120 800 6 la_data_in[40]
port 62 nsew signal input
rlabel metal2 s 383712 0 383824 800 6 la_data_in[41]
port 63 nsew signal input
rlabel metal2 s 388416 0 388528 800 6 la_data_in[42]
port 64 nsew signal input
rlabel metal2 s 393120 0 393232 800 6 la_data_in[43]
port 65 nsew signal input
rlabel metal2 s 397824 0 397936 800 6 la_data_in[44]
port 66 nsew signal input
rlabel metal2 s 402528 0 402640 800 6 la_data_in[45]
port 67 nsew signal input
rlabel metal2 s 407232 0 407344 800 6 la_data_in[46]
port 68 nsew signal input
rlabel metal2 s 411936 0 412048 800 6 la_data_in[47]
port 69 nsew signal input
rlabel metal2 s 416640 0 416752 800 6 la_data_in[48]
port 70 nsew signal input
rlabel metal2 s 421344 0 421456 800 6 la_data_in[49]
port 71 nsew signal input
rlabel metal2 s 209664 0 209776 800 6 la_data_in[4]
port 72 nsew signal input
rlabel metal2 s 426048 0 426160 800 6 la_data_in[50]
port 73 nsew signal input
rlabel metal2 s 430752 0 430864 800 6 la_data_in[51]
port 74 nsew signal input
rlabel metal2 s 435456 0 435568 800 6 la_data_in[52]
port 75 nsew signal input
rlabel metal2 s 440160 0 440272 800 6 la_data_in[53]
port 76 nsew signal input
rlabel metal2 s 444864 0 444976 800 6 la_data_in[54]
port 77 nsew signal input
rlabel metal2 s 449568 0 449680 800 6 la_data_in[55]
port 78 nsew signal input
rlabel metal2 s 454272 0 454384 800 6 la_data_in[56]
port 79 nsew signal input
rlabel metal2 s 458976 0 459088 800 6 la_data_in[57]
port 80 nsew signal input
rlabel metal2 s 463680 0 463792 800 6 la_data_in[58]
port 81 nsew signal input
rlabel metal2 s 468384 0 468496 800 6 la_data_in[59]
port 82 nsew signal input
rlabel metal2 s 214368 0 214480 800 6 la_data_in[5]
port 83 nsew signal input
rlabel metal2 s 473088 0 473200 800 6 la_data_in[60]
port 84 nsew signal input
rlabel metal2 s 477792 0 477904 800 6 la_data_in[61]
port 85 nsew signal input
rlabel metal2 s 482496 0 482608 800 6 la_data_in[62]
port 86 nsew signal input
rlabel metal2 s 487200 0 487312 800 6 la_data_in[63]
port 87 nsew signal input
rlabel metal2 s 219072 0 219184 800 6 la_data_in[6]
port 88 nsew signal input
rlabel metal2 s 223776 0 223888 800 6 la_data_in[7]
port 89 nsew signal input
rlabel metal2 s 228480 0 228592 800 6 la_data_in[8]
port 90 nsew signal input
rlabel metal2 s 233184 0 233296 800 6 la_data_in[9]
port 91 nsew signal input
rlabel metal2 s 192416 0 192528 800 6 la_data_out[0]
port 92 nsew signal output
rlabel metal2 s 239456 0 239568 800 6 la_data_out[10]
port 93 nsew signal output
rlabel metal2 s 244160 0 244272 800 6 la_data_out[11]
port 94 nsew signal output
rlabel metal2 s 248864 0 248976 800 6 la_data_out[12]
port 95 nsew signal output
rlabel metal2 s 253568 0 253680 800 6 la_data_out[13]
port 96 nsew signal output
rlabel metal2 s 258272 0 258384 800 6 la_data_out[14]
port 97 nsew signal output
rlabel metal2 s 262976 0 263088 800 6 la_data_out[15]
port 98 nsew signal output
rlabel metal2 s 267680 0 267792 800 6 la_data_out[16]
port 99 nsew signal output
rlabel metal2 s 272384 0 272496 800 6 la_data_out[17]
port 100 nsew signal output
rlabel metal2 s 277088 0 277200 800 6 la_data_out[18]
port 101 nsew signal output
rlabel metal2 s 281792 0 281904 800 6 la_data_out[19]
port 102 nsew signal output
rlabel metal2 s 197120 0 197232 800 6 la_data_out[1]
port 103 nsew signal output
rlabel metal2 s 286496 0 286608 800 6 la_data_out[20]
port 104 nsew signal output
rlabel metal2 s 291200 0 291312 800 6 la_data_out[21]
port 105 nsew signal output
rlabel metal2 s 295904 0 296016 800 6 la_data_out[22]
port 106 nsew signal output
rlabel metal2 s 300608 0 300720 800 6 la_data_out[23]
port 107 nsew signal output
rlabel metal2 s 305312 0 305424 800 6 la_data_out[24]
port 108 nsew signal output
rlabel metal2 s 310016 0 310128 800 6 la_data_out[25]
port 109 nsew signal output
rlabel metal2 s 314720 0 314832 800 6 la_data_out[26]
port 110 nsew signal output
rlabel metal2 s 319424 0 319536 800 6 la_data_out[27]
port 111 nsew signal output
rlabel metal2 s 324128 0 324240 800 6 la_data_out[28]
port 112 nsew signal output
rlabel metal2 s 328832 0 328944 800 6 la_data_out[29]
port 113 nsew signal output
rlabel metal2 s 201824 0 201936 800 6 la_data_out[2]
port 114 nsew signal output
rlabel metal2 s 333536 0 333648 800 6 la_data_out[30]
port 115 nsew signal output
rlabel metal2 s 338240 0 338352 800 6 la_data_out[31]
port 116 nsew signal output
rlabel metal2 s 342944 0 343056 800 6 la_data_out[32]
port 117 nsew signal output
rlabel metal2 s 347648 0 347760 800 6 la_data_out[33]
port 118 nsew signal output
rlabel metal2 s 352352 0 352464 800 6 la_data_out[34]
port 119 nsew signal output
rlabel metal2 s 357056 0 357168 800 6 la_data_out[35]
port 120 nsew signal output
rlabel metal2 s 361760 0 361872 800 6 la_data_out[36]
port 121 nsew signal output
rlabel metal2 s 366464 0 366576 800 6 la_data_out[37]
port 122 nsew signal output
rlabel metal2 s 371168 0 371280 800 6 la_data_out[38]
port 123 nsew signal output
rlabel metal2 s 375872 0 375984 800 6 la_data_out[39]
port 124 nsew signal output
rlabel metal2 s 206528 0 206640 800 6 la_data_out[3]
port 125 nsew signal output
rlabel metal2 s 380576 0 380688 800 6 la_data_out[40]
port 126 nsew signal output
rlabel metal2 s 385280 0 385392 800 6 la_data_out[41]
port 127 nsew signal output
rlabel metal2 s 389984 0 390096 800 6 la_data_out[42]
port 128 nsew signal output
rlabel metal2 s 394688 0 394800 800 6 la_data_out[43]
port 129 nsew signal output
rlabel metal2 s 399392 0 399504 800 6 la_data_out[44]
port 130 nsew signal output
rlabel metal2 s 404096 0 404208 800 6 la_data_out[45]
port 131 nsew signal output
rlabel metal2 s 408800 0 408912 800 6 la_data_out[46]
port 132 nsew signal output
rlabel metal2 s 413504 0 413616 800 6 la_data_out[47]
port 133 nsew signal output
rlabel metal2 s 418208 0 418320 800 6 la_data_out[48]
port 134 nsew signal output
rlabel metal2 s 422912 0 423024 800 6 la_data_out[49]
port 135 nsew signal output
rlabel metal2 s 211232 0 211344 800 6 la_data_out[4]
port 136 nsew signal output
rlabel metal2 s 427616 0 427728 800 6 la_data_out[50]
port 137 nsew signal output
rlabel metal2 s 432320 0 432432 800 6 la_data_out[51]
port 138 nsew signal output
rlabel metal2 s 437024 0 437136 800 6 la_data_out[52]
port 139 nsew signal output
rlabel metal2 s 441728 0 441840 800 6 la_data_out[53]
port 140 nsew signal output
rlabel metal2 s 446432 0 446544 800 6 la_data_out[54]
port 141 nsew signal output
rlabel metal2 s 451136 0 451248 800 6 la_data_out[55]
port 142 nsew signal output
rlabel metal2 s 455840 0 455952 800 6 la_data_out[56]
port 143 nsew signal output
rlabel metal2 s 460544 0 460656 800 6 la_data_out[57]
port 144 nsew signal output
rlabel metal2 s 465248 0 465360 800 6 la_data_out[58]
port 145 nsew signal output
rlabel metal2 s 469952 0 470064 800 6 la_data_out[59]
port 146 nsew signal output
rlabel metal2 s 215936 0 216048 800 6 la_data_out[5]
port 147 nsew signal output
rlabel metal2 s 474656 0 474768 800 6 la_data_out[60]
port 148 nsew signal output
rlabel metal2 s 479360 0 479472 800 6 la_data_out[61]
port 149 nsew signal output
rlabel metal2 s 484064 0 484176 800 6 la_data_out[62]
port 150 nsew signal output
rlabel metal2 s 488768 0 488880 800 6 la_data_out[63]
port 151 nsew signal output
rlabel metal2 s 220640 0 220752 800 6 la_data_out[6]
port 152 nsew signal output
rlabel metal2 s 225344 0 225456 800 6 la_data_out[7]
port 153 nsew signal output
rlabel metal2 s 230048 0 230160 800 6 la_data_out[8]
port 154 nsew signal output
rlabel metal2 s 234752 0 234864 800 6 la_data_out[9]
port 155 nsew signal output
rlabel metal2 s 193984 0 194096 800 6 la_oenb[0]
port 156 nsew signal input
rlabel metal2 s 241024 0 241136 800 6 la_oenb[10]
port 157 nsew signal input
rlabel metal2 s 245728 0 245840 800 6 la_oenb[11]
port 158 nsew signal input
rlabel metal2 s 250432 0 250544 800 6 la_oenb[12]
port 159 nsew signal input
rlabel metal2 s 255136 0 255248 800 6 la_oenb[13]
port 160 nsew signal input
rlabel metal2 s 259840 0 259952 800 6 la_oenb[14]
port 161 nsew signal input
rlabel metal2 s 264544 0 264656 800 6 la_oenb[15]
port 162 nsew signal input
rlabel metal2 s 269248 0 269360 800 6 la_oenb[16]
port 163 nsew signal input
rlabel metal2 s 273952 0 274064 800 6 la_oenb[17]
port 164 nsew signal input
rlabel metal2 s 278656 0 278768 800 6 la_oenb[18]
port 165 nsew signal input
rlabel metal2 s 283360 0 283472 800 6 la_oenb[19]
port 166 nsew signal input
rlabel metal2 s 198688 0 198800 800 6 la_oenb[1]
port 167 nsew signal input
rlabel metal2 s 288064 0 288176 800 6 la_oenb[20]
port 168 nsew signal input
rlabel metal2 s 292768 0 292880 800 6 la_oenb[21]
port 169 nsew signal input
rlabel metal2 s 297472 0 297584 800 6 la_oenb[22]
port 170 nsew signal input
rlabel metal2 s 302176 0 302288 800 6 la_oenb[23]
port 171 nsew signal input
rlabel metal2 s 306880 0 306992 800 6 la_oenb[24]
port 172 nsew signal input
rlabel metal2 s 311584 0 311696 800 6 la_oenb[25]
port 173 nsew signal input
rlabel metal2 s 316288 0 316400 800 6 la_oenb[26]
port 174 nsew signal input
rlabel metal2 s 320992 0 321104 800 6 la_oenb[27]
port 175 nsew signal input
rlabel metal2 s 325696 0 325808 800 6 la_oenb[28]
port 176 nsew signal input
rlabel metal2 s 330400 0 330512 800 6 la_oenb[29]
port 177 nsew signal input
rlabel metal2 s 203392 0 203504 800 6 la_oenb[2]
port 178 nsew signal input
rlabel metal2 s 335104 0 335216 800 6 la_oenb[30]
port 179 nsew signal input
rlabel metal2 s 339808 0 339920 800 6 la_oenb[31]
port 180 nsew signal input
rlabel metal2 s 344512 0 344624 800 6 la_oenb[32]
port 181 nsew signal input
rlabel metal2 s 349216 0 349328 800 6 la_oenb[33]
port 182 nsew signal input
rlabel metal2 s 353920 0 354032 800 6 la_oenb[34]
port 183 nsew signal input
rlabel metal2 s 358624 0 358736 800 6 la_oenb[35]
port 184 nsew signal input
rlabel metal2 s 363328 0 363440 800 6 la_oenb[36]
port 185 nsew signal input
rlabel metal2 s 368032 0 368144 800 6 la_oenb[37]
port 186 nsew signal input
rlabel metal2 s 372736 0 372848 800 6 la_oenb[38]
port 187 nsew signal input
rlabel metal2 s 377440 0 377552 800 6 la_oenb[39]
port 188 nsew signal input
rlabel metal2 s 208096 0 208208 800 6 la_oenb[3]
port 189 nsew signal input
rlabel metal2 s 382144 0 382256 800 6 la_oenb[40]
port 190 nsew signal input
rlabel metal2 s 386848 0 386960 800 6 la_oenb[41]
port 191 nsew signal input
rlabel metal2 s 391552 0 391664 800 6 la_oenb[42]
port 192 nsew signal input
rlabel metal2 s 396256 0 396368 800 6 la_oenb[43]
port 193 nsew signal input
rlabel metal2 s 400960 0 401072 800 6 la_oenb[44]
port 194 nsew signal input
rlabel metal2 s 405664 0 405776 800 6 la_oenb[45]
port 195 nsew signal input
rlabel metal2 s 410368 0 410480 800 6 la_oenb[46]
port 196 nsew signal input
rlabel metal2 s 415072 0 415184 800 6 la_oenb[47]
port 197 nsew signal input
rlabel metal2 s 419776 0 419888 800 6 la_oenb[48]
port 198 nsew signal input
rlabel metal2 s 424480 0 424592 800 6 la_oenb[49]
port 199 nsew signal input
rlabel metal2 s 212800 0 212912 800 6 la_oenb[4]
port 200 nsew signal input
rlabel metal2 s 429184 0 429296 800 6 la_oenb[50]
port 201 nsew signal input
rlabel metal2 s 433888 0 434000 800 6 la_oenb[51]
port 202 nsew signal input
rlabel metal2 s 438592 0 438704 800 6 la_oenb[52]
port 203 nsew signal input
rlabel metal2 s 443296 0 443408 800 6 la_oenb[53]
port 204 nsew signal input
rlabel metal2 s 448000 0 448112 800 6 la_oenb[54]
port 205 nsew signal input
rlabel metal2 s 452704 0 452816 800 6 la_oenb[55]
port 206 nsew signal input
rlabel metal2 s 457408 0 457520 800 6 la_oenb[56]
port 207 nsew signal input
rlabel metal2 s 462112 0 462224 800 6 la_oenb[57]
port 208 nsew signal input
rlabel metal2 s 466816 0 466928 800 6 la_oenb[58]
port 209 nsew signal input
rlabel metal2 s 471520 0 471632 800 6 la_oenb[59]
port 210 nsew signal input
rlabel metal2 s 217504 0 217616 800 6 la_oenb[5]
port 211 nsew signal input
rlabel metal2 s 476224 0 476336 800 6 la_oenb[60]
port 212 nsew signal input
rlabel metal2 s 480928 0 481040 800 6 la_oenb[61]
port 213 nsew signal input
rlabel metal2 s 485632 0 485744 800 6 la_oenb[62]
port 214 nsew signal input
rlabel metal2 s 490336 0 490448 800 6 la_oenb[63]
port 215 nsew signal input
rlabel metal2 s 222208 0 222320 800 6 la_oenb[6]
port 216 nsew signal input
rlabel metal2 s 226912 0 227024 800 6 la_oenb[7]
port 217 nsew signal input
rlabel metal2 s 231616 0 231728 800 6 la_oenb[8]
port 218 nsew signal input
rlabel metal2 s 236320 0 236432 800 6 la_oenb[9]
port 219 nsew signal input
rlabel metal4 s 65836 3076 66156 26716 6 vdd
port 220 nsew power bidirectional
rlabel metal4 s 195140 3076 195460 26716 6 vdd
port 220 nsew power bidirectional
rlabel metal4 s 324444 3076 324764 26716 6 vdd
port 220 nsew power bidirectional
rlabel metal4 s 453748 3076 454068 26716 6 vdd
port 220 nsew power bidirectional
rlabel metal4 s 130488 3076 130808 26716 6 vss
port 221 nsew ground bidirectional
rlabel metal4 s 259792 3076 260112 26716 6 vss
port 221 nsew ground bidirectional
rlabel metal4 s 389096 3076 389416 26716 6 vss
port 221 nsew ground bidirectional
rlabel metal4 s 518400 3076 518720 26716 6 vss
port 221 nsew ground bidirectional
rlabel metal2 s 24640 0 24752 800 6 wb_clk_i
port 222 nsew signal input
rlabel metal2 s 26208 0 26320 800 6 wb_rst_i
port 223 nsew signal input
rlabel metal2 s 27776 0 27888 800 6 wbs_ack_o
port 224 nsew signal output
rlabel metal2 s 34048 0 34160 800 6 wbs_adr_i[0]
port 225 nsew signal input
rlabel metal2 s 87360 0 87472 800 6 wbs_adr_i[10]
port 226 nsew signal input
rlabel metal2 s 92064 0 92176 800 6 wbs_adr_i[11]
port 227 nsew signal input
rlabel metal2 s 96768 0 96880 800 6 wbs_adr_i[12]
port 228 nsew signal input
rlabel metal2 s 101472 0 101584 800 6 wbs_adr_i[13]
port 229 nsew signal input
rlabel metal2 s 106176 0 106288 800 6 wbs_adr_i[14]
port 230 nsew signal input
rlabel metal2 s 110880 0 110992 800 6 wbs_adr_i[15]
port 231 nsew signal input
rlabel metal2 s 115584 0 115696 800 6 wbs_adr_i[16]
port 232 nsew signal input
rlabel metal2 s 120288 0 120400 800 6 wbs_adr_i[17]
port 233 nsew signal input
rlabel metal2 s 124992 0 125104 800 6 wbs_adr_i[18]
port 234 nsew signal input
rlabel metal2 s 129696 0 129808 800 6 wbs_adr_i[19]
port 235 nsew signal input
rlabel metal2 s 40320 0 40432 800 6 wbs_adr_i[1]
port 236 nsew signal input
rlabel metal2 s 134400 0 134512 800 6 wbs_adr_i[20]
port 237 nsew signal input
rlabel metal2 s 139104 0 139216 800 6 wbs_adr_i[21]
port 238 nsew signal input
rlabel metal2 s 143808 0 143920 800 6 wbs_adr_i[22]
port 239 nsew signal input
rlabel metal2 s 148512 0 148624 800 6 wbs_adr_i[23]
port 240 nsew signal input
rlabel metal2 s 153216 0 153328 800 6 wbs_adr_i[24]
port 241 nsew signal input
rlabel metal2 s 157920 0 158032 800 6 wbs_adr_i[25]
port 242 nsew signal input
rlabel metal2 s 162624 0 162736 800 6 wbs_adr_i[26]
port 243 nsew signal input
rlabel metal2 s 167328 0 167440 800 6 wbs_adr_i[27]
port 244 nsew signal input
rlabel metal2 s 172032 0 172144 800 6 wbs_adr_i[28]
port 245 nsew signal input
rlabel metal2 s 176736 0 176848 800 6 wbs_adr_i[29]
port 246 nsew signal input
rlabel metal2 s 46592 0 46704 800 6 wbs_adr_i[2]
port 247 nsew signal input
rlabel metal2 s 181440 0 181552 800 6 wbs_adr_i[30]
port 248 nsew signal input
rlabel metal2 s 186144 0 186256 800 6 wbs_adr_i[31]
port 249 nsew signal input
rlabel metal2 s 52864 0 52976 800 6 wbs_adr_i[3]
port 250 nsew signal input
rlabel metal2 s 59136 0 59248 800 6 wbs_adr_i[4]
port 251 nsew signal input
rlabel metal2 s 63840 0 63952 800 6 wbs_adr_i[5]
port 252 nsew signal input
rlabel metal2 s 68544 0 68656 800 6 wbs_adr_i[6]
port 253 nsew signal input
rlabel metal2 s 73248 0 73360 800 6 wbs_adr_i[7]
port 254 nsew signal input
rlabel metal2 s 77952 0 78064 800 6 wbs_adr_i[8]
port 255 nsew signal input
rlabel metal2 s 82656 0 82768 800 6 wbs_adr_i[9]
port 256 nsew signal input
rlabel metal2 s 29344 0 29456 800 6 wbs_cyc_i
port 257 nsew signal input
rlabel metal2 s 35616 0 35728 800 6 wbs_dat_i[0]
port 258 nsew signal input
rlabel metal2 s 88928 0 89040 800 6 wbs_dat_i[10]
port 259 nsew signal input
rlabel metal2 s 93632 0 93744 800 6 wbs_dat_i[11]
port 260 nsew signal input
rlabel metal2 s 98336 0 98448 800 6 wbs_dat_i[12]
port 261 nsew signal input
rlabel metal2 s 103040 0 103152 800 6 wbs_dat_i[13]
port 262 nsew signal input
rlabel metal2 s 107744 0 107856 800 6 wbs_dat_i[14]
port 263 nsew signal input
rlabel metal2 s 112448 0 112560 800 6 wbs_dat_i[15]
port 264 nsew signal input
rlabel metal2 s 117152 0 117264 800 6 wbs_dat_i[16]
port 265 nsew signal input
rlabel metal2 s 121856 0 121968 800 6 wbs_dat_i[17]
port 266 nsew signal input
rlabel metal2 s 126560 0 126672 800 6 wbs_dat_i[18]
port 267 nsew signal input
rlabel metal2 s 131264 0 131376 800 6 wbs_dat_i[19]
port 268 nsew signal input
rlabel metal2 s 41888 0 42000 800 6 wbs_dat_i[1]
port 269 nsew signal input
rlabel metal2 s 135968 0 136080 800 6 wbs_dat_i[20]
port 270 nsew signal input
rlabel metal2 s 140672 0 140784 800 6 wbs_dat_i[21]
port 271 nsew signal input
rlabel metal2 s 145376 0 145488 800 6 wbs_dat_i[22]
port 272 nsew signal input
rlabel metal2 s 150080 0 150192 800 6 wbs_dat_i[23]
port 273 nsew signal input
rlabel metal2 s 154784 0 154896 800 6 wbs_dat_i[24]
port 274 nsew signal input
rlabel metal2 s 159488 0 159600 800 6 wbs_dat_i[25]
port 275 nsew signal input
rlabel metal2 s 164192 0 164304 800 6 wbs_dat_i[26]
port 276 nsew signal input
rlabel metal2 s 168896 0 169008 800 6 wbs_dat_i[27]
port 277 nsew signal input
rlabel metal2 s 173600 0 173712 800 6 wbs_dat_i[28]
port 278 nsew signal input
rlabel metal2 s 178304 0 178416 800 6 wbs_dat_i[29]
port 279 nsew signal input
rlabel metal2 s 48160 0 48272 800 6 wbs_dat_i[2]
port 280 nsew signal input
rlabel metal2 s 183008 0 183120 800 6 wbs_dat_i[30]
port 281 nsew signal input
rlabel metal2 s 187712 0 187824 800 6 wbs_dat_i[31]
port 282 nsew signal input
rlabel metal2 s 54432 0 54544 800 6 wbs_dat_i[3]
port 283 nsew signal input
rlabel metal2 s 60704 0 60816 800 6 wbs_dat_i[4]
port 284 nsew signal input
rlabel metal2 s 65408 0 65520 800 6 wbs_dat_i[5]
port 285 nsew signal input
rlabel metal2 s 70112 0 70224 800 6 wbs_dat_i[6]
port 286 nsew signal input
rlabel metal2 s 74816 0 74928 800 6 wbs_dat_i[7]
port 287 nsew signal input
rlabel metal2 s 79520 0 79632 800 6 wbs_dat_i[8]
port 288 nsew signal input
rlabel metal2 s 84224 0 84336 800 6 wbs_dat_i[9]
port 289 nsew signal input
rlabel metal2 s 37184 0 37296 800 6 wbs_dat_o[0]
port 290 nsew signal output
rlabel metal2 s 90496 0 90608 800 6 wbs_dat_o[10]
port 291 nsew signal output
rlabel metal2 s 95200 0 95312 800 6 wbs_dat_o[11]
port 292 nsew signal output
rlabel metal2 s 99904 0 100016 800 6 wbs_dat_o[12]
port 293 nsew signal output
rlabel metal2 s 104608 0 104720 800 6 wbs_dat_o[13]
port 294 nsew signal output
rlabel metal2 s 109312 0 109424 800 6 wbs_dat_o[14]
port 295 nsew signal output
rlabel metal2 s 114016 0 114128 800 6 wbs_dat_o[15]
port 296 nsew signal output
rlabel metal2 s 118720 0 118832 800 6 wbs_dat_o[16]
port 297 nsew signal output
rlabel metal2 s 123424 0 123536 800 6 wbs_dat_o[17]
port 298 nsew signal output
rlabel metal2 s 128128 0 128240 800 6 wbs_dat_o[18]
port 299 nsew signal output
rlabel metal2 s 132832 0 132944 800 6 wbs_dat_o[19]
port 300 nsew signal output
rlabel metal2 s 43456 0 43568 800 6 wbs_dat_o[1]
port 301 nsew signal output
rlabel metal2 s 137536 0 137648 800 6 wbs_dat_o[20]
port 302 nsew signal output
rlabel metal2 s 142240 0 142352 800 6 wbs_dat_o[21]
port 303 nsew signal output
rlabel metal2 s 146944 0 147056 800 6 wbs_dat_o[22]
port 304 nsew signal output
rlabel metal2 s 151648 0 151760 800 6 wbs_dat_o[23]
port 305 nsew signal output
rlabel metal2 s 156352 0 156464 800 6 wbs_dat_o[24]
port 306 nsew signal output
rlabel metal2 s 161056 0 161168 800 6 wbs_dat_o[25]
port 307 nsew signal output
rlabel metal2 s 165760 0 165872 800 6 wbs_dat_o[26]
port 308 nsew signal output
rlabel metal2 s 170464 0 170576 800 6 wbs_dat_o[27]
port 309 nsew signal output
rlabel metal2 s 175168 0 175280 800 6 wbs_dat_o[28]
port 310 nsew signal output
rlabel metal2 s 179872 0 179984 800 6 wbs_dat_o[29]
port 311 nsew signal output
rlabel metal2 s 49728 0 49840 800 6 wbs_dat_o[2]
port 312 nsew signal output
rlabel metal2 s 184576 0 184688 800 6 wbs_dat_o[30]
port 313 nsew signal output
rlabel metal2 s 189280 0 189392 800 6 wbs_dat_o[31]
port 314 nsew signal output
rlabel metal2 s 56000 0 56112 800 6 wbs_dat_o[3]
port 315 nsew signal output
rlabel metal2 s 62272 0 62384 800 6 wbs_dat_o[4]
port 316 nsew signal output
rlabel metal2 s 66976 0 67088 800 6 wbs_dat_o[5]
port 317 nsew signal output
rlabel metal2 s 71680 0 71792 800 6 wbs_dat_o[6]
port 318 nsew signal output
rlabel metal2 s 76384 0 76496 800 6 wbs_dat_o[7]
port 319 nsew signal output
rlabel metal2 s 81088 0 81200 800 6 wbs_dat_o[8]
port 320 nsew signal output
rlabel metal2 s 85792 0 85904 800 6 wbs_dat_o[9]
port 321 nsew signal output
rlabel metal2 s 38752 0 38864 800 6 wbs_sel_i[0]
port 322 nsew signal input
rlabel metal2 s 45024 0 45136 800 6 wbs_sel_i[1]
port 323 nsew signal input
rlabel metal2 s 51296 0 51408 800 6 wbs_sel_i[2]
port 324 nsew signal input
rlabel metal2 s 57568 0 57680 800 6 wbs_sel_i[3]
port 325 nsew signal input
rlabel metal2 s 30912 0 31024 800 6 wbs_stb_i
port 326 nsew signal input
rlabel metal2 s 32480 0 32592 800 6 wbs_we_i
port 327 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 520000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1346638
string GDS_FILE /home/luke/picosoc-w-approximation/openlane/user_proj_example/runs/23_12_10_12_01/results/signoff/user_proj_example.magic.gds
string GDS_START 187076
<< end >>

